library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"B0",X"4F",X"ED",X"56",X"C3",X"81",X"00",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",
		X"0F",X"0F",X"0F",X"0F",X"C9",X"DF",X"DF",X"DF",X"E1",X"D1",X"C1",X"00",X"00",X"C7",X"DF",X"DF",
		X"E1",X"07",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"EB",X"E9",X"DF",X"DF",X"DF",
		X"E1",X"22",X"5A",X"4C",X"C9",X"DF",X"DF",X"DF",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"D9",X"C5",X"D5",X"E5",X"08",X"F5",X"21",X"01",X"50",X"36",X"00",X"32",X"C0",X"50",X"2E",X"07",
		X"36",X"01",X"CD",X"4D",X"06",X"CD",X"63",X"05",X"CD",X"60",X"04",X"CD",X"E8",X"03",X"CD",X"00",
		X"20",X"CD",X"F2",X"05",X"CD",X"E0",X"03",X"3E",X"FF",X"32",X"22",X"4C",X"21",X"01",X"50",X"36",
		X"01",X"F1",X"08",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"FB",
		X"C9",X"21",X"07",X"50",X"36",X"00",X"2B",X"7C",X"FE",X"3F",X"32",X"C0",X"50",X"20",X"F5",X"16",
		X"00",X"D9",X"21",X"00",X"40",X"36",X"00",X"23",X"7C",X"32",X"C0",X"50",X"FE",X"51",X"20",X"F5",
		X"21",X"00",X"40",X"55",X"5D",X"DD",X"21",X"AC",X"00",X"C3",X"0B",X"01",X"21",X"00",X"44",X"DD",
		X"21",X"B6",X"00",X"C3",X"0B",X"01",X"21",X"00",X"4C",X"DD",X"21",X"C0",X"00",X"C3",X"0B",X"01",
		X"21",X"00",X"40",X"36",X"40",X"23",X"7C",X"FE",X"44",X"20",X"F8",X"36",X"03",X"23",X"7C",X"FE",
		X"48",X"20",X"F8",X"7A",X"B3",X"CA",X"67",X"01",X"01",X"E0",X"FF",X"21",X"A6",X"42",X"36",X"42",
		X"09",X"36",X"41",X"09",X"36",X"44",X"09",X"36",X"40",X"09",X"36",X"52",X"09",X"36",X"41",X"09",
		X"36",X"4D",X"09",X"36",X"40",X"DD",X"21",X"FC",X"00",X"C3",X"4A",X"01",X"09",X"41",X"DD",X"21",
		X"05",X"01",X"C3",X"4A",X"01",X"16",X"FF",X"D9",X"C3",X"67",X"01",X"7E",X"B7",X"FD",X"21",X"13",
		X"01",X"20",X"2E",X"3E",X"01",X"47",X"77",X"AE",X"FD",X"21",X"1E",X"01",X"20",X"23",X"78",X"37",
		X"8F",X"32",X"C0",X"50",X"30",X"EF",X"23",X"7D",X"06",X"4F",X"32",X"07",X"50",X"10",X"FB",X"B7",
		X"20",X"D9",X"7C",X"FE",X"44",X"28",X"08",X"FE",X"48",X"28",X"04",X"FE",X"50",X"20",X"CC",X"DD",
		X"E9",X"B3",X"5F",X"7A",X"B7",X"20",X"01",X"54",X"FD",X"E9",X"09",X"7A",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"37",X"77",X"09",X"7A",X"E6",X"0F",X"FE",X"0A",X"38",
		X"02",X"C6",X"37",X"77",X"09",X"DD",X"E9",X"21",X"00",X"00",X"11",X"08",X"01",X"01",X"00",X"08",
		X"3E",X"FF",X"AE",X"32",X"07",X"50",X"32",X"C0",X"50",X"23",X"0D",X"20",X"F5",X"10",X"F3",X"B7",
		X"FD",X"21",X"86",X"01",X"00",X"00",X"14",X"1D",X"20",X"E3",X"CB",X"7A",X"20",X"08",X"D9",X"7A",
		X"B7",X"20",X"03",X"C3",X"22",X"02",X"21",X"00",X"20",X"10",X"FE",X"32",X"C0",X"50",X"2D",X"20",
		X"F8",X"D9",X"21",X"BA",X"42",X"01",X"E0",X"FF",X"36",X"44",X"09",X"36",X"49",X"09",X"36",X"50",
		X"09",X"09",X"36",X"53",X"09",X"36",X"57",X"09",X"3A",X"00",X"50",X"57",X"DD",X"21",X"C3",X"01",
		X"C3",X"4A",X"01",X"3A",X"40",X"50",X"57",X"DD",X"21",X"CD",X"01",X"18",X"F3",X"3A",X"80",X"50",
		X"57",X"DD",X"21",X"D7",X"01",X"18",X"E9",X"D9",X"25",X"20",X"BE",X"C7",X"25",X"20",X"BA",X"C7",
		X"08",X"7A",X"87",X"CB",X"FA",X"E6",X"3F",X"D9",X"21",X"A8",X"42",X"85",X"6F",X"30",X"01",X"24",
		X"01",X"E0",X"FF",X"36",X"42",X"09",X"36",X"41",X"09",X"36",X"44",X"09",X"09",X"36",X"50",X"09",
		X"36",X"52",X"09",X"36",X"4F",X"09",X"36",X"4D",X"09",X"D9",X"7A",X"D9",X"E6",X"0F",X"57",X"DD",
		X"21",X"16",X"02",X"C3",X"4A",X"01",X"08",X"57",X"DD",X"21",X"1F",X"02",X"C3",X"4A",X"01",X"D9",
		X"FD",X"E9",X"18",X"16",X"C3",X"B6",X"02",X"C3",X"80",X"03",X"C3",X"B3",X"03",X"C3",X"C6",X"03",
		X"C3",X"CB",X"03",X"C3",X"D8",X"05",X"6D",X"06",X"8D",X"06",X"21",X"00",X"4C",X"36",X"00",X"11",
		X"01",X"4C",X"01",X"FF",X"03",X"ED",X"B0",X"CD",X"80",X"03",X"3A",X"00",X"50",X"32",X"12",X"4C",
		X"3A",X"C0",X"50",X"A7",X"20",X"02",X"3E",X"FF",X"32",X"13",X"4C",X"FB",X"3E",X"01",X"32",X"01",
		X"50",X"3A",X"00",X"50",X"CB",X"67",X"C2",X"0C",X"07",X"CD",X"C6",X"03",X"A4",X"42",X"41",X"44",
		X"44",X"52",X"45",X"53",X"53",X"20",X"20",X"44",X"41",X"54",X"41",X"24",X"CD",X"C6",X"03",X"66",
		X"42",X"30",X"30",X"30",X"30",X"24",X"11",X"00",X"00",X"0E",X"00",X"CD",X"33",X"03",X"3A",X"00",
		X"50",X"CB",X"47",X"28",X"41",X"CB",X"5F",X"28",X"41",X"CB",X"4F",X"28",X"70",X"CB",X"57",X"28",
		X"7C",X"3A",X"40",X"50",X"CB",X"6F",X"28",X"1C",X"CB",X"77",X"28",X"1E",X"06",X"14",X"CD",X"B6",
		X"02",X"10",X"FB",X"C3",X"8E",X"02",X"AF",X"32",X"22",X"4C",X"3A",X"22",X"4C",X"B7",X"32",X"C0",
		X"50",X"28",X"F7",X"C9",X"3A",X"FF",X"4F",X"12",X"18",X"E2",X"C5",X"D5",X"21",X"D2",X"02",X"E5",
		X"D5",X"C9",X"D1",X"C1",X"18",X"D6",X"06",X"01",X"18",X"02",X"06",X"FF",X"CB",X"59",X"20",X"1F",
		X"CB",X"49",X"20",X"09",X"7A",X"CD",X"51",X"03",X"57",X"2E",X"66",X"18",X"07",X"7B",X"CD",X"51",
		X"03",X"5F",X"2E",X"26",X"26",X"42",X"CD",X"64",X"03",X"ED",X"53",X"F0",X"4F",X"18",X"A2",X"3A",
		X"FF",X"4F",X"CD",X"51",X"03",X"32",X"FF",X"4F",X"CD",X"66",X"06",X"18",X"94",X"0D",X"F2",X"15",
		X"03",X"0E",X"09",X"18",X"18",X"CB",X"51",X"28",X"14",X"0E",X"03",X"18",X"10",X"0C",X"CB",X"51",
		X"28",X"04",X"0E",X"08",X"18",X"07",X"79",X"FE",X"0A",X"38",X"02",X"0E",X"00",X"CD",X"33",X"03",
		X"C3",X"A1",X"02",X"C5",X"D5",X"79",X"32",X"FE",X"4F",X"0C",X"21",X"47",X"41",X"11",X"20",X"00",
		X"06",X"0A",X"79",X"B8",X"3E",X"FF",X"28",X"02",X"3E",X"20",X"77",X"19",X"10",X"F4",X"D1",X"C1",
		X"C9",X"CB",X"41",X"20",X"01",X"D7",X"F5",X"80",X"E6",X"0F",X"47",X"F1",X"E6",X"F0",X"B0",X"CB",
		X"41",X"C0",X"D7",X"C9",X"C5",X"47",X"D7",X"CD",X"74",X"03",X"78",X"01",X"E0",X"FF",X"09",X"CD",
		X"74",X"03",X"C1",X"C9",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"77",X"C9",
		X"AF",X"32",X"00",X"50",X"CD",X"B3",X"03",X"00",X"80",X"50",X"30",X"01",X"CD",X"B3",X"03",X"00",
		X"D0",X"4F",X"30",X"01",X"CD",X"B3",X"03",X"FC",X"00",X"40",X"00",X"04",X"CD",X"B3",X"03",X"03",
		X"00",X"44",X"00",X"04",X"21",X"01",X"4C",X"CB",X"86",X"21",X"00",X"00",X"22",X"06",X"4D",X"22",
		X"08",X"4D",X"C9",X"E1",X"7E",X"23",X"5E",X"23",X"56",X"23",X"46",X"23",X"4E",X"12",X"13",X"10",
		X"FC",X"0D",X"20",X"F9",X"23",X"E9",X"01",X"E0",X"FF",X"18",X"03",X"01",X"FF",X"FF",X"E1",X"5E",
		X"23",X"56",X"23",X"EB",X"1A",X"13",X"FE",X"24",X"28",X"04",X"77",X"09",X"18",X"F6",X"EB",X"E9",
		X"21",X"10",X"4C",X"34",X"C0",X"23",X"34",X"C9",X"3A",X"01",X"4C",X"0F",X"D0",X"3A",X"16",X"4C",
		X"0E",X"1F",X"FE",X"06",X"30",X"07",X"0E",X"0F",X"3D",X"20",X"02",X"0E",X"07",X"3A",X"10",X"4C",
		X"A1",X"C0",X"2A",X"48",X"4C",X"5E",X"23",X"7E",X"23",X"A7",X"28",X"3A",X"57",X"1A",X"FE",X"F0",
		X"30",X"F3",X"EE",X"01",X"12",X"3A",X"16",X"4C",X"A7",X"28",X"EA",X"FE",X"06",X"30",X"E6",X"E5",
		X"21",X"00",X"04",X"19",X"7E",X"FE",X"0F",X"28",X"08",X"FE",X"15",X"20",X"08",X"36",X"0F",X"18",
		X"12",X"36",X"15",X"18",X"0E",X"FE",X"16",X"28",X"08",X"FE",X"14",X"20",X"06",X"36",X"16",X"18",
		X"02",X"36",X"14",X"E1",X"18",X"BF",X"2A",X"06",X"4D",X"7C",X"A7",X"C8",X"0E",X"2E",X"CD",X"56",
		X"04",X"2A",X"08",X"4D",X"0E",X"03",X"7E",X"FE",X"FC",X"79",X"28",X"02",X"3E",X"FC",X"77",X"C9",
		X"3A",X"1D",X"4C",X"A7",X"C8",X"3A",X"00",X"4C",X"FE",X"50",X"D0",X"E6",X"F0",X"FE",X"40",X"CA",
		X"FA",X"04",X"CD",X"80",X"03",X"AF",X"32",X"04",X"50",X"CD",X"03",X"07",X"4C",X"44",X"1C",X"02",
		X"CD",X"03",X"07",X"51",X"44",X"1C",X"07",X"CD",X"03",X"07",X"58",X"44",X"1C",X"05",X"CD",X"B3",
		X"03",X"00",X"23",X"4C",X"06",X"01",X"CD",X"00",X"07",X"06",X"CD",X"C6",X"03",X"0C",X"43",X"50",
		X"55",X"53",X"48",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"2E",X"24",X"21",X"86",X"90",X"22",X"E6",X"4F",X"21",X"88",X"13",X"22",X"D6",X"4F",X"CD",X"C6",
		X"03",X"98",X"43",X"41",X"44",X"44",X"49",X"54",X"49",X"4F",X"4E",X"41",X"4C",X"20",X"2A",X"2A",
		X"20",X"41",X"54",X"20",X"31",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"2E",X"24",X"21",
		X"60",X"62",X"22",X"17",X"42",X"21",X"66",X"64",X"22",X"37",X"42",X"21",X"02",X"02",X"22",X"17",
		X"46",X"22",X"37",X"46",X"21",X"40",X"00",X"22",X"00",X"4C",X"3A",X"10",X"4C",X"E6",X"0F",X"20",
		X"07",X"21",X"D6",X"4F",X"7E",X"EE",X"04",X"77",X"3A",X"1D",X"4C",X"3D",X"20",X"18",X"CD",X"C6",
		X"03",X"D1",X"42",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"4C",X"59",
		X"24",X"3A",X"40",X"50",X"18",X"25",X"CD",X"C6",X"03",X"D1",X"42",X"31",X"20",X"4F",X"52",X"20",
		X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"24",X"3A",X"40",X"50",X"CB",X"77",X"20",
		X"0A",X"3A",X"1D",X"4C",X"D6",X"02",X"11",X"50",X"80",X"18",X"0B",X"E6",X"20",X"C0",X"3A",X"1D",
		X"4C",X"D6",X"01",X"11",X"50",X"00",X"27",X"32",X"1D",X"4C",X"ED",X"53",X"00",X"4C",X"CD",X"06",
		X"07",X"18",X"75",X"3A",X"80",X"50",X"E6",X"03",X"20",X"07",X"3E",X"99",X"32",X"1D",X"4C",X"18",
		X"67",X"3A",X"00",X"50",X"CB",X"77",X"21",X"1F",X"4C",X"CD",X"8F",X"05",X"3A",X"00",X"50",X"CB",
		X"6F",X"21",X"1E",X"4C",X"CD",X"8F",X"05",X"3A",X"00",X"50",X"CB",X"7F",X"21",X"1E",X"4C",X"7E",
		X"28",X"05",X"E6",X"0F",X"C8",X"35",X"C9",X"E6",X"0F",X"CB",X"D6",X"CB",X"8E",X"C0",X"3A",X"80",
		X"50",X"E6",X"03",X"47",X"3A",X"1D",X"4C",X"05",X"28",X"18",X"05",X"20",X"03",X"3C",X"18",X"12",
		X"7E",X"C6",X"80",X"77",X"21",X"33",X"40",X"38",X"04",X"36",X"25",X"18",X"0F",X"36",X"20",X"3A",
		X"1D",X"4C",X"C6",X"01",X"27",X"30",X"02",X"3E",X"99",X"32",X"1D",X"4C",X"3A",X"00",X"4C",X"FE",
		X"50",X"30",X"05",X"3E",X"01",X"32",X"4A",X"4C",X"11",X"1D",X"4C",X"1A",X"21",X"34",X"40",X"E6",
		X"0F",X"C6",X"30",X"77",X"1A",X"D7",X"23",X"E6",X"0F",X"28",X"04",X"C6",X"30",X"77",X"C9",X"36",
		X"20",X"C9",X"3A",X"01",X"4C",X"E6",X"20",X"20",X"17",X"21",X"D2",X"4F",X"11",X"F2",X"4F",X"01",
		X"0C",X"00",X"ED",X"B0",X"21",X"E2",X"4F",X"11",X"A2",X"50",X"01",X"0C",X"00",X"ED",X"B0",X"C9",
		X"DD",X"21",X"D2",X"4F",X"FD",X"21",X"33",X"50",X"01",X"02",X"06",X"26",X"0C",X"11",X"02",X"00",
		X"DD",X"7E",X"00",X"EE",X"03",X"FD",X"77",X"BF",X"DD",X"7E",X"01",X"FD",X"77",X"C0",X"DD",X"7E",
		X"10",X"ED",X"44",X"84",X"FD",X"77",X"6F",X"DD",X"7E",X"11",X"ED",X"44",X"C6",X"10",X"FD",X"77",
		X"70",X"0D",X"20",X"02",X"26",X"0E",X"DD",X"19",X"FD",X"19",X"10",X"D4",X"C9",X"3A",X"00",X"50",
		X"CB",X"67",X"C0",X"3A",X"FE",X"4F",X"CB",X"5F",X"28",X"05",X"3A",X"FF",X"4F",X"18",X"07",X"2A",
		X"F0",X"4F",X"7E",X"32",X"FF",X"4F",X"21",X"66",X"41",X"CD",X"64",X"03",X"C9",X"ED",X"41",X"EE",
		X"41",X"0D",X"42",X"0E",X"42",X"DF",X"40",X"BF",X"40",X"5F",X"41",X"3F",X"41",X"DF",X"42",X"BF",
		X"42",X"5F",X"43",X"3F",X"43",X"BF",X"41",X"DF",X"41",X"3F",X"42",X"5F",X"42",X"82",X"40",X"83",
		X"40",X"93",X"40",X"94",X"40",X"A5",X"40",X"C5",X"40",X"A8",X"40",X"A9",X"40",X"B6",X"40",X"D6",
		X"40",X"CC",X"40",X"EC",X"40",X"0A",X"41",X"2A",X"41",X"26",X"41",X"27",X"41",X"41",X"41",X"42",
		X"41",X"C3",X"41",X"C4",X"41",X"E1",X"41",X"01",X"42",X"C3",X"42",X"E3",X"42",X"41",X"43",X"42",
		X"43",X"05",X"43",X"25",X"43",X"C7",X"42",X"C8",X"42",X"49",X"43",X"4A",X"43",X"0D",X"43",X"2D",
		X"43",X"73",X"43",X"74",X"43",X"36",X"43",X"56",X"43",X"B4",X"41",X"B5",X"41",X"77",X"41",X"97",
		X"41",X"55",X"42",X"56",X"42",X"78",X"42",X"98",X"42",X"00",X"00",X"72",X"CB",X"68",X"3E",X"DC",
		X"28",X"02",X"3E",X"78",X"77",X"18",X"67",X"18",X"71",X"CD",X"52",X"1D",X"CD",X"60",X"2D",X"CD",
		X"C3",X"44",X"0A",X"C3",X"3F",X"0F",X"C3",X"1C",X"0A",X"C3",X"7D",X"09",X"C3",X"12",X"07",X"C3",
		X"86",X"0E",X"3A",X"80",X"50",X"0F",X"0F",X"E6",X"03",X"3C",X"32",X"1A",X"4C",X"21",X"80",X"50",
		X"CB",X"6E",X"28",X"11",X"11",X"29",X"4C",X"06",X"05",X"C5",X"21",X"3C",X"07",X"01",X"06",X"00",
		X"ED",X"B0",X"C1",X"10",X"F4",X"3E",X"01",X"32",X"03",X"50",X"18",X"06",X"00",X"05",X"00",X"4D",
		X"54",X"50",X"3A",X"00",X"4C",X"D7",X"E6",X"0F",X"28",X"0C",X"CB",X"57",X"20",X"12",X"3D",X"20",
		X"0A",X"CD",X"7A",X"07",X"18",X"1F",X"CD",X"0C",X"27",X"18",X"1A",X"CD",X"0F",X"27",X"18",X"15",
		X"E6",X"03",X"28",X"05",X"CD",X"7A",X"07",X"18",X"0C",X"21",X"00",X"4C",X"CB",X"5E",X"20",X"05",
		X"CB",X"DE",X"CD",X"C6",X"0A",X"CD",X"24",X"02",X"18",X"C8",X"3A",X"01",X"4C",X"0F",X"DA",X"0B",
		X"08",X"21",X"00",X"4C",X"CB",X"76",X"20",X"05",X"CD",X"06",X"07",X"18",X"70",X"CD",X"27",X"02",
		X"CD",X"C6",X"0A",X"21",X"01",X"4C",X"CB",X"AE",X"11",X"78",X"4C",X"3E",X"31",X"CB",X"76",X"28",
		X"11",X"3A",X"80",X"50",X"E6",X"10",X"28",X"07",X"CB",X"EE",X"3E",X"01",X"32",X"00",X"50",X"3E",
		X"32",X"13",X"32",X"8B",X"41",X"1A",X"A7",X"20",X"04",X"CB",X"9E",X"18",X"02",X"CB",X"DE",X"CD",
		X"29",X"0B",X"CD",X"2D",X"02",X"6B",X"42",X"50",X"4C",X"41",X"59",X"45",X"52",X"24",X"CD",X"2D",
		X"02",X"2E",X"42",X"52",X"45",X"41",X"44",X"59",X"24",X"21",X"01",X"4C",X"CB",X"7E",X"20",X"0C",
		X"AF",X"21",X"C5",X"47",X"77",X"23",X"77",X"23",X"77",X"32",X"E3",X"47",X"06",X"64",X"CD",X"24",
		X"02",X"10",X"FB",X"3E",X"02",X"32",X"4C",X"4C",X"3E",X"09",X"32",X"4A",X"4C",X"CD",X"CB",X"0B",
		X"2A",X"36",X"02",X"22",X"48",X"4C",X"21",X"01",X"4C",X"CB",X"C6",X"3A",X"00",X"4C",X"E6",X"07",
		X"E7",X"21",X"08",X"AE",X"08",X"B6",X"08",X"03",X"09",X"4C",X"09",X"51",X"09",X"56",X"09",X"06",
		X"27",X"21",X"00",X"05",X"22",X"18",X"4C",X"3A",X"80",X"50",X"CB",X"6F",X"20",X"05",X"3E",X"01",
		X"32",X"16",X"4C",X"AF",X"32",X"20",X"4C",X"21",X"1B",X"4C",X"3A",X"01",X"4C",X"E6",X"40",X"28",
		X"01",X"23",X"35",X"21",X"01",X"4C",X"28",X"04",X"CB",X"A6",X"18",X"02",X"CB",X"E6",X"CD",X"7D",
		X"09",X"3A",X"7A",X"4C",X"A7",X"4F",X"28",X"0C",X"E6",X"E0",X"3E",X"06",X"20",X"06",X"79",X"0F",
		X"0F",X"E6",X"07",X"3C",X"4F",X"5F",X"16",X"00",X"21",X"84",X"08",X"19",X"7E",X"32",X"14",X"4C",
		X"79",X"07",X"07",X"81",X"5F",X"21",X"8B",X"08",X"19",X"11",X"7B",X"4C",X"01",X"05",X"00",X"ED",
		X"B0",X"C3",X"58",X"09",X"00",X"02",X"00",X"05",X"02",X"84",X"FF",X"05",X"09",X"07",X"10",X"15",
		X"07",X"12",X"09",X"13",X"20",X"09",X"16",X"13",X"18",X"27",X"12",X"22",X"17",X"24",X"36",X"15",
		X"27",X"21",X"30",X"45",X"20",X"36",X"28",X"40",X"60",X"25",X"45",X"35",X"50",X"75",X"CD",X"B4",
		X"09",X"CD",X"00",X"10",X"18",X"30",X"3A",X"7A",X"4C",X"E6",X"FC",X"28",X"06",X"CD",X"0C",X"10",
		X"CD",X"06",X"10",X"CD",X"0C",X"10",X"CD",X"06",X"10",X"3A",X"14",X"4C",X"4F",X"A7",X"28",X"19",
		X"21",X"15",X"4C",X"07",X"79",X"30",X"08",X"35",X"20",X"09",X"E6",X"7F",X"77",X"18",X"0A",X"35",
		X"20",X"07",X"77",X"CD",X"0C",X"10",X"CD",X"06",X"10",X"21",X"20",X"4C",X"7E",X"A7",X"28",X"6C",
		X"35",X"20",X"69",X"CD",X"03",X"07",X"AA",X"41",X"07",X"FB",X"CD",X"03",X"07",X"AA",X"45",X"07",
		X"1C",X"18",X"59",X"21",X"00",X"4C",X"CB",X"5E",X"20",X"08",X"CB",X"DE",X"21",X"00",X"00",X"22",
		X"10",X"4C",X"3A",X"10",X"4C",X"47",X"E6",X"0F",X"20",X"42",X"CB",X"60",X"28",X"14",X"CD",X"C9",
		X"0E",X"CD",X"B3",X"0B",X"3A",X"10",X"4C",X"FE",X"80",X"38",X"31",X"21",X"00",X"4C",X"CB",X"9E",
		X"18",X"26",X"3E",X"0C",X"32",X"4A",X"4C",X"CD",X"2A",X"02",X"03",X"40",X"44",X"80",X"04",X"21",
		X"D3",X"4F",X"01",X"03",X"06",X"71",X"23",X"23",X"10",X"FB",X"18",X"10",X"CD",X"00",X"27",X"18",
		X"0B",X"CD",X"03",X"27",X"18",X"06",X"18",X"00",X"21",X"00",X"4C",X"34",X"3A",X"00",X"4C",X"CB",
		X"77",X"C8",X"3A",X"10",X"4C",X"E6",X"0F",X"C0",X"3A",X"01",X"4C",X"21",X"C5",X"47",X"CB",X"77",
		X"20",X"02",X"2E",X"D8",X"7E",X"EE",X"03",X"77",X"23",X"77",X"23",X"77",X"C9",X"11",X"1B",X"4C",
		X"3A",X"01",X"4C",X"CB",X"77",X"28",X"01",X"13",X"21",X"90",X"91",X"01",X"93",X"92",X"1A",X"A7",
		X"C8",X"22",X"CF",X"41",X"ED",X"43",X"EF",X"41",X"3D",X"C8",X"22",X"0F",X"42",X"ED",X"43",X"2F",
		X"42",X"3D",X"C8",X"22",X"8F",X"41",X"ED",X"43",X"AF",X"41",X"3D",X"C8",X"22",X"4F",X"42",X"ED",
		X"43",X"6F",X"42",X"C9",X"21",X"00",X"4C",X"CB",X"5E",X"20",X"1B",X"CB",X"DE",X"3E",X"03",X"32",
		X"18",X"4C",X"21",X"00",X"00",X"22",X"10",X"4C",X"21",X"86",X"98",X"01",X"04",X"02",X"22",X"E4",
		X"4F",X"ED",X"43",X"D4",X"4F",X"C9",X"3A",X"10",X"4C",X"E6",X"0F",X"C0",X"21",X"D4",X"4F",X"7E",
		X"FE",X"20",X"28",X"04",X"C6",X"04",X"77",X"C9",X"D6",X"04",X"77",X"21",X"18",X"4C",X"35",X"C0",
		X"21",X"00",X"00",X"22",X"E4",X"4F",X"22",X"D4",X"4F",X"21",X"60",X"62",X"22",X"ED",X"41",X"21",
		X"66",X"64",X"22",X"0D",X"42",X"21",X"00",X"4C",X"7E",X"E6",X"F0",X"F6",X"02",X"77",X"3E",X"03",
		X"32",X"08",X"4C",X"3E",X"01",X"32",X"0D",X"4C",X"32",X"04",X"4C",X"C9",X"3A",X"1A",X"4C",X"67",
		X"6F",X"22",X"1B",X"4C",X"21",X"00",X"00",X"22",X"78",X"4C",X"AF",X"32",X"7A",X"4C",X"21",X"29",
		X"4C",X"11",X"03",X"4D",X"01",X"03",X"00",X"ED",X"B0",X"21",X"0A",X"4D",X"06",X"08",X"36",X"00",
		X"23",X"10",X"FB",X"C9",X"E1",X"7E",X"23",X"E5",X"06",X"1C",X"21",X"43",X"44",X"11",X"20",X"00",
		X"E5",X"C5",X"06",X"07",X"77",X"23",X"10",X"FC",X"C1",X"E1",X"19",X"10",X"F3",X"CD",X"2D",X"02",
		X"E3",X"42",X"10",X"FF",X"FF",X"11",X"12",X"24",X"CD",X"2D",X"02",X"C4",X"42",X"13",X"18",X"19",
		X"1A",X"24",X"CD",X"2D",X"02",X"E5",X"42",X"1B",X"1C",X"FF",X"FF",X"1E",X"03",X"20",X"20",X"20",
		X"20",X"1B",X"F0",X"03",X"24",X"CD",X"2D",X"02",X"E6",X"42",X"1F",X"00",X"20",X"19",X"1A",X"04",
		X"06",X"08",X"0A",X"0C",X"0E",X"00",X"04",X"1B",X"F0",X"04",X"17",X"24",X"CD",X"2D",X"02",X"07",
		X"43",X"10",X"FF",X"FF",X"FF",X"01",X"02",X"05",X"07",X"09",X"0B",X"0D",X"0F",X"F1",X"05",X"F2",
		X"F4",X"14",X"1D",X"24",X"CD",X"2D",X"02",X"48",X"41",X"F3",X"F5",X"15",X"24",X"CD",X"2D",X"02",
		X"49",X"41",X"0D",X"0F",X"16",X"24",X"CD",X"30",X"02",X"DA",X"43",X"31",X"55",X"50",X"20",X"20",
		X"20",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"20",X"20",X"32",X"55",
		X"50",X"24",X"3E",X"30",X"32",X"F7",X"43",X"32",X"ED",X"43",X"32",X"E3",X"43",X"21",X"FD",X"43",
		X"11",X"25",X"4C",X"CD",X"09",X"10",X"2E",X"E9",X"11",X"28",X"4C",X"CD",X"09",X"10",X"2E",X"F3",
		X"11",X"05",X"4D",X"CD",X"09",X"10",X"CD",X"30",X"02",X"3C",X"40",X"43",X"52",X"45",X"44",X"49",
		X"54",X"20",X"20",X"30",X"20",X"20",X"20",X"40",X"4D",X"41",X"4D",X"41",X"20",X"54",X"4F",X"50",
		X"20",X"31",X"39",X"38",X"33",X"24",X"C3",X"33",X"02",X"32",X"7A",X"4C",X"F5",X"3E",X"FC",X"06",
		X"0A",X"21",X"3C",X"40",X"77",X"2B",X"10",X"FC",X"F1",X"F5",X"0F",X"0F",X"E6",X"07",X"16",X"00",
		X"5F",X"21",X"AE",X"0B",X"19",X"7E",X"21",X"13",X"44",X"11",X"33",X"44",X"06",X"08",X"77",X"12",
		X"23",X"13",X"10",X"FA",X"CD",X"30",X"02",X"1D",X"40",X"41",X"43",X"54",X"24",X"F1",X"F5",X"4F",
		X"E6",X"1F",X"FE",X"0A",X"79",X"38",X"02",X"C6",X"06",X"C6",X"01",X"27",X"4F",X"E6",X"0F",X"C6",
		X"30",X"32",X"3B",X"40",X"79",X"D7",X"E6",X"0F",X"28",X"04",X"C6",X"30",X"18",X"02",X"3E",X"20",
		X"32",X"3C",X"40",X"F1",X"21",X"60",X"66",X"11",X"62",X"64",X"22",X"19",X"40",X"ED",X"53",X"39",
		X"40",X"E6",X"03",X"C8",X"22",X"17",X"40",X"ED",X"53",X"37",X"40",X"3D",X"C8",X"22",X"15",X"40",
		X"ED",X"53",X"35",X"40",X"3D",X"C8",X"22",X"13",X"40",X"ED",X"53",X"33",X"40",X"C9",X"02",X"07",
		X"04",X"01",X"06",X"3E",X"07",X"32",X"D3",X"4F",X"3E",X"13",X"32",X"D7",X"4F",X"32",X"D9",X"4F",
		X"3E",X"01",X"32",X"DB",X"4F",X"3E",X"05",X"32",X"DD",X"4F",X"C9",X"CD",X"B3",X"0B",X"21",X"68",
		X"88",X"22",X"02",X"4C",X"21",X"30",X"00",X"22",X"06",X"4C",X"2E",X"A0",X"22",X"0B",X"4C",X"3E",
		X"02",X"32",X"08",X"4C",X"AF",X"32",X"0D",X"4C",X"32",X"04",X"4C",X"32",X"00",X"4D",X"3D",X"32",
		X"14",X"4D",X"3E",X"20",X"32",X"E3",X"4F",X"21",X"01",X"00",X"22",X"10",X"4C",X"CD",X"2A",X"02",
		X"FC",X"40",X"40",X"80",X"04",X"CD",X"2D",X"02",X"5F",X"43",X"72",X"70",X"FC",X"FC",X"77",X"75",
		X"FC",X"FC",X"72",X"70",X"FC",X"FC",X"76",X"74",X"FC",X"FC",X"73",X"71",X"FC",X"FC",X"76",X"74",
		X"24",X"CD",X"03",X"07",X"5E",X"40",X"1C",X"84",X"CD",X"03",X"07",X"72",X"40",X"1A",X"2D",X"3E",
		X"FB",X"21",X"40",X"40",X"06",X"0D",X"C5",X"CD",X"2F",X"0F",X"C1",X"23",X"10",X"F8",X"11",X"40",
		X"40",X"CD",X"86",X"0E",X"FF",X"22",X"FF",X"FF",X"23",X"FF",X"24",X"FF",X"FF",X"26",X"FF",X"FF",
		X"27",X"FF",X"28",X"29",X"2A",X"2B",X"00",X"11",X"52",X"40",X"CD",X"B5",X"0E",X"11",X"A0",X"43",
		X"CD",X"86",X"0E",X"FF",X"FF",X"FF",X"22",X"24",X"FF",X"D7",X"D8",X"D9",X"D3",X"FF",X"3C",X"24",
		X"FF",X"D7",X"D8",X"D9",X"D3",X"FF",X"22",X"FF",X"00",X"11",X"B5",X"43",X"CD",X"A7",X"0E",X"11",
		X"F2",X"41",X"CD",X"86",X"0E",X"3B",X"22",X"3C",X"00",X"11",X"F5",X"41",X"CD",X"A7",X"0E",X"11",
		X"12",X"42",X"CD",X"B5",X"0E",X"21",X"EC",X"ED",X"22",X"D2",X"41",X"21",X"EE",X"EF",X"22",X"32",
		X"42",X"11",X"7B",X"40",X"CD",X"70",X"0E",X"11",X"BB",X"41",X"CD",X"7B",X"0E",X"11",X"3B",X"42",
		X"CD",X"70",X"0E",X"11",X"7B",X"43",X"CD",X"7B",X"0E",X"11",X"72",X"40",X"CD",X"2E",X"0E",X"11",
		X"53",X"41",X"CD",X"4F",X"0E",X"11",X"34",X"42",X"CD",X"2E",X"0E",X"11",X"12",X"43",X"CD",X"4F",
		X"0E",X"3E",X"C7",X"32",X"92",X"40",X"32",X"72",X"43",X"11",X"60",X"40",X"CD",X"86",X"0E",X"02",
		X"9C",X"9D",X"01",X"A0",X"A1",X"A2",X"02",X"87",X"FC",X"E2",X"FF",X"FF",X"E1",X"E0",X"3F",X"20",
		X"01",X"9A",X"81",X"83",X"A3",X"A4",X"02",X"9C",X"9D",X"85",X"E2",X"FF",X"E1",X"E0",X"20",X"02",
		X"9E",X"9F",X"A5",X"7C",X"98",X"9A",X"80",X"82",X"A3",X"FF",X"E3",X"20",X"04",X"97",X"7E",X"99",
		X"01",X"9E",X"9F",X"B0",X"B1",X"78",X"C4",X"20",X"05",X"95",X"03",X"B2",X"A4",X"97",X"7A",X"C5",
		X"20",X"06",X"9C",X"9D",X"01",X"B3",X"7C",X"98",X"C1",X"FC",X"20",X"01",X"9C",X"9D",X"02",X"9A",
		X"81",X"83",X"A3",X"B4",X"7E",X"99",X"85",X"20",X"DA",X"80",X"82",X"9B",X"02",X"9E",X"9F",X"B5",
		X"01",X"95",X"02",X"85",X"20",X"DB",X"9E",X"9F",X"05",X"B6",X"04",X"87",X"20",X"FF",X"B7",X"0B",
		X"85",X"20",X"A9",X"DB",X"01",X"9C",X"9D",X"08",X"86",X"20",X"01",X"DC",X"DD",X"81",X"83",X"9B",
		X"06",X"86",X"FC",X"20",X"96",X"79",X"DE",X"DF",X"9F",X"07",X"85",X"20",X"97",X"7B",X"99",X"09",
		X"87",X"20",X"01",X"95",X"0A",X"85",X"FC",X"20",X"0D",X"85",X"20",X"0D",X"87",X"20",X"09",X"B7",
		X"03",X"85",X"20",X"03",X"94",X"03",X"9C",X"9D",X"B8",X"03",X"FB",X"85",X"FC",X"FC",X"3F",X"20",
		X"02",X"BD",X"78",X"98",X"01",X"9A",X"81",X"83",X"A7",X"B7",X"02",X"FB",X"FB",X"20",X"02",X"BE",
		X"7A",X"99",X"94",X"01",X"9E",X"9F",X"01",X"B8",X"02",X"94",X"FB",X"85",X"20",X"02",X"B9",X"A8",
		X"96",X"78",X"98",X"03",X"B9",X"BA",X"96",X"78",X"98",X"87",X"20",X"00",X"11",X"20",X"43",X"CD",
		X"0B",X"0E",X"11",X"28",X"43",X"CD",X"0B",X"0E",X"11",X"2E",X"43",X"CD",X"86",X"0E",X"01",X"85",
		X"20",X"FB",X"FB",X"FC",X"3F",X"20",X"02",X"85",X"3F",X"20",X"03",X"EB",X"00",X"CD",X"2D",X"02",
		X"6E",X"42",X"8F",X"AE",X"AE",X"FC",X"FC",X"AE",X"AE",X"AF",X"24",X"CD",X"03",X"07",X"91",X"41",
		X"08",X"8B",X"11",X"6E",X"41",X"CD",X"86",X"0E",X"88",X"89",X"AC",X"8A",X"00",X"11",X"8E",X"42",
		X"CD",X"86",X"0E",X"8E",X"8D",X"AD",X"8C",X"00",X"C3",X"C6",X"0E",X"CD",X"86",X"0E",X"01",X"9C",
		X"9D",X"BB",X"BC",X"7A",X"99",X"20",X"9A",X"80",X"82",X"A7",X"FF",X"A8",X"20",X"01",X"9E",X"9F",
		X"01",X"A9",X"FF",X"A6",X"AA",X"20",X"05",X"A9",X"FF",X"FF",X"A6",X"AA",X"00",X"C9",X"CD",X"86",
		X"0E",X"01",X"C8",X"C9",X"01",X"E2",X"E1",X"E0",X"20",X"C6",X"81",X"83",X"E4",X"E3",X"20",X"01",
		X"CA",X"CB",X"E5",X"7D",X"C4",X"20",X"03",X"C3",X"7F",X"C5",X"20",X"04",X"C1",X"00",X"C9",X"CD",
		X"86",X"0E",X"04",X"C0",X"20",X"03",X"C2",X"79",X"C4",X"20",X"01",X"C8",X"C9",X"E6",X"7B",X"C5",
		X"20",X"C6",X"80",X"82",X"E7",X"E8",X"20",X"01",X"CA",X"CB",X"01",X"E9",X"EA",X"EB",X"00",X"C9",
		X"CD",X"86",X"0E",X"D0",X"D1",X"2A",X"20",X"02",X"D2",X"00",X"C9",X"CD",X"86",X"0E",X"02",X"D6",
		X"20",X"D4",X"D5",X"D9",X"00",X"C9",X"E1",X"D5",X"7E",X"23",X"A7",X"20",X"02",X"D1",X"E9",X"47",
		X"FE",X"20",X"28",X"0B",X"38",X"04",X"12",X"13",X"18",X"EE",X"13",X"10",X"FD",X"18",X"E9",X"E3",
		X"11",X"20",X"00",X"19",X"EB",X"18",X"DF",X"CD",X"86",X"0E",X"3D",X"24",X"FF",X"3E",X"5B",X"5C",
		X"5D",X"5E",X"D9",X"00",X"C9",X"CD",X"86",X"0E",X"FF",X"FF",X"26",X"FF",X"FF",X"2B",X"26",X"3A",
		X"FF",X"FF",X"FF",X"FF",X"00",X"C9",X"CD",X"00",X"30",X"CD",X"2A",X"02",X"1C",X"40",X"44",X"80",
		X"04",X"CD",X"03",X"07",X"72",X"44",X"0B",X"0E",X"CD",X"03",X"07",X"52",X"46",X"0B",X"0E",X"21",
		X"5E",X"44",X"3E",X"1F",X"CD",X"2F",X"0F",X"23",X"3E",X"16",X"CD",X"2F",X"0F",X"2A",X"38",X"02",
		X"5E",X"23",X"7E",X"23",X"A7",X"28",X"08",X"C6",X"04",X"57",X"3E",X"0F",X"12",X"18",X"F1",X"3E",
		X"12",X"06",X"04",X"21",X"6E",X"45",X"C5",X"CD",X"33",X"0F",X"23",X"C1",X"10",X"F8",X"11",X"2B",
		X"0F",X"06",X"04",X"21",X"8F",X"45",X"1A",X"13",X"D5",X"CD",X"4C",X"0F",X"19",X"D1",X"10",X"F6",
		X"3E",X"02",X"21",X"ED",X"45",X"CD",X"4C",X"0F",X"C3",X"03",X"30",X"04",X"05",X"07",X"06",X"06",
		X"1C",X"18",X"02",X"06",X"0A",X"E5",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"E1",X"C9",X"E1",
		X"5E",X"23",X"56",X"23",X"46",X"23",X"7E",X"23",X"E5",X"EB",X"18",X"E9",X"77",X"23",X"77",X"11",
		X"20",X"00",X"19",X"77",X"2B",X"77",X"C9",X"10",X"F4",X"C9",X"7B",X"E6",X"0F",X"DD",X"77",X"05",
		X"7B",X"D7",X"E6",X"0F",X"DD",X"77",X"06",X"7A",X"E6",X"0F",X"DD",X"77",X"07",X"7A",X"D7",X"E6",
		X"0F",X"DD",X"77",X"08",X"C9",X"AF",X"06",X"0C",X"DD",X"E5",X"E1",X"77",X"23",X"10",X"FC",X"C9",
		X"27",X"3F",X"44",X"18",X"25",X"4A",X"89",X"91",X"1F",X"00",X"20",X"3F",X"40",X"56",X"1F",X"5C",
		X"1F",X"00",X"27",X"3E",X"40",X"56",X"16",X"30",X"14",X"20",X"3F",X"16",X"30",X"12",X"27",X"3E",
		X"40",X"56",X"16",X"30",X"14",X"20",X"3F",X"16",X"00",X"27",X"3F",X"4C",X"18",X"30",X"18",X"26",
		X"4F",X"9A",X"1F",X"1F",X"00",X"3F",X"61",X"99",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"18",X"C2",X"18",X"C4",X"18",X"C5",X"18",X"C7",X"18",X"C9",X"18",X"CB",X"18",X"D0",X"18",X"00",
		X"00",X"00",X"4F",X"9A",X"1F",X"1F",X"00",X"3F",X"61",X"99",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"18",X"C2",X"18",X"C4",X"18",X"C5",X"18",X"C7",X"18",X"C9",X"18",X"CB",X"18",X"D0",
		X"18",X"00",X"00",X"00",X"50",X"CB",X"7F",X"7E",X"28",X"05",X"E6",X"0F",X"C8",X"35",X"C9",X"67",
		X"C3",X"B8",X"10",X"C3",X"BB",X"10",X"C3",X"59",X"15",X"C3",X"57",X"1A",X"C3",X"12",X"10",X"C3",
		X"85",X"19",X"3A",X"7A",X"4C",X"CB",X"4F",X"C4",X"00",X"1C",X"2A",X"02",X"4C",X"11",X"00",X"00",
		X"7C",X"FE",X"68",X"38",X"30",X"FE",X"B0",X"30",X"2C",X"7D",X"FE",X"38",X"38",X"27",X"FE",X"98",
		X"30",X"23",X"FE",X"68",X"38",X"03",X"11",X"08",X"08",X"3A",X"ED",X"41",X"01",X"01",X"01",X"0F",
		X"38",X"03",X"01",X"00",X"00",X"21",X"60",X"62",X"09",X"19",X"22",X"ED",X"41",X"21",X"66",X"64",
		X"09",X"19",X"22",X"0D",X"42",X"3A",X"19",X"4C",X"FE",X"02",X"28",X"0F",X"30",X"37",X"CD",X"59",
		X"15",X"3E",X"01",X"32",X"4C",X"4C",X"CD",X"A5",X"10",X"18",X"21",X"3A",X"18",X"4C",X"CB",X"67",
		X"20",X"08",X"CD",X"A5",X"10",X"21",X"02",X"02",X"18",X"15",X"CD",X"2D",X"02",X"2C",X"42",X"46",
		X"45",X"45",X"44",X"21",X"24",X"CD",X"03",X"07",X"AC",X"45",X"05",X"05",X"21",X"0D",X"0D",X"22",
		X"ED",X"45",X"22",X"0D",X"46",X"21",X"18",X"4C",X"35",X"20",X"1D",X"23",X"35",X"20",X"19",X"CD",
		X"09",X"27",X"C3",X"44",X"18",X"CD",X"2D",X"02",X"2C",X"42",X"85",X"87",X"85",X"86",X"FB",X"24",
		X"CD",X"03",X"07",X"AC",X"45",X"05",X"1C",X"C9",X"AF",X"18",X"02",X"3E",X"FF",X"21",X"05",X"4C",
		X"34",X"2B",X"CB",X"46",X"CA",X"CB",X"13",X"CB",X"7E",X"28",X"0B",X"CB",X"4E",X"11",X"BA",X"B8",
		X"CA",X"F8",X"13",X"C3",X"06",X"1C",X"A7",X"C2",X"B7",X"12",X"3A",X"00",X"4C",X"CB",X"77",X"C2",
		X"75",X"12",X"3A",X"10",X"4C",X"E6",X"07",X"C2",X"B7",X"12",X"CD",X"85",X"19",X"E6",X"07",X"06",
		X"FF",X"20",X"09",X"3A",X"03",X"4C",X"FE",X"10",X"38",X"02",X"06",X"00",X"78",X"32",X"14",X"4D",
		X"DD",X"21",X"06",X"4C",X"CD",X"61",X"11",X"DD",X"21",X"0B",X"4C",X"CD",X"61",X"11",X"21",X"04",
		X"4C",X"CB",X"66",X"28",X"0C",X"11",X"68",X"78",X"21",X"00",X"00",X"22",X"84",X"4C",X"C3",X"C7",
		X"11",X"ED",X"5B",X"84",X"4C",X"7B",X"B2",X"C2",X"C7",X"11",X"CD",X"85",X"19",X"3A",X"12",X"4C",
		X"E6",X"3E",X"4F",X"06",X"20",X"C5",X"06",X"00",X"21",X"35",X"12",X"09",X"56",X"23",X"5E",X"D5",
		X"EB",X"11",X"07",X"07",X"19",X"CD",X"33",X"15",X"D1",X"C1",X"38",X"08",X"79",X"C6",X"02",X"E6",
		X"3E",X"4F",X"10",X"E1",X"7A",X"FE",X"ED",X"20",X"02",X"16",X"00",X"ED",X"53",X"84",X"4C",X"18",
		X"66",X"DD",X"46",X"02",X"78",X"E6",X"F8",X"C8",X"FE",X"08",X"20",X"3E",X"CB",X"40",X"C0",X"DD",
		X"7E",X"00",X"FE",X"60",X"28",X"2C",X"FE",X"70",X"28",X"28",X"A7",X"3A",X"02",X"4C",X"06",X"88",
		X"28",X"06",X"4F",X"3E",X"D0",X"91",X"06",X"80",X"FE",X"38",X"D0",X"4F",X"3A",X"03",X"4C",X"DD",
		X"96",X"01",X"D0",X"ED",X"44",X"81",X"4F",X"DD",X"7E",X"01",X"B8",X"30",X"19",X"81",X"B8",X"D0",
		X"18",X"14",X"DD",X"7E",X"01",X"FE",X"20",X"D8",X"18",X"0C",X"CB",X"60",X"C8",X"CB",X"68",X"28",
		X"05",X"78",X"0F",X"A8",X"0F",X"D0",X"21",X"00",X"00",X"22",X"84",X"4C",X"DD",X"5E",X"00",X"DD",
		X"56",X"01",X"AF",X"32",X"14",X"4D",X"E1",X"0E",X"00",X"3A",X"03",X"4C",X"A7",X"20",X"02",X"CB",
		X"D9",X"92",X"30",X"04",X"CB",X"C9",X"ED",X"44",X"FE",X"05",X"30",X"02",X"CB",X"C1",X"47",X"3A",
		X"02",X"4C",X"93",X"30",X"04",X"CB",X"E9",X"ED",X"44",X"FE",X"05",X"30",X"02",X"CB",X"E1",X"B8",
		X"30",X"03",X"CB",X"F1",X"3F",X"1F",X"B8",X"38",X"02",X"CB",X"F9",X"3A",X"04",X"4C",X"47",X"79",
		X"E6",X"11",X"28",X"12",X"FE",X"10",X"28",X"1A",X"38",X"1D",X"CB",X"59",X"28",X"04",X"06",X"01",
		X"18",X"1D",X"78",X"2F",X"18",X"08",X"79",X"07",X"38",X"0D",X"07",X"38",X"05",X"78",X"E6",X"04",
		X"20",X"05",X"79",X"E6",X"02",X"18",X"06",X"79",X"D7",X"E6",X"02",X"F6",X"04",X"3C",X"47",X"21",
		X"04",X"4C",X"C3",X"A4",X"12",X"40",X"54",X"A8",X"9C",X"ED",X"98",X"90",X"30",X"C8",X"5C",X"30",
		X"B8",X"B0",X"34",X"ED",X"18",X"30",X"18",X"38",X"7C",X"78",X"B0",X"20",X"88",X"ED",X"38",X"80",
		X"20",X"98",X"BC",X"28",X"48",X"48",X"0C",X"ED",X"B8",X"A0",X"14",X"48",X"C4",X"D8",X"3C",X"B8",
		X"B0",X"B8",X"18",X"C8",X"A0",X"D8",X"68",X"D0",X"0C",X"D8",X"BC",X"40",X"54",X"A8",X"9C",X"90",
		X"30",X"C8",X"5C",X"30",X"B8",X"CD",X"1D",X"15",X"47",X"3A",X"03",X"4C",X"FE",X"10",X"78",X"30",
		X"02",X"3E",X"FF",X"32",X"14",X"4D",X"78",X"21",X"04",X"4C",X"0F",X"30",X"0D",X"0F",X"30",X"0E",
		X"0F",X"30",X"0F",X"0F",X"38",X"21",X"06",X"01",X"18",X"0A",X"06",X"03",X"18",X"06",X"06",X"07",
		X"18",X"02",X"06",X"05",X"7E",X"E6",X"07",X"B8",X"28",X"0D",X"3E",X"01",X"32",X"05",X"4C",X"7E",
		X"E6",X"F8",X"B0",X"77",X"CD",X"85",X"19",X"46",X"E5",X"3A",X"14",X"4D",X"07",X"D2",X"A2",X"13",
		X"2A",X"02",X"4C",X"CB",X"58",X"C2",X"67",X"13",X"CB",X"50",X"20",X"1C",X"7D",X"C6",X"07",X"6F",
		X"7C",X"C6",X"07",X"CB",X"48",X"28",X"02",X"C6",X"08",X"67",X"CD",X"33",X"15",X"38",X"1B",X"2C",
		X"CD",X"33",X"15",X"38",X"15",X"C3",X"A2",X"13",X"7C",X"C6",X"0A",X"67",X"CB",X"48",X"28",X"04",
		X"7D",X"C6",X"0F",X"6F",X"CD",X"33",X"15",X"D2",X"A2",X"13",X"CB",X"60",X"20",X"16",X"FE",X"70",
		X"DA",X"A2",X"13",X"47",X"3E",X"FE",X"CD",X"F3",X"14",X"3A",X"7B",X"4C",X"47",X"3E",X"01",X"0E",
		X"10",X"C3",X"90",X"13",X"FE",X"70",X"D2",X"A2",X"13",X"AF",X"32",X"D4",X"4F",X"21",X"18",X"4C",
		X"77",X"3A",X"7A",X"4C",X"E6",X"02",X"3E",X"05",X"20",X"01",X"3D",X"23",X"77",X"C5",X"CD",X"A5",
		X"10",X"C1",X"21",X"02",X"02",X"22",X"ED",X"45",X"22",X"0D",X"46",X"3E",X"02",X"32",X"4C",X"4C",
		X"0E",X"03",X"CD",X"1D",X"19",X"3A",X"7C",X"4C",X"CB",X"68",X"28",X"03",X"3A",X"7E",X"4C",X"CD",
		X"97",X"19",X"E1",X"7E",X"E6",X"CF",X"77",X"EB",X"21",X"16",X"4C",X"35",X"EB",X"20",X"44",X"21",
		X"01",X"4C",X"0E",X"03",X"C3",X"99",X"18",X"78",X"E6",X"36",X"20",X"36",X"CB",X"70",X"28",X"32",
		X"3A",X"05",X"4C",X"E6",X"E0",X"28",X"2B",X"26",X"F4",X"7D",X"C6",X"07",X"6F",X"CD",X"33",X"15",
		X"30",X"20",X"47",X"3E",X"FC",X"CD",X"F3",X"14",X"3A",X"7D",X"4C",X"47",X"3E",X"16",X"0E",X"30",
		X"32",X"D5",X"4F",X"78",X"CD",X"97",X"19",X"E1",X"7E",X"B1",X"77",X"0E",X"02",X"CD",X"1D",X"19",
		X"18",X"01",X"E1",X"11",X"02",X"4C",X"0E",X"D0",X"CB",X"5E",X"C2",X"3E",X"14",X"CB",X"56",X"20",
		X"03",X"13",X"0E",X"D8",X"1A",X"CB",X"4E",X"28",X"06",X"B9",X"30",X"0F",X"3C",X"18",X"0B",X"A7",
		X"20",X"07",X"CB",X"56",X"CA",X"28",X"14",X"18",X"02",X"3D",X"12",X"7E",X"0F",X"E6",X"03",X"28",
		X"0B",X"3D",X"28",X"1C",X"3D",X"28",X"1E",X"11",X"AA",X"A2",X"18",X"1C",X"11",X"92",X"90",X"3A",
		X"14",X"4D",X"07",X"38",X"13",X"11",X"9B",X"99",X"E5",X"21",X"03",X"4C",X"35",X"E1",X"18",X"08",
		X"11",X"9A",X"98",X"18",X"03",X"11",X"A0",X"A8",X"CB",X"76",X"28",X"07",X"E5",X"21",X"04",X"04",
		X"19",X"EB",X"E1",X"CD",X"D3",X"14",X"7A",X"32",X"D6",X"4F",X"7B",X"32",X"D8",X"4F",X"3A",X"02",
		X"4C",X"C6",X"17",X"32",X"E8",X"4F",X"C6",X"10",X"32",X"E6",X"4F",X"3A",X"03",X"4C",X"C6",X"20",
		X"32",X"E9",X"4F",X"32",X"E7",X"4F",X"18",X"5C",X"7E",X"C6",X"08",X"77",X"AF",X"32",X"D8",X"4F",
		X"3C",X"32",X"05",X"4C",X"3A",X"02",X"4C",X"C6",X"1F",X"32",X"E6",X"4F",X"18",X"2A",X"CB",X"56",
		X"28",X"21",X"23",X"34",X"CB",X"86",X"2B",X"1A",X"CB",X"4E",X"28",X"08",X"B9",X"0E",X"82",X"28",
		X"0F",X"3C",X"18",X"06",X"0E",X"80",X"A7",X"28",X"07",X"3D",X"12",X"C6",X"1F",X"32",X"E6",X"4F",
		X"79",X"18",X"15",X"CB",X"4E",X"C2",X"EC",X"14",X"CB",X"66",X"28",X"0A",X"3E",X"B0",X"CB",X"76",
		X"28",X"0C",X"C6",X"02",X"18",X"08",X"3E",X"88",X"CB",X"76",X"28",X"02",X"C6",X"04",X"32",X"D6",
		X"4F",X"CD",X"D3",X"14",X"CB",X"66",X"C8",X"46",X"EB",X"2A",X"02",X"4C",X"CB",X"50",X"20",X"1C",
		X"0E",X"60",X"CB",X"48",X"28",X"08",X"7C",X"C6",X"08",X"67",X"0E",X"64",X"18",X"1D",X"3A",X"14",
		X"4D",X"07",X"38",X"17",X"7C",X"D6",X"08",X"67",X"0E",X"65",X"18",X"0F",X"7D",X"D6",X"08",X"6F",
		X"0E",X"68",X"CB",X"48",X"28",X"05",X"C6",X"10",X"6F",X"0E",X"6C",X"7D",X"C6",X"1E",X"32",X"E4",
		X"4F",X"7C",X"C6",X"20",X"32",X"E5",X"4F",X"EB",X"79",X"CB",X"6E",X"28",X"02",X"C6",X"10",X"32",
		X"D4",X"4F",X"C9",X"06",X"0F",X"3A",X"14",X"4D",X"07",X"38",X"07",X"7E",X"E6",X"06",X"28",X"02",
		X"06",X"03",X"3A",X"05",X"4C",X"A0",X"C0",X"7E",X"EE",X"40",X"77",X"C9",X"7E",X"EE",X"08",X"77",
		X"C3",X"CB",X"13",X"ED",X"53",X"12",X"4D",X"12",X"CB",X"78",X"20",X"13",X"CB",X"48",X"01",X"20",
		X"00",X"28",X"03",X"01",X"E0",X"FF",X"EB",X"09",X"77",X"EB",X"CB",X"48",X"C8",X"18",X"09",X"CB",
		X"48",X"20",X"03",X"13",X"12",X"C9",X"1B",X"12",X"ED",X"53",X"12",X"4D",X"C9",X"3A",X"40",X"50",
		X"21",X"01",X"4C",X"CB",X"76",X"C0",X"07",X"07",X"07",X"E6",X"80",X"47",X"3A",X"00",X"50",X"E6",
		X"7F",X"B0",X"C9",X"E5",X"3E",X"EF",X"94",X"0F",X"0F",X"0F",X"E6",X"1F",X"5F",X"7D",X"07",X"07",
		X"57",X"E6",X"E0",X"B3",X"5F",X"7A",X"E6",X"03",X"57",X"21",X"40",X"40",X"19",X"EB",X"1A",X"E1",
		X"FE",X"60",X"30",X"02",X"3F",X"C9",X"FE",X"84",X"C9",X"DD",X"21",X"06",X"4C",X"21",X"DA",X"4F",
		X"CD",X"6A",X"15",X"DD",X"21",X"0B",X"4C",X"21",X"DC",X"4F",X"DD",X"34",X"04",X"DD",X"CB",X"02",
		X"76",X"C2",X"CF",X"18",X"E5",X"21",X"82",X"4C",X"36",X"00",X"3A",X"02",X"4C",X"DD",X"96",X"00",
		X"30",X"04",X"CB",X"CE",X"ED",X"44",X"47",X"5F",X"3A",X"03",X"4C",X"DD",X"96",X"01",X"30",X"04",
		X"CB",X"C6",X"ED",X"44",X"6F",X"4F",X"AF",X"67",X"57",X"19",X"22",X"80",X"4C",X"E1",X"3A",X"14",
		X"4D",X"07",X"38",X"0B",X"79",X"FE",X"09",X"30",X"06",X"78",X"FE",X"11",X"DA",X"A4",X"18",X"DD",
		X"7E",X"02",X"D7",X"E6",X"0F",X"28",X"0C",X"3D",X"CA",X"98",X"17",X"3D",X"CA",X"29",X"18",X"3D",
		X"CA",X"FA",X"16",X"DD",X"7E",X"02",X"CB",X"5F",X"C2",X"1F",X"16",X"0F",X"30",X"3E",X"0F",X"30",
		X"1F",X"CD",X"32",X"19",X"30",X"09",X"3A",X"02",X"4C",X"DD",X"BE",X"00",X"D2",X"B4",X"16",X"DD",
		X"7E",X"00",X"FE",X"D0",X"30",X"32",X"CD",X"3F",X"19",X"38",X"2D",X"DD",X"34",X"00",X"18",X"1C",
		X"CD",X"32",X"19",X"30",X"09",X"3A",X"02",X"4C",X"DD",X"BE",X"00",X"DA",X"AD",X"16",X"DD",X"7E",
		X"00",X"A7",X"28",X"14",X"CD",X"3F",X"19",X"38",X"0F",X"DD",X"35",X"00",X"DD",X"46",X"02",X"78",
		X"E6",X"06",X"C6",X"C0",X"77",X"C3",X"FE",X"18",X"DD",X"36",X"02",X"08",X"C3",X"BB",X"16",X"DD",
		X"7E",X"00",X"A7",X"20",X"0D",X"DD",X"7E",X"01",X"FE",X"88",X"20",X"17",X"CD",X"49",X"19",X"DA",
		X"EA",X"16",X"FE",X"D0",X"20",X"0D",X"DD",X"7E",X"01",X"FE",X"80",X"20",X"06",X"CD",X"49",X"19",
		X"DA",X"F0",X"16",X"DD",X"46",X"02",X"CB",X"40",X"20",X"37",X"CD",X"32",X"19",X"30",X"08",X"3A",
		X"03",X"4C",X"DD",X"BE",X"01",X"30",X"24",X"DD",X"7E",X"01",X"FE",X"58",X"20",X"0D",X"DD",X"7E",
		X"00",X"FE",X"60",X"CA",X"79",X"17",X"FE",X"70",X"CA",X"7F",X"17",X"DD",X"7E",X"01",X"CB",X"48",
		X"20",X"49",X"FE",X"E0",X"30",X"05",X"DD",X"34",X"01",X"18",X"40",X"DD",X"36",X"02",X"09",X"18",
		X"3A",X"CD",X"32",X"19",X"30",X"08",X"3A",X"03",X"4C",X"DD",X"BE",X"01",X"38",X"8A",X"DD",X"7E",
		X"01",X"A7",X"28",X"0A",X"DD",X"35",X"01",X"28",X"05",X"DD",X"35",X"01",X"20",X"1D",X"DD",X"7E",
		X"00",X"A7",X"28",X"09",X"FE",X"D0",X"28",X"0C",X"CD",X"85",X"19",X"38",X"07",X"DD",X"36",X"02",
		X"03",X"C3",X"0C",X"16",X"DD",X"36",X"02",X"01",X"C3",X"0C",X"16",X"DD",X"46",X"02",X"78",X"0F",
		X"E6",X"03",X"E5",X"21",X"E6",X"16",X"16",X"00",X"5F",X"19",X"56",X"78",X"E6",X"01",X"82",X"E1",
		X"77",X"DD",X"7E",X"04",X"E6",X"07",X"C2",X"0B",X"19",X"78",X"C6",X"02",X"E6",X"07",X"C6",X"08",
		X"DD",X"77",X"02",X"C3",X"0B",X"19",X"C8",X"CC",X"CE",X"CA",X"DD",X"36",X"02",X"32",X"18",X"04",
		X"DD",X"36",X"02",X"31",X"DD",X"36",X"03",X"00",X"18",X"61",X"DD",X"7E",X"02",X"CB",X"4F",X"20",
		X"1E",X"CD",X"32",X"19",X"30",X"08",X"3A",X"02",X"4C",X"DD",X"BE",X"00",X"38",X"45",X"DD",X"7E",
		X"00",X"A7",X"CA",X"7B",X"16",X"FE",X"90",X"CA",X"85",X"17",X"DD",X"35",X"00",X"18",X"1D",X"CD",
		X"32",X"19",X"30",X"08",X"3A",X"02",X"4C",X"DD",X"BE",X"00",X"30",X"27",X"DD",X"7E",X"00",X"FE",
		X"D0",X"CA",X"7B",X"16",X"FE",X"40",X"CA",X"8B",X"17",X"DD",X"34",X"00",X"DD",X"7E",X"02",X"CB",
		X"5F",X"28",X"18",X"47",X"0F",X"A8",X"0F",X"38",X"05",X"DD",X"35",X"01",X"18",X"0D",X"DD",X"34",
		X"01",X"18",X"08",X"DD",X"7E",X"02",X"EE",X"02",X"DD",X"77",X"02",X"DD",X"7E",X"02",X"E6",X"06",
		X"C6",X"C0",X"77",X"DD",X"7E",X"02",X"EE",X"08",X"47",X"DD",X"7E",X"04",X"E6",X"07",X"78",X"20",
		X"02",X"EE",X"04",X"DD",X"77",X"02",X"C3",X"0B",X"19",X"DD",X"36",X"02",X"10",X"18",X"10",X"DD",
		X"36",X"02",X"12",X"18",X"0A",X"DD",X"36",X"02",X"11",X"18",X"04",X"DD",X"36",X"02",X"13",X"DD",
		X"36",X"03",X"00",X"0E",X"50",X"CD",X"21",X"19",X"DD",X"7E",X"02",X"E6",X"03",X"07",X"5F",X"16",
		X"00",X"E5",X"21",X"D7",X"17",X"19",X"5E",X"23",X"56",X"EB",X"DD",X"5E",X"03",X"DD",X"34",X"03",
		X"16",X"00",X"19",X"7E",X"E1",X"A7",X"CA",X"07",X"18",X"DD",X"77",X"00",X"DD",X"7E",X"01",X"C6",
		X"04",X"DD",X"CB",X"02",X"46",X"28",X"02",X"D6",X"08",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"E6",
		X"03",X"C6",X"F0",X"77",X"C3",X"0B",X"19",X"DF",X"17",X"FC",X"17",X"E7",X"17",X"EF",X"17",X"60",
		X"60",X"61",X"63",X"65",X"67",X"68",X"00",X"70",X"70",X"6F",X"6D",X"6B",X"69",X"68",X"00",X"48",
		X"50",X"56",X"58",X"5B",X"5E",X"60",X"62",X"64",X"66",X"67",X"68",X"00",X"88",X"7E",X"78",X"74",
		X"70",X"6D",X"6B",X"6A",X"69",X"68",X"00",X"DD",X"7E",X"02",X"E6",X"03",X"F6",X"20",X"DD",X"77",
		X"02",X"DD",X"36",X"03",X"00",X"3A",X"04",X"4C",X"E6",X"70",X"F6",X"81",X"32",X"04",X"4C",X"3E",
		X"FF",X"32",X"14",X"4D",X"0E",X"70",X"C3",X"21",X"19",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"E6",
		X"0F",X"C0",X"DD",X"7E",X"02",X"C6",X"04",X"CB",X"67",X"20",X"09",X"DD",X"77",X"02",X"E6",X"0F",
		X"C6",X"F0",X"77",X"C9",X"21",X"FC",X"FC",X"22",X"ED",X"41",X"22",X"0D",X"42",X"21",X"01",X"4C",
		X"CB",X"66",X"28",X"17",X"CD",X"2D",X"02",X"8B",X"42",X"47",X"41",X"4D",X"45",X"20",X"20",X"4F",
		X"56",X"45",X"52",X"24",X"CD",X"03",X"07",X"6B",X"45",X"0A",X"01",X"06",X"64",X"CD",X"24",X"02",
		X"10",X"FB",X"CD",X"06",X"30",X"21",X"00",X"4C",X"CB",X"76",X"20",X"07",X"21",X"20",X"00",X"22",
		X"00",X"4C",X"C9",X"23",X"CB",X"66",X"C2",X"06",X"27",X"CB",X"7E",X"28",X"08",X"CB",X"56",X"20",
		X"04",X"7E",X"EE",X"40",X"77",X"0E",X"00",X"CB",X"86",X"2B",X"7E",X"E6",X"F0",X"B1",X"77",X"AF",
		X"32",X"14",X"4C",X"C9",X"DD",X"7E",X"01",X"FE",X"08",X"38",X"0B",X"0E",X"40",X"CD",X"21",X"19",
		X"3A",X"7F",X"4C",X"CD",X"97",X"19",X"06",X"49",X"DD",X"7E",X"00",X"FE",X"68",X"30",X"02",X"06",
		X"4B",X"DD",X"70",X"02",X"DD",X"7E",X"01",X"0F",X"E6",X"7F",X"C6",X"50",X"DD",X"77",X"03",X"DD",
		X"46",X"02",X"CB",X"58",X"28",X"17",X"DD",X"7E",X"01",X"D6",X"04",X"38",X"05",X"DD",X"77",X"01",
		X"18",X"18",X"AF",X"DD",X"77",X"01",X"78",X"EE",X"09",X"DD",X"77",X"02",X"47",X"DD",X"35",X"03",
		X"20",X"08",X"CB",X"48",X"CA",X"B4",X"16",X"C3",X"AD",X"16",X"78",X"F6",X"D0",X"77",X"3A",X"10",
		X"4C",X"E6",X"07",X"20",X"06",X"78",X"EE",X"04",X"DD",X"77",X"02",X"11",X"10",X"00",X"19",X"DD",
		X"7E",X"00",X"C6",X"1F",X"77",X"DD",X"7E",X"01",X"23",X"C6",X"20",X"77",X"C9",X"16",X"F0",X"18",
		X"02",X"16",X"0F",X"3A",X"00",X"4C",X"FE",X"50",X"D8",X"3A",X"4A",X"4C",X"A2",X"B1",X"32",X"4A",
		X"4C",X"C9",X"3A",X"81",X"4C",X"A7",X"C0",X"3A",X"80",X"4C",X"FE",X"48",X"D0",X"18",X"46",X"FE",
		X"60",X"28",X"06",X"FE",X"70",X"28",X"02",X"A7",X"C9",X"3A",X"7A",X"4C",X"E6",X"FC",X"20",X"12",
		X"3A",X"01",X"4C",X"E6",X"08",X"28",X"2E",X"CD",X"85",X"19",X"CD",X"85",X"19",X"E6",X"03",X"C8",
		X"37",X"C9",X"3A",X"81",X"4C",X"A7",X"37",X"C0",X"3A",X"80",X"4C",X"FE",X"78",X"3F",X"D8",X"FE",
		X"48",X"30",X"E4",X"3A",X"04",X"4C",X"4F",X"3A",X"82",X"4C",X"CB",X"51",X"20",X"01",X"07",X"A9",
		X"E6",X"02",X"C0",X"37",X"C9",X"E5",X"21",X"13",X"4C",X"7E",X"07",X"2B",X"AE",X"0F",X"7E",X"17",
		X"77",X"23",X"7E",X"17",X"77",X"E1",X"C9",X"E5",X"57",X"E6",X"0F",X"C6",X"30",X"32",X"4A",X"42",
		X"7A",X"D7",X"E6",X"0F",X"20",X"02",X"3E",X"F0",X"C6",X"30",X"32",X"6A",X"42",X"C5",X"D5",X"CD",
		X"03",X"07",X"AA",X"45",X"07",X"07",X"CD",X"2D",X"02",X"2A",X"42",X"30",X"20",X"50",X"54",X"53",
		X"24",X"3E",X"32",X"32",X"20",X"4C",X"D1",X"C1",X"7A",X"21",X"00",X"4C",X"CB",X"76",X"CA",X"55",
		X"1A",X"23",X"CB",X"76",X"21",X"24",X"4C",X"28",X"03",X"21",X"27",X"4C",X"56",X"E5",X"2B",X"06",
		X"03",X"86",X"27",X"77",X"30",X"06",X"23",X"7E",X"C6",X"01",X"10",X"F6",X"21",X"01",X"4C",X"CB",
		X"76",X"21",X"FD",X"43",X"28",X"02",X"2E",X"E9",X"7A",X"D1",X"E6",X"F0",X"20",X"2A",X"1A",X"E6",
		X"F0",X"28",X"25",X"13",X"1A",X"A7",X"20",X"21",X"1B",X"E5",X"21",X"1B",X"4C",X"3A",X"01",X"4C",
		X"E6",X"40",X"28",X"01",X"23",X"34",X"D5",X"C5",X"CD",X"09",X"07",X"0E",X"60",X"CD",X"21",X"19",
		X"21",X"01",X"4C",X"CB",X"A6",X"C1",X"D1",X"E1",X"13",X"D5",X"CD",X"57",X"1A",X"E1",X"E5",X"11",
		X"05",X"4D",X"06",X"03",X"1A",X"BE",X"38",X"09",X"20",X"04",X"2B",X"1B",X"10",X"F6",X"E1",X"18",
		X"14",X"E1",X"11",X"05",X"4D",X"C5",X"01",X"03",X"00",X"ED",X"B8",X"C1",X"11",X"05",X"4D",X"21",
		X"F3",X"43",X"CD",X"57",X"1A",X"E1",X"C9",X"C5",X"01",X"00",X"03",X"1A",X"D7",X"CD",X"69",X"1A",
		X"1A",X"CD",X"69",X"1A",X"1B",X"10",X"F4",X"C1",X"C9",X"E6",X"0F",X"20",X"08",X"CB",X"41",X"20",
		X"06",X"3E",X"20",X"18",X"04",X"CB",X"C1",X"C6",X"30",X"77",X"2B",X"C9",X"18",X"4C",X"69",X"88",
		X"86",X"84",X"88",X"0A",X"82",X"80",X"86",X"D1",X"0A",X"80",X"C4",X"C6",X"82",X"02",X"88",X"82",
		X"86",X"C0",X"02",X"C2",X"C1",X"C6",X"12",X"C6",X"42",X"02",X"4A",X"CA",X"82",X"42",X"82",X"8A",
		X"22",X"02",X"20",X"10",X"80",X"12",X"20",X"00",X"08",X"10",X"00",X"08",X"50",X"20",X"08",X"08",
		X"00",X"40",X"00",X"00",X"08",X"00",X"40",X"40",X"80",X"00",X"80",X"28",X"28",X"02",X"42",X"50",
		X"85",X"17",X"85",X"14",X"05",X"23",X"05",X"07",X"13",X"01",X"25",X"05",X"24",X"24",X"81",X"05",
		X"00",X"23",X"05",X"05",X"05",X"05",X"04",X"14",X"85",X"85",X"0E",X"05",X"15",X"8F",X"AC",X"AE",
		X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"01",X"08",X"00",X"20",
		X"00",X"00",X"00",X"10",X"20",X"00",X"40",X"00",X"20",X"18",X"20",X"00",X"08",X"44",X"01",X"70",
		X"8F",X"86",X"83",X"D6",X"86",X"C7",X"02",X"82",X"82",X"83",X"CA",X"42",X"08",X"82",X"82",X"82",
		X"8A",X"87",X"03",X"C6",X"82",X"43",X"CB",X"83",X"86",X"20",X"83",X"06",X"80",X"98",X"80",X"C2",
		X"40",X"80",X"00",X"30",X"40",X"02",X"00",X"00",X"98",X"00",X"20",X"00",X"00",X"08",X"10",X"00",
		X"40",X"00",X"00",X"E0",X"5A",X"00",X"80",X"00",X"02",X"08",X"58",X"C0",X"00",X"00",X"00",X"02",
		X"07",X"05",X"05",X"50",X"57",X"07",X"0C",X"B0",X"05",X"05",X"45",X"17",X"A5",X"04",X"21",X"85",
		X"07",X"27",X"A5",X"0D",X"25",X"2D",X"26",X"20",X"01",X"06",X"87",X"84",X"85",X"8C",X"03",X"37",
		X"48",X"08",X"00",X"20",X"08",X"00",X"00",X"00",X"00",X"28",X"08",X"00",X"01",X"00",X"00",X"30",
		X"20",X"08",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"53",X"20",X"40",X"48",
		X"86",X"CA",X"86",X"EC",X"98",X"83",X"00",X"CE",X"81",X"80",X"9E",X"C2",X"03",X"02",X"8A",X"26",
		X"C2",X"96",X"CA",X"06",X"A3",X"C2",X"01",X"82",X"82",X"02",X"82",X"82",X"86",X"83",X"02",X"C2",
		X"40",X"08",X"82",X"28",X"00",X"20",X"08",X"10",X"20",X"00",X"C8",X"00",X"08",X"02",X"08",X"48",
		X"00",X"08",X"08",X"00",X"60",X"20",X"40",X"00",X"40",X"88",X"42",X"00",X"00",X"00",X"08",X"04",
		X"24",X"05",X"05",X"10",X"B5",X"11",X"A1",X"01",X"05",X"01",X"85",X"15",X"05",X"74",X"31",X"35",
		X"04",X"0C",X"44",X"07",X"07",X"8C",X"0D",X"0C",X"61",X"A5",X"04",X"15",X"1D",X"A7",X"27",X"05",
		X"00",X"08",X"40",X"20",X"00",X"12",X"00",X"20",X"08",X"09",X"80",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"40",X"10",X"20",X"00",X"08",X"00",X"3C",X"00",X"02",X"88",X"20",X"04",X"40",
		X"C3",X"09",X"1C",X"C3",X"0E",X"1D",X"C3",X"5B",X"1E",X"DD",X"21",X"00",X"4D",X"DD",X"CB",X"00",
		X"46",X"20",X"3C",X"3A",X"04",X"4C",X"07",X"D8",X"0E",X"3F",X"3A",X"16",X"4C",X"CB",X"67",X"20",
		X"0C",X"0E",X"0F",X"CB",X"5F",X"20",X"06",X"0E",X"03",X"CB",X"57",X"28",X"05",X"CD",X"0F",X"10",
		X"A1",X"C0",X"3A",X"02",X"4C",X"FE",X"68",X"21",X"50",X"01",X"3E",X"DF",X"38",X"05",X"21",X"52",
		X"03",X"3E",X"F1",X"DD",X"74",X"00",X"26",X"07",X"22",X"D2",X"4F",X"DD",X"77",X"01",X"C9",X"DD",
		X"CB",X"00",X"7E",X"28",X"1C",X"DD",X"35",X"02",X"C0",X"2A",X"D0",X"4F",X"22",X"D4",X"4F",X"2A",
		X"E0",X"4F",X"22",X"E4",X"4F",X"DD",X"CB",X"00",X"BE",X"21",X"D2",X"4F",X"CB",X"9E",X"C3",X"ED",
		X"1C",X"3A",X"03",X"4C",X"FE",X"08",X"30",X"63",X"DD",X"7E",X"01",X"FE",X"D1",X"30",X"5C",X"3A",
		X"02",X"4C",X"01",X"58",X"81",X"DD",X"96",X"01",X"30",X"05",X"ED",X"44",X"01",X"5A",X"83",X"FE",
		X"14",X"30",X"48",X"DD",X"70",X"00",X"79",X"32",X"D2",X"4F",X"2A",X"D4",X"4F",X"22",X"D0",X"4F",
		X"2A",X"E4",X"4F",X"22",X"E0",X"4F",X"E6",X"02",X"F6",X"5C",X"6F",X"26",X"03",X"22",X"D4",X"4F",
		X"3A",X"02",X"4C",X"C6",X"1E",X"6F",X"26",X"20",X"22",X"E4",X"4F",X"DD",X"36",X"02",X"08",X"21",
		X"4A",X"4C",X"7E",X"E6",X"F0",X"F6",X"0D",X"77",X"AF",X"32",X"05",X"4C",X"3A",X"04",X"4C",X"E6",
		X"30",X"F6",X"83",X"32",X"04",X"4C",X"AF",X"32",X"03",X"4C",X"C9",X"DD",X"34",X"02",X"DD",X"7E",
		X"02",X"E6",X"07",X"20",X"08",X"3A",X"D2",X"4F",X"EE",X"04",X"32",X"D2",X"4F",X"DD",X"7E",X"01",
		X"C6",X"02",X"DD",X"CB",X"00",X"4E",X"20",X"02",X"D6",X"04",X"DD",X"77",X"01",X"4F",X"C6",X"1E",
		X"32",X"E2",X"4F",X"79",X"E6",X"F0",X"FE",X"E0",X"C0",X"DD",X"36",X"00",X"00",X"C9",X"D9",X"21",
		X"01",X"4C",X"CB",X"86",X"CD",X"2A",X"02",X"FC",X"40",X"40",X"80",X"04",X"AF",X"32",X"07",X"4D",
		X"CD",X"2A",X"02",X"00",X"C0",X"4F",X"40",X"01",X"CD",X"03",X"07",X"48",X"44",X"1C",X"05",X"CD",
		X"03",X"07",X"4B",X"44",X"1C",X"05",X"CD",X"03",X"07",X"4E",X"44",X"1C",X"02",X"CD",X"03",X"07",
		X"4E",X"46",X"05",X"07",X"21",X"68",X"1D",X"01",X"E0",X"FF",X"7E",X"23",X"A7",X"20",X"06",X"5E",
		X"23",X"56",X"23",X"18",X"08",X"FE",X"24",X"28",X"2F",X"12",X"EB",X"09",X"EB",X"C5",X"06",X"06",
		X"CD",X"24",X"02",X"10",X"FB",X"C1",X"18",X"E2",X"00",X"48",X"42",X"42",X"45",X"57",X"41",X"52",
		X"45",X"00",X"0B",X"42",X"4F",X"46",X"00",X"CE",X"42",X"53",X"4B",X"55",X"4E",X"4B",X"2F",X"53",
		X"20",X"53",X"50",X"52",X"41",X"59",X"21",X"24",X"21",X"68",X"60",X"22",X"02",X"4C",X"3E",X"01",
		X"32",X"04",X"4C",X"3E",X"FF",X"32",X"14",X"4D",X"3E",X"13",X"32",X"D7",X"4F",X"32",X"D9",X"4F",
		X"3E",X"07",X"32",X"D3",X"4F",X"CD",X"03",X"07",X"5E",X"44",X"1C",X"1F",X"CD",X"03",X"07",X"5E",
		X"40",X"1C",X"84",X"CD",X"03",X"07",X"5F",X"44",X"1C",X"16",X"CD",X"2D",X"02",X"5F",X"43",X"72",
		X"70",X"FC",X"FC",X"77",X"75",X"FC",X"FC",X"72",X"70",X"FC",X"FC",X"76",X"74",X"FC",X"FC",X"73",
		X"71",X"FC",X"FC",X"76",X"74",X"24",X"3E",X"1D",X"32",X"16",X"4C",X"21",X"01",X"4C",X"CB",X"C6",
		X"21",X"E8",X"1D",X"22",X"48",X"4C",X"18",X"1A",X"BF",X"40",X"DF",X"40",X"3F",X"41",X"5F",X"41",
		X"BF",X"41",X"DF",X"41",X"3F",X"42",X"5F",X"42",X"BF",X"42",X"DF",X"42",X"3F",X"43",X"5F",X"43",
		X"00",X"00",X"06",X"20",X"CD",X"52",X"1E",X"10",X"FB",X"3E",X"05",X"32",X"04",X"4C",X"06",X"20",
		X"CD",X"52",X"1E",X"10",X"FB",X"3E",X"01",X"32",X"04",X"4C",X"3A",X"03",X"4C",X"FE",X"08",X"38",
		X"05",X"CD",X"52",X"1E",X"18",X"F4",X"AF",X"32",X"00",X"4D",X"32",X"16",X"4C",X"4F",X"3E",X"20",
		X"32",X"E3",X"4F",X"3A",X"04",X"4C",X"07",X"38",X"06",X"CB",X"41",X"20",X"0E",X"18",X"02",X"0E",
		X"FF",X"C5",X"CD",X"09",X"1C",X"CD",X"52",X"1E",X"C1",X"18",X"E8",X"21",X"01",X"4C",X"CB",X"86",
		X"D9",X"C9",X"C5",X"CD",X"03",X"10",X"CD",X"24",X"02",X"C1",X"C9",X"3A",X"05",X"4C",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"4F",X"06",X"00",X"21",X"C1",X"1E",X"09",X"7E",X"A7",X"28",X"48",X"32",X"D6",
		X"4F",X"AF",X"32",X"D8",X"4F",X"2A",X"02",X"4C",X"7C",X"C6",X"20",X"67",X"7D",X"C6",X"1F",X"6F",
		X"22",X"E6",X"4F",X"3A",X"04",X"4C",X"CB",X"67",X"C8",X"3A",X"D0",X"4F",X"E6",X"F0",X"47",X"79",
		X"A7",X"C8",X"FE",X"04",X"38",X"17",X"20",X"0C",X"7C",X"C6",X"05",X"67",X"78",X"F6",X"06",X"32",
		X"D4",X"4F",X"18",X"0D",X"FE",X"08",X"30",X"05",X"AF",X"32",X"D4",X"4F",X"C9",X"78",X"32",X"D4",
		X"4F",X"2D",X"22",X"E4",X"4F",X"C9",X"3A",X"04",X"4C",X"E6",X"30",X"F6",X"09",X"32",X"04",X"4C",
		X"C9",X"B4",X"B6",X"B4",X"B6",X"48",X"4C",X"4C",X"4C",X"B0",X"B2",X"00",X"05",X"20",X"0C",X"01",
		X"01",X"05",X"15",X"21",X"2D",X"00",X"41",X"04",X"20",X"01",X"04",X"01",X"69",X"76",X"65",X"0D",
		X"00",X"84",X"08",X"21",X"00",X"25",X"10",X"11",X"00",X"3D",X"30",X"10",X"4D",X"10",X"21",X"19",
		X"01",X"24",X"3C",X"54",X"01",X"00",X"41",X"05",X"2D",X"9C",X"20",X"80",X"47",X"7F",X"5C",X"75",
		X"9A",X"C0",X"AA",X"8A",X"82",X"D2",X"02",X"A0",X"DA",X"40",X"80",X"02",X"5A",X"0A",X"92",X"42",
		X"86",X"A2",X"E2",X"0A",X"82",X"82",X"80",X"C8",X"02",X"00",X"82",X"42",X"42",X"22",X"0A",X"C0",
		X"E0",X"D4",X"D6",X"0A",X"92",X"82",X"80",X"80",X"80",X"22",X"28",X"02",X"12",X"08",X"A0",X"B2",
		X"12",X"40",X"80",X"9A",X"F0",X"82",X"42",X"8A",X"40",X"82",X"12",X"A0",X"22",X"10",X"82",X"82",
		X"81",X"45",X"0C",X"21",X"21",X"01",X"21",X"04",X"05",X"00",X"61",X"0C",X"20",X"00",X"04",X"04",
		X"0C",X"51",X"21",X"25",X"45",X"09",X"28",X"15",X"29",X"04",X"05",X"0C",X"19",X"01",X"34",X"76",
		X"12",X"09",X"19",X"02",X"21",X"2C",X"01",X"01",X"01",X"05",X"31",X"00",X"00",X"25",X"01",X"05",
		X"30",X"01",X"24",X"01",X"00",X"00",X"25",X"11",X"05",X"00",X"85",X"60",X"55",X"75",X"75",X"4D",
		X"88",X"92",X"80",X"08",X"28",X"A8",X"00",X"58",X"DA",X"02",X"EA",X"02",X"02",X"00",X"42",X"00",
		X"02",X"50",X"42",X"40",X"42",X"80",X"C8",X"00",X"02",X"4A",X"C6",X"02",X"92",X"02",X"32",X"10",
		X"9A",X"80",X"D3",X"24",X"80",X"C0",X"C2",X"C8",X"0A",X"00",X"8A",X"A3",X"23",X"D8",X"88",X"D0",
		X"82",X"12",X"82",X"A0",X"92",X"D0",X"02",X"02",X"E8",X"E2",X"92",X"A2",X"02",X"F2",X"7B",X"40",
		X"40",X"05",X"05",X"00",X"04",X"3D",X"01",X"05",X"01",X"09",X"24",X"60",X"75",X"11",X"27",X"81",
		X"1C",X"15",X"25",X"05",X"01",X"65",X"2D",X"45",X"01",X"01",X"00",X"A9",X"29",X"65",X"65",X"6D",
		X"70",X"27",X"39",X"39",X"15",X"09",X"05",X"01",X"05",X"08",X"0D",X"25",X"21",X"14",X"05",X"0F",
		X"04",X"60",X"14",X"04",X"25",X"11",X"23",X"25",X"19",X"C1",X"08",X"60",X"DF",X"53",X"65",X"59",
		X"3A",X"4A",X"4C",X"CD",X"32",X"20",X"3A",X"4A",X"4C",X"D7",X"CD",X"32",X"20",X"AF",X"32",X"4A",
		X"4C",X"DD",X"21",X"50",X"4C",X"FD",X"21",X"81",X"50",X"CD",X"FD",X"20",X"DD",X"21",X"5C",X"4C",
		X"FD",X"21",X"86",X"50",X"CD",X"FD",X"20",X"DD",X"21",X"68",X"4C",X"FD",X"21",X"8B",X"50",X"C3",
		X"FD",X"20",X"E6",X"0F",X"C8",X"E7",X"5F",X"22",X"56",X"20",X"5B",X"20",X"60",X"20",X"65",X"20",
		X"77",X"20",X"7C",X"20",X"89",X"20",X"9C",X"20",X"A5",X"20",X"C0",X"20",X"C9",X"20",X"CE",X"20",
		X"72",X"20",X"AE",X"20",X"B7",X"20",X"11",X"B0",X"22",X"18",X"0D",X"11",X"B9",X"22",X"18",X"08",
		X"11",X"B9",X"22",X"18",X"03",X"11",X"C4",X"22",X"DD",X"21",X"5C",X"4C",X"FD",X"21",X"86",X"50",
		X"18",X"67",X"11",X"95",X"24",X"18",X"08",X"11",X"D2",X"22",X"18",X"03",X"11",X"D7",X"22",X"DD",
		X"21",X"68",X"4C",X"FD",X"21",X"8B",X"50",X"18",X"50",X"11",X"F8",X"22",X"CD",X"7F",X"20",X"11",
		X"EC",X"22",X"DD",X"21",X"50",X"4C",X"FD",X"21",X"81",X"50",X"18",X"3D",X"CD",X"E5",X"20",X"02",
		X"23",X"28",X"23",X"58",X"23",X"CD",X"E5",X"20",X"87",X"23",X"BE",X"23",X"EA",X"23",X"CD",X"E5",
		X"20",X"B8",X"24",X"E4",X"24",X"08",X"25",X"CD",X"E5",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"E5",X"20",X"00",X"00",X"00",X"00",X"64",X"24",X"11",X"7B",X"24",X"18",X"B1",X"11",X"88",
		X"24",X"CD",X"68",X"20",X"11",X"00",X"00",X"18",X"B9",X"CD",X"7B",X"22",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"C3",X"77",X"21",X"E1",X"5E",X"23",X"56",X"23",X"E5",X"CD",X"92",X"20",X"E1",X"5E",
		X"23",X"56",X"23",X"E5",X"CD",X"68",X"20",X"E1",X"5E",X"23",X"56",X"18",X"82",X"DD",X"7E",X"02",
		X"A7",X"C8",X"DD",X"7E",X"09",X"A7",X"28",X"27",X"3D",X"47",X"E6",X"0F",X"20",X"1E",X"DD",X"7E",
		X"04",X"CB",X"78",X"20",X"0B",X"E6",X"0F",X"FE",X"0F",X"28",X"0B",X"DD",X"34",X"04",X"18",X"06",
		X"A7",X"28",X"03",X"DD",X"35",X"04",X"78",X"D7",X"E6",X"07",X"B0",X"47",X"DD",X"70",X"09",X"DD",
		X"7E",X"0A",X"A7",X"28",X"3C",X"3D",X"47",X"E6",X"0F",X"20",X"33",X"DD",X"5E",X"05",X"DD",X"7E",
		X"06",X"D7",X"B3",X"5F",X"DD",X"56",X"07",X"DD",X"7E",X"08",X"D7",X"B2",X"57",X"62",X"6B",X"CB",
		X"78",X"20",X"04",X"CB",X"23",X"CB",X"12",X"CB",X"23",X"CB",X"12",X"19",X"EB",X"CB",X"2A",X"CB",
		X"1B",X"CB",X"2A",X"CB",X"1B",X"CD",X"60",X"22",X"78",X"D7",X"E6",X"07",X"B0",X"47",X"DD",X"70",
		X"0A",X"DD",X"35",X"02",X"C2",X"3B",X"22",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7E",X"23",X"47",
		X"D7",X"E6",X"0F",X"20",X"1B",X"78",X"E6",X"0F",X"20",X"06",X"CD",X"7B",X"22",X"C3",X"3B",X"22",
		X"3D",X"20",X"05",X"7E",X"23",X"66",X"6F",X"E9",X"78",X"E6",X"01",X"DD",X"77",X"0B",X"18",X"DD",
		X"3D",X"20",X"1D",X"78",X"E6",X"0F",X"47",X"3A",X"4C",X"4C",X"DD",X"AE",X"0B",X"E6",X"03",X"FE",
		X"03",X"20",X"02",X"CB",X"00",X"DD",X"70",X"02",X"DD",X"75",X"00",X"DD",X"74",X"01",X"18",X"7B",
		X"CB",X"78",X"20",X"11",X"E5",X"DD",X"E5",X"E1",X"23",X"23",X"16",X"00",X"5F",X"19",X"78",X"E6",
		X"0F",X"77",X"E1",X"18",X"A8",X"CB",X"70",X"20",X"28",X"78",X"E6",X"0F",X"D7",X"4F",X"CB",X"68",
		X"20",X"13",X"78",X"E6",X"07",X"B1",X"CB",X"60",X"20",X"05",X"DD",X"77",X"09",X"18",X"8E",X"DD",
		X"77",X"0A",X"C3",X"7D",X"21",X"DD",X"7E",X"0B",X"E6",X"0F",X"B1",X"DD",X"77",X"0B",X"C3",X"7D",
		X"21",X"E5",X"21",X"2F",X"22",X"78",X"E6",X"0F",X"5F",X"16",X"00",X"19",X"5E",X"16",X"00",X"78",
		X"D7",X"E6",X"03",X"28",X"07",X"47",X"CB",X"23",X"CB",X"12",X"10",X"FA",X"CD",X"60",X"22",X"E1",
		X"DD",X"7E",X"0B",X"D7",X"E6",X"0F",X"CA",X"7D",X"21",X"DD",X"77",X"04",X"C3",X"7D",X"21",X"78",
		X"80",X"87",X"90",X"96",X"A0",X"AA",X"B4",X"C0",X"C8",X"D8",X"E1",X"DD",X"7E",X"03",X"FD",X"77",
		X"04",X"DD",X"7E",X"04",X"FD",X"77",X"14",X"DD",X"E5",X"D1",X"7B",X"FE",X"50",X"20",X"02",X"FD",
		X"2B",X"06",X"04",X"DD",X"7E",X"08",X"FD",X"77",X"13",X"DD",X"2B",X"FD",X"2B",X"10",X"F4",X"C9",
		X"7B",X"E6",X"0F",X"DD",X"77",X"05",X"7B",X"D7",X"E6",X"0F",X"DD",X"77",X"06",X"7A",X"E6",X"0F",
		X"DD",X"77",X"07",X"7A",X"D7",X"E6",X"0F",X"DD",X"77",X"08",X"C9",X"AF",X"06",X"0C",X"DD",X"E5",
		X"E1",X"77",X"23",X"10",X"FC",X"C9",X"AF",X"32",X"4F",X"4C",X"21",X"14",X"24",X"22",X"50",X"4C",
		X"C3",X"77",X"21",X"21",X"4F",X"4C",X"7E",X"34",X"07",X"5F",X"16",X"00",X"21",X"AA",X"22",X"19",
		X"5E",X"23",X"56",X"ED",X"53",X"50",X"4C",X"C3",X"77",X"21",X"24",X"24",X"33",X"24",X"42",X"24",
		X"27",X"3F",X"51",X"18",X"25",X"89",X"91",X"1F",X"00",X"3F",X"61",X"99",X"16",X"30",X"12",X"61",
		X"91",X"3F",X"1A",X"00",X"27",X"3F",X"58",X"99",X"16",X"30",X"12",X"26",X"3F",X"68",X"9A",X"1F",
		X"1F",X"00",X"3F",X"6D",X"99",X"18",X"00",X"52",X"89",X"25",X"3C",X"1C",X"24",X"3C",X"1C",X"25",
		X"3C",X"1C",X"24",X"3C",X"1C",X"25",X"3C",X"1C",X"24",X"3C",X"1C",X"00",X"25",X"38",X"6A",X"9A",
		X"18",X"18",X"6A",X"50",X"40",X"18",X"18",X"00",X"27",X"3F",X"4E",X"14",X"24",X"40",X"54",X"91",
		X"1F",X"00",X"03",X"22",X"89",X"AB",X"E7",X"14",X"E7",X"1C",X"E7",X"14",X"E9",X"1C",X"EB",X"18",
		X"30",X"14",X"E7",X"14",X"F0",X"14",X"EB",X"18",X"E7",X"14",X"E7",X"14",X"E2",X"18",X"E0",X"14",
		X"E2",X"14",X"E6",X"1C",X"E7",X"18",X"18",X"00",X"03",X"27",X"89",X"AC",X"C7",X"14",X"C5",X"14",
		X"30",X"14",X"C4",X"14",X"C7",X"14",X"C9",X"14",X"CB",X"14",X"D0",X"14",X"CB",X"14",X"D2",X"14",
		X"30",X"14",X"D4",X"14",X"C7",X"14",X"D2",X"18",X"D7",X"14",X"DB",X"18",X"E0",X"18",X"DB",X"14",
		X"D9",X"14",X"30",X"18",X"D7",X"18",X"18",X"00",X"03",X"89",X"AC",X"C4",X"14",X"C2",X"14",X"30",
		X"14",X"C0",X"14",X"C7",X"14",X"C5",X"14",X"C2",X"14",X"C0",X"14",X"C2",X"14",X"C2",X"14",X"30",
		X"14",X"C4",X"14",X"C4",X"14",X"CB",X"18",X"D0",X"14",X"D2",X"18",X"D4",X"18",X"C7",X"14",X"C7",
		X"14",X"30",X"18",X"C7",X"18",X"18",X"00",X"03",X"22",X"89",X"AB",X"F0",X"14",X"F0",X"14",X"E7",
		X"14",X"E7",X"14",X"F0",X"1C",X"F2",X"14",X"F4",X"14",X"F2",X"14",X"F0",X"14",X"EA",X"14",X"E7",
		X"18",X"E7",X"13",X"E5",X"12",X"E4",X"13",X"E7",X"14",X"EB",X"14",X"F2",X"14",X"30",X"14",X"E9",
		X"18",X"E2",X"18",X"E4",X"14",X"E7",X"14",X"F0",X"18",X"18",X"18",X"01",X"86",X"22",X"03",X"21",
		X"AC",X"D7",X"14",X"D5",X"14",X"D4",X"14",X"D2",X"14",X"D4",X"1C",X"D5",X"14",X"D7",X"14",X"D9",
		X"14",X"30",X"14",X"D7",X"18",X"E0",X"14",X"30",X"18",X"E2",X"1C",X"E4",X"14",X"E5",X"18",X"30",
		X"14",X"EB",X"14",X"F0",X"18",X"18",X"30",X"18",X"18",X"00",X"03",X"27",X"8A",X"AC",X"D0",X"14",
		X"CA",X"14",X"30",X"18",X"C7",X"1C",X"CA",X"14",X"D2",X"14",X"D2",X"14",X"30",X"14",X"C7",X"18",
		X"CA",X"14",X"D0",X"14",X"30",X"14",X"C7",X"14",X"C9",X"14",X"CB",X"14",X"C5",X"18",X"CB",X"18",
		X"D0",X"18",X"18",X"00",X"03",X"8A",X"A9",X"23",X"E0",X"18",X"E0",X"18",X"F0",X"14",X"E7",X"14",
		X"18",X"01",X"93",X"22",X"30",X"14",X"E5",X"14",X"E6",X"14",X"E7",X"14",X"EA",X"18",X"EA",X"18",
		X"01",X"8A",X"22",X"30",X"14",X"F4",X"14",X"F2",X"14",X"F0",X"14",X"EA",X"18",X"F0",X"18",X"01",
		X"8A",X"22",X"30",X"14",X"EA",X"14",X"E9",X"14",X"E7",X"14",X"E5",X"14",X"E7",X"14",X"E4",X"14",
		X"E0",X"14",X"E0",X"14",X"E4",X"18",X"E5",X"1C",X"E7",X"1C",X"EB",X"18",X"F4",X"14",X"F0",X"18",
		X"18",X"01",X"86",X"22",X"26",X"3F",X"6B",X"99",X"18",X"6A",X"58",X"18",X"6A",X"50",X"18",X"69",
		X"58",X"18",X"69",X"50",X"18",X"68",X"58",X"18",X"68",X"18",X"00",X"26",X"3F",X"58",X"99",X"89",
		X"18",X"24",X"3F",X"58",X"80",X"92",X"18",X"00",X"27",X"AF",X"91",X"89",X"C0",X"18",X"D0",X"18",
		X"E0",X"18",X"F0",X"18",X"00",X"27",X"3F",X"52",X"92",X"18",X"24",X"1C",X"00",X"21",X"B8",X"24",
		X"22",X"50",X"4C",X"C3",X"77",X"21",X"21",X"E4",X"24",X"22",X"5C",X"4C",X"C3",X"77",X"21",X"21",
		X"08",X"25",X"22",X"68",X"4C",X"C3",X"77",X"21",X"03",X"22",X"89",X"AA",X"F0",X"14",X"F0",X"14",
		X"30",X"18",X"18",X"E0",X"18",X"E4",X"14",X"E5",X"14",X"8A",X"E7",X"18",X"18",X"18",X"89",X"F0",
		X"14",X"F0",X"14",X"30",X"18",X"18",X"E0",X"18",X"E7",X"14",X"F0",X"14",X"8A",X"F7",X"18",X"18",
		X"18",X"01",X"9D",X"24",X"03",X"89",X"AC",X"E0",X"14",X"DB",X"14",X"D9",X"14",X"D7",X"1C",X"18",
		X"E0",X"18",X"E0",X"18",X"18",X"18",X"E7",X"14",X"E4",X"14",X"E0",X"14",X"D7",X"1C",X"18",X"E7",
		X"18",X"E7",X"18",X"18",X"18",X"01",X"A6",X"24",X"03",X"26",X"89",X"AF",X"99",X"14",X"C0",X"14",
		X"18",X"18",X"C0",X"18",X"C0",X"18",X"18",X"18",X"14",X"C0",X"14",X"01",X"AF",X"24",X"C2",X"80",
		X"80",X"00",X"80",X"24",X"00",X"40",X"10",X"00",X"00",X"00",X"42",X"12",X"00",X"82",X"00",X"B0",
		X"90",X"00",X"28",X"00",X"00",X"80",X"82",X"A2",X"00",X"08",X"00",X"12",X"00",X"00",X"10",X"10",
		X"08",X"05",X"04",X"0F",X"04",X"45",X"05",X"01",X"05",X"0D",X"45",X"49",X"04",X"19",X"05",X"01",
		X"11",X"05",X"A5",X"05",X"05",X"0C",X"85",X"5D",X"09",X"49",X"05",X"05",X"05",X"07",X"97",X"5C",
		X"00",X"01",X"00",X"01",X"21",X"04",X"01",X"10",X"01",X"00",X"00",X"40",X"01",X"01",X"48",X"00",
		X"00",X"00",X"1C",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"10",X"00",X"44",X"45",X"50",X"44",
		X"83",X"A2",X"92",X"AA",X"A2",X"86",X"82",X"B0",X"AA",X"E0",X"A6",X"90",X"92",X"02",X"22",X"92",
		X"80",X"02",X"82",X"81",X"C2",X"42",X"02",X"86",X"92",X"00",X"86",X"A2",X"40",X"42",X"80",X"92",
		X"A0",X"A2",X"A0",X"22",X"00",X"00",X"00",X"02",X"82",X"30",X"20",X"00",X"10",X"00",X"10",X"20",
		X"00",X"22",X"00",X"A0",X"80",X"00",X"02",X"00",X"00",X"02",X"00",X"A2",X"92",X"A0",X"00",X"10",
		X"01",X"01",X"04",X"20",X"04",X"E5",X"26",X"04",X"05",X"05",X"05",X"05",X"25",X"0C",X"C0",X"0D",
		X"05",X"05",X"04",X"06",X"05",X"00",X"44",X"41",X"11",X"05",X"08",X"84",X"91",X"CF",X"8D",X"DD",
		X"00",X"04",X"00",X"00",X"01",X"00",X"01",X"41",X"0C",X"40",X"48",X"00",X"00",X"00",X"00",X"01",
		X"00",X"01",X"01",X"04",X"00",X"09",X"09",X"40",X"00",X"00",X"85",X"01",X"01",X"4C",X"0E",X"49",
		X"82",X"50",X"32",X"BA",X"A2",X"82",X"B0",X"B2",X"D2",X"80",X"82",X"B1",X"92",X"88",X"D2",X"C2",
		X"1A",X"02",X"8B",X"82",X"68",X"C2",X"8A",X"8A",X"A6",X"82",X"82",X"02",X"82",X"B2",X"6A",X"96",
		X"A8",X"68",X"00",X"01",X"10",X"00",X"02",X"00",X"90",X"10",X"00",X"40",X"A2",X"10",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"02",X"00",X"10",X"08",X"60",X"08",X"18",X"00",
		X"14",X"3D",X"C5",X"8C",X"01",X"05",X"54",X"01",X"47",X"05",X"89",X"11",X"03",X"06",X"05",X"0C",
		X"07",X"05",X"05",X"01",X"11",X"25",X"05",X"85",X"B4",X"09",X"21",X"85",X"4D",X"37",X"13",X"0C",
		X"29",X"40",X"00",X"08",X"40",X"00",X"01",X"00",X"41",X"00",X"00",X"00",X"01",X"00",X"21",X"00",
		X"04",X"00",X"08",X"01",X"28",X"01",X"04",X"01",X"00",X"01",X"00",X"04",X"01",X"04",X"08",X"04",
		X"E3",X"83",X"A2",X"8A",X"B2",X"2A",X"98",X"C2",X"A2",X"9A",X"CE",X"02",X"82",X"A2",X"83",X"82",
		X"82",X"22",X"92",X"82",X"83",X"80",X"E0",X"82",X"92",X"8A",X"82",X"92",X"12",X"80",X"B2",X"82",
		X"14",X"B0",X"02",X"30",X"20",X"80",X"02",X"00",X"00",X"C2",X"22",X"00",X"82",X"30",X"00",X"A2",
		X"00",X"00",X"00",X"02",X"10",X"82",X"00",X"00",X"00",X"10",X"80",X"00",X"00",X"10",X"00",X"08",
		X"01",X"15",X"05",X"25",X"14",X"80",X"04",X"09",X"15",X"25",X"5D",X"35",X"40",X"4B",X"25",X"00",
		X"04",X"0C",X"5D",X"45",X"25",X"09",X"0D",X"05",X"45",X"05",X"40",X"14",X"17",X"94",X"11",X"81",
		X"08",X"08",X"00",X"01",X"40",X"00",X"14",X"00",X"01",X"00",X"00",X"00",X"30",X"00",X"04",X"18",
		X"00",X"40",X"08",X"04",X"00",X"00",X"00",X"05",X"08",X"04",X"00",X"44",X"05",X"09",X"08",X"08",
		X"C3",X"F7",X"29",X"C3",X"91",X"2A",X"C3",X"7D",X"2B",X"C3",X"E0",X"2A",X"C3",X"33",X"27",X"21",
		X"00",X"4C",X"CB",X"5E",X"20",X"10",X"CB",X"DE",X"21",X"00",X"00",X"22",X"10",X"4C",X"CD",X"58",
		X"2E",X"CD",X"00",X"07",X"04",X"C9",X"3A",X"11",X"4C",X"FE",X"02",X"C0",X"21",X"00",X"00",X"22",
		X"00",X"4C",X"C9",X"3A",X"00",X"4C",X"E6",X"07",X"E7",X"43",X"27",X"AE",X"27",X"C6",X"27",X"2A",
		X"28",X"0C",X"30",X"CD",X"27",X"02",X"3E",X"1D",X"32",X"16",X"4C",X"3E",X"FF",X"32",X"14",X"4D",
		X"CD",X"00",X"07",X"00",X"21",X"00",X"00",X"22",X"10",X"4C",X"21",X"E0",X"B8",X"22",X"02",X"4C",
		X"21",X"0D",X"00",X"22",X"04",X"4C",X"3E",X"08",X"32",X"D7",X"4F",X"32",X"D9",X"4F",X"3E",X"06",
		X"32",X"DB",X"4F",X"32",X"DD",X"4F",X"3E",X"D8",X"21",X"E7",X"4F",X"06",X"04",X"77",X"23",X"23",
		X"10",X"FB",X"CD",X"03",X"07",X"4C",X"44",X"1C",X"06",X"CD",X"03",X"07",X"4F",X"44",X"1C",X"06",
		X"CD",X"03",X"07",X"52",X"44",X"1C",X"07",X"CD",X"03",X"07",X"55",X"44",X"1C",X"07",X"CD",X"03",
		X"07",X"58",X"44",X"1C",X"05",X"CD",X"03",X"07",X"5B",X"44",X"1C",X"05",X"18",X"13",X"CD",X"03",
		X"10",X"CD",X"14",X"28",X"C6",X"EF",X"32",X"EA",X"4F",X"FE",X"87",X"C0",X"3E",X"05",X"32",X"04",
		X"4C",X"21",X"00",X"4C",X"34",X"C9",X"CD",X"03",X"10",X"CD",X"14",X"28",X"20",X"04",X"21",X"02",
		X"4C",X"35",X"C6",X"E7",X"32",X"EA",X"4F",X"C6",X"10",X"32",X"EC",X"4F",X"FE",X"0F",X"28",X"E1",
		X"3A",X"02",X"4C",X"FE",X"18",X"D8",X"47",X"07",X"D8",X"E6",X"0E",X"C0",X"CD",X"F7",X"27",X"3A",
		X"02",X"4C",X"ED",X"44",X"C6",X"C8",X"47",X"78",X"07",X"07",X"57",X"E6",X"E0",X"5F",X"7A",X"E6",
		X"03",X"57",X"21",X"63",X"44",X"19",X"78",X"0F",X"0F",X"0F",X"E6",X"07",X"3C",X"06",X"07",X"77",
		X"23",X"10",X"FC",X"C9",X"3A",X"D6",X"4F",X"EE",X"02",X"32",X"DA",X"4F",X"3A",X"D8",X"4F",X"EE",
		X"02",X"32",X"DC",X"4F",X"3A",X"02",X"4C",X"ED",X"44",X"C9",X"3A",X"01",X"4C",X"CB",X"47",X"20",
		X"15",X"21",X"9C",X"29",X"22",X"48",X"4C",X"3C",X"32",X"01",X"4C",X"21",X"D6",X"4F",X"06",X"08",
		X"0E",X"00",X"71",X"23",X"10",X"FC",X"CB",X"67",X"C2",X"28",X"29",X"47",X"E6",X"0E",X"4F",X"0F",
		X"81",X"4F",X"78",X"0F",X"E6",X"07",X"E7",X"65",X"28",X"81",X"28",X"9B",X"28",X"AC",X"28",X"BD",
		X"28",X"F3",X"28",X"6E",X"29",X"21",X"90",X"13",X"22",X"D6",X"4F",X"2E",X"92",X"22",X"D8",X"4F",
		X"21",X"C7",X"A8",X"22",X"E6",X"4F",X"2E",X"B7",X"22",X"E8",X"4F",X"21",X"AE",X"29",X"C3",X"15",
		X"29",X"21",X"60",X"62",X"22",X"CE",X"42",X"21",X"66",X"64",X"22",X"EE",X"42",X"21",X"02",X"02",
		X"22",X"CE",X"46",X"22",X"EE",X"46",X"21",X"BA",X"29",X"18",X"7A",X"21",X"C0",X"01",X"22",X"DA",
		X"4F",X"21",X"BF",X"78",X"22",X"EA",X"4F",X"21",X"C4",X"29",X"18",X"69",X"21",X"C0",X"05",X"22",
		X"DC",X"4F",X"21",X"BF",X"60",X"22",X"EC",X"4F",X"21",X"D2",X"29",X"18",X"58",X"C5",X"CD",X"2D",
		X"02",X"F7",X"42",X"C3",X"C2",X"24",X"CD",X"2D",X"02",X"18",X"43",X"C1",X"7A",X"78",X"C0",X"24",
		X"CD",X"2D",X"02",X"F9",X"42",X"C5",X"C4",X"24",X"CD",X"03",X"07",X"D7",X"46",X"02",X"0F",X"CD",
		X"03",X"07",X"D9",X"46",X"02",X"0F",X"CD",X"03",X"07",X"B8",X"46",X"04",X"0F",X"C1",X"21",X"E0",
		X"29",X"18",X"22",X"C5",X"CD",X"2D",X"02",X"FB",X"42",X"72",X"70",X"24",X"CD",X"03",X"07",X"DB",
		X"46",X"02",X"16",X"CD",X"03",X"07",X"BA",X"42",X"04",X"84",X"CD",X"03",X"07",X"BA",X"46",X"04",
		X"1F",X"C1",X"21",X"EC",X"29",X"22",X"02",X"4C",X"21",X"01",X"4C",X"CB",X"E6",X"21",X"2C",X"42",
		X"06",X"00",X"09",X"22",X"04",X"4C",X"18",X"2D",X"3A",X"10",X"4C",X"E6",X"03",X"C0",X"2A",X"02",
		X"4C",X"7E",X"FE",X"24",X"28",X"11",X"23",X"22",X"02",X"4C",X"2A",X"04",X"4C",X"77",X"11",X"E0",
		X"FF",X"19",X"22",X"04",X"4C",X"18",X"0E",X"3A",X"01",X"4C",X"E6",X"EF",X"C6",X"02",X"32",X"01",
		X"4C",X"FE",X"0D",X"30",X"14",X"3A",X"10",X"4C",X"E6",X"0F",X"C0",X"21",X"D6",X"4F",X"06",X"04",
		X"7E",X"EE",X"04",X"77",X"23",X"23",X"10",X"F8",X"C9",X"3E",X"60",X"32",X"02",X"4C",X"3A",X"10",
		X"4C",X"E6",X"03",X"C0",X"11",X"20",X"00",X"06",X"12",X"21",X"E3",X"44",X"C5",X"06",X"07",X"E5",
		X"7E",X"E6",X"07",X"3C",X"77",X"23",X"10",X"FC",X"E1",X"19",X"C1",X"10",X"EF",X"CD",X"55",X"29",
		X"21",X"02",X"4C",X"35",X"C0",X"21",X"04",X"00",X"22",X"00",X"4C",X"C9",X"CE",X"42",X"CF",X"42",
		X"EE",X"42",X"EF",X"42",X"D8",X"42",X"DB",X"42",X"F8",X"42",X"FB",X"42",X"00",X"00",X"42",X"49",
		X"52",X"44",X"49",X"59",X"20",X"4D",X"41",X"4D",X"41",X"24",X"42",X"41",X"42",X"59",X"20",X"42",
		X"49",X"52",X"44",X"24",X"4D",X"4F",X"4E",X"53",X"54",X"45",X"52",X"20",X"52",X"41",X"54",X"20",
		X"41",X"24",X"4D",X"4F",X"4E",X"53",X"54",X"45",X"52",X"20",X"52",X"41",X"54",X"20",X"42",X"24",
		X"43",X"41",X"54",X"45",X"52",X"50",X"49",X"4C",X"4C",X"45",X"52",X"24",X"45",X"41",X"52",X"54",
		X"48",X"20",X"57",X"4F",X"52",X"4D",X"24",X"21",X"00",X"4C",X"CB",X"5E",X"20",X"36",X"CB",X"DE",
		X"21",X"FC",X"FC",X"22",X"ED",X"41",X"22",X"0D",X"42",X"21",X"87",X"98",X"22",X"E6",X"4F",X"2E",
		X"7F",X"22",X"E8",X"4F",X"3E",X"02",X"32",X"D7",X"4F",X"32",X"D9",X"4F",X"3E",X"1C",X"32",X"D6",
		X"4F",X"AF",X"32",X"D8",X"4F",X"32",X"18",X"4C",X"21",X"00",X"00",X"22",X"10",X"4C",X"3E",X"08",
		X"32",X"4A",X"4C",X"C9",X"3A",X"10",X"4C",X"E6",X"0F",X"C0",X"21",X"18",X"4C",X"7E",X"34",X"FE",
		X"0D",X"28",X"36",X"5F",X"16",X"00",X"21",X"80",X"2A",X"19",X"7E",X"32",X"D6",X"4F",X"FE",X"34",
		X"D8",X"20",X"08",X"3E",X"8F",X"32",X"E6",X"4F",X"7E",X"18",X"18",X"47",X"7B",X"FE",X"06",X"38",
		X"11",X"D6",X"06",X"0F",X"38",X"0C",X"5F",X"21",X"8D",X"2A",X"19",X"7E",X"32",X"D7",X"4F",X"32",
		X"D9",X"4F",X"78",X"C6",X"02",X"32",X"D8",X"4F",X"C9",X"21",X"00",X"4C",X"CB",X"9E",X"34",X"C9",
		X"20",X"34",X"38",X"3C",X"40",X"3C",X"40",X"94",X"90",X"94",X"90",X"94",X"90",X"04",X"07",X"06",
		X"13",X"3A",X"00",X"4C",X"FE",X"50",X"30",X"07",X"21",X"20",X"00",X"22",X"00",X"4C",X"C9",X"21",
		X"1B",X"4C",X"11",X"78",X"4C",X"DD",X"21",X"0A",X"4D",X"3A",X"01",X"4C",X"E6",X"40",X"28",X"06",
		X"23",X"13",X"DD",X"21",X"0E",X"4D",X"AF",X"06",X"04",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F9",
		X"34",X"1A",X"3C",X"47",X"E6",X"1C",X"FE",X"14",X"38",X"04",X"78",X"C6",X"0C",X"47",X"78",X"12",
		X"E6",X"03",X"FE",X"02",X"CC",X"03",X"1C",X"21",X"00",X"4C",X"36",X"50",X"23",X"CB",X"86",X"C9",
		X"3A",X"00",X"4C",X"FE",X"50",X"38",X"05",X"3E",X"0A",X"32",X"4A",X"4C",X"3E",X"02",X"32",X"4C",
		X"4C",X"CD",X"2D",X"02",X"6B",X"42",X"54",X"49",X"4D",X"45",X"20",X"4F",X"55",X"54",X"24",X"CD",
		X"03",X"07",X"8B",X"45",X"08",X"05",X"21",X"FC",X"FC",X"22",X"ED",X"41",X"22",X"0D",X"42",X"21",
		X"28",X"0D",X"22",X"DC",X"4F",X"21",X"86",X"98",X"22",X"EC",X"4F",X"21",X"04",X"4C",X"7E",X"E6",
		X"30",X"F6",X"81",X"77",X"21",X"DC",X"4F",X"06",X"08",X"C5",X"06",X"10",X"CD",X"72",X"2B",X"10",
		X"FB",X"7E",X"EE",X"04",X"77",X"C1",X"10",X"F1",X"3E",X"24",X"32",X"DC",X"4F",X"3E",X"97",X"32",
		X"ED",X"4F",X"06",X"20",X"CD",X"72",X"2B",X"10",X"FB",X"3E",X"30",X"32",X"DC",X"4F",X"0E",X"94",
		X"79",X"32",X"ED",X"4F",X"FE",X"20",X"38",X"08",X"D6",X"04",X"4F",X"CD",X"72",X"2B",X"18",X"F0",
		X"3E",X"24",X"32",X"DC",X"4F",X"3E",X"0B",X"32",X"4A",X"4C",X"06",X"64",X"CD",X"72",X"2B",X"10",
		X"FB",X"C9",X"E5",X"C5",X"CD",X"03",X"10",X"CD",X"24",X"02",X"C1",X"E1",X"C9",X"11",X"25",X"4C",
		X"21",X"01",X"4C",X"CB",X"76",X"28",X"03",X"11",X"28",X"4C",X"21",X"43",X"4C",X"06",X"05",X"D5",
		X"E5",X"1A",X"BE",X"38",X"1A",X"20",X"0E",X"1B",X"2B",X"1A",X"BE",X"38",X"12",X"20",X"06",X"1B",
		X"2B",X"1A",X"BE",X"38",X"0A",X"E1",X"11",X"FA",X"FF",X"19",X"D1",X"10",X"E2",X"18",X"02",X"E1",
		X"D1",X"78",X"FE",X"05",X"CA",X"51",X"2D",X"32",X"02",X"4C",X"D5",X"E5",X"ED",X"44",X"C6",X"04",
		X"28",X"0F",X"07",X"4F",X"07",X"81",X"4F",X"06",X"00",X"21",X"40",X"4C",X"11",X"46",X"4C",X"ED",
		X"B8",X"E1",X"11",X"07",X"00",X"19",X"22",X"06",X"4C",X"2B",X"D1",X"D5",X"EB",X"01",X"03",X"00",
		X"ED",X"B8",X"2A",X"06",X"4C",X"36",X"59",X"23",X"36",X"4F",X"23",X"36",X"55",X"CD",X"58",X"2E",
		X"D1",X"21",X"C9",X"42",X"CD",X"17",X"2F",X"CD",X"03",X"07",X"42",X"44",X"1C",X"05",X"CD",X"03",
		X"07",X"44",X"44",X"1C",X"05",X"CD",X"03",X"07",X"47",X"44",X"1C",X"03",X"CD",X"03",X"07",X"09",
		X"45",X"03",X"07",X"CD",X"03",X"07",X"09",X"46",X"07",X"02",X"CD",X"03",X"07",X"EB",X"45",X"07",
		X"04",X"21",X"10",X"10",X"22",X"07",X"45",X"22",X"27",X"45",X"22",X"47",X"45",X"22",X"0A",X"45",
		X"22",X"2A",X"45",X"22",X"4A",X"45",X"CD",X"2D",X"02",X"22",X"43",X"45",X"4E",X"54",X"45",X"52",
		X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"2E",X"24",
		X"CD",X"2D",X"02",X"84",X"43",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"57",X"49",X"54",X"48",
		X"20",X"54",X"48",X"45",X"20",X"4A",X"4F",X"59",X"20",X"53",X"54",X"49",X"43",X"4B",X"2E",X"24",
		X"CD",X"2D",X"02",X"E7",X"42",X"59",X"4F",X"55",X"52",X"20",X"53",X"43",X"4F",X"52",X"45",X"24",
		X"CD",X"2D",X"02",X"49",X"41",X"59",X"4F",X"55",X"24",X"CD",X"2D",X"02",X"AB",X"42",X"54",X"49",
		X"4D",X"45",X"20",X"34",X"30",X"24",X"21",X"E4",X"07",X"22",X"D4",X"4F",X"21",X"3F",X"C0",X"22",
		X"E4",X"4F",X"21",X"E0",X"03",X"22",X"D2",X"4F",X"3E",X"BC",X"32",X"E3",X"4F",X"3E",X"20",X"32",
		X"03",X"4C",X"CD",X"BE",X"2D",X"3E",X"40",X"32",X"05",X"4C",X"3E",X"02",X"32",X"4C",X"4C",X"3E",
		X"0E",X"32",X"4A",X"4C",X"06",X"03",X"C5",X"21",X"01",X"4C",X"3A",X"00",X"50",X"CB",X"76",X"28",
		X"03",X"3A",X"40",X"50",X"0F",X"D4",X"6E",X"2D",X"0F",X"D4",X"BE",X"2D",X"0F",X"D4",X"D0",X"2D",
		X"0F",X"D4",X"83",X"2D",X"3A",X"02",X"4C",X"07",X"5F",X"16",X"00",X"21",X"14",X"45",X"19",X"11",
		X"20",X"00",X"06",X"13",X"7E",X"FE",X"01",X"0E",X"01",X"20",X"02",X"0E",X"03",X"71",X"19",X"10",
		X"FC",X"3A",X"03",X"4C",X"C6",X"09",X"6F",X"26",X"45",X"71",X"06",X"14",X"CD",X"24",X"02",X"10",
		X"FB",X"C1",X"10",X"B2",X"3A",X"05",X"4C",X"D6",X"01",X"28",X"27",X"27",X"32",X"05",X"4C",X"4F",
		X"FE",X"10",X"20",X"06",X"3E",X"01",X"32",X"4C",X"4C",X"79",X"E6",X"0F",X"C6",X"30",X"32",X"EB",
		X"41",X"79",X"D7",X"E6",X"0F",X"20",X"04",X"3E",X"20",X"18",X"02",X"C6",X"30",X"32",X"0B",X"42",
		X"18",X"82",X"3E",X"0F",X"32",X"4A",X"4C",X"CD",X"1E",X"27",X"06",X"00",X"CD",X"24",X"02",X"10",
		X"FB",X"3A",X"01",X"4C",X"CB",X"7F",X"28",X"0F",X"CB",X"57",X"20",X"0B",X"21",X"50",X"C4",X"CB",
		X"77",X"28",X"07",X"26",X"84",X"18",X"03",X"21",X"00",X"00",X"22",X"00",X"4C",X"C9",X"F5",X"3A",
		X"03",X"4C",X"C6",X"07",X"5F",X"16",X"41",X"06",X"05",X"1A",X"CD",X"16",X"2E",X"12",X"13",X"10",
		X"F8",X"18",X"13",X"F5",X"3A",X"03",X"4C",X"C6",X"07",X"5F",X"16",X"41",X"06",X"05",X"1A",X"CD",
		X"2C",X"2E",X"12",X"13",X"10",X"F8",X"3A",X"03",X"4C",X"C6",X"09",X"5F",X"16",X"41",X"3A",X"02",
		X"4C",X"07",X"83",X"C6",X"0B",X"6F",X"62",X"1A",X"77",X"7B",X"07",X"07",X"07",X"E6",X"03",X"ED",
		X"44",X"C6",X"02",X"4F",X"06",X"00",X"2A",X"06",X"4C",X"09",X"1A",X"77",X"F1",X"C9",X"F5",X"3A",
		X"03",X"4C",X"FE",X"40",X"28",X"4E",X"CD",X"42",X"2E",X"3A",X"03",X"4C",X"C6",X"20",X"18",X"1B",
		X"F5",X"3A",X"03",X"4C",X"A7",X"20",X"0C",X"3E",X"43",X"32",X"E2",X"4F",X"3E",X"01",X"32",X"05",
		X"4C",X"18",X"31",X"CD",X"42",X"2E",X"3A",X"03",X"4C",X"D6",X"20",X"32",X"03",X"4C",X"5F",X"0F",
		X"0F",X"C6",X"4B",X"32",X"E2",X"4F",X"7B",X"C6",X"09",X"5F",X"16",X"41",X"1A",X"D5",X"CD",X"16",
		X"2E",X"1B",X"12",X"CD",X"16",X"2E",X"1B",X"12",X"D1",X"1A",X"CD",X"2C",X"2E",X"13",X"12",X"CD",
		X"2C",X"2E",X"13",X"12",X"F1",X"C9",X"FE",X"41",X"0E",X"2C",X"28",X"0E",X"FE",X"2C",X"0E",X"2E",
		X"28",X"08",X"FE",X"2E",X"0E",X"5A",X"28",X"02",X"3D",X"4F",X"79",X"C9",X"FE",X"5A",X"0E",X"2E",
		X"28",X"0E",X"FE",X"2E",X"0E",X"2C",X"28",X"08",X"FE",X"2C",X"0E",X"41",X"28",X"02",X"3C",X"4F",
		X"79",X"C9",X"C6",X"07",X"6F",X"26",X"41",X"3E",X"FC",X"77",X"23",X"77",X"23",X"26",X"45",X"36",
		X"07",X"26",X"41",X"23",X"77",X"23",X"77",X"C9",X"21",X"01",X"4C",X"CB",X"86",X"CD",X"2A",X"02",
		X"FC",X"40",X"40",X"80",X"04",X"CD",X"2A",X"02",X"00",X"D0",X"4F",X"20",X"01",X"CD",X"2A",X"02",
		X"07",X"00",X"45",X"60",X"01",X"CD",X"2A",X"02",X"05",X"00",X"46",X"E0",X"01",X"CD",X"2A",X"02",
		X"02",X"00",X"47",X"60",X"01",X"CD",X"03",X"07",X"4D",X"44",X"1C",X"06",X"CD",X"03",X"07",X"51",
		X"44",X"1C",X"03",X"CD",X"2D",X"02",X"91",X"42",X"53",X"43",X"4F",X"52",X"45",X"20",X"20",X"20",
		X"20",X"20",X"4E",X"41",X"4D",X"45",X"24",X"CD",X"2D",X"02",X"CD",X"42",X"54",X"4F",X"44",X"41",
		X"59",X"2F",X"53",X"20",X"42",X"45",X"53",X"54",X"20",X"35",X"24",X"21",X"54",X"43",X"06",X"05",
		X"DD",X"21",X"29",X"4C",X"E5",X"78",X"C5",X"01",X"E0",X"FF",X"ED",X"44",X"C6",X"05",X"5F",X"C6",
		X"31",X"77",X"09",X"E5",X"7B",X"07",X"5F",X"16",X"00",X"21",X"0D",X"2F",X"19",X"EB",X"E1",X"1A",
		X"77",X"13",X"09",X"1A",X"77",X"09",X"09",X"DD",X"E5",X"D1",X"13",X"13",X"CD",X"17",X"2F",X"11",
		X"40",X"FF",X"19",X"DD",X"7E",X"03",X"77",X"09",X"DD",X"7E",X"04",X"77",X"09",X"DD",X"7E",X"05",
		X"77",X"01",X"06",X"00",X"DD",X"09",X"C1",X"E1",X"23",X"23",X"10",X"B8",X"C9",X"53",X"54",X"4E",
		X"44",X"52",X"44",X"54",X"48",X"54",X"48",X"C5",X"01",X"00",X"03",X"1A",X"D7",X"CD",X"2B",X"2F",
		X"1A",X"CD",X"2B",X"2F",X"1B",X"10",X"F4",X"36",X"30",X"C1",X"C9",X"D5",X"E6",X"0F",X"5F",X"B1",
		X"3E",X"20",X"28",X"05",X"0E",X"FF",X"7B",X"C6",X"30",X"77",X"11",X"E0",X"FF",X"19",X"D1",X"C9",
		X"80",X"45",X"0C",X"21",X"20",X"01",X"21",X"40",X"05",X"00",X"41",X"2C",X"20",X"01",X"44",X"04",
		X"4C",X"51",X"21",X"20",X"45",X"09",X"08",X"1D",X"28",X"04",X"85",X"04",X"19",X"00",X"30",X"76",
		X"12",X"09",X"09",X"02",X"21",X"2C",X"01",X"01",X"01",X"05",X"31",X"08",X"00",X"25",X"01",X"05",
		X"10",X"05",X"24",X"01",X"00",X"02",X"25",X"10",X"05",X"00",X"A5",X"60",X"54",X"75",X"75",X"4D",
		X"88",X"92",X"80",X"08",X"20",X"A8",X"00",X"1A",X"DA",X"02",X"EA",X"02",X"02",X"00",X"42",X"00",
		X"02",X"50",X"42",X"00",X"C2",X"80",X"C8",X"00",X"02",X"4A",X"C6",X"02",X"90",X"00",X"32",X"10",
		X"9A",X"80",X"D3",X"A4",X"82",X"C0",X"C2",X"C8",X"00",X"02",X"80",X"23",X"23",X"D8",X"08",X"D0",
		X"82",X"12",X"82",X"20",X"42",X"70",X"02",X"02",X"E8",X"E2",X"90",X"A2",X"02",X"E2",X"22",X"40",
		X"60",X"05",X"0D",X"00",X"08",X"1D",X"01",X"05",X"01",X"09",X"24",X"60",X"75",X"11",X"27",X"81",
		X"1C",X"15",X"25",X"05",X"00",X"65",X"25",X"45",X"01",X"11",X"00",X"E9",X"09",X"65",X"25",X"2D",
		X"50",X"03",X"19",X"3B",X"15",X"08",X"05",X"01",X"05",X"08",X"1D",X"21",X"21",X"14",X"09",X"0D",
		X"00",X"60",X"04",X"04",X"25",X"11",X"33",X"25",X"19",X"C0",X"00",X"40",X"9F",X"13",X"65",X"59",
		X"C3",X"16",X"30",X"C3",X"8C",X"30",X"C3",X"CE",X"30",X"C3",X"18",X"31",X"C3",X"0F",X"30",X"21",
		X"10",X"00",X"22",X"00",X"4C",X"C9",X"21",X"16",X"4C",X"36",X"1D",X"3A",X"00",X"4C",X"E6",X"40",
		X"C4",X"18",X"31",X"CD",X"03",X"07",X"B2",X"40",X"09",X"BF",X"CD",X"03",X"07",X"52",X"42",X"09",
		X"BF",X"3E",X"BF",X"32",X"72",X"40",X"32",X"92",X"43",X"3A",X"7A",X"4C",X"E6",X"02",X"C0",X"11",
		X"8D",X"40",X"CD",X"0F",X"07",X"02",X"FC",X"CD",X"FF",X"20",X"FC",X"FC",X"CD",X"FF",X"FF",X"20",
		X"01",X"FC",X"CC",X"CF",X"FF",X"20",X"01",X"FC",X"FD",X"CC",X"FF",X"20",X"FC",X"FC",X"FD",X"FD",
		X"FF",X"20",X"2E",X"FF",X"CC",X"FD",X"CF",X"20",X"01",X"FC",X"FC",X"CE",X"FF",X"00",X"21",X"2D",
		X"41",X"22",X"06",X"4D",X"2E",X"0D",X"22",X"08",X"4D",X"11",X"D0",X"42",X"CD",X"0F",X"07",X"CD",
		X"FF",X"20",X"CC",X"FF",X"20",X"FD",X"FF",X"20",X"CE",X"CF",X"00",X"C9",X"3A",X"7A",X"4C",X"E6",
		X"02",X"C0",X"11",X"8D",X"44",X"CD",X"0F",X"07",X"03",X"85",X"85",X"20",X"02",X"85",X"85",X"85",
		X"20",X"02",X"8A",X"85",X"85",X"20",X"02",X"8F",X"8A",X"85",X"20",X"83",X"01",X"8F",X"8F",X"87",
		X"20",X"83",X"83",X"8F",X"8F",X"87",X"20",X"03",X"81",X"87",X"00",X"11",X"D0",X"46",X"CD",X"0F",
		X"07",X"86",X"86",X"20",X"91",X"86",X"20",X"83",X"98",X"20",X"83",X"98",X"00",X"C9",X"21",X"7E",
		X"31",X"11",X"0A",X"4D",X"3A",X"01",X"4C",X"CB",X"77",X"28",X"03",X"11",X"0E",X"4D",X"06",X"04",
		X"C5",X"06",X"08",X"0E",X"01",X"AF",X"12",X"C5",X"4E",X"23",X"7E",X"23",X"A7",X"28",X"1F",X"47",
		X"0A",X"FE",X"F0",X"38",X"19",X"3A",X"04",X"4C",X"E6",X"30",X"28",X"0C",X"3A",X"12",X"4D",X"B9",
		X"20",X"06",X"3A",X"13",X"4D",X"B8",X"28",X"06",X"C1",X"1A",X"B1",X"12",X"18",X"01",X"C1",X"CB",
		X"01",X"10",X"D4",X"13",X"C1",X"10",X"C9",X"C9",X"21",X"7E",X"31",X"11",X"0A",X"4D",X"3A",X"01",
		X"4C",X"CB",X"77",X"28",X"03",X"11",X"0E",X"4D",X"DD",X"21",X"BE",X"31",X"3A",X"7A",X"4C",X"0F",
		X"30",X"04",X"DD",X"21",X"C2",X"31",X"06",X"04",X"C5",X"06",X"08",X"1A",X"13",X"DD",X"4E",X"00",
		X"DD",X"23",X"B1",X"C5",X"F5",X"4E",X"23",X"7E",X"23",X"A7",X"20",X"03",X"F1",X"18",X"28",X"47",
		X"F1",X"0F",X"30",X"23",X"F5",X"E5",X"0A",X"67",X"79",X"E6",X"1F",X"FE",X"1F",X"3E",X"FE",X"20",
		X"02",X"3E",X"FC",X"02",X"CB",X"7C",X"20",X"07",X"21",X"20",X"00",X"09",X"77",X"18",X"02",X"03",
		X"02",X"21",X"16",X"4C",X"35",X"E1",X"F1",X"C1",X"10",X"C9",X"C1",X"10",X"BB",X"C9",X"BF",X"40",
		X"3F",X"41",X"BF",X"42",X"3F",X"43",X"BF",X"41",X"3F",X"42",X"82",X"40",X"93",X"40",X"A5",X"40",
		X"A8",X"40",X"B6",X"40",X"CC",X"40",X"0A",X"41",X"26",X"41",X"41",X"41",X"C3",X"41",X"E1",X"41",
		X"C3",X"42",X"41",X"43",X"05",X"43",X"C7",X"42",X"49",X"43",X"0D",X"43",X"73",X"43",X"36",X"43",
		X"B4",X"41",X"77",X"41",X"55",X"42",X"78",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"68",
		X"16",X"00",X"00",X"16",X"C9",X"12",X"00",X"02",X"00",X"00",X"20",X"C0",X"12",X"10",X"00",X"40",
		X"00",X"22",X"90",X"32",X"00",X"20",X"00",X"30",X"80",X"80",X"00",X"00",X"92",X"02",X"00",X"80",
		X"A3",X"3E",X"C2",X"A2",X"82",X"9B",X"A2",X"32",X"9A",X"BA",X"AA",X"B0",X"A2",X"8A",X"AA",X"82",
		X"82",X"92",X"F6",X"92",X"A2",X"32",X"92",X"A2",X"82",X"82",X"00",X"92",X"B2",X"B3",X"F2",X"F6",
		X"50",X"08",X"40",X"55",X"00",X"00",X"00",X"49",X"00",X"04",X"08",X"44",X"04",X"48",X"0C",X"00",
		X"08",X"01",X"08",X"00",X"00",X"00",X"41",X"40",X"00",X"00",X"44",X"40",X"40",X"0C",X"04",X"44",
		X"5D",X"7D",X"47",X"EB",X"4D",X"CD",X"CD",X"25",X"47",X"4F",X"0D",X"4D",X"4D",X"05",X"4D",X"5D",
		X"0D",X"0D",X"05",X"5D",X"4D",X"1D",X"6D",X"4D",X"0D",X"0D",X"C5",X"81",X"44",X"4D",X"0D",X"69",
		X"02",X"20",X"00",X"92",X"80",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"80",X"00",X"20",X"00",
		X"20",X"28",X"A0",X"10",X"10",X"00",X"20",X"00",X"02",X"90",X"82",X"02",X"72",X"22",X"40",X"A0",
		X"82",X"C2",X"D6",X"82",X"A0",X"92",X"82",X"82",X"82",X"82",X"A7",X"B2",X"9E",X"F2",X"B2",X"E2",
		X"B0",X"8A",X"32",X"9A",X"32",X"86",X"91",X"B2",X"AA",X"B3",X"86",X"B2",X"B6",X"B2",X"D3",X"A6",
		X"0D",X"0C",X"61",X"05",X"00",X"00",X"04",X"00",X"40",X"21",X"40",X"04",X"01",X"04",X"00",X"00",
		X"00",X"44",X"40",X"41",X"40",X"40",X"49",X"00",X"08",X"41",X"01",X"40",X"44",X"48",X"00",X"24",
		X"0F",X"6D",X"2D",X"57",X"0D",X"1D",X"9D",X"05",X"45",X"4F",X"4D",X"8D",X"05",X"5D",X"65",X"C5",
		X"45",X"4D",X"4F",X"05",X"05",X"85",X"2D",X"5D",X"1F",X"45",X"45",X"4D",X"5D",X"D5",X"6D",X"1D",
		X"00",X"00",X"00",X"00",X"02",X"00",X"22",X"B8",X"02",X"02",X"02",X"00",X"00",X"02",X"12",X"10",
		X"02",X"00",X"20",X"00",X"C2",X"00",X"00",X"20",X"20",X"82",X"20",X"20",X"A2",X"60",X"82",X"80",
		X"A2",X"92",X"A0",X"9A",X"A2",X"92",X"B6",X"AA",X"D3",X"B2",X"92",X"BA",X"B2",X"F8",X"F2",X"B2",
		X"82",X"A2",X"EA",X"E2",X"E2",X"B2",X"98",X"80",X"B0",X"82",X"A2",X"B2",X"F2",X"A9",X"B2",X"B2",
		X"01",X"15",X"00",X"40",X"00",X"00",X"01",X"08",X"00",X"09",X"08",X"04",X"49",X"41",X"00",X"08",
		X"20",X"00",X"44",X"08",X"04",X"64",X"40",X"44",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",
		X"7D",X"6D",X"6F",X"6D",X"05",X"0D",X"44",X"4D",X"45",X"05",X"55",X"45",X"2D",X"0D",X"65",X"4C",
		X"75",X"55",X"4C",X"25",X"5D",X"05",X"45",X"1D",X"1D",X"B6",X"75",X"15",X"6D",X"45",X"85",X"5D",
		X"00",X"00",X"00",X"02",X"80",X"00",X"00",X"12",X"00",X"40",X"22",X"00",X"10",X"B0",X"02",X"00",
		X"80",X"10",X"80",X"00",X"C0",X"02",X"00",X"90",X"00",X"20",X"00",X"82",X"9A",X"12",X"20",X"22",
		X"DE",X"89",X"92",X"8A",X"9A",X"94",X"A2",X"92",X"A2",X"A2",X"A2",X"92",X"22",X"B3",X"B2",X"86",
		X"BA",X"92",X"82",X"A2",X"82",X"20",X"B6",X"82",X"BA",X"B2",X"A0",X"A3",X"A6",X"EE",X"B6",X"12",
		X"0D",X"0D",X"04",X"08",X"18",X"00",X"04",X"00",X"00",X"00",X"45",X"04",X"28",X"10",X"48",X"00",
		X"00",X"00",X"40",X"05",X"40",X"41",X"40",X"00",X"44",X"00",X"0C",X"11",X"45",X"44",X"04",X"00",
		X"4D",X"6D",X"65",X"05",X"7D",X"45",X"55",X"4D",X"07",X"65",X"06",X"2D",X"44",X"4D",X"0D",X"0D",
		X"DD",X"4C",X"4D",X"C7",X"45",X"4D",X"A5",X"15",X"4D",X"8D",X"05",X"05",X"25",X"25",X"45",X"05",
		X"80",X"28",X"00",X"E0",X"00",X"00",X"02",X"00",X"00",X"02",X"30",X"A2",X"20",X"90",X"42",X"40",
		X"80",X"02",X"10",X"20",X"00",X"00",X"88",X"A0",X"00",X"02",X"20",X"10",X"00",X"9A",X"30",X"00",
		X"92",X"82",X"A2",X"A2",X"B2",X"92",X"8A",X"12",X"B2",X"92",X"92",X"83",X"82",X"92",X"9A",X"B4",
		X"B2",X"B2",X"BA",X"B2",X"A2",X"F8",X"B2",X"B2",X"D2",X"82",X"B1",X"B2",X"B6",X"A3",X"B6",X"EE",
		X"EA",X"80",X"8A",X"10",X"92",X"80",X"82",X"02",X"80",X"A2",X"8C",X"16",X"02",X"F2",X"A2",X"80",
		X"82",X"8A",X"80",X"92",X"A3",X"02",X"02",X"A2",X"30",X"0A",X"DA",X"9A",X"9A",X"82",X"80",X"C2",
		X"42",X"22",X"B2",X"90",X"00",X"00",X"08",X"90",X"80",X"10",X"00",X"90",X"00",X"70",X"1A",X"10",
		X"00",X"40",X"08",X"80",X"A0",X"02",X"10",X"82",X"00",X"12",X"00",X"00",X"80",X"80",X"A0",X"00",
		X"25",X"05",X"05",X"05",X"11",X"05",X"27",X"05",X"15",X"05",X"05",X"41",X"07",X"75",X"35",X"24",
		X"24",X"01",X"87",X"0D",X"08",X"45",X"41",X"06",X"0D",X"0C",X"05",X"08",X"95",X"45",X"DC",X"2B",
		X"04",X"00",X"00",X"04",X"00",X"04",X"01",X"20",X"00",X"00",X"40",X"01",X"84",X"09",X"0D",X"00",
		X"01",X"01",X"05",X"08",X"44",X"04",X"00",X"04",X"01",X"04",X"04",X"24",X"41",X"00",X"44",X"42",
		X"A3",X"93",X"A2",X"82",X"04",X"D2",X"A2",X"C0",X"82",X"12",X"A2",X"86",X"8A",X"A2",X"82",X"82",
		X"B2",X"AE",X"F2",X"9A",X"82",X"82",X"8A",X"D1",X"CA",X"00",X"82",X"92",X"02",X"A2",X"06",X"92",
		X"82",X"E0",X"00",X"80",X"10",X"80",X"22",X"90",X"20",X"00",X"80",X"80",X"00",X"40",X"10",X"1A",
		X"C0",X"00",X"80",X"40",X"00",X"90",X"80",X"80",X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"80",
		X"0C",X"2D",X"05",X"0D",X"B1",X"14",X"21",X"45",X"04",X"45",X"24",X"00",X"05",X"31",X"6C",X"35",
		X"05",X"25",X"79",X"45",X"04",X"05",X"45",X"45",X"25",X"85",X"05",X"04",X"65",X"09",X"2D",X"25",
		X"00",X"01",X"00",X"0D",X"04",X"08",X"05",X"01",X"00",X"04",X"08",X"04",X"01",X"20",X"20",X"05",
		X"00",X"04",X"10",X"00",X"44",X"01",X"05",X"04",X"24",X"04",X"00",X"8C",X"48",X"49",X"4C",X"45",
		X"8A",X"B6",X"82",X"88",X"82",X"82",X"82",X"8A",X"A2",X"32",X"A2",X"88",X"A0",X"C2",X"B2",X"C2",
		X"90",X"98",X"A2",X"C0",X"06",X"82",X"22",X"40",X"A2",X"C6",X"C2",X"C1",X"82",X"31",X"C2",X"80",
		X"80",X"10",X"80",X"30",X"00",X"40",X"10",X"00",X"00",X"00",X"42",X"10",X"20",X"82",X"00",X"B0",
		X"90",X"00",X"28",X"00",X"00",X"00",X"82",X"A2",X"00",X"08",X"00",X"12",X"00",X"02",X"10",X"90",
		X"0C",X"05",X"04",X"0D",X"04",X"45",X"05",X"05",X"05",X"0D",X"45",X"4D",X"04",X"19",X"05",X"05",
		X"11",X"05",X"A5",X"05",X"05",X"1D",X"85",X"5D",X"09",X"49",X"05",X"05",X"05",X"07",X"9F",X"DC",
		X"01",X"41",X"40",X"01",X"21",X"04",X"01",X"00",X"01",X"00",X"00",X"40",X"01",X"01",X"48",X"00",
		X"00",X"00",X"1C",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"00",X"44",X"44",X"40",X"44",
		X"83",X"A2",X"92",X"8A",X"A2",X"82",X"82",X"B0",X"AA",X"E0",X"A6",X"90",X"92",X"02",X"22",X"92",
		X"80",X"02",X"82",X"81",X"C2",X"42",X"82",X"86",X"92",X"80",X"86",X"A2",X"00",X"42",X"80",X"92",
		X"A1",X"A2",X"A0",X"22",X"00",X"00",X"80",X"02",X"82",X"30",X"20",X"00",X"10",X"00",X"10",X"20",
		X"00",X"20",X"00",X"A0",X"80",X"00",X"82",X"00",X"00",X"12",X"00",X"A2",X"92",X"80",X"00",X"10",
		X"01",X"01",X"05",X"00",X"04",X"25",X"26",X"04",X"05",X"05",X"05",X"05",X"25",X"4C",X"C4",X"4D",
		X"05",X"05",X"04",X"07",X"05",X"80",X"44",X"01",X"1D",X"05",X"09",X"04",X"91",X"CF",X"8D",X"DD",
		X"00",X"04",X"00",X"00",X"01",X"00",X"01",X"01",X"0C",X"40",X"48",X"00",X"00",X"00",X"01",X"01",
		X"00",X"01",X"01",X"05",X"00",X"09",X"09",X"40",X"00",X"00",X"85",X"01",X"01",X"4C",X"0E",X"48",
		X"82",X"D2",X"92",X"BA",X"A2",X"82",X"B0",X"B2",X"D2",X"80",X"82",X"B1",X"92",X"88",X"D2",X"EA",
		X"1A",X"02",X"8B",X"82",X"68",X"C2",X"8A",X"8A",X"A6",X"82",X"82",X"02",X"82",X"B2",X"6A",X"96",
		X"A8",X"6A",X"00",X"01",X"10",X"00",X"02",X"00",X"90",X"10",X"00",X"40",X"A2",X"10",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"02",X"20",X"10",X"08",X"40",X"08",X"18",X"00",
		X"14",X"3D",X"C5",X"8C",X"01",X"05",X"54",X"01",X"47",X"05",X"89",X"11",X"07",X"06",X"05",X"0C",
		X"07",X"05",X"05",X"01",X"11",X"25",X"05",X"05",X"14",X"09",X"21",X"85",X"4D",X"37",X"13",X"4C",
		X"29",X"40",X"00",X"08",X"40",X"00",X"01",X"00",X"61",X"00",X"00",X"00",X"01",X"00",X"21",X"00",
		X"04",X"00",X"08",X"01",X"28",X"01",X"04",X"01",X"00",X"01",X"00",X"04",X"01",X"0C",X"08",X"04",
		X"E3",X"83",X"A2",X"8A",X"B2",X"22",X"98",X"C6",X"A2",X"9A",X"CE",X"02",X"82",X"A2",X"83",X"82",
		X"8A",X"22",X"92",X"82",X"83",X"80",X"E2",X"82",X"92",X"8A",X"82",X"92",X"92",X"80",X"B2",X"82",
		X"14",X"A0",X"02",X"32",X"20",X"00",X"02",X"00",X"00",X"C2",X"22",X"00",X"82",X"30",X"00",X"A2",
		X"00",X"00",X"00",X"02",X"10",X"02",X"00",X"00",X"00",X"10",X"80",X"00",X"10",X"10",X"00",X"08",
		X"01",X"15",X"05",X"25",X"14",X"80",X"04",X"0D",X"15",X"65",X"5D",X"25",X"40",X"49",X"25",X"00",
		X"04",X"0C",X"5D",X"45",X"25",X"09",X"0D",X"05",X"45",X"05",X"40",X"14",X"17",X"94",X"35",X"91",
		X"00",X"08",X"00",X"01",X"40",X"00",X"14",X"00",X"01",X"00",X"00",X"00",X"30",X"00",X"04",X"18",
		X"00",X"40",X"08",X"04",X"00",X"00",X"00",X"05",X"08",X"00",X"00",X"44",X"05",X"09",X"08",X"08",
		X"A2",X"82",X"AA",X"30",X"A2",X"82",X"92",X"A2",X"02",X"02",X"CA",X"82",X"88",X"87",X"82",X"38",
		X"C3",X"92",X"B8",X"B2",X"90",X"02",X"80",X"C2",X"00",X"02",X"53",X"C2",X"C2",X"92",X"8A",X"A3",
		X"82",X"22",X"A0",X"12",X"00",X"06",X"00",X"00",X"80",X"08",X"00",X"20",X"20",X"00",X"42",X"00",
		X"08",X"02",X"80",X"00",X"80",X"40",X"00",X"10",X"02",X"10",X"10",X"00",X"30",X"00",X"80",X"00",
		X"55",X"01",X"04",X"48",X"1D",X"09",X"00",X"05",X"09",X"45",X"05",X"0C",X"05",X"25",X"0C",X"14",
		X"14",X"00",X"09",X"07",X"64",X"41",X"7C",X"84",X"81",X"05",X"05",X"05",X"6D",X"47",X"26",X"45",
		X"00",X"00",X"00",X"45",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"48",X"01",X"01",X"04",X"04",X"05",X"00",X"0C",X"00",X"00",X"08",X"40",X"4C",X"00",X"09",X"00",
		X"9E",X"A1",X"92",X"F0",X"02",X"82",X"12",X"90",X"8A",X"9A",X"02",X"A1",X"82",X"02",X"82",X"A4",
		X"90",X"82",X"02",X"02",X"D0",X"42",X"22",X"A0",X"42",X"92",X"82",X"B2",X"E2",X"B2",X"90",X"92",
		X"90",X"84",X"28",X"30",X"80",X"A0",X"10",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"02",X"00",
		X"02",X"10",X"80",X"A0",X"00",X"00",X"20",X"10",X"80",X"02",X"00",X"80",X"00",X"10",X"20",X"00",
		X"25",X"01",X"04",X"04",X"45",X"45",X"05",X"85",X"09",X"05",X"29",X"45",X"05",X"25",X"05",X"05",
		X"15",X"41",X"0C",X"00",X"1D",X"04",X"45",X"07",X"91",X"C4",X"41",X"0D",X"1E",X"04",X"61",X"1F",
		X"19",X"01",X"0C",X"08",X"6C",X"05",X"00",X"04",X"01",X"00",X"01",X"0D",X"08",X"00",X"04",X"41",
		X"0C",X"14",X"08",X"00",X"00",X"00",X"0C",X"01",X"00",X"04",X"40",X"00",X"41",X"41",X"45",X"4D",
		X"9A",X"02",X"8C",X"02",X"02",X"84",X"80",X"00",X"A2",X"42",X"82",X"E2",X"80",X"0E",X"84",X"02",
		X"80",X"02",X"C0",X"0A",X"82",X"86",X"82",X"CF",X"00",X"C2",X"42",X"88",X"40",X"42",X"82",X"80",
		X"40",X"10",X"08",X"00",X"00",X"10",X"04",X"40",X"00",X"40",X"00",X"02",X"60",X"00",X"12",X"00",
		X"C0",X"00",X"00",X"58",X"10",X"40",X"08",X"10",X"10",X"00",X"82",X"40",X"00",X"00",X"00",X"80",
		X"02",X"20",X"01",X"05",X"01",X"07",X"05",X"11",X"00",X"25",X"05",X"05",X"05",X"05",X"05",X"00",
		X"05",X"05",X"00",X"07",X"04",X"04",X"00",X"05",X"21",X"20",X"05",X"09",X"0D",X"00",X"05",X"35",
		X"30",X"10",X"80",X"18",X"00",X"24",X"40",X"08",X"10",X"01",X"08",X"20",X"10",X"00",X"43",X"08",
		X"40",X"20",X"00",X"14",X"20",X"10",X"20",X"00",X"00",X"09",X"00",X"00",X"00",X"68",X"28",X"09",
		X"0A",X"B6",X"CA",X"02",X"82",X"0A",X"83",X"00",X"83",X"42",X"82",X"C2",X"88",X"40",X"00",X"20",
		X"C0",X"03",X"86",X"42",X"9B",X"8A",X"8A",X"02",X"82",X"46",X"02",X"82",X"86",X"02",X"8A",X"04",
		X"00",X"50",X"40",X"20",X"00",X"02",X"22",X"00",X"20",X"80",X"28",X"00",X"02",X"42",X"00",X"20",
		X"00",X"02",X"00",X"20",X"00",X"00",X"02",X"12",X"08",X"00",X"00",X"48",X"01",X"02",X"40",X"00",
		X"04",X"00",X"04",X"85",X"05",X"85",X"05",X"11",X"15",X"80",X"0D",X"84",X"05",X"11",X"85",X"00",
		X"05",X"05",X"05",X"05",X"05",X"02",X"00",X"07",X"01",X"80",X"25",X"94",X"05",X"49",X"05",X"8D",
		X"00",X"00",X"40",X"00",X"00",X"60",X"20",X"18",X"60",X"00",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"20",X"00",X"20",X"4C",X"61",X"08",X"50",
		X"C5",X"3B",X"82",X"85",X"90",X"06",X"80",X"82",X"83",X"97",X"82",X"02",X"04",X"02",X"0A",X"C0",
		X"C2",X"96",X"02",X"C7",X"02",X"86",X"82",X"E3",X"8A",X"02",X"43",X"42",X"82",X"47",X"D2",X"22",
		X"0A",X"30",X"60",X"40",X"00",X"40",X"10",X"80",X"00",X"40",X"00",X"08",X"00",X"00",X"48",X"20",
		X"E0",X"28",X"00",X"08",X"00",X"00",X"12",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"28",X"08",
		X"02",X"05",X"07",X"00",X"84",X"45",X"1D",X"02",X"01",X"55",X"05",X"81",X"20",X"23",X"0C",X"B5",
		X"00",X"60",X"05",X"04",X"01",X"01",X"15",X"02",X"05",X"22",X"01",X"07",X"85",X"07",X"75",X"0D",
		X"00",X"08",X"00",X"08",X"04",X"00",X"00",X"00",X"04",X"11",X"40",X"00",X"00",X"00",X"04",X"00",
		X"04",X"08",X"10",X"00",X"05",X"08",X"00",X"09",X"20",X"40",X"2C",X"00",X"40",X"30",X"08",X"10",
		X"00",X"84",X"E6",X"82",X"84",X"82",X"83",X"04",X"81",X"90",X"82",X"00",X"02",X"80",X"82",X"80",
		X"88",X"44",X"82",X"12",X"80",X"8A",X"82",X"62",X"56",X"46",X"05",X"32",X"CA",X"1A",X"04",X"50",
		X"52",X"F0",X"40",X"40",X"00",X"08",X"00",X"00",X"00",X"00",X"50",X"00",X"20",X"00",X"00",X"00",
		X"48",X"00",X"00",X"02",X"00",X"00",X"40",X"22",X"00",X"20",X"00",X"00",X"00",X"0A",X"08",X"00",
		X"27",X"0D",X"01",X"2E",X"05",X"00",X"25",X"05",X"00",X"01",X"01",X"01",X"01",X"25",X"0D",X"2D",
		X"04",X"45",X"89",X"04",X"05",X"95",X"07",X"05",X"27",X"11",X"14",X"11",X"A5",X"65",X"91",X"03",
		X"00",X"48",X"00",X"00",X"28",X"48",X"00",X"01",X"05",X"00",X"08",X"00",X"00",X"00",X"08",X"00",
		X"10",X"10",X"40",X"08",X"10",X"01",X"01",X"10",X"00",X"30",X"00",X"38",X"49",X"60",X"40",X"20",
		X"82",X"83",X"8A",X"82",X"82",X"12",X"92",X"8A",X"80",X"42",X"00",X"C2",X"02",X"84",X"07",X"03",
		X"C2",X"0A",X"86",X"82",X"82",X"06",X"4A",X"02",X"06",X"82",X"42",X"83",X"06",X"02",X"A2",X"08",
		X"02",X"98",X"08",X"00",X"04",X"00",X"00",X"20",X"00",X"00",X"52",X"00",X"20",X"00",X"50",X"40",
		X"00",X"40",X"22",X"00",X"00",X"00",X"A0",X"40",X"40",X"08",X"82",X"00",X"54",X"00",X"00",X"08",
		X"00",X"05",X"45",X"09",X"21",X"04",X"87",X"24",X"05",X"01",X"00",X"01",X"84",X"04",X"09",X"05",
		X"05",X"84",X"04",X"24",X"05",X"04",X"A4",X"14",X"23",X"11",X"00",X"01",X"24",X"07",X"05",X"E5",
		X"24",X"60",X"40",X"00",X"08",X"80",X"34",X"40",X"01",X"84",X"20",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"08",X"00",X"49",X"00",X"04",X"08",X"04",X"04",X"10",X"4C",X"69",X"88",
		X"86",X"84",X"00",X"0A",X"82",X"80",X"86",X"D1",X"08",X"80",X"84",X"84",X"82",X"00",X"88",X"82",
		X"86",X"00",X"02",X"06",X"C1",X"C4",X"02",X"86",X"42",X"02",X"0A",X"C8",X"02",X"02",X"82",X"0A",
		X"22",X"02",X"20",X"10",X"C0",X"12",X"20",X"00",X"08",X"10",X"00",X"08",X"00",X"20",X"00",X"08",
		X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"40",X"80",X"00",X"A0",X"28",X"20",X"02",X"02",X"50",
		X"85",X"17",X"8D",X"14",X"05",X"23",X"05",X"07",X"13",X"01",X"05",X"00",X"04",X"24",X"01",X"25",
		X"00",X"23",X"05",X"05",X"05",X"05",X"04",X"16",X"84",X"84",X"04",X"05",X"05",X"0F",X"AC",X"8C",
		X"08",X"00",X"00",X"40",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"20",
		X"00",X"00",X"00",X"10",X"20",X"00",X"40",X"00",X"20",X"08",X"00",X"00",X"08",X"04",X"01",X"70",
		X"8F",X"04",X"83",X"47",X"86",X"C7",X"42",X"82",X"82",X"83",X"C8",X"42",X"08",X"02",X"82",X"82",
		X"8A",X"87",X"01",X"42",X"82",X"43",X"8A",X"82",X"02",X"00",X"83",X"06",X"00",X"10",X"80",X"42",
		X"40",X"80",X"00",X"30",X"00",X"02",X"00",X"10",X"98",X"00",X"20",X"04",X"00",X"08",X"10",X"00",
		X"40",X"00",X"00",X"E0",X"52",X"00",X"80",X"00",X"02",X"08",X"58",X"C0",X"00",X"00",X"00",X"02",
		X"07",X"05",X"04",X"50",X"57",X"07",X"0C",X"B0",X"05",X"05",X"45",X"17",X"A5",X"04",X"21",X"05",
		X"06",X"05",X"A1",X"09",X"25",X"24",X"22",X"20",X"01",X"02",X"05",X"84",X"80",X"8C",X"03",X"37",
		X"48",X"28",X"00",X"20",X"08",X"00",X"00",X"00",X"00",X"28",X"08",X"00",X"01",X"00",X"00",X"30",
		X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"53",X"20",X"40",X"48",
		X"82",X"CA",X"82",X"E5",X"90",X"02",X"00",X"C6",X"81",X"80",X"92",X"86",X"03",X"02",X"0A",X"26",
		X"80",X"96",X"0B",X"06",X"A3",X"C2",X"01",X"82",X"82",X"06",X"82",X"82",X"84",X"83",X"02",X"C2",
		X"40",X"08",X"82",X"28",X"00",X"28",X"08",X"10",X"00",X"00",X"D8",X"00",X"08",X"0A",X"08",X"40",
		X"00",X"00",X"08",X"04",X"60",X"20",X"00",X"00",X"40",X"80",X"42",X"00",X"00",X"00",X"08",X"04",
		X"20",X"04",X"15",X"10",X"B5",X"11",X"A0",X"11",X"05",X"01",X"85",X"05",X"05",X"6C",X"31",X"21",
		X"04",X"0C",X"04",X"07",X"07",X"84",X"0D",X"04",X"01",X"85",X"00",X"15",X"0D",X"84",X"27",X"25",
		X"00",X"08",X"00",X"00",X"00",X"12",X"00",X"20",X"08",X"09",X"80",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"08",X"00",X"18",X"00",X"00",X"0C",X"08",X"04",X"44",
		X"20",X"4A",X"22",X"06",X"80",X"02",X"1C",X"00",X"50",X"CA",X"02",X"DA",X"10",X"00",X"C2",X"4A",
		X"80",X"C2",X"02",X"8A",X"20",X"02",X"43",X"50",X"08",X"82",X"80",X"00",X"82",X"22",X"C2",X"82",
		X"22",X"A7",X"52",X"06",X"0B",X"00",X"82",X"C2",X"A2",X"02",X"22",X"A2",X"10",X"88",X"C0",X"E0",
		X"8A",X"02",X"82",X"8A",X"82",X"CA",X"0A",X"A0",X"CA",X"22",X"82",X"8E",X"80",X"A2",X"02",X"0A",
		X"01",X"05",X"21",X"00",X"21",X"24",X"08",X"0C",X"04",X"00",X"24",X"11",X"04",X"0D",X"00",X"04",
		X"35",X"10",X"30",X"01",X"05",X"34",X"40",X"00",X"0D",X"01",X"00",X"21",X"05",X"8C",X"2E",X"44",
		X"00",X"01",X"42",X"75",X"40",X"24",X"41",X"15",X"04",X"10",X"05",X"10",X"17",X"47",X"01",X"05",
		X"01",X"05",X"04",X"3D",X"61",X"24",X"04",X"05",X"01",X"00",X"25",X"00",X"51",X"32",X"94",X"85",
		X"02",X"82",X"B4",X"2A",X"82",X"82",X"00",X"08",X"CA",X"02",X"4E",X"92",X"C2",X"B2",X"82",X"82",
		X"E2",X"42",X"CA",X"00",X"62",X"02",X"82",X"C0",X"82",X"80",X"C2",X"02",X"A0",X"02",X"82",X"62",
		X"92",X"63",X"02",X"18",X"08",X"02",X"02",X"38",X"80",X"0E",X"02",X"C2",X"00",X"40",X"D2",X"00",
		X"B2",X"52",X"1A",X"98",X"02",X"00",X"92",X"8A",X"00",X"0A",X"92",X"92",X"A2",X"44",X"80",X"42",
		X"00",X"00",X"10",X"01",X"25",X"05",X"34",X"01",X"0D",X"4C",X"45",X"11",X"10",X"11",X"01",X"21",
		X"35",X"01",X"2C",X"45",X"45",X"64",X"05",X"41",X"25",X"15",X"05",X"28",X"85",X"35",X"25",X"04",
		X"00",X"6D",X"24",X"51",X"40",X"24",X"04",X"05",X"24",X"01",X"21",X"30",X"10",X"25",X"09",X"85",
		X"41",X"71",X"01",X"01",X"00",X"05",X"01",X"21",X"25",X"21",X"00",X"21",X"30",X"0C",X"65",X"5D",
		X"0A",X"C8",X"EA",X"08",X"02",X"24",X"28",X"30",X"C2",X"68",X"80",X"02",X"90",X"02",X"92",X"82",
		X"80",X"42",X"00",X"42",X"42",X"22",X"0A",X"02",X"CA",X"0A",X"62",X"00",X"40",X"00",X"90",X"C2",
		X"92",X"9A",X"06",X"90",X"13",X"92",X"12",X"20",X"18",X"48",X"82",X"20",X"02",X"82",X"90",X"00",
		X"10",X"82",X"02",X"00",X"12",X"00",X"80",X"A0",X"10",X"00",X"A8",X"82",X"10",X"00",X"82",X"08",
		X"28",X"2C",X"25",X"05",X"05",X"A1",X"01",X"01",X"00",X"00",X"1C",X"20",X"14",X"B0",X"21",X"15",
		X"04",X"29",X"31",X"05",X"55",X"11",X"05",X"25",X"34",X"01",X"2D",X"30",X"4D",X"05",X"75",X"45",
		X"41",X"0D",X"01",X"45",X"40",X"05",X"05",X"14",X"05",X"00",X"25",X"25",X"86",X"41",X"00",X"05",
		X"04",X"01",X"01",X"30",X"29",X"21",X"81",X"05",X"11",X"05",X"08",X"05",X"42",X"49",X"51",X"86",
		X"B0",X"B2",X"92",X"92",X"C8",X"12",X"00",X"C2",X"0E",X"48",X"00",X"48",X"0A",X"D0",X"88",X"82",
		X"02",X"00",X"80",X"00",X"8A",X"42",X"00",X"02",X"AA",X"46",X"02",X"42",X"00",X"3A",X"00",X"D0",
		X"42",X"50",X"FF",X"E3",X"80",X"02",X"02",X"92",X"22",X"82",X"02",X"8A",X"00",X"82",X"00",X"C4",
		X"92",X"10",X"00",X"00",X"40",X"C8",X"30",X"2A",X"02",X"92",X"0A",X"00",X"82",X"52",X"00",X"8A",
		X"31",X"0D",X"05",X"60",X"04",X"01",X"00",X"00",X"25",X"11",X"00",X"00",X"01",X"04",X"40",X"01",
		X"40",X"05",X"04",X"01",X"35",X"08",X"10",X"00",X"00",X"09",X"00",X"15",X"27",X"3D",X"49",X"1D",
		X"10",X"01",X"64",X"C5",X"55",X"80",X"00",X"0C",X"05",X"05",X"2C",X"06",X"05",X"09",X"08",X"09",
		X"18",X"14",X"25",X"04",X"24",X"55",X"04",X"01",X"21",X"20",X"05",X"81",X"C5",X"4C",X"5D",X"1D",
		X"A8",X"08",X"C8",X"48",X"84",X"80",X"82",X"82",X"80",X"02",X"63",X"C0",X"02",X"82",X"4A",X"02",
		X"82",X"80",X"8A",X"C2",X"86",X"E0",X"82",X"B2",X"83",X"02",X"E2",X"A2",X"80",X"C2",X"82",X"42",
		X"92",X"02",X"2A",X"62",X"02",X"02",X"C0",X"0A",X"40",X"02",X"C2",X"00",X"06",X"43",X"D2",X"80",
		X"02",X"8A",X"06",X"DA",X"02",X"02",X"22",X"22",X"80",X"02",X"02",X"82",X"8A",X"10",X"58",X"47",
		X"44",X"40",X"00",X"0D",X"00",X"15",X"15",X"00",X"50",X"01",X"01",X"04",X"14",X"00",X"20",X"11",
		X"05",X"01",X"40",X"05",X"21",X"10",X"01",X"15",X"60",X"00",X"15",X"04",X"15",X"ED",X"24",X"15",
		X"16",X"05",X"15",X"02",X"04",X"69",X"10",X"01",X"00",X"05",X"25",X"04",X"15",X"22",X"05",X"41",
		X"01",X"51",X"00",X"14",X"24",X"00",X"11",X"10",X"01",X"15",X"11",X"0C",X"45",X"10",X"3C",X"A6",
		X"F0",X"80",X"88",X"1A",X"82",X"82",X"C0",X"08",X"88",X"80",X"CA",X"CC",X"4A",X"80",X"8A",X"80",
		X"02",X"02",X"02",X"82",X"88",X"8A",X"A2",X"80",X"C0",X"8A",X"02",X"B0",X"83",X"A2",X"00",X"82",
		X"02",X"48",X"02",X"82",X"00",X"92",X"08",X"8A",X"42",X"90",X"80",X"48",X"42",X"C2",X"00",X"C2",
		X"07",X"32",X"22",X"00",X"40",X"80",X"05",X"E8",X"40",X"08",X"A3",X"C2",X"06",X"02",X"4A",X"0A",
		X"21",X"05",X"00",X"05",X"40",X"05",X"04",X"05",X"14",X"15",X"10",X"05",X"01",X"20",X"04",X"01",
		X"01",X"05",X"05",X"01",X"2D",X"00",X"41",X"04",X"20",X"01",X"04",X"01",X"61",X"72",X"65",X"0D",
		X"00",X"80",X"0A",X"21",X"00",X"25",X"10",X"13",X"40",X"34",X"30",X"10",X"4D",X"10",X"20",X"18",
		X"01",X"24",X"3C",X"54",X"01",X"00",X"41",X"05",X"04",X"1C",X"20",X"80",X"17",X"5B",X"5C",X"35",
		X"9A",X"C0",X"AA",X"8A",X"82",X"D2",X"02",X"A0",X"CA",X"40",X"80",X"04",X"5A",X"0A",X"90",X"02",
		X"86",X"A2",X"E2",X"0A",X"84",X"82",X"80",X"C8",X"12",X"08",X"82",X"02",X"02",X"22",X"0A",X"C0",
		X"E0",X"D4",X"D7",X"08",X"92",X"80",X"00",X"00",X"80",X"22",X"20",X"06",X"12",X"00",X"A0",X"32",
		X"12",X"50",X"00",X"82",X"F0",X"82",X"42",X"8A",X"40",X"02",X"1A",X"A0",X"20",X"00",X"C0",X"82",
		X"80",X"45",X"0C",X"21",X"20",X"01",X"21",X"00",X"05",X"00",X"41",X"0C",X"20",X"00",X"44",X"0C",
		X"0C",X"51",X"21",X"21",X"45",X"09",X"08",X"15",X"29",X"04",X"85",X"0C",X"19",X"00",X"30",X"76",
		X"12",X"09",X"09",X"02",X"21",X"2C",X"01",X"01",X"01",X"05",X"21",X"00",X"00",X"25",X"01",X"05",
		X"10",X"05",X"24",X"01",X"00",X"02",X"25",X"10",X"05",X"00",X"A5",X"60",X"55",X"75",X"75",X"4D",
		X"88",X"92",X"80",X"08",X"20",X"A8",X"00",X"1A",X"DA",X"02",X"EA",X"02",X"02",X"00",X"42",X"00",
		X"02",X"50",X"42",X"40",X"C2",X"80",X"C8",X"00",X"02",X"4A",X"C6",X"02",X"90",X"00",X"32",X"10",
		X"9A",X"80",X"D3",X"A4",X"80",X"C0",X"C2",X"C8",X"00",X"02",X"8A",X"23",X"23",X"D8",X"08",X"D0",
		X"82",X"12",X"82",X"20",X"92",X"F0",X"02",X"02",X"E8",X"E2",X"90",X"A2",X"02",X"E0",X"22",X"40",
		X"60",X"05",X"0D",X"00",X"04",X"1D",X"01",X"05",X"01",X"09",X"24",X"60",X"75",X"11",X"27",X"81",
		X"1C",X"15",X"25",X"05",X"00",X"25",X"25",X"45",X"01",X"11",X"00",X"E9",X"09",X"65",X"25",X"2D",
		X"50",X"07",X"19",X"3B",X"15",X"00",X"05",X"01",X"05",X"08",X"1D",X"21",X"21",X"14",X"0D",X"0D",
		X"04",X"60",X"04",X"04",X"25",X"11",X"23",X"25",X"19",X"C0",X"00",X"40",X"9F",X"13",X"65",X"59");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
