library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"A1",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"70",X"B0",X"80",X"C1",X"40",X"41",X"40",X"00",
		X"80",X"90",X"10",X"38",X"20",X"28",X"20",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"41",X"81",X"F0",
		X"00",X"00",X"80",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"A0",X"B0",X"00",X"E0",X"20",X"20",X"20",X"00",
		X"00",X"90",X"10",X"0C",X"20",X"2C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"80",X"03",X"43",X"30",
		X"00",X"00",X"00",X"00",X"00",X"80",X"58",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"60",X"20",X"10",X"10",X"00",X"00",
		X"80",X"00",X"00",X"1C",X"00",X"06",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"00",X"80",X"03",X"21",X"50",
		X"00",X"00",X"00",X"00",X"00",X"10",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"90",X"50",X"20",X"10",X"00",X"00",X"00",
		X"80",X"90",X"02",X"04",X"03",X"80",X"40",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"40",X"00",X"12",X"43",X"70",
		X"00",X"00",X"00",X"00",X"20",X"10",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"B0",X"90",X"70",X"60",X"00",X"00",X"00",
		X"C0",X"82",X"06",X"00",X"C1",X"60",X"00",X"00",X"00",X"80",X"40",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"20",X"30",X"00",X"00",X"00",X"10",X"00",X"00",X"96",X"61",
		X"00",X"00",X"00",X"80",X"60",X"10",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"B0",X"C0",X"70",X"20",X"00",X"00",X"00",
		X"C1",X"83",X"80",X"40",X"B0",X"00",X"00",X"00",X"40",X"00",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"60",X"00",X"00",X"00",X"10",X"00",X"80",X"34",X"43",
		X"00",X"00",X"00",X"C0",X"E0",X"30",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"70",X"D0",X"60",X"10",X"00",X"00",X"00",
		X"C1",X"C1",X"40",X"B0",X"80",X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"34",X"43",
		X"00",X"00",X"00",X"E0",X"20",X"00",X"00",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"0C",
		X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"70",X"50",X"60",X"10",X"00",X"00",X"00",
		X"81",X"C1",X"20",X"90",X"80",X"00",X"00",X"00",X"04",X"04",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"04",
		X"00",X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"61",X"B0",X"20",X"70",X"00",X"00",X"00",X"00",
		X"C1",X"C0",X"10",X"C0",X"80",X"00",X"00",X"00",X"04",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"10",X"60",X"00",X"20",X"43",
		X"00",X"00",X"00",X"80",X"00",X"20",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"00",X"04",X"04",
		X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"61",X"70",X"30",X"70",X"00",X"00",X"00",X"00",
		X"80",X"80",X"10",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"00",X"03",
		X"00",X"00",X"00",X"00",X"30",X"00",X"01",X"01",X"00",X"00",X"00",X"C0",X"00",X"0C",X"04",X"00",
		X"20",X"00",X"00",X"10",X"30",X"00",X"00",X"00",X"07",X"34",X"30",X"80",X"D0",X"00",X"00",X"00",
		X"C0",X"90",X"20",X"60",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"A0",X"80",X"01",
		X"00",X"00",X"00",X"00",X"40",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"08",X"04",X"00",X"20",
		X"10",X"20",X"00",X"00",X"10",X"10",X"00",X"00",X"25",X"70",X"70",X"60",X"B0",X"50",X"00",X"00",
		X"00",X"D0",X"70",X"F0",X"C0",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"30",X"40",X"80",X"00",X"30",
		X"00",X"00",X"40",X"81",X"00",X"86",X"02",X"20",X"00",X"00",X"00",X"00",X"08",X"00",X"40",X"80",
		X"00",X"30",X"10",X"20",X"00",X"00",X"00",X"00",X"C3",X"E1",X"30",X"20",X"30",X"C0",X"00",X"00",
		X"80",X"80",X"80",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"80",X"80",X"B0",
		X"00",X"00",X"00",X"03",X"05",X"02",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"21",X"61",X"70",X"10",X"00",X"00",X"30",X"40",
		X"48",X"90",X"B0",X"60",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"40",X"C0",X"80",
		X"00",X"80",X"06",X"02",X"06",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"83",X"61",X"70",X"90",X"80",X"80",X"30",X"00",
		X"08",X"10",X"30",X"60",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"80",X"B0",
		X"00",X"10",X"1C",X"10",X"1C",X"00",X"10",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"A1",X"30",X"10",X"40",X"40",X"00",X"00",
		X"58",X"58",X"D0",X"A0",X"A0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"00",X"41",X"00",X"80",X"80",
		X"00",X"00",X"08",X"00",X"28",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"A1",X"B0",X"20",X"40",X"20",X"20",X"00",
		X"58",X"58",X"D0",X"C0",X"00",X"40",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"77",X"23",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"44",X"FF",X"77",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"DD",X"BB",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"88",X"08",X"0C",X"08",
		X"03",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"08",X"00",X"88",X"EE",X"FF",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"44",X"EE",X"55",X"33",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"88",X"08",X"0C",
		X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"EE",X"FF",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"00",
		X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",
		X"00",X"00",X"88",X"88",X"11",X"22",X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"44",X"88",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"66",X"88",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"88",X"22",X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"88",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"50",X"00",
		X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"88",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"D0",X"29",
		X"00",X"42",X"43",X"43",X"52",X"24",X"80",X"48",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",
		X"16",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"38",X"D0",X"E0",X"F0",X"F0",X"70",X"00",X"00",
		X"48",X"A0",X"16",X"C3",X"C3",X"C3",X"43",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"70",X"30",X"00",X"00",X"00",X"00",X"08",X"0C",X"1C",X"A1",
		X"00",X"00",X"00",X"00",X"10",X"21",X"92",X"48",X"00",X"00",X"00",X"80",X"0C",X"0C",X"E0",X"00",
		X"30",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"A1",X"D0",X"E0",X"E1",X"E1",X"21",X"21",X"00",
		X"48",X"A0",X"70",X"78",X"2C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"10",X"30",X"30",X"00",X"02",X"0E",X"0E",X"86",X"C2",X"D0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",
		X"30",X"70",X"30",X"10",X"01",X"00",X"00",X"00",X"B0",X"D0",X"86",X"5A",X"D2",X"1E",X"02",X"00",
		X"50",X"80",X"40",X"E0",X"E0",X"C0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"21",X"21",X"21",X"01",X"80",X"D0",X"B0",
		X"00",X"0C",X"0C",X"0C",X"08",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"03",X"03",X"10",X"00",X"00",X"00",X"B0",X"94",X"A4",X"B4",X"78",X"70",X"00",X"00",
		X"C0",X"83",X"61",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"0E",X"0C",X"0C",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"10",
		X"00",X"00",X"00",X"00",X"D0",X"C0",X"00",X"80",X"00",X"00",X"00",X"01",X"81",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"D0",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"81",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"08",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"30",X"01",X"00",X"00",
		X"00",X"00",X"C0",X"D0",X"C0",X"08",X"00",X"00",X"00",X"00",X"01",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"38",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"F0",X"30",X"40",
		X"00",X"00",X"08",X"08",X"00",X"D0",X"C0",X"20",X"00",X"00",X"00",X"00",X"01",X"81",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"70",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"6F",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",X"0C",X"8E",X"CF",X"FE",X"FC",X"F9",X"FF",
		X"00",X"02",X"06",X"0C",X"08",X"00",X"08",X"8D",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0C",
		X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"BB",X"11",X"00",X"11",X"01",X"03",X"06",X"00",
		X"FE",X"FC",X"F9",X"FF",X"FF",X"77",X"33",X"00",X"08",X"0C",X"8E",X"CE",X"CF",X"EF",X"EF",X"CF",
		X"0F",X"6F",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",X"0C",X"8E",X"CF",X"EF",X"FD",X"BD",X"F3",
		X"01",X"03",X"06",X"84",X"08",X"00",X"08",X"8D",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"11",X"00",X"11",X"01",X"03",X"06",X"0C",
		X"EF",X"FC",X"77",X"F7",X"FF",X"77",X"33",X"00",X"80",X"0C",X"8E",X"CE",X"CF",X"EF",X"EF",X"CF",
		X"0F",X"6F",X"FF",X"FF",X"77",X"77",X"33",X"01",X"00",X"0C",X"8E",X"DE",X"EF",X"FF",X"F3",X"7B",
		X"00",X"04",X"84",X"08",X"08",X"00",X"08",X"8D",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"84",
		X"21",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"11",X"00",X"11",X"01",X"21",X"02",X"00",
		X"FE",X"FF",X"FF",X"7B",X"7B",X"77",X"33",X"00",X"08",X"0C",X"8E",X"CE",X"CF",X"EF",X"EF",X"CF",
		X"0F",X"6F",X"FF",X"FF",X"77",X"77",X"33",X"10",X"00",X"0C",X"8E",X"CF",X"EF",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"00",X"08",X"8D",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"84",
		X"03",X"06",X"0C",X"08",X"00",X"00",X"00",X"00",X"BB",X"11",X"00",X"11",X"00",X"00",X"00",X"00",
		X"EF",X"FF",X"BD",X"F3",X"FF",X"77",X"33",X"00",X"08",X"0C",X"8E",X"CE",X"CF",X"EF",X"EF",X"CF",
		X"10",X"10",X"10",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"70",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"10",X"10",X"10",X"70",X"70",X"30",X"00",X"00",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"00",X"00",X"F0",X"F0",X"F0",X"30",X"70",X"70",X"70",X"70",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"70",X"70",X"30",X"00",X"00",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"00",X"00",X"E0",X"E0",X"E0",X"70",X"70",X"70",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"10",X"00",X"00",X"70",X"70",X"70",
		X"80",X"80",X"80",X"00",X"00",X"C0",X"C0",X"C0",X"70",X"70",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"30",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"30",X"00",X"00",X"10",X"10",X"10",
		X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"70",X"70",X"70",X"00",X"00",X"00",X"00",X"70",
		X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"10",X"00",X"00",X"40",X"40",X"40",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"70",
		X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"70",X"70",X"30",X"00",X"00",X"80",X"80",X"80",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"10",
		X"00",X"10",X"30",X"30",X"20",X"80",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"70",X"30",X"00",X"00",X"00",X"10",X"70",X"00",X"F0",X"F0",X"F0",X"70",X"00",
		X"90",X"00",X"00",X"A0",X"F0",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"B0",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"08",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"70",X"30",X"00",X"00",X"00",X"F0",X"60",X"00",X"E0",X"F0",X"F0",X"70",X"10",
		X"F0",X"20",X"00",X"20",X"B0",X"B0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"10",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"70",X"30",X"00",X"00",X"00",X"D0",X"40",X"00",X"C0",X"D0",X"D0",X"B0",X"00",
		X"80",X"E0",X"00",X"E0",X"F0",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"E0",X"20",X"00",X"10",
		X"80",X"80",X"80",X"80",X"00",X"40",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"70",X"10",X"00",X"00",X"00",X"10",X"00",X"80",X"F0",X"F0",X"F0",X"70",X"00",
		X"80",X"00",X"10",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"C0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"21",X"F0",X"E1",X"30",X"30",X"EE",X"00",X"00",
		X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"21",X"F0",X"E1",X"30",X"30",X"00",X"00",X"00",
		X"00",X"30",X"30",X"00",X"00",X"EE",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"00",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"10",X"B0",X"70",X"F0",X"F0",X"E0",X"80",X"C0",X"E0",X"F0",X"F0",X"B0",X"30",X"B0",
		X"10",X"00",X"10",X"30",X"10",X"00",X"00",X"00",X"70",X"F0",X"F0",X"E0",X"D0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"B0",X"30",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"00",X"10",X"00",X"01",X"01",X"43",
		X"F0",X"F0",X"10",X"B0",X"70",X"78",X"78",X"0E",X"80",X"C0",X"E0",X"F0",X"F0",X"B0",X"30",X"B0",
		X"10",X"00",X"10",X"30",X"10",X"00",X"00",X"00",X"70",X"F0",X"F0",X"E0",X"D0",X"80",X"00",X"00",
		X"68",X"08",X"80",X"00",X"80",X"00",X"00",X"00",X"B0",X"30",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"00",X"10",X"20",X"21",X"87",X"43",
		X"F0",X"F0",X"10",X"B0",X"34",X"3C",X"0F",X"0E",X"80",X"C0",X"E0",X"F0",X"F0",X"B0",X"30",X"B0",
		X"10",X"00",X"10",X"30",X"10",X"00",X"00",X"00",X"52",X"E1",X"F0",X"E0",X"D0",X"80",X"00",X"00",
		X"0E",X"3C",X"84",X"40",X"80",X"00",X"00",X"00",X"B0",X"30",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"30",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"E0",X"10",X"30",X"30",X"10",X"60",X"60",X"00",X"00",X"00",X"80",X"C0",X"E0",X"D0",X"10",X"10",
		X"20",X"20",X"20",X"70",X"70",X"30",X"10",X"00",X"70",X"30",X"D0",X"C0",X"80",X"F0",X"80",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"30",X"00",X"00",X"00",X"10",X"10",X"10",X"30",
		X"E0",X"10",X"30",X"30",X"10",X"60",X"60",X"80",X"00",X"00",X"80",X"C0",X"E0",X"D0",X"10",X"10",
		X"30",X"20",X"20",X"70",X"70",X"30",X"10",X"00",X"F0",X"30",X"D0",X"D0",X"90",X"F0",X"80",X"00",
		X"F0",X"80",X"00",X"00",X"00",X"C0",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",
		X"E0",X"10",X"30",X"30",X"D0",X"E0",X"F0",X"F0",X"00",X"00",X"80",X"C0",X"E0",X"D0",X"10",X"10",
		X"30",X"30",X"30",X"70",X"70",X"30",X"10",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"00",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"74",X"44",X"44",X"00",X"00",X"00",X"00",X"D0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"60",
		X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"60",
		X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"70",X"69",X"69",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"4B",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"86",
		X"30",X"12",X"21",X"10",X"00",X"00",X"00",X"00",X"78",X"78",X"F0",X"F0",X"F0",X"70",X"10",X"00",
		X"E1",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"86",X"E0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5A",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",
		X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"84",X"C0",X"E0",X"70",X"00",X"00",
		X"5A",X"F0",X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"08",X"28",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"10",X"10",X"00",X"00",
		X"28",X"28",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"C0",X"60",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"70",X"80",X"70",X"00",X"00",
		X"E0",X"E0",X"A0",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"40",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"D0",X"30",X"00",
		X"20",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"24",X"60",X"00",X"00",X"10",X"10",X"10",
		X"29",X"29",X"B0",X"08",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"01",X"10",X"10",X"10",X"00",X"00",
		X"C0",X"84",X"84",X"C8",X"C8",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"20",X"00",X"00",X"00",
		X"00",X"00",X"80",X"82",X"14",X"50",X"48",X"80",X"00",X"00",X"00",X"00",X"0C",X"08",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"34",X"25",X"46",X"C4",X"88",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"02",X"60",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"08",X"80",X"C2",X"C0",X"80",
		X"00",X"00",X"00",X"10",X"11",X"20",X"00",X"00",X"30",X"3C",X"4A",X"8E",X"80",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"01",X"52",X"30",X"00",X"61",X"84",X"00",X"00",X"08",X"80",X"80",X"08",X"00",X"C0",
		X"01",X"52",X"67",X"C9",X"00",X"00",X"00",X"00",X"70",X"68",X"08",X"00",X"00",X"00",X"00",X"00",
		X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"61",X"70",X"00",
		X"73",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"96",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"70",X"61",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"77",X"44",X"00",X"00",X"00",X"33",X"11",X"11",X"99",X"FF",X"33",X"00",
		X"44",X"44",X"44",X"77",X"77",X"44",X"00",X"00",X"00",X"99",X"99",X"99",X"FF",X"FF",X"33",X"00",
		X"33",X"66",X"44",X"66",X"77",X"44",X"00",X"00",X"88",X"CC",X"44",X"44",X"CC",X"FF",X"33",X"00",
		X"33",X"77",X"44",X"44",X"77",X"44",X"00",X"00",X"00",X"BB",X"FF",X"CC",X"88",X"FF",X"33",X"00",
		X"66",X"11",X"00",X"33",X"77",X"66",X"00",X"00",X"00",X"00",X"CC",X"FF",X"33",X"00",X"00",X"00",
		X"33",X"33",X"66",X"44",X"77",X"44",X"00",X"00",X"CC",X"EE",X"33",X"11",X"99",X"FF",X"33",X"00",
		X"00",X"77",X"77",X"66",X"55",X"00",X"00",X"00",X"11",X"FF",X"FF",X"44",X"44",X"CC",X"77",X"00",
		X"00",X"77",X"77",X"66",X"55",X"00",X"00",X"00",X"11",X"FF",X"FF",X"44",X"44",X"CC",X"77",X"00",
		X"33",X"77",X"44",X"44",X"77",X"44",X"00",X"00",X"00",X"BB",X"FF",X"CC",X"88",X"FF",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"77",X"77",X"44",X"00",X"00",X"00",X"99",X"99",X"99",X"FF",X"FF",X"33",X"00",
		X"66",X"11",X"00",X"33",X"77",X"66",X"00",X"00",X"00",X"00",X"CC",X"FF",X"33",X"00",X"00",X"00",
		X"66",X"11",X"00",X"11",X"77",X"11",X"00",X"00",X"00",X"CC",X"77",X"FF",X"CC",X"88",X"77",X"00",
		X"66",X"11",X"11",X"77",X"00",X"11",X"77",X"00",X"00",X"CC",X"FF",X"88",X"44",X"FF",X"88",X"00",
		X"33",X"77",X"44",X"44",X"66",X"33",X"00",X"00",X"88",X"EE",X"33",X"11",X"11",X"FF",X"EE",X"00",
		X"44",X"44",X"66",X"77",X"55",X"44",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"77",X"77",X"44",X"00",X"00",X"00",X"99",X"99",X"99",X"FF",X"FF",X"33",X"00",
		X"33",X"77",X"44",X"44",X"66",X"33",X"00",X"00",X"88",X"EE",X"33",X"11",X"11",X"FF",X"EE",X"00",
		X"F7",X"FF",X"F0",X"EC",X"EC",X"FD",X"F5",X"70",X"FE",X"EC",X"C0",X"00",X"00",X"EC",X"FE",X"F0",
		X"FF",X"F7",X"F0",X"00",X"70",X"F7",X"FF",X"F0",X"FE",X"FF",X"F0",X"73",X"F3",X"FB",X"FA",X"E0",
		X"70",X"F7",X"FF",X"F0",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"F0",X"00",X"00",X"00",X"00",
		X"70",X"F7",X"FF",X"F0",X"00",X"00",X"00",X"00",X"E0",X"FE",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"F7",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"70",X"FE",X"EC",X"C0",X"00",X"C0",X"EC",X"FE",X"F0",
		X"FF",X"F7",X"70",X"00",X"00",X"F7",X"FF",X"F0",X"FE",X"FF",X"F0",X"73",X"73",X"FB",X"FA",X"A0",
		X"F7",X"FF",X"F0",X"EC",X"EC",X"EC",X"E4",X"60",X"FE",X"FC",X"F1",X"31",X"31",X"10",X"10",X"10",
		X"00",X"80",X"C8",X"C8",X"F8",X"F3",X"FF",X"F0",X"10",X"31",X"73",X"73",X"F3",X"FB",X"FA",X"E0",
		X"F7",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"50",X"FE",X"EC",X"C0",X"00",X"C0",X"EC",X"FE",X"E0",
		X"FF",X"F7",X"70",X"00",X"70",X"F7",X"FF",X"F0",X"EE",X"FF",X"F0",X"73",X"F3",X"FB",X"FA",X"A0",
		X"70",X"F7",X"FF",X"F0",X"EC",X"EC",X"EC",X"E4",X"E0",X"FE",X"EC",X"F1",X"31",X"31",X"10",X"00",
		X"F0",X"FF",X"F3",X"F8",X"C8",X"C8",X"80",X"00",X"E0",X"FE",X"FF",X"F0",X"73",X"73",X"73",X"72",
		X"77",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"50",X"FE",X"EC",X"C0",X"00",X"C0",X"EC",X"FE",X"E0",
		X"FF",X"F7",X"70",X"00",X"70",X"F7",X"FF",X"F0",X"FE",X"FF",X"F0",X"73",X"F3",X"FB",X"FA",X"A0",
		X"00",X"80",X"C8",X"EC",X"EC",X"FC",X"FD",X"F5",X"00",X"10",X"10",X"31",X"31",X"F1",X"FC",X"FE",
		X"00",X"FF",X"F3",X"F8",X"C8",X"C8",X"C8",X"80",X"00",X"EE",X"FF",X"F0",X"73",X"73",X"73",X"72",
		X"F7",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"70",X"FE",X"EC",X"C0",X"00",X"C0",X"EC",X"FE",X"E0",
		X"FF",X"F7",X"70",X"00",X"70",X"F7",X"FF",X"F0",X"FE",X"FF",X"F0",X"73",X"F3",X"FB",X"FA",X"E0",
		X"F7",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"50",X"EC",X"FE",X"F1",X"31",X"F1",X"FE",X"EC",X"E0",
		X"73",X"F7",X"F8",X"C8",X"F8",X"F7",X"73",X"70",X"FE",X"FF",X"F0",X"73",X"F3",X"FB",X"FA",X"A0",
		X"F7",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"70",X"FE",X"EC",X"C0",X"00",X"C0",X"EC",X"FE",X"E0",
		X"FF",X"F7",X"70",X"00",X"70",X"F7",X"FF",X"F0",X"FE",X"FF",X"F0",X"33",X"B3",X"FB",X"FA",X"E0",
		X"F7",X"FF",X"F0",X"EC",X"FC",X"FD",X"F5",X"50",X"FE",X"EC",X"C0",X"00",X"C0",X"EC",X"FE",X"E0",
		X"FF",X"F7",X"70",X"00",X"70",X"F7",X"FF",X"F0",X"FE",X"FF",X"F0",X"73",X"F3",X"FB",X"FA",X"A0",
		X"00",X"00",X"00",X"10",X"21",X"12",X"12",X"71",X"00",X"10",X"61",X"97",X"7B",X"F7",X"F3",X"FF",
		X"00",X"80",X"48",X"A4",X"DA",X"C3",X"C7",X"FE",X"00",X"00",X"00",X"00",X"80",X"48",X"A4",X"2C",
		X"37",X"35",X"12",X"01",X"00",X"00",X"00",X"00",X"FF",X"F3",X"F7",X"FF",X"F7",X"78",X"07",X"00",
		X"FE",X"EF",X"E7",X"C3",X"C3",X"2D",X"48",X"00",X"2C",X"48",X"48",X"48",X"48",X"80",X"00",X"00",
		X"00",X"10",X"21",X"21",X"52",X"3D",X"7B",X"7B",X"F0",X"2D",X"1E",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"3C",X"C3",X"ED",X"FE",X"FF",X"FF",X"FF",X"00",X"80",X"48",X"2C",X"2C",X"96",X"D2",X"96",
		X"7B",X"F7",X"73",X"73",X"35",X"16",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"78",X"07",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"E3",X"0F",X"07",X"DA",X"D2",X"96",X"A4",X"48",X"48",X"48",X"80",
		X"00",X"10",X"03",X"01",X"31",X"7B",X"7B",X"F7",X"94",X"2D",X"0F",X"C3",X"F8",X"FC",X"FE",X"FF",
		X"48",X"2D",X"0F",X"C3",X"E1",X"F4",X"F6",X"F8",X"00",X"80",X"48",X"2C",X"0E",X"3C",X"87",X"2C",
		X"F7",X"F7",X"73",X"71",X"34",X"16",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F0",X"07",
		X"FC",X"FE",X"FE",X"FE",X"FC",X"E1",X"0F",X"16",X"96",X"87",X"1E",X"2C",X"0C",X"0C",X"48",X"00",
		X"20",X"07",X"03",X"03",X"03",X"03",X"16",X"1F",X"10",X"87",X"0F",X"3C",X"7B",X"F1",X"F8",X"FC",
		X"C0",X"1E",X"2D",X"C3",X"F8",X"FC",X"F4",X"E1",X"00",X"80",X"68",X"48",X"0C",X"2C",X"2C",X"0F",
		X"1E",X"12",X"01",X"03",X"03",X"05",X"00",X"00",X"FC",X"F1",X"F5",X"7E",X"3E",X"0F",X"03",X"01",
		X"E9",X"FC",X"FE",X"E9",X"87",X"0F",X"08",X"00",X"1E",X"2C",X"2C",X"0C",X"0C",X"2C",X"E0",X"20",
		X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"07",X"31",X"31",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"01",X"04",X"00",X"00",X"00",X"00",X"00",
		X"8E",X"42",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"64",X"11",X"00",X"C8",X"C0",X"10",X"00",X"40",X"00",
		X"00",X"00",X"31",X"10",X"88",X"A0",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"C4",X"40",
		X"00",X"00",X"22",X"00",X"11",X"00",X"00",X"00",X"64",X"22",X"00",X"00",X"C0",X"88",X"11",X"00",
		X"40",X"10",X"80",X"10",X"31",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"32",X"80",X"00",X"00",X"40",X"00",X"20",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"44",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"44",X"C0",X"00",
		X"30",X"22",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"60",X"44",X"00",X"00",X"10",X"00",X"00",
		X"00",X"40",X"62",X"00",X"00",X"90",X"88",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"32",X"00",X"00",X"11",X"00",X"C8",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"62",X"20",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"C4",X"00",
		X"00",X"00",X"10",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"22",X"00",X"20",X"22",X"00",X"00",
		X"00",X"10",X"00",X"80",X"44",X"00",X"44",X"00",X"00",X"80",X"99",X"00",X"80",X"00",X"00",X"00",
		X"00",X"40",X"02",X"10",X"01",X"00",X"40",X"60",X"00",X"40",X"60",X"00",X"8D",X"4B",X"78",X"72",
		X"00",X"00",X"90",X"C0",X"30",X"08",X"0E",X"84",X"00",X"00",X"80",X"00",X"00",X"00",X"A0",X"80",
		X"00",X"20",X"30",X"00",X"00",X"10",X"10",X"00",X"B3",X"73",X"71",X"12",X"40",X"10",X"80",X"00",
		X"C2",X"CB",X"CA",X"A5",X"93",X"02",X"00",X"30",X"00",X"40",X"60",X"00",X"08",X"84",X"02",X"00",
		X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"21",X"61",X"1E",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"1E",X"E1",X"E1",X"61",X"00",X"80",X"00",X"00",
		X"87",X"68",X"48",X"08",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"02",X"32",X"26",X"26",X"3E",X"AE",X"AE",
		X"00",X"04",X"C4",X"46",X"46",X"C7",X"57",X"57",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"11",X"33",X"23",X"23",X"33",X"11",X"00",X"00",X"BE",X"B7",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",
		X"D7",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"88",X"CC",X"4C",X"4C",X"CC",X"88",X"00",X"00",
		X"00",X"11",X"11",X"01",X"01",X"11",X"11",X"01",X"66",X"F3",X"99",X"99",X"7C",X"4C",X"AE",X"BE",
		X"00",X"00",X"88",X"A6",X"9F",X"FB",X"56",X"F5",X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"C4",
		X"01",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"FF",X"FF",X"BF",X"BF",X"BF",X"FF",X"57",X"11",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"EF",X"88",X"CA",X"EE",X"E6",X"C4",X"88",X"08",X"00",X"00",
		X"00",X"11",X"00",X"44",X"26",X"13",X"13",X"11",X"00",X"08",X"8E",X"75",X"32",X"51",X"88",X"DC",
		X"00",X"00",X"00",X"0C",X"EF",X"F0",X"9F",X"C7",X"00",X"00",X"00",X"00",X"08",X"8C",X"C6",X"EA",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"BE",X"9F",X"AF",X"BF",X"DF",X"67",X"33",X"00",
		X"EF",X"FF",X"FF",X"7F",X"BF",X"DF",X"6F",X"00",X"6C",X"6E",X"AE",X"CE",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"57",X"73",X"40",X"4C",X"37",X"00",X"00",X"00",X"2F",X"F3",X"FC",X"B3",X"90",
		X"00",X"00",X"00",X"4F",X"FC",X"DB",X"E3",X"CF",X"00",X"00",X"00",X"08",X"8C",X"C6",X"CE",X"6E",
		X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"FF",X"DF",X"DF",X"67",X"33",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"9F",X"CC",X"00",X"0F",X"EF",X"CE",X"8E",X"8C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"77",X"20",X"00",X"00",X"00",X"01",X"37",X"78",X"FF",X"40",
		X"00",X"00",X"17",X"FC",X"FB",X"87",X"FF",X"F7",X"00",X"00",X"88",X"C0",X"2E",X"6F",X"EF",X"FF",
		X"20",X"77",X"11",X"00",X"00",X"00",X"00",X"00",X"40",X"FF",X"FF",X"77",X"11",X"00",X"00",X"00",
		X"F7",X"FF",X"4F",X"BF",X"CF",X"77",X"00",X"00",X"FF",X"FF",X"3F",X"CC",X"0C",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"12",X"00",X"23",X"17",X"7E",X"5F",X"FC",X"F3",X"DC",
		X"00",X"CE",X"FB",X"F6",X"F9",X"F7",X"FF",X"FF",X"00",X"00",X"00",X"4C",X"8E",X"CE",X"EE",X"7F",
		X"37",X"CC",X"40",X"73",X"47",X"00",X"00",X"00",X"90",X"B3",X"CF",X"3F",X"FF",X"00",X"00",X"00",
		X"FC",X"7F",X"BF",X"CF",X"FF",X"00",X"00",X"00",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"03",X"16",X"3D",X"AF",X"BE",X"9F",X"AF",
		X"00",X"86",X"2D",X"7B",X"F7",X"FF",X"FF",X"EF",X"00",X"00",X"00",X"08",X"8C",X"EE",X"EE",X"CE",
		X"11",X"23",X"13",X"26",X"54",X"00",X"11",X"00",X"5C",X"88",X"51",X"23",X"57",X"EE",X"88",X"00",
		X"5F",X"FF",X"0F",X"FF",X"CC",X"00",X"00",X"00",X"AE",X"6E",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"01",X"11",X"01",X"01",X"11",X"17",X"4F",X"2F",X"BE",X"BE",X"FD",X"FD",
		X"08",X"4B",X"E7",X"F7",X"FF",X"FF",X"EF",X"EF",X"00",X"00",X"08",X"CC",X"AE",X"6E",X"CE",X"AE",
		X"11",X"11",X"11",X"11",X"01",X"11",X"11",X"00",X"FA",X"AE",X"4C",X"F4",X"99",X"99",X"F3",X"33",
		X"F7",X"77",X"8F",X"BF",X"6E",X"CC",X"88",X"00",X"6E",X"4E",X"8C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"23",X"23",X"23",X"33",X"11",X"17",X"AF",X"BF",X"BF",X"BF",X"BF",X"B7",X"BE",
		X"8E",X"5F",X"DF",X"DF",X"DF",X"DF",X"DE",X"D7",X"00",X"00",X"08",X"4C",X"4C",X"4C",X"CC",X"88",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AE",X"AE",X"BE",X"66",X"66",X"32",X"22",X"00",
		X"57",X"57",X"D7",X"66",X"66",X"C4",X"44",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"13",X"77",X"37",X"00",X"00",X"02",X"37",X"EF",X"BF",X"FF",X"FF",
		X"00",X"00",X"04",X"CE",X"7F",X"DF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"8C",X"EE",X"CE",
		X"77",X"77",X"77",X"77",X"33",X"11",X"00",X"00",X"33",X"11",X"11",X"11",X"11",X"11",X"00",X"00",
		X"CC",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"13",X"77",X"00",X"00",X"99",X"FF",X"9E",X"DE",X"FF",X"7F",
		X"00",X"00",X"0F",X"FF",X"EF",X"7F",X"A6",X"C8",X"00",X"00",X"00",X"4C",X"8C",X"CE",X"CE",X"FF",
		X"77",X"77",X"77",X"33",X"13",X"01",X"00",X"00",X"5F",X"99",X"88",X"88",X"CC",X"CC",X"44",X"00",
		X"8C",X"CC",X"CC",X"EE",X"66",X"00",X"00",X"00",X"77",X"67",X"26",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"77",X"00",X"00",X"9F",X"CF",X"ED",X"FE",X"FF",X"FF",
		X"00",X"06",X"6F",X"FB",X"7D",X"19",X"80",X"88",X"00",X"00",X"00",X"08",X"CC",X"EE",X"EE",X"66",
		X"67",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"DF",X"08",X"88",X"CC",X"EE",X"FF",X"77",X"00",
		X"CC",X"EE",X"77",X"22",X"00",X"00",X"88",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"13",X"11",X"11",X"33",X"00",X"11",X"17",X"BF",X"7F",X"79",X"FE",X"FF",
		X"00",X"0E",X"EF",X"FF",X"3F",X"08",X"80",X"88",X"00",X"00",X"88",X"0C",X"CC",X"EE",X"00",X"00",
		X"33",X"33",X"33",X"11",X"11",X"01",X"00",X"00",X"FF",X"FF",X"EE",X"CC",X"FF",X"FF",X"77",X"11",
		X"EF",X"FF",X"33",X"00",X"08",X"AF",X"EF",X"CC",X"00",X"88",X"88",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"03",X"37",X"FC",X"3F",X"8F",X"8F",X"FF",
		X"00",X"0F",X"FF",X"FF",X"00",X"00",X"08",X"FF",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"CC",
		X"11",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"CF",X"FF",X"77",X"33",X"00",
		X"FF",X"88",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"CC",X"00",X"00",X"00",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"01",X"01",X"11",X"33",X"33",X"23",X"01",X"17",X"7F",X"FF",X"CE",X"AE",X"CF",X"3F",
		X"0C",X"CF",X"EE",X"00",X"00",X"13",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"00",
		X"13",X"11",X"11",X"33",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"EF",X"77",X"37",X"11",X"00",
		X"88",X"88",X"08",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"EE",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"37",X"76",X"77",X"00",X"37",X"7F",X"EE",X"CC",X"80",X"08",X"7D",
		X"00",X"88",X"00",X"00",X"03",X"77",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"67",X"13",X"33",X"33",X"11",X"00",X"00",X"00",X"FB",X"F7",X"FF",X"FF",X"FF",X"FF",X"11",X"00",
		X"88",X"88",X"99",X"BF",X"7F",X"FF",X"EE",X"00",X"66",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"01",X"13",X"13",X"37",X"77",X"67",X"00",X"CC",X"4C",X"8C",X"88",X"88",X"99",X"1F",
		X"00",X"00",X"00",X"46",X"6E",X"AE",X"CE",X"CC",X"00",X"00",X"00",X"00",X"02",X"46",X"67",X"77",
		X"77",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"00",X"00",
		X"8C",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"EE",X"EE",X"CC",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"01",X"13",X"37",X"37",X"77",X"77",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"13",
		X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"8C",X"00",X"00",X"08",X"8C",X"CE",X"CE",X"EE",X"EE",
		X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"BF",X"FF",X"FF",X"FF",X"77",X"22",X"00",X"00",
		X"DF",X"FF",X"FF",X"FF",X"EE",X"44",X"00",X"00",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"00",X"00",X"00",X"44",X"CC",X"CC",X"7F",X"6F",
		X"00",X"00",X"00",X"22",X"33",X"33",X"EF",X"6F",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",
		X"77",X"77",X"77",X"07",X"00",X"00",X"00",X"00",X"4F",X"4F",X"9E",X"3E",X"3F",X"3F",X"77",X"00",
		X"2F",X"2F",X"1F",X"4F",X"CF",X"CF",X"EE",X"00",X"EE",X"EE",X"EE",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"13",X"33",X"33",X"67",X"00",X"01",X"00",X"00",X"00",X"8B",X"8F",X"CF",
		X"00",X"08",X"2E",X"FF",X"5F",X"5F",X"2F",X"2F",X"00",X"00",X"00",X"08",X"8C",X"CE",X"CE",X"EE",
		X"77",X"77",X"77",X"33",X"13",X"00",X"00",X"00",X"4F",X"4F",X"DF",X"DF",X"47",X"33",X"11",X"00",
		X"1F",X"A7",X"2F",X"FF",X"FF",X"CC",X"88",X"00",X"EE",X"08",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"33",X"33",X"00",X"00",X"77",X"33",X"11",X"01",X"03",X"CB",
		X"00",X"00",X"EF",X"FF",X"BF",X"DF",X"6F",X"0F",X"00",X"00",X"08",X"0C",X"8E",X"CE",X"CC",X"08",
		X"33",X"33",X"33",X"33",X"13",X"01",X"00",X"00",X"ED",X"F6",X"FB",X"FD",X"FF",X"EE",X"4C",X"00",
		X"2F",X"97",X"FB",X"FF",X"FF",X"FF",X"22",X"00",X"0C",X"0C",X"8E",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"11",X"77",X"EF",X"77",X"13",X"07",X"07",
		X"00",X"8E",X"EF",X"FF",X"3F",X"EF",X"0F",X"3F",X"00",X"00",X"08",X"08",X"00",X"08",X"0C",X"0E",
		X"77",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"0F",X"CF",X"3F",X"CF",X"FF",X"FF",X"77",X"00",
		X"97",X"5B",X"FF",X"FF",X"FF",X"88",X"88",X"00",X"CE",X"CC",X"CC",X"88",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"33",X"77",X"FC",X"FF",X"03",X"03",
		X"00",X"0F",X"EF",X"EF",X"D2",X"FC",X"3F",X"0F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"EE",X"EE",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"FF",X"CF",X"77",X"33",X"11",X"00",
		X"3C",X"3F",X"CF",X"2F",X"EF",X"EF",X"FF",X"00",X"EE",X"EE",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"11",X"33",X"77",X"00",X"77",X"FF",X"FF",X"DF",X"3F",X"CF",X"0F",
		X"00",X"88",X"88",X"8F",X"1F",X"7F",X"1F",X"79",X"00",X"00",X"00",X"08",X"88",X"CC",X"CC",X"CE",
		X"44",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"07",X"07",X"13",X"FF",X"EF",X"77",X"11",X"00",
		X"3F",X"0F",X"EF",X"3F",X"FF",X"FF",X"EE",X"00",X"8E",X"0C",X"08",X"00",X"88",X"88",X"00",X"00",
		X"00",X"00",X"01",X"03",X"13",X"33",X"33",X"33",X"00",X"0C",X"4E",X"FF",X"CF",X"AF",X"6F",X"CF",
		X"00",X"02",X"1F",X"3F",X"7F",X"BF",X"3D",X"7B",X"00",X"00",X"00",X"88",X"CC",X"EE",X"CC",X"CC",
		X"33",X"33",X"22",X"00",X"00",X"00",X"00",X"00",X"8F",X"03",X"01",X"11",X"33",X"77",X"00",X"00",
		X"3F",X"6F",X"DF",X"BF",X"FF",X"FF",X"00",X"00",X"88",X"8C",X"EE",X"EE",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"03",X"13",X"37",X"37",X"77",X"00",X"01",X"03",X"17",X"5F",X"DF",X"4F",X"4F",
		X"00",X"08",X"EE",X"FF",X"FF",X"2F",X"6B",X"87",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"8E",
		X"67",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"CF",X"8F",X"8B",X"88",X"00",X"00",X"11",X"00",
		X"3F",X"2F",X"5F",X"5F",X"FF",X"EE",X"88",X"00",X"EE",X"EE",X"CE",X"8C",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"37",X"3F",X"3F",X"2F",X"BE",X"4F",X"6F",
		X"00",X"CE",X"CF",X"CF",X"4F",X"D7",X"2F",X"6F",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",
		X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"CC",X"CC",X"44",X"00",X"00",X"00",
		X"EF",X"EF",X"33",X"33",X"22",X"00",X"00",X"00",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"11",X"37",X"77",X"00",X"03",X"7E",X"FF",X"7F",X"7F",X"BF",X"FF",
		X"00",X"0C",X"E7",X"FF",X"EF",X"EF",X"DF",X"FF",X"00",X"00",X"00",X"08",X"00",X"88",X"CE",X"EE",
		X"77",X"77",X"77",X"66",X"66",X"44",X"00",X"00",X"8F",X"06",X"66",X"66",X"00",X"00",X"00",X"00",
		X"1F",X"06",X"66",X"66",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"66",X"66",X"22",X"00",X"00",
		X"00",X"11",X"33",X"13",X"77",X"23",X"23",X"77",X"37",X"97",X"FB",X"FF",X"FF",X"FF",X"FF",X"6F",
		X"8C",X"CE",X"8E",X"BF",X"BF",X"BF",X"9F",X"2E",X"00",X"00",X"00",X"8C",X"CC",X"EE",X"EE",X"FF",
		X"77",X"77",X"77",X"33",X"33",X"11",X"11",X"00",X"0E",X"3F",X"33",X"02",X"00",X"00",X"00",X"00",
		X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"16",X"7F",X"7F",X"BF",X"6F",X"0F",X"DF",X"CF",X"EF",X"EF",X"FF",X"EF",X"CF",
		X"00",X"67",X"FF",X"FF",X"3F",X"0C",X"6E",X"77",X"00",X"00",X"08",X"8C",X"CE",X"EF",X"11",X"00",
		X"33",X"33",X"77",X"77",X"33",X"11",X"00",X"00",X"0E",X"BF",X"BB",X"99",X"CC",X"CC",X"CC",X"66",
		X"23",X"00",X"88",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"13",X"77",X"37",X"1F",X"FB",X"FF",X"00",X"99",X"3F",X"9F",X"CF",X"EF",X"FF",X"EF",
		X"00",X"EE",X"FF",X"FF",X"0C",X"0E",X"7F",X"26",X"00",X"00",X"88",X"EE",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"37",X"11",X"11",X"11",X"00",X"00",X"EF",X"8F",X"DF",X"EE",X"FF",X"FF",X"77",X"00",
		X"00",X"88",X"CC",X"CC",X"00",X"88",X"CC",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"33",X"37",X"17",X"00",X"33",X"33",X"77",X"C3",X"FC",X"FF",X"FF",
		X"00",X"FF",X"FF",X"EE",X"88",X"0F",X"3F",X"08",X"00",X"CC",X"08",X"00",X"00",X"00",X"00",X"00",
		X"71",X"77",X"33",X"13",X"01",X"00",X"00",X"00",X"FF",X"FF",X"DF",X"7F",X"77",X"33",X"33",X"00",
		X"08",X"7F",X"7F",X"88",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"CC",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
