library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity LLANDER_VEC_ROM_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of LLANDER_VEC_ROM_2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"30",X"60",X"00",X"94",X"58",X"C6",X"58",X"FA",X"58",X"2E",X"59",X"48",X"59",X"79",X"59",
		X"9C",X"59",X"10",X"5A",X"36",X"5A",X"86",X"5A",X"D2",X"5A",X"0C",X"5B",X"4E",X"5B",X"82",X"5B",
		X"EA",X"5B",X"36",X"5C",X"8D",X"5C",X"A6",X"5C",X"EC",X"5C",X"6A",X"5D",X"AA",X"5D",X"ED",X"5D",
		X"02",X"5E",X"23",X"5E",X"A5",X"58",X"D7",X"58",X"0B",X"59",X"35",X"59",X"5D",X"59",X"82",X"59",
		X"C5",X"59",X"1D",X"5A",X"55",X"5A",X"9C",X"5A",X"E4",X"5A",X"21",X"5B",X"5F",X"5B",X"A3",X"5B",
		X"06",X"5C",X"47",X"5C",X"AD",X"5C",X"C5",X"5C",X"18",X"5D",X"7C",X"5D",X"C4",X"5D",X"F4",X"5D",
		X"0E",X"5E",X"38",X"5E",X"B1",X"58",X"E7",X"58",X"1A",X"59",X"3D",X"59",X"6B",X"59",X"8B",X"59",
		X"F1",X"59",X"2B",X"5A",X"70",X"5A",X"B1",X"5A",X"FA",X"5A",X"39",X"5B",X"71",X"5B",X"C4",X"5B",
		X"22",X"5C",X"6C",X"5C",X"CE",X"5C",X"E3",X"5C",X"3C",X"5D",X"83",X"5D",X"DA",X"5D",X"FB",X"5D",
		X"1A",X"5E",X"51",X"5E",X"16",X"34",X"34",X"3E",X"46",X"1E",X"38",X"00",X"3A",X"3E",X"38",X"00",
		X"3A",X"3C",X"16",X"38",X"BC",X"34",X"3E",X"2C",X"3A",X"16",X"38",X"00",X"3A",X"3C",X"16",X"38",
		X"BC",X"3A",X"3C",X"16",X"38",X"3C",X"2A",X"30",X"32",X"1E",X"34",X"20",X"1E",X"00",X"1C",X"38",
		X"3E",X"1E",X"1A",X"2A",X"1E",X"B0",X"1A",X"16",X"38",X"18",X"3E",X"38",X"16",X"30",X"3C",X"00",
		X"1C",X"26",X"2E",X"26",X"30",X"3E",X"9E",X"34",X"32",X"1A",X"32",X"00",X"1A",X"32",X"2E",X"18",
		X"3E",X"3A",X"3C",X"26",X"18",X"2C",X"9E",X"3C",X"38",X"1E",X"26",X"18",X"3A",X"3C",X"32",X"20",
		X"20",X"00",X"22",X"1E",X"24",X"3C",X"00",X"16",X"3E",X"BA",X"34",X"2C",X"3E",X"3A",X"00",X"1C",
		X"1E",X"00",X"1A",X"16",X"38",X"18",X"3E",X"38",X"16",X"30",X"BC",X"3A",X"26",X"30",X"00",X"1A",
		X"32",X"2E",X"18",X"3E",X"3A",X"3C",X"26",X"18",X"2C",X"9E",X"3C",X"38",X"1E",X"26",X"18",X"3A",
		X"3C",X"32",X"20",X"20",X"3C",X"16",X"30",X"2A",X"3A",X"00",X"2C",X"1E",X"1E",X"B8",X"34",X"1E",
		X"38",X"1C",X"3E",X"1E",X"BA",X"34",X"1E",X"38",X"1C",X"26",X"1C",X"16",X"BA",X"3C",X"1E",X"26",
		X"2C",X"40",X"1E",X"38",X"2C",X"3E",X"3A",X"BC",X"26",X"30",X"3C",X"38",X"32",X"1C",X"3E",X"26",
		X"38",X"1E",X"00",X"2C",X"1E",X"3A",X"00",X"34",X"26",X"1E",X"1A",X"1E",X"BA",X"26",X"30",X"3A",
		X"1E",X"38",X"3C",X"1E",X"00",X"20",X"26",X"1A",X"24",X"16",X"BA",X"22",X"1E",X"2C",X"1C",X"00",
		X"16",X"3E",X"3A",X"42",X"1E",X"38",X"20",X"1E",X"B0",X"34",X"16",X"38",X"00",X"34",X"26",X"1E",
		X"1A",X"9E",X"34",X"32",X"38",X"00",X"20",X"26",X"1A",X"24",X"96",X"48",X"3E",X"2A",X"16",X"3E",
		X"20",X"00",X"34",X"38",X"32",X"00",X"2E",X"3E",X"1E",X"30",X"48",X"9E",X"38",X"1E",X"3A",X"1E",
		X"38",X"40",X"32",X"26",X"38",X"00",X"16",X"3E",X"44",X"26",X"2C",X"26",X"16",X"26",X"38",X"1E",
		X"00",X"1C",X"1E",X"00",X"1A",X"16",X"38",X"18",X"3E",X"38",X"16",X"30",X"3C",X"00",X"1C",X"1E",
		X"3C",X"38",X"3E",X"26",X"BC",X"3C",X"16",X"30",X"36",X"3E",X"1E",X"3A",X"00",X"16",X"3E",X"44",
		X"26",X"2C",X"26",X"16",X"38",X"1E",X"3A",X"00",X"1C",X"1E",X"00",X"1A",X"32",X"2E",X"18",X"3E",
		X"3A",X"3C",X"26",X"18",X"2C",X"1E",X"00",X"1C",X"1E",X"3A",X"3C",X"38",X"3E",X"26",X"1C",X"32",
		X"BA",X"48",X"3E",X"3A",X"16",X"3C",X"48",X"3C",X"38",X"1E",X"26",X"18",X"3A",X"3C",X"32",X"20",
		X"20",X"3C",X"16",X"30",X"2A",X"3A",X"00",X"48",X"1E",X"38",X"3A",X"3C",X"32",X"1E",X"38",X"BC",
		X"20",X"1E",X"2C",X"26",X"1A",X"26",X"3C",X"16",X"3C",X"26",X"32",X"30",X"BA",X"20",X"1E",X"2C",
		X"26",X"1A",X"26",X"3C",X"16",X"1A",X"26",X"32",X"30",X"1E",X"BA",X"22",X"38",X"16",X"3C",X"3E",
		X"2C",X"16",X"3C",X"26",X"32",X"B0",X"40",X"32",X"3E",X"3A",X"00",X"16",X"40",X"1E",X"48",X"00",
		X"16",X"3C",X"3C",X"1E",X"38",X"38",X"26",X"00",X"1C",X"26",X"20",X"20",X"26",X"1A",X"26",X"2C",
		X"1E",X"2E",X"1E",X"30",X"BC",X"3E",X"3A",X"3C",X"1E",X"1C",X"00",X"16",X"2C",X"3E",X"30",X"26",
		X"48",X"32",X"00",X"40",X"26",X"32",X"2C",X"1E",X"30",X"3C",X"16",X"2E",X"1E",X"30",X"3C",X"9E",
		X"3A",X"26",X"1E",X"00",X"3A",X"26",X"30",X"1C",X"00",X"24",X"16",X"38",X"3C",X"00",X"22",X"1E",
		X"2C",X"16",X"30",X"1C",X"1E",X"BC",X"3A",X"34",X"2C",X"1E",X"30",X"1C",X"26",X"1C",X"1E",X"00",
		X"16",X"3C",X"3C",X"1E",X"38",X"38",X"26",X"3A",X"3A",X"16",X"22",X"9E",X"20",X"3E",X"1E",X"00",
		X"3E",X"30",X"00",X"22",X"38",X"16",X"30",X"00",X"16",X"2C",X"3E",X"30",X"26",X"48",X"16",X"28",
		X"9E",X"1C",X"26",X"1E",X"3A",X"00",X"42",X"16",X"38",X"00",X"1E",X"26",X"30",X"1E",X"00",X"22",
		X"38",X"32",X"3A",X"3A",X"16",X"38",X"3C",X"26",X"22",X"1E",X"00",X"2C",X"16",X"30",X"1C",X"3E",
		X"30",X"A2",X"2C",X"1E",X"00",X"1E",X"16",X"22",X"2C",X"1E",X"00",X"16",X"00",X"16",X"3C",X"3C",
		X"1E",X"38",X"38",X"A6",X"1E",X"2C",X"00",X"16",X"22",X"3E",X"26",X"2C",X"16",X"00",X"24",X"16",
		X"00",X"16",X"2C",X"3E",X"30",X"26",X"48",X"16",X"1C",X"B2",X"1E",X"16",X"22",X"2C",X"1E",X"00",
		X"26",X"3A",X"3C",X"00",X"22",X"1E",X"2C",X"16",X"30",X"1C",X"1E",X"BC",X"2C",X"1E",X"00",X"1A",
		X"32",X"2C",X"3E",X"2E",X"18",X"26",X"16",X"00",X"16",X"00",X"16",X"3C",X"3C",X"1E",X"38",X"38",
		X"A6",X"1E",X"2C",X"00",X"1A",X"32",X"2C",X"3E",X"2E",X"18",X"26",X"16",X"00",X"24",X"16",X"00",
		X"16",X"2C",X"3E",X"30",X"26",X"48",X"16",X"1C",X"B2",X"1A",X"32",X"2C",X"3E",X"2E",X"18",X"26",
		X"16",X"00",X"26",X"3A",X"3C",X"00",X"22",X"1E",X"2C",X"16",X"30",X"1C",X"1E",X"BC",X"40",X"32",
		X"3E",X"3A",X"00",X"16",X"40",X"1E",X"48",X"00",X"16",X"3C",X"3C",X"1E",X"38",X"38",X"A6",X"3E",
		X"3A",X"3C",X"1E",X"1C",X"00",X"24",X"16",X"00",X"16",X"2C",X"3E",X"30",X"26",X"48",X"16",X"1C",
		X"B2",X"3A",X"26",X"1E",X"00",X"3A",X"26",X"30",X"1C",X"00",X"22",X"1E",X"2C",X"16",X"30",X"1C",
		X"1E",X"BC",X"2C",X"1E",X"00",X"3A",X"3E",X"34",X"34",X"32",X"38",X"3C",X"00",X"1C",X"1E",X"00",
		X"3A",X"16",X"3E",X"40",X"1E",X"3C",X"16",X"22",X"1E",X"00",X"1E",X"3A",X"3C",X"00",X"34",X"16",
		X"38",X"3C",X"A6",X"1E",X"36",X"3E",X"26",X"34",X"32",X"00",X"1C",X"1E",X"00",X"3A",X"3E",X"34",
		X"1E",X"38",X"40",X"26",X"40",X"1E",X"30",X"1A",X"26",X"16",X"00",X"1C",X"1E",X"3A",X"3C",X"38",
		X"3E",X"26",X"1C",X"B2",X"2C",X"1E",X"18",X"1E",X"30",X"3A",X"38",X"1E",X"3C",X"3C",X"3E",X"30",
		X"22",X"3A",X"3A",X"46",X"3A",X"3C",X"1E",X"2E",X"1E",X"00",X"3A",X"26",X"30",X"1C",X"00",X"16",
		X"3E",X"3A",X"22",X"1E",X"20",X"16",X"2C",X"2C",X"1E",X"B0",X"40",X"32",X"3C",X"38",X"1E",X"00",
		X"40",X"32",X"46",X"16",X"22",X"1E",X"00",X"1E",X"3A",X"3C",X"00",X"3A",X"16",X"30",X"3A",X"00",
		X"38",X"1E",X"3C",X"32",X"3E",X"B8",X"3A",X"3E",X"00",X"40",X"26",X"16",X"28",X"1E",X"00",X"1E",
		X"3A",X"00",X"1C",X"1E",X"00",X"26",X"1C",X"16",X"00",X"3A",X"32",X"2C",X"16",X"2E",X"1E",X"30",
		X"3C",X"9E",X"38",X"1E",X"26",X"3A",X"1E",X"00",X"32",X"24",X"30",X"1E",X"00",X"38",X"3E",X"1E",
		X"1A",X"2A",X"2A",X"1E",X"24",X"B8",X"34",X"1E",X"38",X"1C",X"3E",X"00",X"3A",X"16",X"30",X"3A",
		X"00",X"1E",X"3A",X"34",X"32",X"26",X"B8",X"2C",X"16",X"2E",X"1E",X"30",X"3C",X"16",X"18",X"2C",
		X"1E",X"2E",X"1E",X"30",X"3C",X"1E",X"00",X"3E",X"3A",X"3C",X"1E",X"1C",X"00",X"30",X"32",X"00",
		X"34",X"3E",X"1E",X"1C",X"1E",X"00",X"40",X"32",X"2C",X"40",X"1E",X"B8",X"2A",X"1E",X"26",X"30",
		X"00",X"38",X"3E",X"1E",X"1A",X"2A",X"3A",X"3C",X"16",X"38",X"3C",X"00",X"48",X"3E",X"38",X"00",
		X"1E",X"38",X"1C",X"1E",X"00",X"2E",X"32",X"1E",X"22",X"2C",X"26",X"1A",X"A4",X"3A",X"46",X"3A",
		X"3C",X"1E",X"2E",X"1E",X"00",X"1C",X"1E",X"00",X"1A",X"32",X"2E",X"2E",X"3E",X"30",X"26",X"1A",
		X"16",X"3C",X"26",X"32",X"30",X"00",X"1C",X"1E",X"3C",X"38",X"3E",X"26",X"BC",X"3A",X"26",X"3A",
		X"3C",X"1E",X"2E",X"16",X"00",X"1C",X"1E",X"00",X"1A",X"32",X"2E",X"3E",X"30",X"26",X"1A",X"16",
		X"1A",X"26",X"32",X"30",X"00",X"1C",X"1E",X"3A",X"3C",X"38",X"3E",X"26",X"1C",X"B2",X"2A",X"32",
		X"2E",X"2E",X"3E",X"30",X"26",X"2A",X"16",X"3C",X"26",X"32",X"30",X"3A",X"3A",X"46",X"3A",X"3C",
		X"1E",X"2E",X"00",X"48",X"1E",X"38",X"3A",X"3C",X"32",X"1E",X"38",X"BC",X"40",X"32",X"3E",X"3A",
		X"00",X"16",X"40",X"1E",X"48",X"00",X"1A",X"38",X"1E",X"1E",X"00",X"3E",X"30",X"00",X"1A",X"38",
		X"16",X"3C",X"1E",X"38",X"1E",X"00",X"1C",X"1E",X"00",X"1C",X"1E",X"3E",X"44",X"00",X"2A",X"26",
		X"2C",X"32",X"2E",X"1E",X"3C",X"38",X"1E",X"BA",X"3E",X"3A",X"3C",X"1E",X"1C",X"00",X"1A",X"38",
		X"1E",X"32",X"00",X"3E",X"30",X"00",X"1A",X"38",X"16",X"3C",X"1E",X"38",X"00",X"1C",X"1E",X"00",
		X"06",X"00",X"2A",X"26",X"2C",X"32",X"2E",X"1E",X"3C",X"38",X"32",X"BA",X"3A",X"26",X"1E",X"00",
		X"24",X"16",X"18",X"1E",X"30",X"00",X"1E",X"26",X"30",X"1E",X"30",X"00",X"06",X"00",X"2A",X"26",
		X"2C",X"32",X"2E",X"1E",X"3C",X"1E",X"38",X"00",X"2A",X"38",X"16",X"3C",X"1E",X"38",X"00",X"16",
		X"3E",X"20",X"22",X"1E",X"38",X"26",X"3A",X"3A",X"1E",X"B0",X"40",X"32",X"3E",X"3A",X"00",X"16",
		X"40",X"1E",X"48",X"00",X"3E",X"30",X"00",X"1A",X"38",X"16",X"3A",X"A4",X"1C",X"1E",X"2E",X"32",
		X"2C",X"1E",X"B8",X"0C",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"00",X"2E",X"16",
		X"38",X"2A",X"00",X"3A",X"26",X"30",X"1C",X"00",X"26",X"30",X"00",X"1C",X"26",X"1E",X"00",X"2C",
		X"3E",X"20",X"3C",X"00",X"22",X"1E",X"28",X"16",X"22",X"BC",X"26",X"2C",X"00",X"30",X"1E",X"46",
		X"00",X"16",X"00",X"34",X"16",X"3A",X"00",X"1C",X"1E",X"00",X"3A",X"3E",X"38",X"40",X"26",X"40",
		X"16",X"30",X"3C",X"BA",X"30",X"32",X"00",X"24",X"3E",X"18",X"32",X"00",X"3A",X"32",X"18",X"38",
		X"1E",X"40",X"26",X"40",X"26",X"1E",X"30",X"3C",X"1E",X"BA",X"2A",X"1E",X"26",X"30",X"1E",X"00",
		X"3E",X"1E",X"18",X"1E",X"38",X"2C",X"1E",X"18",X"1E",X"30",X"1C",X"1E",X"B0",X"00",X"34",X"32",
		X"26",X"30",X"3C",X"BA",X"00",X"34",X"3E",X"30",X"3C",X"32",X"BA",X"00",X"34",X"3E",X"30",X"2A",
		X"3C",X"9E",X"1A",X"24",X"32",X"26",X"44",X"00",X"1C",X"3E",X"00",X"28",X"1E",X"BE",X"1E",X"2C",
		X"1E",X"22",X"26",X"38",X"00",X"28",X"3E",X"1E",X"22",X"B2",X"3A",X"34",X"26",X"1E",X"2C",X"42",
		X"16",X"24",X"AC",X"00",X"3E",X"30",X"26",X"3C",X"1E",X"3A",X"00",X"1C",X"1E",X"00",X"1A",X"16",
		X"38",X"18",X"3E",X"38",X"16",X"30",X"3C",X"80",X"00",X"3E",X"30",X"26",X"1C",X"16",X"1C",X"1E",
		X"3A",X"00",X"1C",X"1E",X"00",X"1A",X"32",X"2E",X"18",X"3E",X"3A",X"3C",X"26",X"18",X"2C",X"1E",
		X"80",X"00",X"3C",X"38",X"1E",X"26",X"18",X"3A",X"3C",X"32",X"20",X"20",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"5E",X"D5",X"5E",X"33",X"5F",X"EC",
		X"A2",X"28",X"00",X"00",X"70",X"00",X"00",X"3A",X"1A",X"32",X"38",X"9E",X"C0",X"55",X"C0",X"07",
		X"1C",X"3E",X"38",X"1E",X"1E",X"00",X"1C",X"3E",X"00",X"28",X"1E",X"BE",X"70",X"74",X"40",X"06",
		X"1A",X"32",X"2E",X"18",X"3E",X"3A",X"3C",X"26",X"18",X"2C",X"9E",X"70",X"80",X"40",X"03",X"16",
		X"2C",X"3C",X"26",X"3C",X"3E",X"1C",X"9E",X"E0",X"64",X"00",X"07",X"40",X"26",X"3C",X"1E",X"3A",
		X"3A",X"1E",X"00",X"24",X"32",X"38",X"26",X"48",X"32",X"30",X"3C",X"16",X"2C",X"9E",X"70",X"74",
		X"90",X"07",X"40",X"26",X"3C",X"1E",X"3A",X"3A",X"1E",X"00",X"40",X"1E",X"38",X"3C",X"26",X"1A",
		X"16",X"2C",X"9E",X"00",X"D0",X"EC",X"A2",X"64",X"00",X"00",X"70",X"00",X"00",X"34",X"3E",X"30",
		X"3C",X"16",X"28",X"9E",X"E0",X"64",X"A0",X"06",X"3C",X"26",X"1E",X"2E",X"34",X"B2",X"E0",X"64",
		X"40",X"06",X"34",X"1E",X"3C",X"38",X"32",X"AC",X"70",X"80",X"10",X"03",X"16",X"2C",X"3C",X"26",
		X"3C",X"3E",X"9C",X"E0",X"64",X"A0",X"06",X"40",X"1E",X"2C",X"32",X"1A",X"26",X"1C",X"16",X"1C",
		X"00",X"24",X"32",X"38",X"26",X"48",X"32",X"30",X"3C",X"16",X"AC",X"70",X"74",X"C0",X"07",X"40",
		X"1E",X"2C",X"32",X"1A",X"26",X"1C",X"16",X"1C",X"00",X"40",X"1E",X"38",X"3C",X"26",X"1A",X"16",
		X"AC",X"00",X"D0",X"EC",X"A2",X"4C",X"00",X"00",X"70",X"00",X"00",X"34",X"3E",X"30",X"2A",X"3C",
		X"48",X"16",X"24",X"AC",X"E0",X"64",X"60",X"07",X"38",X"1E",X"3A",X"3C",X"48",X"1E",X"26",X"BC",
		X"E0",X"64",X"00",X"07",X"34",X"1E",X"3C",X"38",X"32",X"AC",X"70",X"80",X"B0",X"02",X"24",X"32",
		X"1E",X"24",X"9E",X"C0",X"55",X"C0",X"07",X"24",X"32",X"38",X"26",X"48",X"32",X"30",X"3C",X"16",
		X"2C",X"1E",X"00",X"22",X"1E",X"3A",X"1A",X"24",X"42",X"26",X"30",X"1C",X"26",X"22",X"2A",X"1E",
		X"26",X"BC",X"38",X"84",X"88",X"06",X"40",X"1E",X"38",X"3C",X"26",X"2A",X"16",X"2C",X"1E",X"00",
		X"22",X"1E",X"3A",X"1A",X"24",X"42",X"26",X"30",X"1C",X"26",X"22",X"2A",X"1E",X"26",X"BC",X"00",
		X"D0",X"00",X"1D",X"3A",X"EB",X"EE",X"EE",X"F7",X"E5",X"FD",X"DF",X"06",X"D0",X"06",X"12",X"09",
		X"15",X"F7",X"06",X"27",X"FA",X"63",X"F4",X"42",X"2A",X"00",X"03",X"E5",X"00",X"00",X"00",X"00",
		X"00",X"FA",X"F1",X"F4",X"F4",X"FA",X"FD",X"D6",X"03",X"DC",X"09",X"06",X"00",X"12",X"F7",X"06",
		X"EB",X"F7",X"5D",X"0C",X"63",X"36",X"00",X"03",X"D9",X"00",X"00",X"00",X"00",X"00",X"DF",X"E8",
		X"E5",X"EB",X"FA",X"E5",X"FD",X"0C",X"EB",X"E5",X"12",X"09",X"15",X"E8",X"1E",X"F7",X"00",X"5D",
		X"EE",X"03",X"3F",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
