library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MRDONIGHTMARE_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MRDONIGHTMARE_ROM_PGM_0 is
	type rom is array(0 to  10239) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"70",X"C3",X"D0",X"00",X"3A",X"36",X"40",X"3C",X"E6",X"07",X"32",X"36",X"40",
		X"20",X"1A",X"06",X"1A",X"11",X"09",X"58",X"1A",X"FE",X"05",X"28",X"09",X"FE",X"06",X"20",X"08",
		X"3E",X"05",X"12",X"18",X"03",X"3E",X"06",X"12",X"13",X"13",X"10",X"EB",X"C9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"01",X"70",X"3A",X"00",X"40",X"3C",X"32",X"00",X"40",X"3A",X"35",X"40",X"3C",X"32",X"35",X"40",
		X"CD",X"07",X"00",X"CD",X"FB",X"1B",X"AF",X"32",X"05",X"68",X"3A",X"00",X"60",X"CB",X"47",X"20",
		X"06",X"AF",X"32",X"02",X"40",X"18",X"18",X"3A",X"02",X"40",X"B7",X"20",X"12",X"3E",X"01",X"32",
		X"02",X"40",X"3A",X"01",X"40",X"37",X"3F",X"3C",X"27",X"32",X"01",X"40",X"CD",X"1D",X"17",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3A",X"00",X"78",X"3E",X"01",X"32",X"01",X"70",X"F1",X"C9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"00",X"50",X"06",X"04",X"3E",X"10",X"77",X"2C",X"20",X"FC",X"24",X"3A",X"00",X"78",X"10",
		X"F4",X"21",X"00",X"58",X"AF",X"77",X"2C",X"20",X"FC",X"3E",X"01",X"21",X"00",X"60",X"06",X"08",
		X"77",X"23",X"10",X"FC",X"AF",X"21",X"00",X"68",X"06",X"08",X"77",X"23",X"10",X"FC",X"06",X"08",
		X"21",X"01",X"70",X"77",X"23",X"10",X"FC",X"3D",X"32",X"00",X"78",X"3A",X"00",X"78",X"06",X"04",
		X"21",X"00",X"40",X"AF",X"77",X"2C",X"20",X"FC",X"24",X"3A",X"00",X"78",X"10",X"F5",X"31",X"00",
		X"44",X"18",X"1D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"64",X"14",X"3E",X"01",X"32",X"07",X"68",X"3E",X"01",X"32",X"01",X"70",X"CD",X"70",X"14",
		X"AF",X"32",X"06",X"70",X"32",X"07",X"70",X"CD",X"6B",X"15",X"CD",X"AD",X"14",X"AF",X"32",X"30",
		X"40",X"3E",X"03",X"32",X"37",X"40",X"3E",X"01",X"32",X"32",X"40",X"AF",X"CD",X"B8",X"0E",X"CD",
		X"C5",X"02",X"CD",X"F5",X"12",X"3A",X"00",X"78",X"CD",X"B9",X"14",X"3A",X"33",X"40",X"CD",X"B8",
		X"0E",X"CD",X"93",X"0F",X"CD",X"87",X"13",X"CD",X"B4",X"0F",X"CD",X"5F",X"13",X"AF",X"32",X"35",
		X"40",X"3A",X"40",X"40",X"32",X"40",X"58",X"3A",X"41",X"40",X"32",X"43",X"58",X"AF",X"32",X"4A",
		X"40",X"32",X"42",X"40",X"32",X"43",X"40",X"32",X"57",X"40",X"32",X"59",X"40",X"32",X"5B",X"40",
		X"32",X"44",X"58",X"32",X"48",X"58",X"32",X"4C",X"58",X"CD",X"E2",X"0F",X"CD",X"74",X"0C",X"21",
		X"9C",X"1C",X"3A",X"45",X"40",X"B7",X"28",X"03",X"21",X"8B",X"1D",X"AF",X"CD",X"70",X"1C",X"3A",
		X"40",X"58",X"E6",X"0F",X"20",X"1B",X"3A",X"43",X"58",X"E6",X"0F",X"20",X"14",X"CD",X"74",X"02",
		X"B7",X"20",X"1A",X"3A",X"43",X"40",X"B7",X"28",X"11",X"47",X"AF",X"32",X"43",X"40",X"78",X"18",
		X"0C",X"CD",X"74",X"02",X"B7",X"28",X"03",X"32",X"43",X"40",X"3A",X"42",X"40",X"CB",X"57",X"C2",
		X"20",X"03",X"CB",X"5F",X"C2",X"4B",X"03",X"CB",X"47",X"C2",X"76",X"03",X"CB",X"4F",X"C2",X"A1",
		X"03",X"CD",X"83",X"05",X"CD",X"98",X"07",X"CD",X"BC",X"13",X"CD",X"B6",X"11",X"3A",X"3A",X"40",
		X"FE",X"1F",X"CA",X"B9",X"10",X"3A",X"2E",X"40",X"B7",X"28",X"07",X"3A",X"00",X"68",X"CB",X"4F",
		X"20",X"17",X"3A",X"44",X"40",X"B7",X"20",X"34",X"CD",X"7F",X"12",X"3A",X"4A",X"40",X"FE",X"04",
		X"20",X"2A",X"3A",X"45",X"40",X"B7",X"C2",X"2F",X"11",X"3A",X"32",X"40",X"37",X"3F",X"3C",X"27",
		X"32",X"32",X"40",X"3A",X"33",X"40",X"3C",X"32",X"33",X"40",X"FE",X"0C",X"20",X"0B",X"AF",X"32",
		X"33",X"40",X"3A",X"34",X"40",X"3C",X"32",X"34",X"40",X"C3",X"75",X"01",X"3E",X"01",X"CD",X"D5",
		X"0C",X"C3",X"CF",X"01",X"C5",X"AF",X"4F",X"3A",X"00",X"60",X"CB",X"57",X"28",X"04",X"79",X"C6",
		X"04",X"4F",X"3A",X"00",X"60",X"CB",X"5F",X"28",X"04",X"79",X"C6",X"08",X"4F",X"3A",X"00",X"60",
		X"CB",X"67",X"28",X"04",X"79",X"C6",X"10",X"4F",X"3A",X"00",X"68",X"CB",X"57",X"28",X"04",X"79",
		X"C6",X"01",X"4F",X"3A",X"00",X"68",X"CB",X"5F",X"28",X"04",X"79",X"C6",X"02",X"4F",X"79",X"C1",
		X"C9",X"3A",X"30",X"40",X"B7",X"28",X"02",X"18",X"0C",X"01",X"0D",X"01",X"21",X"32",X"40",X"11",
		X"3F",X"41",X"ED",X"B0",X"C9",X"01",X"0D",X"01",X"21",X"32",X"40",X"11",X"4C",X"42",X"ED",X"B0",
		X"C9",X"3A",X"30",X"40",X"B7",X"28",X"02",X"18",X"0C",X"01",X"0D",X"01",X"21",X"3F",X"41",X"11",
		X"32",X"40",X"ED",X"B0",X"C9",X"01",X"0D",X"01",X"21",X"4C",X"42",X"11",X"32",X"40",X"ED",X"B0",
		X"C9",X"3A",X"2F",X"40",X"B7",X"C8",X"3A",X"30",X"40",X"EE",X"01",X"32",X"30",X"40",X"CD",X"D1",
		X"02",X"3A",X"37",X"40",X"B7",X"28",X"EF",X"CD",X"87",X"13",X"CD",X"DC",X"13",X"CD",X"5F",X"13",
		X"3A",X"2D",X"40",X"B7",X"28",X"09",X"3A",X"30",X"40",X"32",X"06",X"70",X"32",X"07",X"70",X"C9",
		X"32",X"42",X"40",X"CD",X"DC",X"03",X"38",X"20",X"CD",X"61",X"04",X"3A",X"40",X"58",X"3D",X"32",
		X"40",X"58",X"E6",X"0F",X"01",X"00",X"00",X"DD",X"21",X"CC",X"03",X"4F",X"DD",X"09",X"DD",X"7E",
		X"00",X"4F",X"3E",X"14",X"81",X"32",X"41",X"58",X"C3",X"11",X"02",X"32",X"42",X"40",X"CD",X"1C",
		X"04",X"38",X"20",X"CD",X"C3",X"04",X"3A",X"40",X"58",X"3C",X"32",X"40",X"58",X"E6",X"0F",X"01",
		X"00",X"00",X"DD",X"21",X"CC",X"03",X"4F",X"DD",X"09",X"DD",X"7E",X"00",X"4F",X"3E",X"94",X"81",
		X"32",X"41",X"58",X"C3",X"11",X"02",X"32",X"42",X"40",X"CD",X"30",X"04",X"38",X"20",X"CD",X"E0",
		X"04",X"3A",X"43",X"58",X"3D",X"32",X"43",X"58",X"E6",X"0F",X"01",X"00",X"00",X"DD",X"21",X"CC",
		X"03",X"4F",X"DD",X"09",X"DD",X"7E",X"00",X"4F",X"3E",X"17",X"81",X"32",X"41",X"58",X"C3",X"11",
		X"02",X"32",X"42",X"40",X"CD",X"4A",X"04",X"38",X"20",X"CD",X"04",X"05",X"3A",X"43",X"58",X"3C",
		X"32",X"43",X"58",X"E6",X"0F",X"01",X"00",X"00",X"DD",X"21",X"CC",X"03",X"4F",X"DD",X"09",X"DD",
		X"7E",X"00",X"4F",X"3E",X"57",X"81",X"32",X"41",X"58",X"C3",X"11",X"02",X"01",X"01",X"01",X"01",
		X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"3A",X"40",X"58",X"E6",
		X"0F",X"20",X"2D",X"3A",X"40",X"58",X"FE",X"20",X"28",X"24",X"CD",X"25",X"05",X"2B",X"7E",X"FE",
		X"00",X"28",X"1B",X"FE",X"02",X"28",X"17",X"FE",X"06",X"CA",X"1B",X"0C",X"FE",X"07",X"28",X"0E",
		X"FE",X"0D",X"28",X"0A",X"FE",X"0E",X"28",X"06",X"FE",X"0F",X"28",X"07",X"18",X"02",X"37",X"C9",
		X"37",X"3F",X"C9",X"3A",X"4A",X"40",X"FE",X"03",X"20",X"F4",X"18",X"F4",X"3A",X"40",X"58",X"E6",
		X"0F",X"20",X"ED",X"3A",X"40",X"58",X"FE",X"D0",X"28",X"E4",X"CD",X"25",X"05",X"23",X"18",X"BE",
		X"3A",X"43",X"58",X"E6",X"0F",X"20",X"D9",X"3A",X"43",X"58",X"FE",X"20",X"28",X"D0",X"CD",X"25",
		X"05",X"11",X"10",X"00",X"37",X"3F",X"ED",X"52",X"18",X"A4",X"3A",X"43",X"58",X"E6",X"0F",X"20",
		X"BF",X"3A",X"43",X"58",X"FE",X"E0",X"28",X"B6",X"CD",X"25",X"05",X"11",X"10",X"00",X"19",X"18",
		X"8D",X"3A",X"40",X"58",X"E6",X"0F",X"FE",X"08",X"20",X"58",X"3A",X"40",X"58",X"C6",X"08",X"32",
		X"2C",X"41",X"3A",X"43",X"58",X"32",X"2D",X"41",X"CD",X"31",X"05",X"2B",X"7E",X"FE",X"03",X"28",
		X"1C",X"FE",X"04",X"28",X"13",X"FE",X"05",X"20",X"39",X"3E",X"20",X"CD",X"BC",X"0D",X"3A",X"4D",
		X"40",X"B7",X"20",X"0E",X"3C",X"32",X"4D",X"40",X"3E",X"20",X"CD",X"BC",X"0D",X"3E",X"10",X"CD",
		X"BC",X"0D",X"3A",X"44",X"40",X"3D",X"32",X"44",X"40",X"3E",X"01",X"E5",X"21",X"64",X"1F",X"CD",
		X"70",X"1C",X"E1",X"3E",X"01",X"77",X"CD",X"4D",X"05",X"3E",X"01",X"CD",X"04",X"0E",X"CD",X"7D",
		X"0D",X"C9",X"C9",X"3A",X"40",X"58",X"E6",X"0F",X"FE",X"08",X"20",X"F6",X"3A",X"40",X"58",X"D6",
		X"08",X"32",X"2C",X"41",X"3A",X"43",X"58",X"32",X"2D",X"41",X"CD",X"31",X"05",X"23",X"18",X"9C",
		X"3A",X"43",X"58",X"E6",X"0F",X"FE",X"08",X"20",X"D9",X"3A",X"43",X"58",X"C6",X"08",X"32",X"2D",
		X"41",X"3A",X"40",X"58",X"32",X"2C",X"41",X"CD",X"31",X"05",X"11",X"10",X"00",X"37",X"3F",X"ED",
		X"52",X"C3",X"7C",X"04",X"3A",X"43",X"58",X"E6",X"0F",X"FE",X"08",X"20",X"B5",X"3A",X"43",X"58",
		X"D6",X"08",X"32",X"2D",X"41",X"3A",X"40",X"58",X"32",X"2C",X"41",X"CD",X"31",X"05",X"11",X"10",
		X"00",X"19",X"C3",X"7C",X"04",X"3A",X"40",X"58",X"32",X"2C",X"41",X"3A",X"43",X"58",X"32",X"2D",
		X"41",X"3A",X"2C",X"41",X"D6",X"20",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"3A",
		X"2D",X"41",X"D6",X"20",X"85",X"6F",X"26",X"00",X"11",X"5C",X"40",X"19",X"C9",X"D5",X"E5",X"11",
		X"5C",X"40",X"37",X"3F",X"ED",X"52",X"7D",X"E6",X"0F",X"CB",X"27",X"C6",X"02",X"47",X"7D",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"27",X"C6",X"04",X"4F",X"E1",X"D1",X"C9",X"79",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"B0",X"06",X"00",X"4F",X"DD",X"21",X"5C",X"40",
		X"DD",X"09",X"C9",X"3A",X"55",X"40",X"3C",X"32",X"55",X"40",X"47",X"3A",X"54",X"40",X"B8",X"30",
		X"22",X"AF",X"32",X"55",X"40",X"3A",X"53",X"40",X"E6",X"01",X"28",X"03",X"CD",X"E7",X"05",X"3A",
		X"53",X"40",X"E6",X"02",X"28",X"03",X"CD",X"4C",X"06",X"3A",X"53",X"40",X"E6",X"04",X"28",X"03",
		X"CD",X"B1",X"06",X"CD",X"16",X"07",X"CD",X"30",X"07",X"CD",X"4A",X"07",X"3A",X"50",X"58",X"57",
		X"3A",X"53",X"58",X"5F",X"CD",X"64",X"07",X"DA",X"1B",X"0C",X"3A",X"54",X"58",X"57",X"3A",X"57",
		X"58",X"5F",X"CD",X"64",X"07",X"DA",X"1B",X"0C",X"3A",X"58",X"58",X"57",X"3A",X"5B",X"58",X"5F",
		X"CD",X"64",X"07",X"DA",X"1B",X"0C",X"C9",X"3A",X"57",X"40",X"B7",X"20",X"47",X"3A",X"56",X"40",
		X"47",X"3A",X"47",X"58",X"80",X"32",X"47",X"58",X"FE",X"20",X"28",X"04",X"FE",X"E0",X"20",X"06",
		X"78",X"ED",X"44",X"32",X"56",X"40",X"3A",X"47",X"58",X"E6",X"0F",X"20",X"27",X"3A",X"47",X"58",
		X"E6",X"F0",X"47",X"3A",X"43",X"58",X"E6",X"F0",X"B8",X"20",X"19",X"3E",X"01",X"32",X"05",X"68",
		X"32",X"57",X"40",X"3E",X"1E",X"32",X"45",X"58",X"3A",X"44",X"58",X"32",X"50",X"58",X"3A",X"47",
		X"58",X"32",X"53",X"58",X"3A",X"57",X"40",X"B7",X"28",X"11",X"FE",X"10",X"30",X"0D",X"3C",X"32",
		X"57",X"40",X"FE",X"10",X"20",X"05",X"3E",X"1D",X"32",X"45",X"58",X"C9",X"3A",X"59",X"40",X"B7",
		X"20",X"47",X"3A",X"58",X"40",X"47",X"3A",X"4B",X"58",X"80",X"32",X"4B",X"58",X"FE",X"20",X"28",
		X"04",X"FE",X"E0",X"20",X"06",X"78",X"ED",X"44",X"32",X"58",X"40",X"3A",X"4B",X"58",X"E6",X"0F",
		X"20",X"27",X"3A",X"4B",X"58",X"E6",X"F0",X"47",X"3A",X"43",X"58",X"E6",X"F0",X"B8",X"20",X"19",
		X"3E",X"01",X"32",X"05",X"68",X"32",X"59",X"40",X"3E",X"9E",X"32",X"49",X"58",X"3A",X"48",X"58",
		X"32",X"54",X"58",X"3A",X"4B",X"58",X"32",X"57",X"58",X"3A",X"59",X"40",X"B7",X"28",X"11",X"FE",
		X"10",X"30",X"0D",X"3C",X"32",X"59",X"40",X"FE",X"10",X"20",X"05",X"3E",X"9D",X"32",X"49",X"58",
		X"C9",X"3A",X"5B",X"40",X"B7",X"20",X"47",X"3A",X"5A",X"40",X"47",X"3A",X"4C",X"58",X"80",X"32",
		X"4C",X"58",X"FE",X"20",X"28",X"04",X"FE",X"D0",X"20",X"06",X"78",X"ED",X"44",X"32",X"5A",X"40",
		X"3A",X"4C",X"58",X"E6",X"0F",X"20",X"27",X"3A",X"4C",X"58",X"E6",X"F0",X"47",X"3A",X"40",X"58",
		X"E6",X"F0",X"B8",X"20",X"19",X"3E",X"01",X"32",X"05",X"68",X"32",X"5B",X"40",X"3E",X"62",X"32",
		X"4D",X"58",X"3A",X"4C",X"58",X"32",X"58",X"58",X"3A",X"4F",X"58",X"32",X"5B",X"58",X"3A",X"5B",
		X"40",X"B7",X"28",X"11",X"FE",X"10",X"30",X"0D",X"3C",X"32",X"5B",X"40",X"FE",X"10",X"20",X"05",
		X"3E",X"61",X"32",X"4D",X"58",X"C9",X"3A",X"57",X"40",X"B7",X"28",X"13",X"3A",X"50",X"58",X"3C",
		X"3C",X"32",X"50",X"58",X"FE",X"D8",X"20",X"07",X"AF",X"32",X"50",X"58",X"32",X"57",X"40",X"C9",
		X"3A",X"59",X"40",X"B7",X"28",X"13",X"3A",X"54",X"58",X"3D",X"3D",X"32",X"54",X"58",X"FE",X"18",
		X"20",X"07",X"AF",X"32",X"54",X"58",X"32",X"59",X"40",X"C9",X"3A",X"5B",X"40",X"B7",X"28",X"13",
		X"3A",X"5B",X"58",X"3C",X"3C",X"32",X"5B",X"58",X"FE",X"E8",X"20",X"07",X"AF",X"32",X"58",X"58",
		X"32",X"5B",X"40",X"C9",X"7A",X"C6",X"04",X"4F",X"3A",X"40",X"58",X"C6",X"04",X"CD",X"7F",X"07",
		X"30",X"0C",X"7B",X"C6",X"04",X"4F",X"3A",X"43",X"58",X"C6",X"04",X"CD",X"7F",X"07",X"C9",X"47",
		X"B8",X"38",X"08",X"79",X"90",X"FE",X"08",X"38",X"0D",X"18",X"08",X"78",X"91",X"FE",X"08",X"38",
		X"05",X"18",X"00",X"37",X"3F",X"C9",X"37",X"C9",X"3A",X"45",X"40",X"B7",X"C0",X"3A",X"4D",X"40",
		X"B7",X"20",X"4C",X"3A",X"4B",X"40",X"3C",X"32",X"4B",X"40",X"FE",X"3C",X"38",X"40",X"AF",X"32",
		X"4B",X"40",X"3A",X"4C",X"40",X"FE",X"01",X"20",X"12",X"3A",X"5C",X"58",X"C6",X"10",X"32",X"5C",
		X"58",X"3A",X"3B",X"40",X"CB",X"27",X"32",X"3B",X"40",X"18",X"10",X"3A",X"5C",X"58",X"D6",X"10",
		X"32",X"5C",X"58",X"3A",X"3B",X"40",X"CB",X"3F",X"32",X"3B",X"40",X"3A",X"5C",X"58",X"FE",X"58",
		X"28",X"04",X"FE",X"98",X"20",X"08",X"3A",X"4C",X"40",X"ED",X"44",X"32",X"4C",X"40",X"C9",X"3A",
		X"4D",X"40",X"FE",X"01",X"20",X"1C",X"CD",X"FA",X"09",X"30",X"12",X"3A",X"4D",X"40",X"3C",X"32",
		X"4D",X"40",X"AF",X"32",X"4B",X"40",X"32",X"51",X"40",X"32",X"50",X"40",X"C9",X"AF",X"32",X"4D",
		X"40",X"C9",X"FE",X"02",X"20",X"55",X"3A",X"4B",X"40",X"3C",X"32",X"4B",X"40",X"FE",X"0A",X"C0",
		X"AF",X"32",X"4B",X"40",X"3A",X"5C",X"58",X"47",X"3A",X"50",X"40",X"32",X"5C",X"58",X"78",X"32",
		X"50",X"40",X"3A",X"51",X"40",X"3C",X"32",X"51",X"40",X"FE",X"08",X"C0",X"3E",X"03",X"32",X"4D",
		X"40",X"AF",X"32",X"51",X"40",X"3A",X"4E",X"40",X"C6",X"02",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"CB",X"27",X"32",X"5C",X"58",X"3A",X"4F",X"40",X"C6",X"02",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"CB",X"27",X"32",X"5F",X"58",X"3E",X"39",X"32",X"5D",X"58",X"C9",X"FE",X"03",X"20",X"77",X"3A",
		X"4B",X"40",X"3C",X"32",X"4B",X"40",X"FE",X"0A",X"C0",X"AF",X"32",X"4B",X"40",X"3A",X"5C",X"58",
		X"47",X"3A",X"50",X"40",X"32",X"5C",X"58",X"78",X"32",X"50",X"40",X"3A",X"4E",X"40",X"3C",X"CB",
		X"27",X"47",X"3A",X"4F",X"40",X"3C",X"3C",X"CB",X"27",X"4F",X"3A",X"5C",X"58",X"B7",X"20",X"07",
		X"3E",X"06",X"CD",X"04",X"0E",X"18",X"05",X"3E",X"01",X"CD",X"04",X"0E",X"3A",X"51",X"40",X"3C",
		X"32",X"51",X"40",X"FE",X"08",X"C0",X"3E",X"04",X"32",X"4D",X"40",X"AF",X"32",X"4B",X"40",X"32",
		X"51",X"40",X"32",X"4C",X"40",X"32",X"52",X"40",X"AF",X"21",X"9E",X"1E",X"CD",X"70",X"1C",X"3A",
		X"4E",X"40",X"47",X"3A",X"4F",X"40",X"4F",X"CD",X"6F",X"05",X"3E",X"01",X"DD",X"77",X"00",X"CD",
		X"E4",X"14",X"CD",X"79",X"0A",X"C9",X"3A",X"4B",X"40",X"3C",X"E6",X"3F",X"32",X"4B",X"40",X"3A",
		X"52",X"40",X"B7",X"20",X"16",X"3A",X"4B",X"40",X"B7",X"20",X"4B",X"3A",X"51",X"40",X"3C",X"32",
		X"51",X"40",X"FE",X"0A",X"20",X"40",X"3E",X"01",X"32",X"52",X"40",X"CD",X"7C",X"09",X"30",X"36",
		X"AF",X"32",X"52",X"40",X"32",X"4D",X"40",X"3A",X"4E",X"40",X"3C",X"CB",X"27",X"47",X"3A",X"4F",
		X"40",X"3C",X"3C",X"CB",X"27",X"4F",X"3E",X"06",X"CD",X"04",X"0E",X"3A",X"4E",X"40",X"47",X"3A",
		X"4F",X"40",X"4F",X"CD",X"6F",X"05",X"3E",X"06",X"DD",X"77",X"00",X"CD",X"7B",X"10",X"AF",X"21",
		X"9C",X"1C",X"CD",X"70",X"1C",X"C9",X"CD",X"E3",X"09",X"38",X"6B",X"3A",X"4B",X"40",X"E6",X"01",
		X"C8",X"3A",X"4B",X"40",X"E6",X"10",X"28",X"04",X"3E",X"39",X"18",X"02",X"3E",X"3A",X"32",X"5D",
		X"58",X"3A",X"4C",X"40",X"CB",X"57",X"C2",X"35",X"0A",X"CB",X"5F",X"C2",X"46",X"0A",X"CB",X"47",
		X"C2",X"57",X"0A",X"CB",X"4F",X"C2",X"68",X"0A",X"CD",X"79",X"0A",X"C9",X"3A",X"5C",X"58",X"E6",
		X"0F",X"20",X"2E",X"3A",X"5F",X"58",X"E6",X"0F",X"20",X"27",X"3A",X"5C",X"58",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"D6",X"02",X"32",X"4E",X"40",X"4F",X"3A",X"5F",X"58",X"D6",X"20",
		X"81",X"06",X"00",X"4F",X"DD",X"21",X"5C",X"40",X"DD",X"09",X"DD",X"7E",X"00",X"FE",X"01",X"28",
		X"03",X"37",X"3F",X"C9",X"37",X"C9",X"AF",X"32",X"4D",X"40",X"3A",X"3B",X"40",X"47",X"3A",X"3A",
		X"40",X"B0",X"32",X"3A",X"40",X"CD",X"DC",X"13",X"CD",X"7B",X"10",X"3E",X"50",X"CD",X"BC",X"0D",
		X"CD",X"7D",X"0D",X"AF",X"21",X"9C",X"1C",X"CD",X"70",X"1C",X"3E",X"01",X"21",X"6D",X"1F",X"CD",
		X"70",X"1C",X"C9",X"3A",X"40",X"58",X"4F",X"3A",X"5C",X"58",X"CD",X"7F",X"07",X"30",X"0A",X"3A",
		X"43",X"58",X"4F",X"3A",X"5F",X"58",X"CD",X"7F",X"07",X"C9",X"AF",X"32",X"4F",X"40",X"0E",X"0D",
		X"DD",X"21",X"5C",X"40",X"AF",X"32",X"4E",X"40",X"06",X"0C",X"DD",X"7E",X"00",X"FE",X"06",X"28",
		X"22",X"DD",X"23",X"3A",X"4E",X"40",X"3C",X"32",X"4E",X"40",X"10",X"EE",X"DD",X"23",X"DD",X"23",
		X"DD",X"23",X"DD",X"23",X"3A",X"4F",X"40",X"3C",X"32",X"4F",X"40",X"0D",X"79",X"B7",X"20",X"D4",
		X"37",X"3F",X"C9",X"37",X"C9",X"3A",X"5C",X"58",X"3D",X"32",X"5C",X"58",X"E6",X"0F",X"20",X"03",
		X"CD",X"79",X"0A",X"C3",X"7B",X"09",X"3A",X"5C",X"58",X"3C",X"32",X"5C",X"58",X"E6",X"0F",X"20",
		X"03",X"CD",X"79",X"0A",X"C3",X"7B",X"09",X"3A",X"5F",X"58",X"3D",X"32",X"5F",X"58",X"E6",X"0F",
		X"20",X"03",X"CD",X"79",X"0A",X"C3",X"7B",X"09",X"3A",X"5F",X"58",X"3C",X"32",X"5F",X"58",X"E6",
		X"0F",X"20",X"03",X"CD",X"79",X"0A",X"C3",X"7B",X"09",X"06",X"10",X"AF",X"DD",X"21",X"2F",X"41",
		X"DD",X"77",X"00",X"DD",X"23",X"10",X"F5",X"3A",X"5C",X"58",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"D6",X"02",X"32",X"4E",X"40",X"47",X"3A",X"5F",X"58",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"D6",X"02",X"32",X"4F",X"40",X"4F",X"CD",X"9B",X"0B",X"DD",X"21",X"2F",X"41",
		X"1E",X"00",X"3A",X"2E",X"41",X"CB",X"57",X"28",X"07",X"DD",X"36",X"00",X"04",X"DD",X"23",X"1C",
		X"CB",X"5F",X"28",X"07",X"DD",X"36",X"00",X"08",X"DD",X"23",X"1C",X"CB",X"47",X"28",X"07",X"DD",
		X"36",X"00",X"01",X"DD",X"23",X"1C",X"CB",X"4F",X"28",X"07",X"DD",X"36",X"00",X"02",X"DD",X"23",
		X"1C",X"3A",X"4C",X"40",X"B7",X"28",X"19",X"47",X"3A",X"2E",X"41",X"A0",X"28",X"12",X"DD",X"77",
		X"00",X"DD",X"23",X"1C",X"DD",X"77",X"00",X"DD",X"23",X"1C",X"DD",X"77",X"00",X"DD",X"23",X"1C",
		X"3A",X"40",X"58",X"47",X"3A",X"5C",X"58",X"B8",X"38",X"1E",X"3A",X"2E",X"41",X"CB",X"5F",X"28",
		X"33",X"DD",X"36",X"00",X"08",X"DD",X"23",X"1C",X"DD",X"36",X"00",X"08",X"DD",X"23",X"1C",X"DD",
		X"36",X"00",X"08",X"DD",X"23",X"1C",X"18",X"1C",X"3A",X"2E",X"41",X"CB",X"57",X"28",X"15",X"DD",
		X"36",X"00",X"04",X"DD",X"23",X"1C",X"DD",X"36",X"00",X"04",X"DD",X"23",X"1C",X"DD",X"36",X"00",
		X"04",X"DD",X"23",X"1C",X"3A",X"43",X"58",X"47",X"3A",X"5F",X"58",X"B8",X"38",X"1E",X"3A",X"2E",
		X"41",X"CB",X"4F",X"28",X"33",X"DD",X"36",X"00",X"02",X"DD",X"23",X"1C",X"DD",X"36",X"00",X"02",
		X"DD",X"23",X"1C",X"DD",X"36",X"00",X"02",X"DD",X"23",X"1C",X"18",X"1C",X"3A",X"2E",X"41",X"CB",
		X"47",X"28",X"15",X"DD",X"36",X"00",X"01",X"DD",X"23",X"1C",X"DD",X"36",X"00",X"01",X"DD",X"23",
		X"1C",X"DD",X"36",X"00",X"01",X"DD",X"23",X"1C",X"CD",X"ED",X"14",X"DD",X"21",X"2F",X"41",X"4F",
		X"06",X"00",X"DD",X"09",X"DD",X"7E",X"00",X"32",X"4C",X"40",X"C9",X"AF",X"32",X"2E",X"41",X"C5",
		X"D1",X"79",X"FE",X"00",X"28",X"0F",X"0D",X"CD",X"F8",X"0B",X"30",X"09",X"06",X"01",X"3A",X"2E",
		X"41",X"B0",X"32",X"2E",X"41",X"D5",X"C1",X"79",X"FE",X"0C",X"28",X"0F",X"0C",X"CD",X"F8",X"0B",
		X"30",X"09",X"06",X"02",X"3A",X"2E",X"41",X"B0",X"32",X"2E",X"41",X"D5",X"C1",X"78",X"FE",X"00",
		X"28",X"0F",X"05",X"CD",X"F8",X"0B",X"30",X"09",X"06",X"04",X"3A",X"2E",X"41",X"B0",X"32",X"2E",
		X"41",X"D5",X"C1",X"78",X"FE",X"0B",X"28",X"0F",X"04",X"CD",X"F8",X"0B",X"30",X"09",X"06",X"08",
		X"3A",X"2E",X"41",X"B0",X"32",X"2E",X"41",X"C9",X"CD",X"6F",X"05",X"DD",X"7E",X"00",X"FE",X"01",
		X"28",X"17",X"FE",X"09",X"28",X"13",X"FE",X"0A",X"28",X"0F",X"FE",X"08",X"28",X"0B",X"FE",X"0B",
		X"28",X"07",X"FE",X"0C",X"28",X"03",X"37",X"3F",X"C9",X"37",X"C9",X"AF",X"32",X"50",X"58",X"32",
		X"54",X"58",X"32",X"58",X"58",X"3E",X"00",X"21",X"5A",X"1E",X"CD",X"70",X"1C",X"3A",X"4D",X"40",
		X"B7",X"28",X"07",X"AF",X"32",X"5C",X"58",X"32",X"4D",X"40",X"06",X"04",X"0E",X"24",X"79",X"32",
		X"41",X"58",X"3E",X"1C",X"CD",X"D5",X"0C",X"0C",X"10",X"F4",X"AF",X"32",X"40",X"58",X"3E",X"1E",
		X"CD",X"D5",X"0C",X"3A",X"45",X"40",X"B7",X"C2",X"2F",X"11",X"3A",X"37",X"40",X"3D",X"32",X"37",
		X"40",X"CD",X"B1",X"02",X"CD",X"87",X"13",X"3A",X"37",X"40",X"B7",X"CA",X"57",X"1B",X"CD",X"F1",
		X"02",X"C3",X"84",X"01",X"06",X"0A",X"3A",X"40",X"58",X"32",X"50",X"40",X"78",X"E6",X"01",X"28",
		X"0B",X"3A",X"50",X"40",X"32",X"40",X"58",X"CD",X"A1",X"0C",X"18",X"07",X"AF",X"32",X"40",X"58",
		X"CD",X"BD",X"0C",X"3E",X"0F",X"CD",X"D5",X"0C",X"10",X"E2",X"3A",X"50",X"40",X"32",X"40",X"58",
		X"C9",X"C5",X"3A",X"30",X"40",X"B7",X"28",X"09",X"01",X"00",X"18",X"DD",X"21",X"CB",X"14",X"18",
		X"07",X"01",X"00",X"01",X"DD",X"21",X"C7",X"14",X"CD",X"0D",X"0D",X"C1",X"C9",X"C5",X"3A",X"30",
		X"40",X"B7",X"28",X"05",X"01",X"00",X"18",X"18",X"03",X"01",X"00",X"01",X"DD",X"21",X"CF",X"14",
		X"CD",X"0D",X"0D",X"C1",X"C9",X"C5",X"47",X"AF",X"32",X"35",X"40",X"3A",X"00",X"78",X"3A",X"35",
		X"40",X"B8",X"38",X"F7",X"C1",X"C9",X"21",X"00",X"50",X"06",X"04",X"3E",X"10",X"77",X"2C",X"20",
		X"FC",X"24",X"10",X"F7",X"C9",X"21",X"00",X"50",X"06",X"04",X"7D",X"E6",X"1F",X"28",X"07",X"FE",
		X"01",X"28",X"03",X"3E",X"10",X"77",X"2C",X"20",X"F1",X"24",X"10",X"EE",X"C9",X"21",X"A0",X"53",
		X"11",X"E0",X"FF",X"78",X"FE",X"00",X"28",X"03",X"19",X"10",X"FD",X"09",X"DD",X"7E",X"00",X"B7",
		X"C8",X"FE",X"20",X"20",X"04",X"3E",X"10",X"18",X"0E",X"FE",X"30",X"38",X"08",X"FE",X"39",X"30",
		X"04",X"D6",X"30",X"18",X"02",X"D6",X"30",X"77",X"19",X"DD",X"23",X"18",X"DF",X"C5",X"F5",X"21",
		X"A0",X"53",X"11",X"E0",X"FF",X"78",X"FE",X"00",X"28",X"03",X"19",X"10",X"FD",X"09",X"F1",X"FE",
		X"20",X"20",X"04",X"3E",X"10",X"18",X"0E",X"FE",X"30",X"38",X"08",X"FE",X"39",X"30",X"04",X"D6",
		X"30",X"18",X"02",X"D6",X"30",X"77",X"C1",X"C9",X"C5",X"F5",X"21",X"A0",X"53",X"11",X"E0",X"FF",
		X"78",X"FE",X"00",X"28",X"03",X"19",X"10",X"FD",X"09",X"F1",X"77",X"C1",X"C9",X"01",X"01",X"00",
		X"3A",X"30",X"40",X"B7",X"28",X"03",X"01",X"01",X"16",X"3A",X"3F",X"40",X"CD",X"DE",X"0D",X"04",
		X"04",X"3A",X"3E",X"40",X"CD",X"DE",X"0D",X"04",X"04",X"3A",X"3D",X"40",X"CD",X"DE",X"0D",X"C9",
		X"3A",X"06",X"40",X"01",X"01",X"0B",X"CD",X"DE",X"0D",X"01",X"01",X"0D",X"3A",X"05",X"40",X"CD",
		X"DE",X"0D",X"01",X"01",X"0F",X"3A",X"04",X"40",X"CD",X"DE",X"0D",X"C9",X"F5",X"C5",X"37",X"3F",
		X"47",X"3A",X"3D",X"40",X"80",X"27",X"32",X"3D",X"40",X"3A",X"3E",X"40",X"CE",X"00",X"27",X"32",
		X"3E",X"40",X"3A",X"3F",X"40",X"CE",X"00",X"27",X"32",X"3F",X"40",X"C1",X"F1",X"C9",X"C5",X"F5",
		X"21",X"A0",X"53",X"11",X"E0",X"FF",X"78",X"FE",X"00",X"28",X"03",X"19",X"10",X"FD",X"09",X"F1",
		X"F5",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"77",X"11",X"E0",X"FF",X"19",X"F1",X"E6",
		X"0F",X"77",X"C1",X"C9",X"F5",X"21",X"A0",X"53",X"11",X"E0",X"FF",X"78",X"FE",X"00",X"28",X"03",
		X"19",X"10",X"FD",X"09",X"F1",X"DD",X"21",X"3C",X"0E",X"CB",X"27",X"CB",X"27",X"4F",X"06",X"00",
		X"DD",X"09",X"DD",X"7E",X"00",X"77",X"23",X"DD",X"23",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",
		X"DD",X"7E",X"00",X"77",X"2B",X"DD",X"23",X"DD",X"7E",X"00",X"77",X"C9",X"10",X"10",X"10",X"10",
		X"2E",X"2F",X"2D",X"2C",X"A0",X"A3",X"A0",X"A3",X"36",X"37",X"35",X"34",X"3A",X"3B",X"39",X"38",
		X"3E",X"3F",X"3D",X"3C",X"42",X"43",X"41",X"40",X"46",X"47",X"45",X"44",X"4A",X"4B",X"49",X"48",
		X"4E",X"2F",X"2D",X"4C",X"2E",X"4F",X"4D",X"2C",X"6A",X"2F",X"2D",X"68",X"2E",X"6B",X"69",X"2C",
		X"6E",X"6F",X"6D",X"6C",X"72",X"73",X"71",X"70",X"72",X"73",X"71",X"70",X"52",X"53",X"51",X"50",
		X"56",X"57",X"55",X"54",X"5A",X"5B",X"59",X"58",X"BA",X"BB",X"B9",X"B8",X"BE",X"BF",X"BD",X"BC",
		X"C2",X"C3",X"D5",X"C0",X"C6",X"C7",X"C5",X"C4",X"CA",X"CB",X"C9",X"C8",X"CE",X"CF",X"CD",X"CC",
		X"D2",X"D3",X"D1",X"D0",X"D6",X"D7",X"D5",X"D4",X"DA",X"DB",X"D9",X"D8",X"DE",X"DF",X"DD",X"DC",
		X"32",X"33",X"31",X"30",X"FA",X"FB",X"F9",X"F8",X"21",X"B8",X"23",X"B7",X"28",X"07",X"47",X"11",
		X"52",X"00",X"19",X"10",X"FD",X"7E",X"32",X"53",X"40",X"23",X"7E",X"32",X"54",X"40",X"23",X"7E",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"C6",X"20",X"32",X"40",X"40",X"23",X"7E",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"C6",X"20",X"32",X"41",X"40",X"23",X"06",X"0D",X"11",
		X"5C",X"40",X"C5",X"06",X"06",X"7E",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"12",X"13",
		X"7E",X"E6",X"0F",X"12",X"13",X"23",X"10",X"ED",X"C1",X"13",X"13",X"13",X"13",X"10",X"E3",X"06",
		X"1A",X"AF",X"11",X"09",X"58",X"12",X"13",X"13",X"10",X"FB",X"11",X"10",X"00",X"DD",X"21",X"5C",
		X"40",X"FD",X"21",X"09",X"58",X"06",X"0D",X"DD",X"7E",X"00",X"FE",X"07",X"20",X"12",X"3E",X"05",
		X"FD",X"77",X"00",X"FD",X"23",X"FD",X"23",X"FD",X"77",X"00",X"FD",X"23",X"FD",X"23",X"18",X"08",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"DD",X"19",X"10",X"DB",X"AF",X"32",X"44",X"40",
		X"06",X"D0",X"DD",X"21",X"5C",X"40",X"DD",X"7E",X"00",X"FE",X"0F",X"CC",X"76",X"0F",X"FE",X"03",
		X"28",X"08",X"FE",X"04",X"28",X"04",X"FE",X"05",X"20",X"07",X"3A",X"44",X"40",X"3C",X"32",X"44",
		X"40",X"DD",X"23",X"10",X"E1",X"C9",X"3E",X"D0",X"90",X"4F",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"C6",X"04",X"32",X"48",X"40",X"79",X"E6",X"0F",X"CB",X"27",X"C6",X"02",X"32",X"47",
		X"40",X"AF",X"C9",X"3A",X"34",X"40",X"B7",X"28",X"08",X"47",X"C5",X"CD",X"A2",X"0F",X"C1",X"10",
		X"F9",X"C9",X"3A",X"54",X"40",X"B7",X"28",X"06",X"3D",X"32",X"54",X"40",X"18",X"05",X"3E",X"07",
		X"32",X"53",X"40",X"C9",X"DD",X"21",X"5C",X"40",X"01",X"04",X"02",X"DD",X"7E",X"00",X"C5",X"DD",
		X"E5",X"CD",X"04",X"0E",X"DD",X"E1",X"C1",X"DD",X"23",X"04",X"04",X"78",X"FE",X"1A",X"20",X"EB",
		X"06",X"02",X"0C",X"0C",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"79",X"FE",X"1E",X"20",
		X"DA",X"C9",X"3E",X"94",X"32",X"41",X"58",X"3E",X"01",X"32",X"42",X"58",X"3A",X"45",X"40",X"B7",
		X"28",X"05",X"CD",X"98",X"10",X"18",X"03",X"CD",X"7B",X"10",X"3A",X"53",X"40",X"E6",X"01",X"28",
		X"19",X"3E",X"10",X"32",X"44",X"58",X"3E",X"1D",X"32",X"45",X"58",X"3E",X"01",X"32",X"46",X"58",
		X"3E",X"20",X"32",X"47",X"58",X"3E",X"01",X"32",X"56",X"40",X"3A",X"53",X"40",X"E6",X"02",X"28",
		X"19",X"3E",X"E0",X"32",X"48",X"58",X"3E",X"9D",X"32",X"49",X"58",X"3E",X"01",X"32",X"4A",X"58",
		X"3E",X"E0",X"32",X"4B",X"58",X"3E",X"FF",X"32",X"58",X"40",X"3A",X"53",X"40",X"E6",X"04",X"28",
		X"19",X"3E",X"D0",X"32",X"4C",X"58",X"3E",X"61",X"32",X"4D",X"58",X"3E",X"01",X"32",X"4E",X"58",
		X"3E",X"10",X"32",X"4F",X"58",X"3E",X"FF",X"32",X"5A",X"40",X"AF",X"32",X"50",X"58",X"32",X"54",
		X"58",X"32",X"58",X"58",X"3E",X"02",X"32",X"52",X"58",X"32",X"56",X"58",X"32",X"5A",X"58",X"3E",
		X"23",X"32",X"51",X"58",X"32",X"55",X"58",X"32",X"59",X"58",X"C9",X"3E",X"58",X"32",X"5C",X"58",
		X"3E",X"EF",X"32",X"5F",X"58",X"3E",X"38",X"32",X"5D",X"58",X"3E",X"04",X"32",X"5E",X"58",X"3E",
		X"01",X"32",X"4C",X"40",X"32",X"3B",X"40",X"C9",X"3E",X"90",X"32",X"5C",X"58",X"21",X"B6",X"10",
		X"3A",X"3C",X"40",X"4F",X"06",X"00",X"09",X"7E",X"32",X"5F",X"58",X"3E",X"14",X"32",X"5D",X"58",
		X"3E",X"01",X"32",X"5E",X"58",X"C9",X"B0",X"70",X"30",X"AF",X"32",X"5C",X"58",X"CD",X"94",X"1C",
		X"06",X"04",X"C5",X"AF",X"32",X"3A",X"40",X"CD",X"DC",X"13",X"3E",X"14",X"CD",X"D5",X"0C",X"3E",
		X"1F",X"32",X"3A",X"40",X"CD",X"DC",X"13",X"3E",X"14",X"CD",X"D5",X"0C",X"C1",X"10",X"E3",X"CD",
		X"ED",X"11",X"CD",X"D3",X"11",X"01",X"0B",X"08",X"DD",X"21",X"FB",X"11",X"CD",X"0D",X"0D",X"01",
		X"0E",X"04",X"DD",X"21",X"07",X"12",X"CD",X"0D",X"0D",X"3E",X"04",X"32",X"1D",X"58",X"01",X"12",
		X"09",X"DD",X"21",X"1C",X"12",X"CD",X"0D",X"0D",X"3E",X"C8",X"CD",X"D5",X"0C",X"AF",X"32",X"1D",
		X"58",X"32",X"35",X"40",X"32",X"3A",X"40",X"CD",X"DC",X"13",X"3E",X"01",X"32",X"45",X"40",X"AF",
		X"32",X"46",X"40",X"21",X"90",X"27",X"CD",X"C5",X"0E",X"CD",X"B4",X"0F",X"C3",X"84",X"01",X"CD",
		X"D3",X"11",X"CD",X"ED",X"11",X"01",X"0B",X"05",X"DD",X"21",X"26",X"12",X"CD",X"0D",X"0D",X"3A",
		X"44",X"40",X"B7",X"28",X"1A",X"47",X"AF",X"37",X"3F",X"3C",X"27",X"10",X"FC",X"01",X"0E",X"04",
		X"CD",X"DE",X"0D",X"01",X"0E",X"07",X"DD",X"21",X"38",X"12",X"CD",X"0D",X"0D",X"18",X"21",X"01",
		X"0E",X"04",X"DD",X"21",X"4A",X"12",X"CD",X"0D",X"0D",X"3A",X"3E",X"40",X"37",X"3F",X"C6",X"10",
		X"27",X"32",X"3E",X"40",X"3A",X"3F",X"40",X"CE",X"00",X"27",X"32",X"3F",X"40",X"CD",X"7D",X"0D",
		X"3A",X"46",X"40",X"B7",X"20",X"0C",X"01",X"12",X"07",X"DD",X"21",X"71",X"12",X"CD",X"0D",X"0D",
		X"18",X"0A",X"01",X"12",X"05",X"DD",X"21",X"5E",X"12",X"CD",X"0D",X"0D",X"3E",X"F0",X"CD",X"D5",
		X"0C",X"AF",X"32",X"45",X"40",X"32",X"46",X"40",X"3A",X"3C",X"40",X"FE",X"02",X"28",X"04",X"3C",
		X"32",X"3C",X"40",X"C3",X"49",X"02",X"3A",X"45",X"40",X"B7",X"C8",X"CD",X"E3",X"09",X"D0",X"3E",
		X"01",X"32",X"46",X"40",X"AF",X"32",X"5C",X"58",X"3A",X"37",X"40",X"3C",X"32",X"37",X"40",X"CD",
		X"87",X"13",X"C9",X"01",X"04",X"02",X"AF",X"C5",X"CD",X"04",X"0E",X"C1",X"04",X"04",X"78",X"FE",
		X"1A",X"20",X"F3",X"06",X"02",X"0C",X"0C",X"79",X"FE",X"1E",X"20",X"EA",X"C9",X"AF",X"01",X"1F",
		X"00",X"21",X"40",X"58",X"11",X"41",X"58",X"77",X"ED",X"B0",X"C9",X"42",X"4F",X"4E",X"55",X"53",
		X"20",X"52",X"4F",X"55",X"4E",X"44",X"00",X"45",X"58",X"54",X"52",X"41",X"20",X"4C",X"49",X"46",
		X"45",X"20",X"43",X"48",X"41",X"4C",X"4C",X"45",X"4E",X"47",X"45",X"00",X"47",X"45",X"54",X"20",
		X"52",X"45",X"41",X"44",X"59",X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",X"52",X"4F",X"55",X"4E",
		X"44",X"20",X"53",X"54",X"41",X"54",X"53",X"00",X"43",X"48",X"45",X"52",X"52",X"49",X"45",X"53",
		X"20",X"52",X"45",X"4D",X"41",X"49",X"4E",X"45",X"44",X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",
		X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",X"20",X"31",X"30",X"30",X"30",X"00",X"52",X"45",
		X"43",X"45",X"49",X"56",X"45",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4C",X"49",X"46",X"45",
		X"00",X"4E",X"4F",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4C",X"49",X"46",X"45",X"00",X"3A",
		X"4A",X"40",X"B7",X"28",X"0D",X"FE",X"01",X"28",X"20",X"FE",X"02",X"28",X"2E",X"FE",X"03",X"28",
		X"3E",X"C9",X"3A",X"47",X"40",X"47",X"3A",X"48",X"40",X"4F",X"3E",X"1D",X"CD",X"04",X"0E",X"AF",
		X"32",X"49",X"40",X"3C",X"32",X"4A",X"40",X"18",X"E8",X"3A",X"49",X"40",X"3C",X"32",X"49",X"40",
		X"FE",X"3C",X"20",X"DD",X"3E",X"02",X"32",X"4A",X"40",X"18",X"D6",X"3A",X"47",X"40",X"47",X"3A",
		X"48",X"40",X"4F",X"3E",X"1E",X"CD",X"04",X"0E",X"3E",X"03",X"32",X"4A",X"40",X"18",X"C2",X"3A",
		X"40",X"58",X"E6",X"0F",X"20",X"BB",X"3A",X"43",X"58",X"E6",X"0F",X"20",X"B4",X"CD",X"25",X"05",
		X"7E",X"FE",X"0F",X"20",X"AC",X"AF",X"CD",X"94",X"1C",X"3E",X"3C",X"CD",X"D5",X"0C",X"3E",X"04",
		X"32",X"4A",X"40",X"18",X"9C",X"CD",X"E6",X"0C",X"DD",X"21",X"3F",X"13",X"CD",X"73",X"13",X"01",
		X"00",X"01",X"DD",X"21",X"C7",X"14",X"CD",X"0D",X"0D",X"01",X"00",X"09",X"DD",X"21",X"D3",X"14",
		X"CD",X"0D",X"0D",X"3A",X"2F",X"40",X"B7",X"28",X"16",X"01",X"00",X"18",X"DD",X"21",X"CB",X"14",
		X"CD",X"0D",X"0D",X"3E",X"01",X"32",X"30",X"40",X"CD",X"7D",X"0D",X"AF",X"32",X"30",X"40",X"CD",
		X"7D",X"0D",X"CD",X"A0",X"0D",X"CD",X"DC",X"13",X"CD",X"87",X"13",X"CD",X"5F",X"13",X"C9",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"1E",X"17",X"DD",X"21",X"DE",X"14",X"CD",X"0D",X"0D",X"01",X"1F",X"1A",X"3A",X"32",X"40",X"CD",
		X"DE",X"0D",X"C9",X"C5",X"E5",X"21",X"01",X"58",X"06",X"20",X"DD",X"7E",X"00",X"77",X"23",X"23",
		X"DD",X"23",X"10",X"F6",X"E1",X"C1",X"C9",X"16",X"00",X"D5",X"7A",X"CB",X"27",X"47",X"0E",X"1E",
		X"3A",X"37",X"40",X"B7",X"28",X"08",X"3D",X"BA",X"28",X"04",X"38",X"02",X"18",X"04",X"3E",X"00",
		X"18",X"0F",X"3A",X"38",X"40",X"DD",X"21",X"D8",X"13",X"16",X"00",X"5F",X"DD",X"19",X"DD",X"7E",
		X"00",X"CD",X"04",X"0E",X"D1",X"14",X"7A",X"FE",X"04",X"20",X"CE",X"C9",X"3A",X"39",X"40",X"3C",
		X"32",X"39",X"40",X"FE",X"0F",X"38",X"10",X"AF",X"32",X"39",X"40",X"3A",X"38",X"40",X"3C",X"E6",
		X"03",X"32",X"38",X"40",X"CD",X"87",X"13",X"C9",X"11",X"12",X"11",X"10",X"3A",X"3A",X"40",X"CB",
		X"47",X"20",X"04",X"3E",X"13",X"18",X"02",X"3E",X"18",X"01",X"1E",X"09",X"CD",X"04",X"0E",X"3A",
		X"3A",X"40",X"CB",X"4F",X"20",X"04",X"3E",X"14",X"18",X"02",X"3E",X"19",X"01",X"1E",X"0B",X"CD",
		X"04",X"0E",X"3A",X"3A",X"40",X"CB",X"57",X"20",X"04",X"3E",X"15",X"18",X"02",X"3E",X"1A",X"01",
		X"1E",X"0D",X"CD",X"04",X"0E",X"3A",X"3A",X"40",X"CB",X"5F",X"20",X"04",X"3E",X"16",X"18",X"02",
		X"3E",X"1B",X"01",X"1E",X"0F",X"CD",X"04",X"0E",X"3A",X"3A",X"40",X"CB",X"67",X"20",X"04",X"3E",
		X"17",X"18",X"02",X"3E",X"1C",X"01",X"1E",X"11",X"CD",X"04",X"0E",X"C9",X"00",X"50",X"00",X"49",
		X"56",X"41",X"4E",X"20",X"00",X"30",X"00",X"4D",X"49",X"4B",X"45",X"20",X"00",X"20",X"00",X"4D",
		X"52",X"20",X"44",X"4F",X"00",X"10",X"00",X"4D",X"52",X"20",X"58",X"20",X"00",X"00",X"00",X"48",
		X"45",X"4E",X"43",X"48",X"01",X"28",X"00",X"21",X"3C",X"14",X"11",X"04",X"40",X"ED",X"B0",X"C9",
		X"3A",X"00",X"60",X"E6",X"20",X"FE",X"20",X"20",X"05",X"3E",X"01",X"32",X"2D",X"40",X"3A",X"00",
		X"68",X"E6",X"C0",X"FE",X"C0",X"20",X"05",X"3E",X"01",X"32",X"2C",X"40",X"3A",X"00",X"70",X"E6",
		X"01",X"FE",X"01",X"20",X"05",X"3E",X"01",X"32",X"2E",X"40",X"C9",X"AF",X"DD",X"77",X"00",X"DD",
		X"23",X"DD",X"E5",X"C1",X"3A",X"00",X"78",X"78",X"FE",X"43",X"20",X"EF",X"C9",X"DD",X"21",X"30",
		X"40",X"18",X"E8",X"DD",X"21",X"00",X"40",X"18",X"E2",X"AF",X"01",X"EF",X"00",X"21",X"40",X"40",
		X"11",X"41",X"40",X"77",X"ED",X"B0",X"C9",X"31",X"53",X"54",X"00",X"32",X"4E",X"44",X"00",X"20",
		X"20",X"20",X"00",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"00",X"53",X"43",
		X"45",X"4E",X"45",X"00",X"3A",X"00",X"40",X"E6",X"3F",X"32",X"59",X"43",X"C9",X"DD",X"21",X"0B",
		X"15",X"3A",X"59",X"43",X"06",X"00",X"4F",X"DD",X"09",X"DD",X"7E",X"00",X"47",X"93",X"30",X"FC",
		X"3A",X"59",X"43",X"3C",X"E6",X"3F",X"32",X"59",X"43",X"78",X"C9",X"44",X"41",X"6A",X"B1",X"8D",
		X"5F",X"AF",X"C5",X"CE",X"DB",X"2C",X"13",X"B7",X"39",X"A3",X"4C",X"D2",X"8E",X"B4",X"90",X"17",
		X"8C",X"3E",X"89",X"09",X"5A",X"20",X"C6",X"EF",X"5A",X"A0",X"BC",X"80",X"22",X"0A",X"5B",X"19",
		X"97",X"D6",X"A7",X"74",X"D9",X"C8",X"B3",X"49",X"13",X"CC",X"0C",X"61",X"E9",X"A4",X"DC",X"2E",
		X"49",X"56",X"90",X"84",X"1A",X"9F",X"80",X"00",X"0F",X"D0",X"17",X"00",X"03",X"00",X"00",X"01",
		X"01",X"01",X"01",X"00",X"07",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"06",X"CD",X"E6",X"0C",X"3E",X"00",
		X"32",X"03",X"40",X"AF",X"CD",X"94",X"1C",X"DD",X"21",X"4B",X"15",X"CD",X"73",X"13",X"01",X"00",
		X"09",X"DD",X"21",X"D3",X"14",X"CD",X"0D",X"0D",X"CD",X"A0",X"0D",X"01",X"00",X"01",X"DD",X"21",
		X"C7",X"14",X"CD",X"0D",X"0D",X"AF",X"32",X"30",X"40",X"CD",X"D9",X"02",X"CD",X"7D",X"0D",X"3A",
		X"2F",X"40",X"B7",X"28",X"15",X"01",X"00",X"18",X"DD",X"21",X"CB",X"14",X"CD",X"0D",X"0D",X"3E",
		X"01",X"32",X"30",X"40",X"CD",X"E5",X"02",X"CD",X"7D",X"0D",X"01",X"04",X"08",X"DD",X"21",X"E3",
		X"16",X"DD",X"7E",X"00",X"CD",X"68",X"0D",X"04",X"DD",X"23",X"78",X"FE",X"14",X"20",X"F2",X"06",
		X"08",X"0C",X"79",X"FE",X"08",X"20",X"EA",X"01",X"09",X"0A",X"DD",X"21",X"13",X"17",X"CD",X"0D",
		X"0D",X"01",X"1F",X"00",X"DD",X"21",X"8D",X"16",X"3A",X"2C",X"40",X"B7",X"28",X"04",X"DD",X"21",
		X"95",X"16",X"CD",X"0D",X"0D",X"CD",X"1D",X"17",X"01",X"1D",X"02",X"DD",X"21",X"B6",X"16",X"CD",
		X"0D",X"0D",X"AF",X"32",X"5A",X"43",X"32",X"5B",X"43",X"3A",X"00",X"68",X"CB",X"47",X"28",X"17",
		X"3A",X"2C",X"40",X"B7",X"20",X"0B",X"3A",X"01",X"40",X"B7",X"28",X"2A",X"3D",X"27",X"32",X"01",
		X"40",X"AF",X"32",X"2F",X"40",X"18",X"2C",X"CB",X"4F",X"28",X"1B",X"3A",X"2C",X"40",X"B7",X"20",
		X"0E",X"3A",X"01",X"40",X"FE",X"02",X"38",X"0E",X"3D",X"27",X"3D",X"27",X"32",X"01",X"40",X"3E",
		X"01",X"32",X"2F",X"40",X"18",X"0D",X"3E",X"01",X"CD",X"D5",X"0C",X"CD",X"34",X"17",X"CD",X"72",
		X"17",X"18",X"B6",X"3E",X"01",X"32",X"03",X"40",X"C9",X"50",X"52",X"45",X"53",X"53",X"20",X"31",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"4F",X"4E",
		X"4C",X"59",X"00",X"50",X"52",X"45",X"53",X"53",X"20",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"00",X"43",X"52",X"45",
		X"44",X"49",X"54",X"53",X"00",X"46",X"52",X"45",X"45",X"50",X"4C",X"41",X"59",X"00",X"49",X"4E",
		X"53",X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"00",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"00",X"41",X"20",X"4B",X"52",X"41",X"5A",X"59",X"20",X"49",X"56",
		X"41",X"4E",X"20",X"50",X"52",X"4F",X"44",X"55",X"43",X"54",X"49",X"4F",X"4E",X"00",X"48",X"20",
		X"49",X"20",X"47",X"20",X"48",X"20",X"20",X"53",X"20",X"43",X"20",X"4F",X"20",X"52",X"20",X"45",
		X"20",X"53",X"00",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"10",X"A1",X"A2",X"10",X"A4",
		X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",
		X"B5",X"B6",X"B7",X"EC",X"ED",X"EE",X"EF",X"10",X"10",X"10",X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",
		X"F6",X"F7",X"C1",X"4E",X"49",X"47",X"48",X"54",X"4D",X"41",X"52",X"45",X"00",X"3A",X"2C",X"40",
		X"B7",X"20",X"10",X"3A",X"03",X"40",X"FE",X"00",X"20",X"09",X"3A",X"01",X"40",X"01",X"1F",X"08",
		X"CD",X"DE",X"0D",X"C9",X"3A",X"5A",X"43",X"3C",X"32",X"5A",X"43",X"3A",X"2C",X"40",X"B7",X"3E",
		X"02",X"20",X"1C",X"3A",X"01",X"40",X"B7",X"20",X"16",X"DD",X"21",X"9E",X"16",X"3A",X"5A",X"43",
		X"E6",X"20",X"28",X"04",X"DD",X"21",X"AA",X"16",X"01",X"0B",X"09",X"CD",X"0D",X"0D",X"C9",X"DD",
		X"21",X"59",X"16",X"FE",X"01",X"28",X"04",X"DD",X"21",X"73",X"16",X"01",X"0B",X"02",X"CD",X"0D",
		X"0D",X"C9",X"3A",X"5B",X"43",X"B7",X"CA",X"FC",X"18",X"FE",X"01",X"CA",X"65",X"19",X"FE",X"02",
		X"CA",X"7C",X"19",X"FE",X"03",X"CA",X"CB",X"19",X"FE",X"04",X"CA",X"65",X"19",X"FE",X"05",X"CA",
		X"7C",X"19",X"FE",X"06",X"CA",X"E4",X"19",X"FE",X"07",X"CA",X"65",X"19",X"FE",X"08",X"CA",X"7C",
		X"19",X"FE",X"09",X"CA",X"FD",X"19",X"FE",X"0A",X"CA",X"16",X"1A",X"FE",X"0B",X"CA",X"7C",X"19",
		X"FE",X"0C",X"CA",X"56",X"1A",X"FE",X"0D",X"CA",X"65",X"19",X"FE",X"0E",X"CA",X"7C",X"19",X"FE",
		X"0F",X"CA",X"71",X"1A",X"FE",X"10",X"CA",X"65",X"19",X"FE",X"11",X"CA",X"7E",X"1A",X"FE",X"12",
		X"CA",X"65",X"19",X"FE",X"13",X"CA",X"7E",X"1A",X"FE",X"14",X"CA",X"65",X"19",X"FE",X"15",X"CA",
		X"7E",X"1A",X"FE",X"16",X"CA",X"65",X"19",X"FE",X"17",X"CA",X"91",X"1A",X"FE",X"18",X"CA",X"65",
		X"19",X"FE",X"19",X"CA",X"C1",X"1A",X"FE",X"1A",X"CA",X"99",X"1A",X"FE",X"1B",X"CA",X"65",X"19",
		X"FE",X"1C",X"CA",X"E2",X"1A",X"C9",X"49",X"4E",X"53",X"54",X"52",X"55",X"43",X"54",X"49",X"4F",
		X"4E",X"53",X"00",X"43",X"4F",X"4C",X"4C",X"45",X"43",X"54",X"20",X"43",X"48",X"45",X"52",X"52",
		X"49",X"45",X"53",X"20",X"46",X"4F",X"52",X"20",X"32",X"30",X"20",X"00",X"20",X"43",X"4F",X"4C",
		X"4C",X"45",X"43",X"54",X"20",X"41",X"50",X"50",X"4C",X"45",X"53",X"20",X"46",X"4F",X"52",X"20",
		X"33",X"30",X"20",X"20",X"00",X"20",X"44",X"49",X"41",X"4D",X"4F",X"4E",X"44",X"53",X"20",X"52",
		X"45",X"4C",X"45",X"41",X"53",X"45",X"20",X"4D",X"52",X"20",X"58",X"20",X"20",X"00",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"43",X"41",X"54",X"43",X"48",X"20",X"4D",X"52",X"20",X"58",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"41",X"56",X"4F",
		X"49",X"44",X"20",X"44",X"45",X"41",X"54",X"48",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"0D",X"0D",X"0D",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"03",X"01",X"04",X"01",X"05",X"01",X"06",X"01",X"06",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"0E",X"0E",X"0E",X"01",X"0E",X"02",X"DD",X"21",X"90",X"18",X"DD",X"E5",X"C5",X"CD",
		X"0D",X"0D",X"C1",X"DD",X"E1",X"0C",X"79",X"FE",X"1C",X"20",X"F1",X"C9",X"3E",X"01",X"32",X"5B",
		X"43",X"DD",X"21",X"4B",X"15",X"CD",X"73",X"13",X"CD",X"E5",X"18",X"DD",X"21",X"06",X"18",X"01",
		X"0E",X"08",X"CD",X"0D",X"0D",X"01",X"12",X"02",X"DD",X"21",X"A9",X"18",X"C5",X"DD",X"E5",X"DD",
		X"7E",X"00",X"CD",X"04",X"0E",X"DD",X"E1",X"C1",X"DD",X"23",X"04",X"04",X"78",X"FE",X"1A",X"20",
		X"EB",X"06",X"02",X"0C",X"0C",X"79",X"FE",X"1C",X"20",X"E2",X"DD",X"21",X"13",X"18",X"01",X"10",
		X"02",X"CD",X"0D",X"0D",X"3E",X"20",X"32",X"40",X"58",X"3E",X"B0",X"32",X"43",X"58",X"3E",X"01",
		X"32",X"42",X"58",X"3E",X"94",X"32",X"41",X"58",X"3E",X"20",X"32",X"5C",X"43",X"3E",X"3C",X"32",
		X"5D",X"43",X"C3",X"05",X"18",X"3A",X"5D",X"43",X"B7",X"28",X"07",X"3D",X"32",X"5D",X"43",X"C3",
		X"05",X"18",X"3A",X"5B",X"43",X"3C",X"32",X"5B",X"43",X"C3",X"05",X"18",X"3A",X"5C",X"43",X"B7",
		X"28",X"23",X"3D",X"32",X"5C",X"43",X"3A",X"40",X"58",X"3C",X"32",X"40",X"58",X"E6",X"0F",X"DD",
		X"21",X"CC",X"03",X"4F",X"06",X"00",X"DD",X"09",X"DD",X"7E",X"00",X"4F",X"3E",X"94",X"81",X"32",
		X"41",X"58",X"C3",X"05",X"18",X"3A",X"5B",X"43",X"3C",X"32",X"5B",X"43",X"C3",X"05",X"18",X"3A",
		X"40",X"58",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"D6",X"02",X"47",X"3A",X"43",X"58",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"4F",X"3E",X"01",X"CD",X"04",X"0E",X"C9",X"CD",X"AF",X"19",X"DD",X"21",
		X"2C",X"18",X"01",X"10",X"02",X"CD",X"0D",X"0D",X"3E",X"20",X"32",X"5C",X"43",X"3E",X"78",X"32",
		X"5D",X"43",X"18",X"C1",X"CD",X"AF",X"19",X"DD",X"21",X"45",X"18",X"01",X"10",X"02",X"CD",X"0D",
		X"0D",X"3E",X"20",X"32",X"5C",X"43",X"3E",X"78",X"32",X"5D",X"43",X"18",X"A8",X"CD",X"AF",X"19",
		X"DD",X"21",X"5E",X"18",X"01",X"10",X"02",X"CD",X"0D",X"0D",X"3E",X"18",X"32",X"5C",X"43",X"3E",
		X"20",X"32",X"5D",X"43",X"18",X"8F",X"3A",X"5A",X"43",X"E6",X"08",X"28",X"0F",X"3E",X"06",X"01",
		X"16",X"12",X"CD",X"04",X"0E",X"AF",X"32",X"5C",X"58",X"C3",X"05",X"18",X"3E",X"01",X"01",X"16",
		X"12",X"CD",X"04",X"0E",X"3E",X"A0",X"32",X"5C",X"58",X"3E",X"B0",X"32",X"5F",X"58",X"3E",X"39",
		X"32",X"5D",X"58",X"3E",X"04",X"32",X"5E",X"58",X"3A",X"5D",X"43",X"B7",X"CA",X"A5",X"19",X"3D",
		X"32",X"5D",X"43",X"C3",X"05",X"18",X"AF",X"32",X"5C",X"58",X"DD",X"21",X"77",X"18",X"01",X"10",
		X"02",X"CD",X"0D",X"0D",X"3E",X"18",X"32",X"5C",X"43",X"3E",X"3C",X"32",X"5D",X"43",X"C3",X"A5",
		X"19",X"3E",X"24",X"32",X"41",X"58",X"3E",X"1E",X"32",X"5D",X"43",X"C3",X"A5",X"19",X"3A",X"41",
		X"58",X"FE",X"27",X"28",X"04",X"3C",X"32",X"41",X"58",X"3E",X"1E",X"32",X"5D",X"43",X"C3",X"A5",
		X"19",X"3E",X"78",X"32",X"5D",X"43",X"C3",X"A5",X"19",X"3E",X"FF",X"32",X"5D",X"43",X"C3",X"A5",
		X"19",X"00",X"03",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"07",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"02",X"00",
		X"06",X"AF",X"32",X"40",X"58",X"DD",X"21",X"A1",X"1A",X"CD",X"73",X"13",X"CD",X"E5",X"18",X"DD",
		X"21",X"CE",X"16",X"01",X"0E",X"04",X"CD",X"0D",X"0D",X"01",X"11",X"06",X"CD",X"E9",X"1A",X"C3",
		X"A5",X"19",X"AF",X"32",X"5B",X"43",X"C3",X"05",X"18",X"DD",X"21",X"04",X"40",X"16",X"01",X"D5",
		X"7A",X"CD",X"68",X"0D",X"DD",X"23",X"DD",X"23",X"DD",X"7E",X"00",X"04",X"04",X"04",X"CD",X"DE",
		X"0D",X"DD",X"2B",X"DD",X"7E",X"00",X"04",X"04",X"CD",X"DE",X"0D",X"DD",X"2B",X"DD",X"7E",X"00",
		X"04",X"04",X"CD",X"DE",X"0D",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"04",X"04",X"04",X"04",X"DD",
		X"7E",X"00",X"CD",X"3D",X"0D",X"DD",X"23",X"04",X"DD",X"7E",X"00",X"CD",X"3D",X"0D",X"DD",X"23",
		X"04",X"DD",X"7E",X"00",X"CD",X"3D",X"0D",X"DD",X"23",X"04",X"DD",X"7E",X"00",X"CD",X"3D",X"0D",
		X"DD",X"23",X"04",X"DD",X"7E",X"00",X"CD",X"3D",X"0D",X"DD",X"23",X"0C",X"0C",X"06",X"06",X"D1",
		X"14",X"7A",X"FE",X"06",X"20",X"99",X"C9",X"3A",X"31",X"40",X"3C",X"32",X"31",X"40",X"AF",X"01",
		X"1F",X"00",X"21",X"40",X"58",X"11",X"41",X"58",X"77",X"ED",X"B0",X"3E",X"00",X"21",X"79",X"1E",
		X"CD",X"70",X"1C",X"01",X"0E",X"05",X"DD",X"21",X"E7",X"1B",X"CD",X"0D",X"0D",X"01",X"0F",X"05",
		X"DD",X"21",X"E7",X"1B",X"CD",X"0D",X"0D",X"01",X"10",X"05",X"DD",X"21",X"E7",X"1B",X"CD",X"0D",
		X"0D",X"DD",X"21",X"D6",X"1B",X"01",X"0F",X"06",X"DD",X"7E",X"00",X"B7",X"28",X"13",X"DD",X"E5",
		X"C5",X"CD",X"3D",X"0D",X"3E",X"0F",X"CD",X"D5",X"0C",X"C1",X"DD",X"E1",X"DD",X"23",X"04",X"18",
		X"E7",X"3E",X"3C",X"CD",X"D5",X"0C",X"CD",X"8A",X"1F",X"3A",X"2F",X"40",X"B7",X"28",X"14",X"3A",
		X"31",X"40",X"FE",X"01",X"20",X"0D",X"CD",X"F1",X"02",X"DD",X"21",X"3F",X"13",X"CD",X"73",X"13",
		X"C3",X"84",X"01",X"C3",X"50",X"01",X"47",X"20",X"41",X"20",X"4D",X"20",X"45",X"20",X"20",X"4F",
		X"20",X"56",X"20",X"45",X"20",X"52",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"DD",X"21",X"5E",X"43",X"CD",
		X"21",X"1C",X"B7",X"20",X"02",X"06",X"FF",X"3A",X"65",X"43",X"B7",X"28",X"07",X"DD",X"21",X"65",
		X"43",X"CD",X"21",X"1C",X"3A",X"6C",X"43",X"B8",X"C8",X"78",X"32",X"00",X"78",X"32",X"6C",X"43",
		X"C9",X"DD",X"7E",X"00",X"B7",X"28",X"40",X"DD",X"7E",X"05",X"B7",X"28",X"06",X"3D",X"DD",X"77",
		X"05",X"18",X"39",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"7E",X"DD",X"77",X"06",X"23",X"7E",X"23",
		X"DD",X"74",X"03",X"DD",X"75",X"04",X"B7",X"28",X"05",X"DD",X"77",X"05",X"18",X"1E",X"DD",X"7E",
		X"00",X"FE",X"FF",X"28",X"04",X"3D",X"DD",X"77",X"00",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"DD",
		X"74",X"03",X"DD",X"75",X"04",X"18",X"BA",X"3E",X"FF",X"DD",X"77",X"06",X"DD",X"46",X"06",X"C9",
		X"CD",X"89",X"1C",X"7E",X"DD",X"77",X"00",X"23",X"DD",X"74",X"01",X"DD",X"75",X"02",X"DD",X"74",
		X"03",X"DD",X"75",X"04",X"AF",X"DD",X"77",X"05",X"C9",X"DD",X"21",X"5E",X"43",X"B7",X"C8",X"DD",
		X"21",X"65",X"43",X"C9",X"CD",X"89",X"1C",X"AF",X"DD",X"77",X"00",X"C9",X"FF",X"8E",X"18",X"70",
		X"12",X"40",X"06",X"55",X"06",X"70",X"06",X"FF",X"06",X"70",X"18",X"55",X"06",X"40",X"06",X"FF",
		X"06",X"70",X"06",X"FF",X"06",X"70",X"06",X"FF",X"06",X"A0",X"0C",X"8E",X"12",X"80",X"18",X"40",
		X"06",X"8E",X"18",X"70",X"12",X"40",X"06",X"55",X"06",X"70",X"06",X"FF",X"06",X"70",X"18",X"55",
		X"06",X"40",X"06",X"FF",X"06",X"70",X"06",X"FF",X"06",X"96",X"06",X"8E",X"06",X"80",X"06",X"70",
		X"30",X"FF",X"06",X"8E",X"18",X"70",X"12",X"40",X"06",X"55",X"06",X"70",X"06",X"FF",X"06",X"70",
		X"18",X"55",X"06",X"40",X"06",X"FF",X"06",X"70",X"06",X"FF",X"06",X"70",X"06",X"FF",X"06",X"A0",
		X"0C",X"8E",X"12",X"80",X"18",X"40",X"06",X"8E",X"18",X"70",X"12",X"40",X"06",X"55",X"06",X"70",
		X"06",X"FF",X"06",X"70",X"18",X"55",X"06",X"40",X"06",X"FF",X"06",X"70",X"06",X"FF",X"06",X"96",
		X"06",X"8E",X"06",X"80",X"06",X"70",X"30",X"FF",X"06",X"8E",X"12",X"70",X"12",X"40",X"0C",X"8E",
		X"12",X"70",X"18",X"8A",X"06",X"70",X"06",X"40",X"06",X"FF",X"06",X"8A",X"12",X"80",X"18",X"FF",
		X"18",X"8E",X"12",X"70",X"12",X"40",X"0C",X"8E",X"12",X"70",X"18",X"8A",X"06",X"70",X"06",X"40",
		X"0C",X"A0",X"18",X"FF",X"30",X"8E",X"18",X"70",X"12",X"40",X"06",X"55",X"06",X"70",X"06",X"FF",
		X"06",X"70",X"18",X"55",X"06",X"8E",X"06",X"70",X"06",X"40",X"0C",X"55",X"12",X"70",X"18",X"FF",
		X"18",X"55",X"06",X"A0",X"0C",X"AA",X"0C",X"A0",X"0C",X"AA",X"0C",X"A0",X"12",X"40",X"06",X"96",
		X"06",X"8E",X"06",X"80",X"0C",X"70",X"18",X"FF",X"48",X"00",X"00",X"FF",X"9A",X"06",X"80",X"06",
		X"68",X"06",X"9A",X"06",X"80",X"06",X"68",X"06",X"9A",X"06",X"80",X"06",X"68",X"06",X"9A",X"06",
		X"80",X"06",X"68",X"06",X"9A",X"06",X"68",X"06",X"80",X"06",X"9A",X"06",X"A0",X"06",X"80",X"06",
		X"68",X"06",X"A0",X"06",X"80",X"06",X"68",X"06",X"80",X"06",X"A0",X"06",X"8E",X"06",X"78",X"06",
		X"55",X"06",X"8E",X"06",X"78",X"06",X"55",X"06",X"78",X"06",X"8E",X"06",X"9A",X"06",X"80",X"06",
		X"68",X"06",X"9A",X"06",X"80",X"06",X"68",X"06",X"9A",X"06",X"80",X"06",X"68",X"06",X"9A",X"06",
		X"80",X"06",X"68",X"06",X"9A",X"06",X"68",X"06",X"80",X"06",X"9A",X"06",X"A0",X"06",X"80",X"06",
		X"68",X"06",X"A0",X"06",X"80",X"06",X"68",X"06",X"80",X"06",X"A0",X"06",X"8E",X"06",X"78",X"06",
		X"55",X"06",X"8E",X"06",X"78",X"06",X"55",X"06",X"78",X"06",X"8E",X"06",X"B4",X"06",X"B4",X"06",
		X"B4",X"06",X"B4",X"06",X"B4",X"0C",X"B4",X"06",X"C0",X"0C",X"C0",X"06",X"BC",X"0C",X"B4",X"0C",
		X"AA",X"0C",X"B4",X"06",X"B4",X"06",X"B4",X"06",X"B4",X"06",X"B4",X"0C",X"B4",X"06",X"C0",X"0C",
		X"C0",X"06",X"BC",X"0C",X"B4",X"0C",X"AA",X"0C",X"B4",X"06",X"B4",X"06",X"B4",X"06",X"B4",X"06",
		X"B4",X"0C",X"B4",X"06",X"C0",X"0C",X"C0",X"06",X"BC",X"0C",X"B4",X"0C",X"AA",X"0C",X"B4",X"0C",
		X"CD",X"0C",X"C7",X"0C",X"C0",X"06",X"C7",X"30",X"00",X"00",X"01",X"FF",X"02",X"8E",X"08",X"80",
		X"08",X"70",X"08",X"FF",X"08",X"80",X"08",X"70",X"08",X"68",X"08",X"FF",X"08",X"70",X"08",X"68",
		X"08",X"55",X"08",X"FF",X"08",X"40",X"10",X"00",X"00",X"01",X"40",X"10",X"80",X"08",X"80",X"08",
		X"68",X"10",X"40",X"10",X"40",X"10",X"80",X"08",X"80",X"08",X"68",X"10",X"40",X"10",X"40",X"10",
		X"80",X"08",X"80",X"08",X"80",X"20",X"FF",X"08",X"02",X"10",X"40",X"18",X"00",X"00",X"FF",X"40",
		X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",
		X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",
		X"05",X"8E",X"05",X"40",X"05",X"70",X"05",X"40",X"05",X"8E",X"05",X"40",X"05",X"70",X"05",X"40",
		X"05",X"8E",X"05",X"40",X"05",X"70",X"05",X"40",X"05",X"8E",X"05",X"40",X"05",X"70",X"05",X"40",
		X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",
		X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",X"05",X"80",X"05",X"40",X"05",X"68",X"05",X"40",
		X"05",X"70",X"05",X"40",X"05",X"55",X"05",X"40",X"05",X"70",X"05",X"40",X"05",X"55",X"05",X"40",
		X"05",X"70",X"05",X"40",X"05",X"55",X"05",X"40",X"05",X"70",X"05",X"40",X"05",X"55",X"05",X"00",
		X"00",X"FF",X"40",X"06",X"FF",X"06",X"A0",X"04",X"FF",X"08",X"68",X"06",X"FF",X"06",X"A0",X"04",
		X"FF",X"08",X"70",X"06",X"FF",X"06",X"A0",X"04",X"FF",X"08",X"70",X"06",X"68",X"06",X"70",X"06",
		X"FF",X"06",X"55",X"06",X"FF",X"06",X"9A",X"04",X"FF",X"08",X"55",X"06",X"FF",X"06",X"9A",X"04",
		X"FF",X"08",X"68",X"06",X"FF",X"06",X"9A",X"04",X"FF",X"08",X"55",X"06",X"68",X"06",X"55",X"06",
		X"FF",X"06",X"00",X"00",X"01",X"12",X"01",X"18",X"01",X"22",X"01",X"00",X"00",X"01",X"FF",X"04",
		X"40",X"04",X"55",X"04",X"68",X"04",X"70",X"04",X"80",X"08",X"FF",X"04",X"00",X"00",X"06",X"03",
		X"1A",X"BE",X"D8",X"C0",X"1B",X"2B",X"10",X"F8",X"37",X"C9",X"11",X"3F",X"40",X"21",X"26",X"40",
		X"CD",X"7E",X"1F",X"D8",X"01",X"00",X"04",X"21",X"06",X"40",X"11",X"3F",X"40",X"E5",X"D5",X"C5",
		X"CD",X"7E",X"1F",X"C1",X"D1",X"E1",X"30",X"09",X"D5",X"11",X"08",X"00",X"19",X"D1",X"0C",X"10",
		X"EC",X"2B",X"2B",X"E5",X"79",X"32",X"6D",X"43",X"78",X"B7",X"28",X"10",X"AF",X"C6",X"08",X"10",
		X"FC",X"4F",X"06",X"00",X"21",X"23",X"40",X"11",X"2B",X"40",X"ED",X"B8",X"D1",X"21",X"3D",X"40",
		X"01",X"03",X"00",X"ED",X"B0",X"D5",X"E1",X"3E",X"20",X"12",X"13",X"01",X"04",X"00",X"ED",X"B0",
		X"CD",X"F5",X"0C",X"DD",X"21",X"EC",X"22",X"CD",X"73",X"13",X"CD",X"A0",X"0D",X"01",X"06",X"06",
		X"CD",X"E9",X"1A",X"DD",X"21",X"0C",X"23",X"01",X"04",X"06",X"CD",X"0D",X"0D",X"DD",X"21",X"1C",
		X"23",X"01",X"13",X"06",X"CD",X"0D",X"0D",X"DD",X"21",X"2C",X"23",X"01",X"15",X"05",X"CD",X"0D",
		X"0D",X"DD",X"21",X"3E",X"23",X"01",X"17",X"05",X"CD",X"0D",X"0D",X"DD",X"21",X"50",X"23",X"01",
		X"19",X"06",X"CD",X"0D",X"0D",X"DD",X"21",X"60",X"23",X"01",X"1B",X"05",X"CD",X"0D",X"0D",X"3A",
		X"6D",X"43",X"CB",X"27",X"C6",X"06",X"CB",X"27",X"16",X"00",X"5F",X"21",X"01",X"58",X"19",X"3E",
		X"04",X"77",X"3E",X"35",X"32",X"5C",X"58",X"3E",X"A3",X"32",X"5F",X"58",X"3E",X"3F",X"32",X"5D",
		X"58",X"3E",X"04",X"32",X"5E",X"58",X"AF",X"32",X"4E",X"40",X"32",X"4F",X"40",X"32",X"6E",X"43",
		X"32",X"70",X"43",X"21",X"21",X"1F",X"CD",X"70",X"1C",X"3A",X"6D",X"43",X"B7",X"28",X"06",X"47",
		X"AF",X"C6",X"08",X"10",X"FC",X"C6",X"03",X"F5",X"3A",X"6E",X"43",X"47",X"F1",X"80",X"4F",X"06",
		X"00",X"DD",X"21",X"04",X"40",X"DD",X"09",X"AF",X"32",X"42",X"40",X"AF",X"32",X"71",X"43",X"3A",
		X"42",X"40",X"B7",X"20",X"03",X"CD",X"74",X"02",X"CB",X"47",X"C2",X"E3",X"20",X"CB",X"4F",X"C2",
		X"37",X"21",X"CB",X"57",X"C2",X"9B",X"21",X"CB",X"5F",X"C2",X"C4",X"21",X"CB",X"67",X"C2",X"0B",
		X"22",X"CD",X"C7",X"22",X"06",X"0A",X"AF",X"32",X"42",X"40",X"3E",X"01",X"CD",X"D5",X"0C",X"3A",
		X"71",X"43",X"B7",X"20",X"09",X"CD",X"74",X"02",X"B7",X"28",X"03",X"32",X"42",X"40",X"10",X"EA",
		X"3A",X"70",X"43",X"3C",X"32",X"70",X"43",X"FE",X"F0",X"20",X"B0",X"AF",X"32",X"5C",X"58",X"CD",
		X"94",X"1C",X"C9",X"3E",X"01",X"32",X"71",X"43",X"3A",X"5F",X"58",X"FE",X"A3",X"28",X"24",X"D6",
		X"10",X"32",X"5F",X"58",X"3A",X"4F",X"40",X"3D",X"32",X"4F",X"40",X"FE",X"02",X"20",X"0E",X"3A",
		X"4E",X"40",X"4F",X"06",X"00",X"21",X"B5",X"23",X"09",X"7E",X"32",X"4E",X"40",X"CD",X"EF",X"21",
		X"C3",X"B1",X"20",X"3E",X"D3",X"32",X"5F",X"58",X"3E",X"03",X"32",X"4F",X"40",X"3A",X"4E",X"40",
		X"06",X"00",X"4F",X"21",X"AC",X"23",X"09",X"7E",X"32",X"4E",X"40",X"4F",X"21",X"A9",X"23",X"09",
		X"7E",X"32",X"5C",X"58",X"C3",X"B1",X"20",X"3E",X"01",X"32",X"71",X"43",X"3A",X"5F",X"58",X"FE",
		X"D3",X"28",X"35",X"C6",X"10",X"32",X"5F",X"58",X"3A",X"4F",X"40",X"3C",X"32",X"4F",X"40",X"FE",
		X"02",X"20",X"0D",X"3A",X"4E",X"40",X"FE",X"08",X"20",X"18",X"3D",X"32",X"4E",X"40",X"18",X"12",
		X"FE",X"03",X"20",X"0E",X"3A",X"4E",X"40",X"06",X"00",X"4F",X"21",X"AC",X"23",X"09",X"7E",X"32",
		X"4E",X"40",X"CD",X"EF",X"21",X"C3",X"B1",X"20",X"3E",X"A3",X"32",X"5F",X"58",X"AF",X"32",X"4F",
		X"40",X"3A",X"4E",X"40",X"06",X"00",X"4F",X"21",X"B5",X"23",X"09",X"7E",X"32",X"4E",X"40",X"4F",
		X"21",X"79",X"23",X"09",X"7E",X"32",X"5C",X"58",X"C3",X"B1",X"20",X"3E",X"01",X"32",X"71",X"43",
		X"3A",X"4E",X"40",X"B7",X"28",X"0A",X"3D",X"32",X"4E",X"40",X"CD",X"EF",X"21",X"C3",X"B1",X"20",
		X"3A",X"4F",X"40",X"4F",X"06",X"00",X"21",X"72",X"23",X"09",X"7E",X"32",X"4E",X"40",X"CD",X"EF",
		X"21",X"C3",X"B1",X"20",X"3E",X"01",X"32",X"71",X"43",X"3A",X"4F",X"40",X"4F",X"06",X"00",X"21",
		X"72",X"23",X"09",X"7E",X"47",X"3A",X"4E",X"40",X"B8",X"28",X"0A",X"3C",X"32",X"4E",X"40",X"CD",
		X"EF",X"21",X"C3",X"B1",X"20",X"AF",X"32",X"4E",X"40",X"CD",X"EF",X"21",X"C3",X"B1",X"20",X"3A",
		X"4F",X"40",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"06",X"00",X"4F",X"21",X"79",X"23",
		X"09",X"3A",X"4E",X"40",X"4F",X"09",X"7E",X"32",X"5C",X"58",X"C9",X"3A",X"00",X"78",X"CD",X"74",
		X"02",X"CB",X"67",X"20",X"F6",X"3E",X"01",X"21",X"64",X"1F",X"DD",X"E5",X"CD",X"70",X"1C",X"DD",
		X"E1",X"3A",X"4F",X"40",X"FE",X"03",X"28",X"5C",X"4F",X"06",X"00",X"21",X"76",X"23",X"09",X"7E",
		X"4F",X"3A",X"4E",X"40",X"81",X"CD",X"3E",X"22",X"CD",X"55",X"22",X"C3",X"B1",X"20",X"F5",X"3A",
		X"6D",X"43",X"CB",X"27",X"C6",X"06",X"4F",X"3A",X"6E",X"43",X"C6",X"11",X"47",X"F1",X"DD",X"77",
		X"00",X"CD",X"3D",X"0D",X"C9",X"3A",X"6E",X"43",X"FE",X"04",X"28",X"10",X"AF",X"32",X"6F",X"43",
		X"CD",X"C7",X"22",X"3A",X"6E",X"43",X"3C",X"32",X"6E",X"43",X"DD",X"23",X"C9",X"3A",X"6E",X"43",
		X"B7",X"28",X"F9",X"AF",X"32",X"6F",X"43",X"CD",X"C7",X"22",X"3A",X"6E",X"43",X"3D",X"32",X"6E",
		X"43",X"DD",X"2B",X"C9",X"3A",X"4E",X"40",X"FE",X"00",X"20",X"0B",X"3E",X"20",X"CD",X"3E",X"22",
		X"CD",X"55",X"22",X"C3",X"B1",X"20",X"FE",X"01",X"20",X"19",X"3A",X"6E",X"43",X"FE",X"04",X"20",
		X"07",X"DD",X"7E",X"00",X"FE",X"20",X"20",X"03",X"CD",X"6D",X"22",X"3E",X"20",X"CD",X"3E",X"22",
		X"C3",X"B1",X"20",X"AF",X"32",X"6F",X"43",X"CD",X"C7",X"22",X"AF",X"32",X"5C",X"58",X"CD",X"94",
		X"1C",X"3E",X"A0",X"CD",X"D5",X"0C",X"C9",X"3A",X"6F",X"43",X"3C",X"E6",X"01",X"32",X"6F",X"43",
		X"20",X"04",X"3E",X"5B",X"18",X"02",X"3E",X"20",X"F5",X"3A",X"6D",X"43",X"CB",X"27",X"C6",X"07",
		X"4F",X"3A",X"6E",X"43",X"C6",X"11",X"47",X"F1",X"CD",X"3D",X"0D",X"C9",X"00",X"03",X"00",X"00",
		X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"4F",X"4E",X"47",
		X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"00",X"45",X"4E",X"54",X"45",
		X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"4E",X"41",X"4D",X"45",X"00",X"41",X"20",X"42",X"20",
		X"43",X"20",X"44",X"20",X"45",X"20",X"46",X"20",X"47",X"20",X"48",X"20",X"49",X"00",X"4A",X"20",
		X"4B",X"20",X"4C",X"20",X"4D",X"20",X"4E",X"20",X"4F",X"20",X"50",X"20",X"51",X"20",X"52",X"00",
		X"53",X"20",X"54",X"20",X"55",X"20",X"56",X"20",X"57",X"20",X"58",X"20",X"59",X"20",X"5A",X"00",
		X"53",X"50",X"41",X"43",X"45",X"20",X"20",X"45",X"52",X"41",X"53",X"45",X"20",X"20",X"45",X"4E",
		X"44",X"00",X"08",X"08",X"07",X"02",X"41",X"4A",X"53",X"35",X"45",X"55",X"65",X"75",X"85",X"95",
		X"A5",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"45",X"55",X"65",X"75",X"85",X"95",
		X"A5",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"4D",X"5D",X"6D",X"7D",X"8D",X"9D",
		X"AD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"45",X"7D",X"AD",X"00",X"00",X"00",X"01",
		X"01",X"01",X"01",X"02",X"02",X"00",X"04",X"07",X"05",X"02",X"05",X"07",X"DE",X"11",X"11",X"11",
		X"11",X"ED",X"11",X"11",X"11",X"11",X"11",X"11",X"13",X"31",X"13",X"31",X"13",X"31",X"13",X"31",
		X"13",X"31",X"13",X"31",X"13",X"31",X"63",X"36",X"13",X"31",X"13",X"31",X"13",X"31",X"13",X"31",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"AC",X"CA",X"AA",X"AA",
		X"AC",X"CA",X"78",X"87",X"77",X"77",X"78",X"87",X"9B",X"B9",X"99",X"99",X"9B",X"B9",X"11",X"11",
		X"11",X"11",X"11",X"11",X"EF",X"11",X"51",X"15",X"11",X"FD",X"07",X"02",X"00",X"0C",X"11",X"31",
		X"11",X"11",X"31",X"11",X"F1",X"11",X"13",X"11",X"11",X"11",X"DD",X"DD",X"DD",X"DD",X"DD",X"11",
		X"61",X"11",X"11",X"11",X"41",X"11",X"11",X"11",X"14",X"11",X"11",X"11",X"11",X"41",X"11",X"11",
		X"11",X"15",X"11",X"EE",X"EE",X"EE",X"EE",X"EE",X"11",X"41",X"11",X"11",X"11",X"15",X"11",X"11",
		X"14",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"41",X"11",X"DD",X"DD",X"DD",X"DD",X"DD",X"11",
		X"11",X"11",X"13",X"11",X"11",X"11",X"11",X"31",X"11",X"11",X"31",X"16",X"07",X"01",X"00",X"07",
		X"00",X"DD",X"12",X"11",X"DD",X"00",X"0D",X"11",X"11",X"11",X"11",X"D0",X"D1",X"11",X"12",X"11",
		X"16",X"1D",X"D1",X"11",X"42",X"31",X"11",X"1D",X"11",X"14",X"12",X"13",X"11",X"11",X"11",X"41",
		X"42",X"31",X"31",X"11",X"21",X"22",X"22",X"22",X"22",X"12",X"11",X"13",X"13",X"25",X"14",X"11",
		X"11",X"11",X"31",X"21",X"41",X"11",X"E1",X"11",X"13",X"24",X"11",X"1E",X"E1",X"11",X"11",X"21",
		X"11",X"1E",X"0E",X"11",X"11",X"11",X"11",X"F0",X"00",X"EE",X"11",X"21",X"EE",X"00",X"07",X"01",
		X"03",X"09",X"51",X"40",X"00",X"00",X"01",X"15",X"11",X"14",X"00",X"00",X"11",X"11",X"11",X"11",
		X"40",X"01",X"11",X"14",X"01",X"11",X"11",X"11",X"11",X"40",X"00",X"11",X"11",X"11",X"14",X"00",
		X"00",X"01",X"16",X"61",X"10",X"00",X"00",X"01",X"1E",X"F1",X"10",X"00",X"00",X"01",X"16",X"61",
		X"10",X"00",X"00",X"11",X"11",X"11",X"14",X"00",X"01",X"11",X"11",X"11",X"11",X"40",X"11",X"11",
		X"40",X"01",X"11",X"14",X"11",X"14",X"00",X"00",X"11",X"11",X"51",X"40",X"00",X"00",X"01",X"15",
		X"07",X"01",X"05",X"04",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"14",X"61",X"11",X"11",
		X"11",X"11",X"41",X"14",X"11",X"11",X"11",X"14",X"11",X"11",X"41",X"11",X"11",X"41",X"11",X"11",
		X"14",X"11",X"16",X"11",X"1D",X"E1",X"11",X"41",X"14",X"11",X"1F",X"D1",X"11",X"61",X"11",X"41",
		X"11",X"11",X"14",X"11",X"11",X"14",X"11",X"11",X"41",X"11",X"11",X"11",X"41",X"14",X"11",X"11",
		X"11",X"11",X"16",X"41",X"11",X"11",X"15",X"11",X"11",X"11",X"11",X"51",X"11",X"11",X"11",X"11",
		X"11",X"11",X"06",X"01",X"00",X"0C",X"11",X"12",X"44",X"61",X"21",X"11",X"12",X"12",X"44",X"11",
		X"21",X"21",X"12",X"11",X"11",X"11",X"11",X"21",X"12",X"22",X"11",X"33",X"22",X"21",X"11",X"12",
		X"11",X"33",X"21",X"11",X"11",X"12",X"11",X"11",X"21",X"11",X"12",X"22",X"11",X"D1",X"22",X"21",
		X"12",X"11",X"11",X"D1",X"11",X"21",X"12",X"1D",X"EF",X"EE",X"D1",X"21",X"12",X"11",X"D1",X"11",
		X"11",X"21",X"12",X"21",X"D1",X"33",X"12",X"21",X"11",X"21",X"11",X"33",X"12",X"51",X"11",X"21",
		X"11",X"33",X"12",X"55",X"07",X"01",X"01",X"0C",X"DD",X"11",X"21",X"33",X"21",X"33",X"D1",X"11",
		X"11",X"13",X"21",X"13",X"11",X"11",X"21",X"11",X"21",X"11",X"AC",X"AA",X"2C",X"AA",X"2C",X"AA",
		X"78",X"77",X"78",X"77",X"78",X"77",X"9B",X"99",X"2B",X"99",X"2B",X"99",X"51",X"11",X"26",X"11",
		X"21",X"11",X"AA",X"CA",X"2A",X"1A",X"2A",X"CA",X"77",X"87",X"77",X"87",X"77",X"87",X"99",X"B9",
		X"29",X"B9",X"29",X"B9",X"11",X"11",X"21",X"11",X"21",X"11",X"11",X"1F",X"23",X"11",X"11",X"13",
		X"11",X"EE",X"23",X"31",X"21",X"33",X"06",X"00",X"01",X"01",X"01",X"11",X"13",X"10",X"00",X"00",
		X"11",X"13",X"11",X"13",X"00",X"00",X"11",X"FD",X"ED",X"E1",X"00",X"00",X"01",X"11",X"C1",X"10",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"B1",X"11",X"60",X"00",X"00",X"3E",
		X"DE",X"D1",X"11",X"00",X"00",X"11",X"31",X"31",X"11",X"00",X"00",X"01",X"11",X"C1",X"10",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"B1",X"11",X"10",X"00",X"00",X"5E",X"DE",
		X"D1",X"11",X"00",X"00",X"13",X"13",X"13",X"16",X"07",X"01",X"05",X"04",X"00",X"11",X"11",X"11",
		X"11",X"00",X"01",X"3D",X"F1",X"1D",X"E3",X"10",X"13",X"DE",X"31",X"1E",X"DE",X"31",X"1D",X"E3",
		X"11",X"11",X"3D",X"E1",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"12",X"22",X"22",X"21",X"D1",
		X"1D",X"11",X"31",X"13",X"11",X"D1",X"4D",X"1D",X"DD",X"DD",X"D1",X"D4",X"1D",X"11",X"16",X"61",
		X"11",X"D1",X"4D",X"1E",X"EE",X"EE",X"E1",X"D4",X"1D",X"11",X"31",X"13",X"11",X"D1",X"1D",X"12",
		X"22",X"22",X"21",X"D1",X"11",X"11",X"15",X"51",X"11",X"11",X"07",X"01",X"05",X"08",X"11",X"11",
		X"11",X"11",X"11",X"15",X"1D",X"DD",X"D1",X"1E",X"EE",X"F1",X"1D",X"33",X"31",X"13",X"33",X"E1",
		X"1D",X"32",X"21",X"12",X"23",X"E1",X"1D",X"12",X"41",X"61",X"21",X"E1",X"AA",X"CA",X"AA",X"AA",
		X"AC",X"AA",X"77",X"87",X"77",X"77",X"78",X"77",X"99",X"B9",X"99",X"99",X"9B",X"99",X"1E",X"12",
		X"11",X"14",X"21",X"D1",X"1E",X"32",X"21",X"12",X"23",X"D1",X"1E",X"33",X"31",X"13",X"33",X"D1",
		X"1E",X"EE",X"E1",X"1D",X"DD",X"D1",X"51",X"11",X"11",X"11",X"11",X"11",X"07",X"01",X"02",X"0C",
		X"00",X"25",X"11",X"11",X"12",X"00",X"02",X"55",X"11",X"11",X"11",X"20",X"22",X"22",X"22",X"22",
		X"21",X"22",X"24",X"44",X"11",X"21",X"44",X"42",X"24",X"14",X"21",X"21",X"41",X"42",X"24",X"44",
		X"21",X"21",X"44",X"42",X"21",X"11",X"21",X"11",X"11",X"12",X"22",X"21",X"22",X"22",X"22",X"22",
		X"E1",X"E1",X"11",X"11",X"1E",X"1F",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"77",X"77",X"77",X"77",
		X"77",X"87",X"99",X"99",X"99",X"99",X"99",X"B9",X"11",X"16",X"16",X"16",X"11",X"11",X"07",X"01",
		X"02",X"06",X"EE",X"11",X"11",X"D1",X"11",X"11",X"F1",X"11",X"11",X"D1",X"11",X"11",X"11",X"11",
		X"D1",X"D1",X"11",X"61",X"11",X"11",X"D1",X"D1",X"11",X"11",X"DD",X"D1",X"D1",X"D1",X"61",X"11",
		X"11",X"11",X"D1",X"D1",X"11",X"11",X"11",X"11",X"D1",X"D1",X"11",X"61",X"11",X"11",X"D1",X"D1",
		X"11",X"11",X"1D",X"DD",X"D1",X"D1",X"61",X"11",X"11",X"11",X"D1",X"D1",X"11",X"11",X"15",X"55",
		X"D1",X"D1",X"11",X"61",X"11",X"55",X"D1",X"11",X"11",X"11",X"11",X"11",X"D1",X"11",X"11",X"11",
		X"07",X"00",X"00",X"0C",X"33",X"33",X"33",X"33",X"33",X"3F",X"30",X"00",X"00",X"01",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"10",X"00",X"00",X"03",X"33",X"33",X"33",X"33",
		X"33",X"33",X"30",X"00",X"00",X"01",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",
		X"10",X"00",X"00",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"00",X"00",X"01",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"10",X"00",X"00",X"03",X"13",X"33",X"33",X"33",
		X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
