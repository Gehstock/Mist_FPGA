library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity egs7 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of egs7 is
	type rom is array(0 to  1023) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"05",X"28",X"10",X"10",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"0E",X"00",X"00",X"00",X"00",X"40",X"00",X"FE",X"0F",X"40",X"00",X"F0",X"A1",X"08",X"43",
		X"84",X"FF",X"82",X"3F",X"C2",X"0F",X"FC",X"03",X"F9",X"01",X"62",X"00",X"FE",X"07",X"02",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0E",X"E0",X"0F",X"30",X"0C",X"20",X"4F",
		X"F8",X"3F",X"24",X"49",X"4A",X"95",X"52",X"A5",X"A4",X"49",X"18",X"30",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"3E",X"FF",X"7F",X"80",X"7F",X"00",X"1F",X"F8",X"7F",
		X"FC",X"FF",X"54",X"55",X"FE",X"FF",X"FC",X"7F",X"A8",X"2A",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"02",X"F0",X"7F",X"00",X"02",X"85",X"0F",X"C2",X"10",X"FF",X"21",X"FC",X"41",X"F0",X"43",
		X"C0",X"3F",X"80",X"9F",X"00",X"46",X"E0",X"7F",X"02",X"0E",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"C0",X"00",X"70",X"00",X"F0",X"07",X"30",X"0C",X"F2",X"04",X"FC",X"1B",X"92",X"24",X"A9",X"52",
		X"A5",X"4A",X"92",X"25",X"0C",X"18",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",
		X"7C",X"00",X"FE",X"FF",X"FE",X"01",X"F8",X"00",X"FE",X"3F",X"FF",X"7F",X"AA",X"2A",X"FF",X"7F",
		X"FE",X"3F",X"54",X"15",X"06",X"0E",X"00",X"40",X"01",X"80",X"07",X"00",X"00",X"78",X"03",X"D8",
		X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"DF",X"07",X"F4",X"FD",X"05",X"B8",X"DF",
		X"0F",X"F6",X"FD",X"0D",X"BC",X"DF",X"0F",X"F7",X"FD",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"7E",X"9F",X"DF",X"EF",X"37",X"FC",X"7E",X"BF",X"DF",X"EF",X"37",X"FC",X"7E",X"BF",X"DF",
		X"EF",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"DF",X"EF",X"F7",X"FB",X"3D",X"BF",X"DF",
		X"EF",X"F7",X"FB",X"3D",X"BF",X"DF",X"EF",X"F7",X"FB",X"3D",X"04",X"14",X"40",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"30",X"00",X"00",X"E0",X"30",X"46",X"00",
		X"E0",X"20",X"46",X"00",X"F0",X"3D",X"62",X"00",X"F8",X"B3",X"5E",X"00",X"5A",X"BB",X"C6",X"0F",
		X"FE",X"FF",X"EE",X"1F",X"1E",X"FF",X"3F",X"0E",X"4E",X"FE",X"9F",X"1C",X"54",X"FD",X"AF",X"1A",
		X"E0",X"00",X"C0",X"01",X"50",X"01",X"A0",X"02",X"40",X"00",X"80",X"00",X"04",X"07",X"9E",X"E3",
		X"3C",X"1F",X"41",X"14",X"45",X"01",X"41",X"10",X"45",X"01",X"4E",X"10",X"3D",X"0F",X"50",X"10",
		X"15",X"01",X"50",X"14",X"25",X"01",X"8F",X"E3",X"44",X"1F",X"02",X"07",X"44",X"0E",X"44",X"04",
		X"44",X"04",X"7C",X"64",X"44",X"04",X"44",X"04",X"44",X"0E",X"07",X"07",X"E0",X"39",X"D1",X"07",
		X"27",X"FA",X"1E",X"10",X"44",X"5B",X"80",X"28",X"0A",X"22",X"10",X"44",X"55",X"80",X"28",X"0A",
		X"22",X"90",X"7D",X"D5",X"83",X"28",X"7A",X"1E",X"10",X"45",X"51",X"80",X"28",X"0A",X"0A",X"10",
		X"45",X"51",X"80",X"48",X"09",X"12",X"E0",X"45",X"D1",X"07",X"87",X"F8",X"22",X"08",X"07",X"17",
		X"79",X"DF",X"F3",X"C1",X"71",X"2E",X"02",X"12",X"05",X"41",X"44",X"20",X"8A",X"24",X"02",X"32",
		X"05",X"41",X"44",X"20",X"88",X"64",X"02",X"52",X"39",X"CF",X"43",X"20",X"88",X"A4",X"02",X"92",
		X"41",X"41",X"41",X"20",X"88",X"24",X"03",X"12",X"41",X"41",X"42",X"20",X"8A",X"24",X"02",X"17",
		X"3D",X"5F",X"44",X"C0",X"71",X"2E",X"02",X"04",X"14",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"30",X"00",X"00",X"E0",X"30",X"46",X"00",X"E0",X"20",X"46",
		X"00",X"F0",X"3D",X"62",X"00",X"F8",X"B3",X"5E",X"00",X"5A",X"BB",X"C6",X"0F",X"FE",X"FF",X"EE",
		X"1F",X"1E",X"FF",X"3F",X"0E",X"AE",X"FE",X"5F",X"1D",X"44",X"FC",X"8F",X"18",X"F0",X"01",X"E0",
		X"03",X"40",X"00",X"80",X"00",X"A0",X"00",X"40",X"01",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"02",X"C0",X"1F",X"00",X"02",X"82",X"0F",X"C5",X"10",X"FE",X"21",X"FC",X"41",X"F0",X"43",X"C0",
		X"3F",X"80",X"9F",X"00",X"46",X"E0",X"7F",X"02",X"0E",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",
		X"00",X"70",X"00",X"F0",X"07",X"30",X"0C",X"F2",X"04",X"FC",X"1B",X"92",X"24",X"A5",X"4A",X"A9",
		X"52",X"92",X"25",X"0C",X"18",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"7C",
		X"00",X"FE",X"FF",X"FE",X"01",X"F8",X"00",X"FE",X"3F",X"FF",X"7F",X"54",X"15",X"FE",X"3F",X"FF",
		X"7F",X"AA",X"2A",X"02",X"0E",X"00",X"00",X"00",X"00",X"40",X"00",X"F8",X"03",X"40",X"00",X"F0",
		X"41",X"08",X"A3",X"84",X"7F",X"82",X"3F",X"C2",X"0F",X"FC",X"03",X"F9",X"01",X"62",X"00",X"FE",
		X"07",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0E",X"E0",X"0F",X"30",
		X"0C",X"20",X"4F",X"F8",X"3F",X"24",X"49",X"52",X"A5",X"4A",X"95",X"A4",X"49",X"18",X"30",X"02",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"3E",X"FF",X"7F",X"80",X"7F",X"00",
		X"1F",X"F8",X"7F",X"FC",X"FF",X"A8",X"2A",X"FC",X"7F",X"FE",X"FF",X"54",X"55",X"00",X"01",X"0E",
		X"38",X"38",X"44",X"44",X"64",X"64",X"54",X"54",X"4C",X"4C",X"44",X"44",X"38",X"38",X"01",X"01",
		X"0E",X"10",X"10",X"18",X"18",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"38",X"38",X"02",
		X"01",X"0E",X"38",X"38",X"44",X"44",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"7C",X"7C",
		X"03",X"01",X"0E",X"7C",X"7C",X"20",X"20",X"10",X"10",X"20",X"20",X"40",X"40",X"44",X"44",X"38",
		X"38",X"04",X"01",X"0E",X"30",X"30",X"28",X"28",X"24",X"24",X"7C",X"7C",X"20",X"20",X"20",X"20",
		X"20",X"20",X"05",X"01",X"0E",X"7C",X"7C",X"04",X"04",X"3C",X"3C",X"40",X"40",X"40",X"40",X"44",
		X"44",X"38",X"38",X"06",X"01",X"0E",X"30",X"30",X"08",X"08",X"04",X"04",X"3C",X"3C",X"44",X"44",
		X"44",X"44",X"38",X"38",X"07",X"01",X"0E",X"7C",X"7C",X"40",X"40",X"20",X"20",X"10",X"10",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"01",X"0E",X"38",X"38",X"44",X"44",X"44",X"44",X"38",X"38",
		X"44",X"44",X"44",X"44",X"38",X"38",X"09",X"01",X"0E",X"38",X"38",X"44",X"44",X"44",X"44",X"78",
		X"78",X"40",X"40",X"20",X"20",X"18",X"18",X"10",X"01",X"6A",X"1C",X"59",X"1E",X"10",X"1C",X"B3",
		X"1E",X"1C",X"02",X"A6",X"1C",X"95",X"1E",X"4C",X"1C",X"EF",X"1E",X"28",X"03",X"88",X"1C",X"77",
		X"1E",X"2E",X"1C",X"D1",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
