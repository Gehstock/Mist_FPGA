library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"11",X"11",X"11",X"77",X"6F",X"9F",X"00",X"77",X"FF",X"FF",X"CE",X"8F",X"0F",X"CF",
		X"EE",X"CC",X"88",X"00",X"0C",X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"BF",X"3D",X"73",X"77",X"13",X"00",X"00",X"EF",X"EF",X"EF",X"DF",X"BF",X"7F",X"19",X"00",
		X"27",X"3F",X"0C",X"8C",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",X"88",X"00",X"00",
		X"00",X"00",X"11",X"33",X"77",X"77",X"77",X"23",X"66",X"CC",X"CC",X"CC",X"99",X"BB",X"1F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"BF",X"7F",X"7F",X"47",X"21",X"11",X"00",X"CF",X"EF",X"FF",X"EF",X"EF",X"EF",X"DF",X"6F",
		X"77",X"2E",X"0C",X"7F",X"FF",X"FF",X"33",X"00",X"00",X"11",X"FF",X"EE",X"CC",X"88",X"00",X"00",
		X"00",X"11",X"11",X"33",X"33",X"37",X"77",X"77",X"00",X"00",X"00",X"00",X"02",X"BB",X"8F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"08",X"23",X"67",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",
		X"77",X"23",X"23",X"57",X"33",X"13",X"11",X"00",X"0F",X"7F",X"FF",X"FF",X"FF",X"BF",X"97",X"73",
		X"4E",X"1F",X"BF",X"BF",X"FF",X"EE",X"CE",X"8C",X"FF",X"EE",X"EE",X"CC",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"44",X"46",X"66",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"66",X"66",X"06",X"8F",
		X"00",X"00",X"00",X"00",X"66",X"66",X"06",X"1F",X"00",X"00",X"22",X"26",X"66",X"EE",X"EE",X"EE",
		X"77",X"77",X"11",X"00",X"01",X"00",X"00",X"00",X"8F",X"BF",X"7F",X"7F",X"FF",X"6F",X"32",X"00",
		X"1F",X"DF",X"EF",X"EF",X"FF",X"6F",X"C4",X"00",X"EE",X"EE",X"88",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"36",X"6F",X"EB",X"AB",X"EE",X"EE",
		X"00",X"04",X"C6",X"6F",X"7D",X"5D",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"33",X"22",X"33",X"33",X"00",X"00",X"FF",X"FF",X"FF",X"13",X"13",X"11",X"00",X"00",
		X"FF",X"FF",X"7F",X"4C",X"0C",X"08",X"00",X"00",X"44",X"44",X"CC",X"44",X"CC",X"CC",X"00",X"00",
		X"00",X"00",X"11",X"13",X"13",X"13",X"13",X"01",X"22",X"BB",X"F9",X"9F",X"CF",X"C7",X"46",X"EE",
		X"00",X"0C",X"0E",X"86",X"8A",X"EE",X"6F",X"6F",X"00",X"00",X"00",X"00",X"00",X"CC",X"44",X"44",
		X"02",X"00",X"22",X"11",X"11",X"01",X"00",X"00",X"DF",X"6F",X"37",X"1D",X"88",X"CC",X"CC",X"00",
		X"2F",X"AF",X"AE",X"CE",X"4E",X"00",X"00",X"00",X"EE",X"66",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"54",X"67",X"75",X"66",X"33",X"00",X"EE",X"FB",X"5D",X"3F",X"0B",X"8D",X"DF",
		X"00",X"00",X"00",X"99",X"CC",X"EF",X"7F",X"2E",X"00",X"00",X"00",X"00",X"88",X"4C",X"66",X"77",
		X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"EF",X"FF",X"37",X"26",X"8C",X"77",X"33",X"11",
		X"8E",X"4F",X"AF",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"77",X"21",X"ED",X"77",X"00",X"00",X"0C",X"EF",X"D9",X"FF",X"0F",X"0C",
		X"00",X"08",X"22",X"11",X"0D",X"8F",X"4E",X"8F",X"00",X"00",X"00",X"CC",X"EE",X"66",X"00",X"00",
		X"76",X"77",X"11",X"00",X"00",X"00",X"00",X"00",X"DF",X"67",X"FF",X"33",X"66",X"77",X"00",X"00",
		X"EF",X"3F",X"CF",X"08",X"08",X"EE",X"EE",X"22",X"08",X"88",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"77",X"21",X"00",X"00",X"00",X"00",X"0F",X"4B",X"FF",X"0F",
		X"00",X"00",X"FF",X"02",X"0E",X"0E",X"0F",X"0F",X"00",X"00",X"CC",X"4C",X"00",X"00",X"08",X"0C",
		X"30",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"C0",X"FF",X"B3",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"8F",X"EE",X"CE",X"02",X"FF",X"00",X"00",X"CC",X"08",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"37",X"76",X"00",X"00",X"77",X"44",X"13",X"FF",X"67",X"9F",
		X"22",X"EE",X"EE",X"08",X"0C",X"0F",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"08",
		X"7F",X"ED",X"21",X"77",X"33",X"00",X"00",X"00",X"0C",X"1F",X"FF",X"D9",X"FF",X"CC",X"00",X"00",
		X"AF",X"EF",X"CF",X"CD",X"11",X"2A",X"00",X"00",X"00",X"00",X"66",X"EE",X"8C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"33",X"67",X"8C",X"06",X"27",X"CF",X"8F",
		X"00",X"00",X"00",X"00",X"06",X"2F",X"4F",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"66",X"75",X"67",X"54",X"00",X"11",X"00",X"9F",X"8D",X"1B",X"3F",X"5D",X"FB",X"EE",X"00",
		X"6E",X"FF",X"FF",X"CC",X"99",X"00",X"00",X"00",X"77",X"66",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"22",X"00",X"02",X"00",X"CC",X"CC",X"88",X"0D",X"27",X"6F",X"DF",
		X"00",X"00",X"00",X"4E",X"CE",X"CE",X"8E",X"AF",X"00",X"00",X"00",X"00",X"00",X"37",X"26",X"6E",
		X"01",X"11",X"13",X"33",X"11",X"11",X"00",X"00",X"CF",X"46",X"C6",X"CF",X"9F",X"F9",X"BB",X"33",
		X"AF",X"6F",X"EE",X"AA",X"C6",X"CC",X"8C",X"00",X"44",X"44",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"23",X"22",X"23",X"22",X"22",X"00",X"00",X"11",X"13",X"13",X"5F",X"DF",X"FF",
		X"00",X"00",X"08",X"0C",X"4C",X"6F",X"7F",X"7F",X"00",X"00",X"CC",X"4C",X"44",X"4C",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"AB",X"EB",X"EF",X"76",X"22",X"00",
		X"7F",X"7F",X"5D",X"7D",X"7F",X"E6",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"99",X"99",X"19",
		X"00",X"08",X"88",X"88",X"88",X"99",X"99",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"57",X"57",X"57",X"44",X"00",X"00",X"00",X"5F",X"DF",X"DF",X"BF",X"37",X"37",X"01",X"33",
		X"AF",X"BF",X"BF",X"DF",X"CE",X"CE",X"08",X"CC",X"22",X"AE",X"AE",X"AE",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"01",X"04",X"CE",X"CE",X"67",X"67",X"33",X"33",X"BB",
		X"00",X"00",X"00",X"46",X"22",X"03",X"7F",X"BF",X"00",X"00",X"00",X"00",X"44",X"66",X"2E",X"AE",
		X"00",X"44",X"47",X"23",X"23",X"11",X"00",X"00",X"5F",X"DF",X"DF",X"5F",X"19",X"00",X"00",X"00",
		X"BF",X"DF",X"CF",X"EF",X"8E",X"37",X"CC",X"00",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"27",X"33",X"11",X"00",X"00",X"22",X"00",X"00",X"11",X"08",X"8C",X"CE",X"67",X"33",
		X"00",X"00",X"11",X"99",X"27",X"FF",X"3F",X"1F",X"00",X"00",X"00",X"88",X"CC",X"0E",X"88",X"00",
		X"11",X"00",X"02",X"23",X"11",X"00",X"00",X"00",X"57",X"5F",X"EF",X"7F",X"2E",X"8C",X"44",X"00",
		X"CF",X"EF",X"EF",X"4F",X"19",X"22",X"00",X"00",X"08",X"00",X"04",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"7F",X"77",X"01",X"00",X"00",X"00",X"23",X"11",X"08",X"EF",X"FF",
		X"00",X"66",X"33",X"03",X"7F",X"7F",X"0F",X"8F",X"00",X"00",X"88",X"4C",X"08",X"00",X"00",X"08",
		X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"13",X"33",X"BF",X"37",X"03",X"CF",X"77",X"00",
		X"FF",X"FF",X"BF",X"CF",X"88",X"08",X"80",X"88",X"8A",X"2E",X"4C",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"00",X"67",X"00",X"00",X"FF",
		X"00",X"FF",X"07",X"77",X"7F",X"EF",X"8F",X"9F",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"CF",
		X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"77",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EF",X"7F",X"77",X"07",X"FF",X"00",X"DF",X"CD",X"0C",X"00",X"00",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"77",X"8F",X"13",X"37",X"BF",X"23",X"03",
		X"88",X"08",X"08",X"88",X"8F",X"1F",X"7F",X"FF",X"00",X"00",X"00",X"08",X"04",X"4C",X"2E",X"8A",
		X"01",X"77",X"7F",X"06",X"00",X"00",X"00",X"00",X"FF",X"CF",X"08",X"01",X"77",X"44",X"00",X"00",
		X"EF",X"3F",X"FF",X"6F",X"03",X"13",X"66",X"00",X"08",X"00",X"00",X"08",X"0C",X"88",X"00",X"00",
		X"00",X"00",X"00",X"11",X"23",X"00",X"00",X"11",X"00",X"04",X"8C",X"2E",X"7F",X"EF",X"6F",X"57",
		X"00",X"00",X"02",X"19",X"0F",X"6F",X"FF",X"EF",X"00",X"00",X"00",X"00",X"88",X"04",X"00",X"08",
		X"22",X"00",X"00",X"01",X"13",X"37",X"02",X"00",X"33",X"37",X"6E",X"CC",X"88",X"11",X"00",X"00",
		X"DF",X"BF",X"FF",X"27",X"89",X"11",X"00",X"00",X"00",X"88",X"2E",X"4C",X"88",X"00",X"00",X"00",
		X"00",X"00",X"01",X"23",X"23",X"47",X"44",X"00",X"00",X"00",X"00",X"0D",X"CF",X"DF",X"DF",X"7F",
		X"00",X"CC",X"73",X"AC",X"EF",X"EF",X"DF",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",
		X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"33",X"37",X"37",X"6F",X"6E",X"CE",X"04",
		X"BF",X"7F",X"03",X"22",X"46",X"04",X"00",X"00",X"2E",X"2E",X"66",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"57",X"57",X"57",X"44",X"13",X"01",X"37",X"37",X"BF",X"DF",X"DF",X"7F",
		X"8C",X"08",X"CE",X"CE",X"DF",X"BF",X"BF",X"AF",X"00",X"00",X"00",X"02",X"AE",X"AE",X"AE",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"99",X"99",X"11",X"11",X"11",X"11",X"00",
		X"89",X"99",X"99",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"00",X"70",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"70",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"10",X"00",X"30",X"B0",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"30",X"00",X"10",X"00",X"70",X"00",X"00",
		X"D0",X"C0",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"80",X"00",X"20",X"10",X"03",X"12",
		X"00",X"00",X"80",X"40",X"E0",X"E0",X"78",X"1C",X"40",X"20",X"30",X"30",X"A0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"21",X"20",X"20",X"20",X"10",X"00",X"00",
		X"A4",X"08",X"80",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"00",X"E0",X"10",X"03",X"12",
		X"00",X"00",X"80",X"40",X"E0",X"E0",X"78",X"1C",X"40",X"20",X"30",X"30",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"21",X"20",X"20",X"30",X"10",X"00",X"00",
		X"A4",X"08",X"80",X"E0",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"70",X"F0",X"30",X"00",X"C0",X"03",X"12",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"68",X"3C",X"C0",X"60",X"70",X"70",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"21",X"20",X"30",X"30",X"10",X"00",X"00",
		X"A4",X"48",X"E0",X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"70",X"F0",X"30",X"10",X"00",X"D0",X"03",
		X"00",X"00",X"80",X"C0",X"E0",X"60",X"48",X"0C",X"C0",X"E0",X"70",X"70",X"20",X"20",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"30",X"30",X"30",X"30",X"10",X"00",X"00",
		X"94",X"68",X"F0",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"70",X"F0",X"30",X"10",X"00",X"D0",X"03",
		X"10",X"10",X"80",X"80",X"C0",X"C0",X"48",X"0C",X"C0",X"E0",X"F0",X"70",X"30",X"30",X"60",X"C0",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"30",X"30",X"30",X"30",X"10",X"00",X"00",
		X"94",X"78",X"70",X"C0",X"C0",X"80",X"00",X"00",X"80",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"20",X"40",X"40",X"10",X"30",X"10",X"C0",X"E0",X"30",X"10",X"00",X"D0",X"E1",
		X"F0",X"30",X"00",X"00",X"80",X"C0",X"80",X"48",X"00",X"80",X"C0",X"40",X"20",X"20",X"40",X"E0",
		X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"F0",X"B0",X"B0",X"B0",X"30",X"10",X"00",X"00",
		X"58",X"F0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"E0",X"80",X"20",X"20",X"40",X"80",X"00",X"00",
		X"00",X"00",X"10",X"20",X"00",X"40",X"10",X"30",X"30",X"C0",X"00",X"E0",X"10",X"00",X"D0",X"E1",
		X"F0",X"30",X"00",X"00",X"80",X"40",X"C0",X"48",X"00",X"C0",X"E0",X"60",X"30",X"30",X"10",X"10",
		X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"B0",X"B0",X"B0",X"B0",X"D0",X"10",X"00",X"00",
		X"48",X"80",X"C0",X"C0",X"C0",X"80",X"20",X"00",X"10",X"10",X"20",X"20",X"40",X"80",X"00",X"00",
		X"00",X"00",X"10",X"20",X"00",X"40",X"10",X"30",X"30",X"C0",X"00",X"70",X"00",X"10",X"E1",X"D2",
		X"F0",X"30",X"00",X"00",X"80",X"C0",X"48",X"2C",X"00",X"C0",X"E0",X"60",X"30",X"30",X"10",X"10",
		X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"52",X"61",X"70",X"B0",X"B0",X"10",X"00",X"00",
		X"A4",X"48",X"80",X"C0",X"C0",X"80",X"20",X"00",X"10",X"10",X"20",X"20",X"40",X"80",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"C0",X"30",X"00",X"00",X"C0",X"D0",X"D0",X"00",X"E0",X"F0",
		X"70",X"70",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"30",X"30",X"80",X"C0",X"F0",X"F0",X"70",X"80",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",
		X"80",X"C0",X"D0",X"D0",X"B0",X"B0",X"F0",X"70",X"80",X"00",X"C0",X"C0",X"C0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"10",X"00",X"30",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"60",
		X"00",X"00",X"C0",X"F0",X"F0",X"00",X"E0",X"E0",X"10",X"20",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"30",X"30",X"00",X"00",X"80",X"60",X"70",X"70",X"70",X"00",X"00",X"00",X"30",X"30",X"30",X"21",
		X"F0",X"F0",X"00",X"00",X"C0",X"E0",X"E0",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"C0",X"80",
		X"60",X"E0",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"E0",X"90",X"00",X"20",X"20",X"40",X"40",X"80",X"80",X"40",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"10",X"10",X"30",X"F0",X"F0",X"F0",X"78",X"10",X"00",X"80",X"F0",X"E0",X"90",X"10",X"10",
		X"00",X"80",X"40",X"B0",X"00",X"30",X"20",X"60",X"00",X"30",X"C0",X"00",X"00",X"F0",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"C0",X"30",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"E0",X"F0",
		X"70",X"70",X"70",X"30",X"10",X"00",X"30",X"10",X"30",X"30",X"80",X"C0",X"F0",X"F0",X"70",X"40",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",
		X"80",X"C0",X"D0",X"D0",X"B0",X"B0",X"F0",X"70",X"00",X"00",X"C0",X"C0",X"C0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"10",X"00",X"30",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"60",
		X"00",X"00",X"C0",X"F0",X"F0",X"00",X"E0",X"E0",X"10",X"20",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"80",X"40",X"00",X"60",X"70",X"70",X"70",X"00",X"00",X"00",X"30",X"30",X"30",X"21",
		X"F0",X"F0",X"00",X"00",X"C0",X"E0",X"E0",X"00",X"10",X"10",X"10",X"00",X"30",X"10",X"00",X"00",
		X"60",X"E0",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"E0",X"90",X"10",X"20",X"20",X"40",X"40",X"80",X"80",X"40",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"10",X"10",X"30",X"F0",X"F0",X"F0",X"78",X"D0",X"80",X"80",X"C0",X"E0",X"90",X"10",X"10",
		X"00",X"80",X"40",X"30",X"C0",X"30",X"20",X"60",X"00",X"30",X"C0",X"00",X"00",X"F0",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"C0",X"30",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"E0",X"F0",
		X"70",X"70",X"70",X"30",X"50",X"60",X"20",X"00",X"30",X"30",X"80",X"C0",X"F0",X"F0",X"70",X"00",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",
		X"80",X"C0",X"D0",X"D0",X"B0",X"B0",X"F0",X"70",X"00",X"00",X"C0",X"C0",X"C0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"10",X"00",X"30",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"60",
		X"00",X"00",X"C0",X"F0",X"F0",X"00",X"E0",X"E0",X"10",X"20",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"60",X"E0",X"40",X"00",X"60",X"70",X"70",X"70",X"00",X"00",X"00",X"30",X"30",X"30",X"21",
		X"F0",X"F0",X"00",X"00",X"C0",X"E0",X"E0",X"00",X"10",X"10",X"10",X"00",X"00",X"20",X"60",X"40",
		X"60",X"E0",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"E0",X"90",X"10",X"20",X"20",X"40",X"40",X"80",X"80",X"40",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"10",X"10",X"30",X"F0",X"F0",X"F0",X"78",X"10",X"20",X"80",X"C0",X"E0",X"90",X"10",X"10",
		X"00",X"80",X"40",X"30",X"C0",X"30",X"20",X"60",X"00",X"30",X"C0",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"F0",
		X"00",X"00",X"00",X"30",X"78",X"70",X"F0",X"78",X"00",X"00",X"00",X"00",X"04",X"00",X"80",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"D0",X"28",X"70",X"70",X"68",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"10",X"00",X"00",X"01",X"00",X"00",X"12",X"D0",X"E0",X"D0",X"10",X"10",X"00",X"00",
		X"49",X"F0",X"F0",X"F0",X"40",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"20",X"A0",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"30",X"11",X"10",X"00",X"00",X"00",
		X"A0",X"10",X"00",X"A0",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"00",X"20",X"00",X"00",X"70",X"10",X"00",X"00",X"90",
		X"00",X"C0",X"F0",X"10",X"00",X"30",X"31",X"BA",X"00",X"00",X"00",X"00",X"00",X"20",X"90",X"80",
		X"10",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"D8",X"E8",X"CC",X"F1",X"73",X"30",X"00",X"00",
		X"60",X"44",X"00",X"CC",X"C0",X"A0",X"10",X"00",X"00",X"00",X"40",X"C0",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"51",X"40",X"00",X"70",X"72",X"30",X"00",X"00",X"00",X"10",X"30",X"73",X"72",
		X"00",X"00",X"10",X"40",X"74",X"E4",X"C0",X"72",X"80",X"40",X"20",X"20",X"30",X"90",X"10",X"A0",
		X"72",X"31",X"B0",X"11",X"20",X"30",X"00",X"00",X"F6",X"E0",X"40",X"FC",X"F9",X"B1",X"D0",X"10",
		X"75",X"73",X"60",X"C4",X"D9",X"C8",X"D0",X"80",X"20",X"00",X"00",X"C8",X"C8",X"80",X"00",X"00",
		X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"20",X"10",X"00",X"40",X"E4",X"99",
		X"D0",X"20",X"20",X"D0",X"40",X"44",X"44",X"88",X"00",X"00",X"10",X"C0",X"00",X"90",X"80",X"80",
		X"00",X"00",X"40",X"00",X"00",X"30",X"40",X"80",X"F1",X"70",X"73",X"50",X"20",X"00",X"00",X"90",
		X"22",X"E4",X"EC",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"90",X"40",X"00",
		X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"E0",X"80",X"00",X"00",X"50",
		X"00",X"00",X"00",X"80",X"40",X"00",X"10",X"88",X"00",X"00",X"00",X"20",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"73",X"50",X"B0",X"00",X"20",X"11",X"10",X"80",
		X"C0",X"80",X"00",X"22",X"64",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"51",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B3",X"51",X"31",X"30",X"10",X"40",X"00",X"00",
		X"88",X"00",X"44",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"70",X"10",X"00",X"20",X"10",X"20",X"00",X"B0",X"90",X"50",X"40",X"C0",X"E6",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"10",X"50",X"70",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E6",X"F7",X"20",X"00",X"00",X"C0",X"F0",X"E0",X"C0",X"B0",
		X"90",X"FE",X"E4",X"E0",X"E0",X"80",X"10",X"FB",X"80",X"C0",X"70",X"72",X"F7",X"70",X"80",X"80",
		X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"A0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"70",X"72",X"60",X"00",X"00",X"00",X"60",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"30",X"30",X"00",X"22",X"11",X"00",X"00",X"F6",X"FC",X"64",X"00",X"11",X"11",X"32",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"10",X"30",X"73",X"F7",X"F7",X"00",X"30",X"00",X"00",X"E0",X"C8",X"E8",X"88",
		X"EC",X"FE",X"F4",X"E0",X"00",X"80",X"80",X"D8",X"00",X"10",X"10",X"31",X"72",X"20",X"00",X"A0",
		X"00",X"44",X"A8",X"10",X"D0",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"B1",X"10",X"00",X"00",X"00",X"00",X"00",X"40",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"30",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"88",
		X"00",X"00",X"00",X"70",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"00",
		X"88",X"80",X"00",X"10",X"30",X"31",X"30",X"00",X"00",X"10",X"10",X"80",X"CC",X"CC",X"C4",X"C4",
		X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F7",X"71",X"10",X"30",X"00",X"00",X"60",
		X"C8",X"A0",X"A0",X"88",X"62",X"D0",X"30",X"E0",X"73",X"F1",X"71",X"30",X"00",X"00",X"32",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"20",X"70",X"00",X"00",X"00",X"00",X"00",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"E0",X"CC",X"88",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"30",X"00",X"00",X"20",X"60",X"70",
		X"C0",X"E8",X"88",X"00",X"00",X"10",X"90",X"30",X"00",X"00",X"10",X"70",X"F0",X"F4",X"FF",X"F7",
		X"FF",X"F9",X"90",X"80",X"C0",X"80",X"00",X"D8",X"80",X"90",X"10",X"31",X"72",X"20",X"00",X"A0",
		X"70",X"60",X"80",X"10",X"D0",X"71",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"B1",X"90",X"70",X"00",X"00",X"00",X"00",X"70",X"E8",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"A0",X"00",X"00",X"40",X"40",X"00",
		X"00",X"C0",X"30",X"00",X"00",X"00",X"40",X"60",X"00",X"00",X"00",X"C0",X"20",X"20",X"20",X"20",
		X"00",X"00",X"E0",X"F0",X"F6",X"F7",X"F7",X"F3",X"00",X"00",X"00",X"80",X"D0",X"C8",X"C8",X"C8",
		X"E0",X"C0",X"00",X"00",X"C0",X"E0",X"F4",X"F6",X"60",X"20",X"10",X"10",X"10",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F7",X"F1",X"30",X"30",X"00",X"00",X"20",
		X"D8",X"A0",X"A0",X"88",X"62",X"D0",X"30",X"F0",X"F7",X"F7",X"F3",X"70",X"30",X"30",X"32",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"FC",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",X"70",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"20",X"00",X"10",X"88",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"73",X"E0",X"40",X"00",X"20",X"60",X"70",
		X"80",X"00",X"00",X"00",X"70",X"30",X"B1",X"30",X"00",X"00",X"00",X"C0",X"EC",X"FC",X"FE",X"F6",
		X"88",X"CC",X"E8",X"E4",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"10",X"31",X"72",X"20",X"80",X"80",
		X"30",X"70",X"F0",X"80",X"00",X"11",X"D5",X"F7",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"40",
		X"10",X"33",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"40",X"C8",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"E2",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"80",X"00",X"00",X"80",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"80",X"00",X"00",X"00",X"90",X"F1",X"F3",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"C8",X"C8",
		X"00",X"00",X"00",X"40",X"E0",X"F0",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"30",X"10",X"00",X"00",X"00",X"00",X"10",X"20",X"F6",X"F6",X"F3",X"73",X"70",X"10",X"A0",X"20",
		X"10",X"90",X"80",X"E0",X"B0",X"80",X"00",X"F0",X"FF",X"F3",X"F0",X"30",X"00",X"80",X"90",X"F0",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F7",X"F2",X"10",X"00",X"00",X"00",X"00",X"F6",X"FF",X"F0",X"30",X"10",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"30",X"20",X"00",X"00",X"00",X"30",X"D0",X"10",X"40",X"60",X"70",X"E4",
		X"80",X"70",X"E0",X"E0",X"60",X"00",X"80",X"20",X"F0",X"80",X"00",X"30",X"73",X"70",X"40",X"40",
		X"10",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"C0",X"E4",X"E0",X"80",X"90",X"80",X"C0",X"E4",
		X"20",X"00",X"00",X"00",X"80",X"00",X"00",X"10",X"00",X"80",X"00",X"00",X"00",X"60",X"F0",X"FE",
		X"F0",X"F9",X"FF",X"FC",X"E8",X"C0",X"00",X"F0",X"80",X"A0",X"F0",X"A0",X"10",X"30",X"40",X"00",
		X"F6",X"E0",X"00",X"00",X"00",X"00",X"60",X"F4",X"10",X"30",X"20",X"20",X"10",X"20",X"00",X"80",
		X"FE",X"FF",X"FF",X"E0",X"C0",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"E0",X"80",X"00",X"00",X"30",X"00",
		X"00",X"E0",X"10",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"20",X"20",X"60",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"40",X"40",X"40",X"C0",X"E0",
		X"00",X"00",X"00",X"60",X"10",X"10",X"10",X"30",X"70",X"60",X"70",X"00",X"00",X"80",X"90",X"A0",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F7",X"F1",X"30",X"30",X"00",X"00",X"20",
		X"D8",X"A0",X"A0",X"88",X"62",X"D0",X"30",X"F0",X"F7",X"F7",X"F3",X"70",X"30",X"30",X"32",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"20",X"00",X"10",X"88",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"76",X"73",X"E0",X"40",X"00",X"20",X"60",X"70",
		X"80",X"00",X"00",X"00",X"00",X"10",X"90",X"30",X"00",X"00",X"00",X"00",X"E0",X"F4",X"FE",X"F6",
		X"88",X"CC",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"10",X"31",X"72",X"20",X"00",X"80",
		X"30",X"70",X"F0",X"80",X"00",X"11",X"D5",X"F7",X"90",X"80",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"10",X"33",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"40",X"C8",X"C0",X"00",X"10",X"10",X"00",X"00",
		X"73",X"70",X"00",X"60",X"10",X"00",X"80",X"40",X"C8",X"80",X"00",X"00",X"00",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"10",X"20",X"80",X"00",X"00",X"80",X"C0",X"80",
		X"10",X"10",X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",
		X"C8",X"80",X"00",X"00",X"00",X"90",X"F1",X"F3",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"C8",X"C8",
		X"00",X"00",X"00",X"40",X"E0",X"F0",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F7",X"71",X"10",X"30",X"00",X"00",X"60",
		X"C8",X"A0",X"A0",X"88",X"62",X"D0",X"30",X"E0",X"73",X"71",X"70",X"30",X"00",X"00",X"32",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"20",X"00",X"00",
		X"F1",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"E0",X"CC",X"88",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"30",X"33",X"30",X"00",X"00",X"20",X"60",X"70",
		X"C0",X"E8",X"CC",X"00",X"00",X"10",X"90",X"30",X"00",X"00",X"10",X"70",X"F0",X"F4",X"FF",X"F7",
		X"FF",X"F9",X"90",X"80",X"C0",X"80",X"00",X"D8",X"80",X"90",X"10",X"31",X"72",X"20",X"00",X"A0",
		X"70",X"60",X"80",X"10",X"D0",X"71",X"10",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"B1",X"90",X"70",X"00",X"00",X"00",X"00",X"70",X"E8",X"C0",X"80",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"60",X"10",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"10",X"20",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"F6",X"F7",X"F7",X"F3",X"00",X"00",X"00",X"80",X"D0",X"C8",X"C8",X"C8",
		X"C0",X"C0",X"00",X"00",X"C0",X"E0",X"F4",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"73",X"72",X"30",X"00",X"00",X"00",X"00",
		X"C8",X"A0",X"20",X"00",X"62",X"30",X"30",X"60",X"73",X"71",X"30",X"10",X"00",X"00",X"32",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"20",X"00",X"00",
		X"F1",X"E0",X"30",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",
		X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"E0",X"CC",X"88",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"30",X"73",X"F0",X"40",X"20",X"40",X"80",X"30",
		X"80",X"C8",X"EC",X"70",X"10",X"40",X"C4",X"80",X"00",X"30",X"00",X"80",X"00",X"30",X"F0",X"F0",
		X"FC",X"F2",X"70",X"20",X"00",X"80",X"80",X"D8",X"80",X"90",X"10",X"31",X"72",X"20",X"00",X"A0",
		X"70",X"60",X"80",X"10",X"D0",X"71",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"D0",X"B1",X"90",X"70",X"00",X"00",X"00",X"00",X"70",X"E8",X"C0",X"80",X"10",X"10",X"00",X"00",
		X"00",X"00",X"20",X"60",X"10",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"30",X"10",X"20",X"F0",X"80",X"10",X"30",X"00",X"88",
		X"10",X"20",X"00",X"70",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"E0",X"C0",X"C0",X"00",
		X"88",X"80",X"00",X"10",X"30",X"71",X"F3",X"F7",X"00",X"00",X"00",X"80",X"D0",X"C8",X"C8",X"C8",
		X"40",X"C0",X"00",X"00",X"C0",X"E0",X"F4",X"F6",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"B0",X"30",X"00",X"62",X"31",X"30",X"00",X"F6",X"FC",X"64",X"00",X"51",X"11",X"32",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"40",X"80",
		X"00",X"40",X"F0",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"F0",
		X"20",X"10",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"20",X"20",X"00",X"00",X"00",X"40",X"80",X"00",
		X"00",X"20",X"10",X"10",X"30",X"73",X"F7",X"F7",X"00",X"30",X"00",X"00",X"E0",X"C8",X"E8",X"88",
		X"EC",X"FE",X"F4",X"E0",X"00",X"80",X"80",X"D8",X"00",X"10",X"10",X"31",X"72",X"20",X"00",X"A0",
		X"00",X"44",X"A8",X"10",X"D0",X"71",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"D0",X"B1",X"90",X"70",X"00",X"00",X"00",X"00",X"60",X"C8",X"90",X"B0",X"30",X"10",X"00",X"00",
		X"00",X"80",X"E0",X"60",X"10",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",
		X"40",X"40",X"00",X"00",X"00",X"00",X"31",X"30",X"10",X"20",X"F0",X"80",X"10",X"30",X"00",X"88",
		X"10",X"20",X"00",X"70",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"E0",X"C0",X"C0",X"00",
		X"88",X"80",X"00",X"10",X"30",X"31",X"30",X"00",X"00",X"00",X"00",X"80",X"CC",X"CC",X"C4",X"C4",
		X"40",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"60",X"60",X"00",X"80",X"C0",X"C0",X"B0",
		X"80",X"00",X"00",X"30",X"60",X"00",X"00",X"00",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"70",X"10",X"00",X"20",X"10",X"20",X"00",X"B0",X"90",X"50",X"40",X"C0",X"E6",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"20",X"20",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"60",X"80",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"10",X"50",X"70",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E6",X"F7",X"20",X"00",X"00",X"80",X"C0",X"E0",X"C0",X"80",
		X"90",X"FE",X"E4",X"E0",X"E0",X"80",X"10",X"FB",X"80",X"C0",X"70",X"72",X"F7",X"70",X"80",X"80",
		X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"70",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"60",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"E0",X"A0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",
		X"00",X"80",X"00",X"00",X"00",X"70",X"72",X"60",X"00",X"00",X"00",X"60",X"20",X"00",X"00",X"00",
		X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"20",X"50",X"80",X"00",X"10",X"00",X"00",X"00",X"30",X"10",X"50",X"70",X"F3",X"F7",X"F0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"30",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"70",X"E0",X"00",X"00",X"10",X"00",X"00",X"00",X"E0",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"10",X"10",X"30",X"30",X"00",X"40",X"20",X"00",X"00",X"00",X"C0",X"C8",X"C0",X"80",
		X"EC",X"FE",X"F4",X"E0",X"00",X"80",X"B0",X"FB",X"00",X"00",X"00",X"20",X"40",X"40",X"90",X"80",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"70",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"60",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"E0",X"A0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"30",X"30",X"30",X"00",X"20",X"20",X"10",X"50",X"00",X"30",X"00",X"30",
		X"20",X"C0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"D4",X"E6",X"F4",X"F0",X"70",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"00",X"00",X"00",X"20",X"22",
		X"00",X"00",X"00",X"30",X"30",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"AA",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"20",X"00",X"C0",X"C0",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"C3",X"34",X"0F",X"0F",X"C3",X"F0",X"F0",X"3C",X"F0",X"F0",
		X"E0",X"A0",X"90",X"90",X"F0",X"E0",X"C0",X"C0",X"F0",X"70",X"E0",X"10",X"80",X"70",X"F0",X"B4",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",
		X"E0",X"F0",X"D2",X"D2",X"B4",X"B4",X"F0",X"70",X"87",X"87",X"C3",X"C3",X"C3",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",
		X"07",X"2D",X"0F",X"1E",X"0F",X"3C",X"4B",X"96",X"3C",X"3C",X"3C",X"0F",X"0F",X"F0",X"F0",X"69",
		X"07",X"C3",X"F0",X"F0",X"F0",X"1E",X"E1",X"E1",X"1E",X"2D",X"0F",X"C2",X"F0",X"87",X"0F",X"0F",
		X"3C",X"58",X"12",X"20",X"D0",X"D0",X"C0",X"90",X"F0",X"30",X"00",X"00",X"00",X"30",X"71",X"73",
		X"90",X"80",X"10",X"30",X"80",X"C0",X"E0",X"F0",X"30",X"30",X"30",X"01",X"80",X"00",X"01",X"87",
		X"69",X"E1",X"E1",X"2D",X"07",X"0F",X"0F",X"0F",X"78",X"78",X"0F",X"0F",X"87",X"2D",X"0F",X"0E",
		X"1E",X"1E",X"0F",X"2D",X"2D",X"E1",X"E1",X"C3",X"87",X"87",X"87",X"C3",X"C3",X"E1",X"E1",X"E0",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"E1",X"E1",X"2D",X"2D",X"E1",X"96",X"01",X"2C",X"3C",X"78",X"78",X"F0",X"F0",X"F0",X"70",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"C0",X"EC",X"D0",X"B0",X"B1",X"B0",X"D0",X"00",X"00",X"00",X"80",X"C0",X"D8",X"EC",X"D0",
		X"F0",X"F0",X"F0",X"34",X"4B",X"3C",X"2D",X"69",X"E0",X"F0",X"C3",X"0F",X"0F",X"F0",X"78",X"78",
		X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"C3",X"34",X"0F",X"0F",X"C3",X"F0",X"F0",X"3C",X"F0",X"F0",
		X"C3",X"F0",X"C1",X"81",X"A1",X"C2",X"C0",X"40",X"B5",X"3E",X"4F",X"9E",X"2D",X"00",X"D0",X"A4",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",
		X"E0",X"F0",X"D2",X"D2",X"B4",X"B4",X"F0",X"70",X"87",X"87",X"C3",X"C3",X"C3",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",
		X"07",X"2D",X"0F",X"1E",X"0F",X"3C",X"4B",X"96",X"3C",X"3C",X"3C",X"0F",X"0F",X"F0",X"F0",X"69",
		X"07",X"C3",X"F0",X"F0",X"F0",X"1E",X"E1",X"E1",X"1E",X"2D",X"0F",X"C2",X"F0",X"87",X"0F",X"0F",
		X"3C",X"38",X"12",X"01",X"C3",X"E1",X"E1",X"F0",X"78",X"F0",X"78",X"3C",X"2D",X"2D",X"E1",X"1F",
		X"9E",X"3C",X"1E",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"A5",X"80",X"80",X"0D",X"0F",
		X"69",X"E1",X"E1",X"2D",X"07",X"0F",X"0F",X"0F",X"78",X"78",X"0F",X"0F",X"87",X"2D",X"0F",X"0E",
		X"1E",X"1E",X"0F",X"2D",X"2D",X"E1",X"E1",X"C3",X"87",X"87",X"87",X"C3",X"C3",X"E1",X"E1",X"E0",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"E1",X"E1",X"2D",X"2D",X"E1",X"96",X"0F",X"2C",X"3C",X"78",X"78",X"F0",X"F0",X"F0",X"60",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"E1",X"E1",X"C0",X"34",X"07",X"A7",X"D6",X"F8",X"30",X"70",X"E0",X"78",X"E1",X"F0",X"B0",X"50",
		X"F0",X"F0",X"F0",X"B4",X"4B",X"3C",X"2D",X"69",X"E0",X"F0",X"C3",X"0F",X"0F",X"F0",X"78",X"78",
		X"03",X"03",X"12",X"78",X"78",X"34",X"34",X"12",X"0F",X"0F",X"F0",X"87",X"F0",X"F0",X"F0",X"F0",
		X"2D",X"5A",X"86",X"1C",X"F0",X"B0",X"D0",X"F0",X"53",X"2F",X"96",X"68",X"B0",X"16",X"D2",X"F0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"78",X"34",X"01",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"78",X"30",X"10",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"12",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"61",X"E1",X"69",
		X"00",X"00",X"10",X"70",X"B4",X"3C",X"3C",X"3C",X"00",X"30",X"D2",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"21",X"07",X"34",X"78",X"78",X"03",X"03",X"03",X"69",X"69",X"E1",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"3C",X"3C",X"3C",X"F0",X"F0",X"78",X"0F",X"1E",X"1E",X"1E",X"3C",X"78",X"C2",X"2D",X"E1",X"C3",
		X"0F",X"3C",X"78",X"85",X"B0",X"86",X"87",X"87",X"70",X"38",X"B0",X"3C",X"E1",X"E1",X"F0",X"F0",
		X"48",X"0C",X"08",X"F0",X"0F",X"0F",X"87",X"87",X"00",X"00",X"00",X"F0",X"1E",X"1E",X"2C",X"2C",
		X"87",X"C3",X"C3",X"E1",X"E1",X"87",X"87",X"80",X"F0",X"F0",X"F0",X"F0",X"E1",X"C0",X"C0",X"00",
		X"C3",X"C3",X"C3",X"0E",X"00",X"00",X"00",X"00",X"48",X"48",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"87",X"87",X"87",X"87",X"87",X"87",X"00",X"C0",X"C0",X"F0",X"E1",X"E1",X"E1",X"E1",
		X"00",X"00",X"00",X"00",X"E0",X"1E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"48",
		X"87",X"07",X"30",X"F0",X"1A",X"0F",X"5E",X"9E",X"F0",X"F0",X"F0",X"D0",X"68",X"B0",X"B4",X"70",
		X"0F",X"0F",X"87",X"87",X"F0",X"08",X"08",X"08",X"2C",X"2C",X"1E",X"1E",X"F0",X"00",X"00",X"00",
		X"00",X"30",X"07",X"70",X"0F",X"87",X"87",X"87",X"00",X"D0",X"0E",X"F0",X"0E",X"C3",X"C3",X"C3",
		X"00",X"A0",X"4A",X"58",X"30",X"78",X"61",X"21",X"71",X"72",X"F0",X"C0",X"83",X"0F",X"30",X"0F",
		X"87",X"87",X"87",X"F0",X"43",X"43",X"30",X"00",X"C3",X"C3",X"F0",X"0F",X"0F",X"0F",X"F0",X"00",
		X"69",X"69",X"4B",X"69",X"69",X"78",X"F0",X"00",X"0F",X"3C",X"0F",X"0F",X"1E",X"F0",X"F0",X"00",
		X"00",X"30",X"07",X"70",X"0F",X"87",X"87",X"87",X"00",X"F0",X"0F",X"F0",X"0F",X"C3",X"C3",X"C3",
		X"00",X"F0",X"5A",X"69",X"69",X"4B",X"69",X"69",X"00",X"F0",X"F0",X"1E",X"0F",X"0F",X"3C",X"0F",
		X"87",X"87",X"87",X"F0",X"43",X"70",X"03",X"00",X"C3",X"C3",X"F0",X"0F",X"0F",X"F0",X"0F",X"00",
		X"69",X"69",X"4B",X"68",X"68",X"F0",X"4B",X"00",X"0F",X"3C",X"0F",X"01",X"08",X"41",X"34",X"31",
		X"E1",X"E1",X"C2",X"F0",X"69",X"E1",X"F0",X"E1",X"69",X"0F",X"F0",X"07",X"0F",X"0F",X"87",X"0F",
		X"3C",X"3C",X"F0",X"3C",X"0F",X"3C",X"3C",X"3C",X"80",X"80",X"80",X"F0",X"1E",X"1E",X"1E",X"1E",
		X"E1",X"F0",X"E1",X"69",X"F0",X"F0",X"C0",X"00",X"0F",X"87",X"0F",X"0F",X"3C",X"C0",X"00",X"00",
		X"3C",X"3C",X"3C",X"0F",X"F0",X"00",X"00",X"00",X"1E",X"1E",X"1E",X"96",X"F0",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F0",X"69",X"E1",X"F0",X"E1",X"00",X"00",X"C0",X"3C",X"0F",X"0F",X"87",X"0E",
		X"00",X"00",X"00",X"F0",X"0F",X"3C",X"3C",X"34",X"00",X"00",X"00",X"F0",X"96",X"1E",X"1E",X"1E",
		X"C1",X"40",X"A0",X"58",X"F1",X"E2",X"E4",X"F8",X"01",X"20",X"C1",X"89",X"03",X"B0",X"05",X"18",
		X"34",X"3C",X"3C",X"3C",X"0F",X"F0",X"3C",X"3C",X"1E",X"1E",X"1E",X"96",X"1E",X"80",X"80",X"80",
		X"02",X"02",X"02",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",X"80",X"F0",X"D0",X"D0",X"D0",
		X"10",X"10",X"00",X"00",X"F0",X"E0",X"E0",X"E0",X"D2",X"E1",X"30",X"00",X"F0",X"90",X"D0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"50",X"30",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"60",X"20",X"10",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"60",X"C0",X"40",
		X"00",X"00",X"10",X"60",X"A0",X"20",X"20",X"20",X"00",X"30",X"D0",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"30",X"70",X"70",X"02",X"02",X"02",X"40",X"40",X"C0",X"D0",X"F0",X"00",X"00",X"00",
		X"20",X"20",X"20",X"E0",X"F0",X"60",X"00",X"10",X"10",X"10",X"00",X"70",X"00",X"30",X"E1",X"C3",
		X"3C",X"78",X"F0",X"00",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"20",X"E0",X"A0",X"B0",X"B0",
		X"48",X"0C",X"08",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"60",X"60",X"00",X"00",X"80",X"B0",X"B0",X"B0",X"B0",X"A0",X"80",X"C0",X"00",
		X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"C0",X"68",X"3C",X"A0",X"B0",X"30",X"F0",X"20",X"30",X"30",X"F0",
		X"00",X"00",X"80",X"80",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"00",X"00",X"30",X"30",X"30",
		X"00",X"00",X"C0",X"F0",X"D0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"F0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"00",X"30",X"30",X"00",X"00",X"F0",X"F0",X"F0",X"00",
		X"F0",X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",X"00",
		X"00",X"00",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"00",X"00",X"30",X"30",X"30",
		X"00",X"00",X"C0",X"F0",X"D0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"F0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"00",X"00",X"30",X"30",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"F0",X"D0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"E0",X"F0",X"F0",X"E0",X"F0",X"F0",X"00",X"00",
		X"00",X"50",X"10",X"F0",X"30",X"60",X"F0",X"70",X"69",X"96",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"B0",X"B0",X"B0",X"00",X"00",X"00",X"00",X"E0",X"60",X"60",X"60",
		X"60",X"F0",X"70",X"20",X"F0",X"F0",X"C0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",
		X"B0",X"B0",X"B0",X"E0",X"F0",X"00",X"00",X"00",X"60",X"20",X"20",X"A0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"20",X"60",X"F0",X"60",X"00",X"00",X"00",X"C0",X"F0",X"70",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"E0",X"B0",X"B0",X"B0",X"00",X"00",X"00",X"00",X"E0",X"60",X"60",X"60",
		X"60",X"F0",X"60",X"20",X"F0",X"00",X"40",X"00",X"70",X"F0",X"F0",X"40",X"80",X"00",X"00",X"06",
		X"B0",X"B0",X"B0",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
