library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity program0x is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of program0x is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"40",X"01",X"00",X"11",X"36",X"00",X"23",X"0B",X"78",
		X"B1",X"20",X"F8",X"21",X"00",X"48",X"01",X"00",X"04",X"36",X"5E",X"23",X"0B",X"78",X"B1",X"20",
		X"F8",X"C3",X"D6",X"81",X"21",X"00",X"04",X"11",X"00",X"41",X"01",X"60",X"00",X"ED",X"B0",X"3E",
		X"01",X"32",X"01",X"70",X"21",X"23",X"50",X"06",X"09",X"36",X"02",X"23",X"23",X"10",X"FA",X"06",
		X"06",X"36",X"04",X"23",X"23",X"10",X"FA",X"21",X"1B",X"50",X"06",X"0A",X"36",X"07",X"2B",X"2B",
		X"10",X"FA",X"21",X"85",X"0E",X"11",X"40",X"50",X"01",X"20",X"00",X"ED",X"B0",X"00",X"00",X"00",
		X"00",X"C3",X"06",X"03",X"00",X"00",X"F5",X"E5",X"D5",X"C5",X"AF",X"32",X"01",X"70",X"3E",X"01",
		X"32",X"01",X"70",X"2A",X"00",X"42",X"23",X"22",X"00",X"42",X"21",X"00",X"40",X"3A",X"00",X"60",
		X"E6",X"10",X"28",X"08",X"CB",X"56",X"28",X"06",X"CB",X"C6",X"18",X"02",X"CB",X"D6",X"3A",X"00",
		X"68",X"E6",X"10",X"28",X"08",X"CB",X"5E",X"28",X"06",X"CB",X"CE",X"18",X"02",X"CB",X"DE",X"CD",
		X"1A",X"A7",X"CD",X"02",X"8E",X"C1",X"D1",X"E1",X"F1",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"78",X"67",X"66",X"66",X"66",X"65",X"65",X"55",X"55",X"55",X"54",X"45",
		X"55",X"54",X"44",X"43",X"44",X"44",X"44",X"43",X"34",X"34",X"34",X"34",X"34",X"43",X"33",X"34",
		X"43",X"33",X"33",X"33",X"33",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"00",
		X"00",X"00",X"EB",X"3A",X"04",X"41",X"6F",X"26",X"01",X"4E",X"21",X"08",X"41",X"7E",X"FE",X"F0",
		X"28",X"0B",X"36",X"F0",X"A1",X"EB",X"94",X"2F",X"C6",X"05",X"67",X"C9",X"00",X"36",X"0F",X"A1",
		X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"04",X"41",X"FE",X"9E",X"28",X"04",X"3C",X"32",X"04",X"41",
		X"78",X"18",X"E2",X"3A",X"04",X"41",X"FE",X"93",X"30",X"04",X"0E",X"00",X"18",X"02",X"0E",X"01",
		X"CD",X"51",X"2C",X"0F",X"38",X"1C",X"3A",X"00",X"60",X"CB",X"5F",X"28",X"01",X"2C",X"CB",X"57",
		X"28",X"01",X"2D",X"CB",X"77",X"28",X"02",X"24",X"24",X"CB",X"7F",X"C8",X"25",X"CB",X"41",X"C0",
		X"25",X"C9",X"3A",X"00",X"60",X"E6",X"02",X"28",X"06",X"25",X"CB",X"41",X"20",X"01",X"25",X"3A",
		X"00",X"68",X"CB",X"5F",X"28",X"01",X"2C",X"CB",X"57",X"28",X"01",X"2D",X"CB",X"7F",X"C8",X"24",
		X"24",X"C9",X"00",X"00",X"00",X"00",X"00",X"7E",X"FE",X"80",X"D8",X"FE",X"83",X"38",X"02",X"37",
		X"C9",X"2B",X"7E",X"23",X"D6",X"8B",X"D0",X"C6",X"0B",X"C9",X"32",X"40",X"50",X"D6",X"10",X"32",
		X"44",X"50",X"7C",X"FE",X"F0",X"38",X"03",X"3E",X"00",X"67",X"32",X"43",X"50",X"32",X"47",X"50",
		X"22",X"02",X"41",X"C9",X"2A",X"02",X"41",X"CD",X"A2",X"01",X"CD",X"E9",X"30",X"E5",X"3A",X"03",
		X"41",X"BC",X"30",X"6C",X"11",X"F3",X"10",X"19",X"CD",X"64",X"08",X"11",X"20",X"00",X"CD",X"18",
		X"19",X"38",X"4A",X"2B",X"1E",X"A0",X"CD",X"3C",X"0E",X"0E",X"08",X"1E",X"20",X"19",X"0D",X"28",
		X"20",X"CD",X"95",X"15",X"38",X"F7",X"0F",X"C6",X"2B",X"4F",X"06",X"03",X"36",X"5E",X"19",X"36",
		X"5E",X"10",X"FB",X"2B",X"36",X"5E",X"CD",X"3C",X"0E",X"36",X"5E",X"06",X"19",X"0A",X"CD",X"4E",
		X"14",X"E1",X"7C",X"3C",X"E6",X"F8",X"67",X"3E",X"73",X"32",X"04",X"41",X"3E",X"0F",X"32",X"08",
		X"41",X"7D",X"FE",X"22",X"30",X"27",X"3E",X"22",X"6F",X"CD",X"3A",X"02",X"C9",X"CD",X"3C",X"0E",
		X"CD",X"18",X"19",X"00",X"00",X"19",X"19",X"00",X"00",X"00",X"00",X"CD",X"18",X"19",X"00",X"00",
		X"C3",X"2E",X"2D",X"E1",X"CD",X"D6",X"14",X"38",X"D8",X"26",X"C7",X"18",X"CA",X"FE",X"E0",X"38",
		X"D8",X"3E",X"E0",X"18",X"D3",X"E1",X"CD",X"3B",X"8B",X"C3",X"D9",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"14",X"0A",X"CD",X"37",X"0A",X"CD",X"E1",X"0A",X"C9",
		X"60",X"0D",X"E5",X"C3",X"C8",X"2E",X"00",X"00",X"CD",X"B2",X"8D",X"CD",X"94",X"08",X"CD",X"A0",
		X"3C",X"CD",X"9C",X"99",X"CD",X"3B",X"0A",X"CD",X"51",X"18",X"CD",X"DB",X"10",X"CD",X"9D",X"9B",
		X"CD",X"B3",X"11",X"CD",X"70",X"84",X"CD",X"A1",X"82",X"CD",X"E8",X"3A",X"CD",X"50",X"26",X"CD",
		X"04",X"17",X"CD",X"E4",X"17",X"CD",X"7F",X"88",X"CD",X"AB",X"32",X"CD",X"B9",X"34",X"CD",X"A9",
		X"3A",X"CD",X"80",X"3E",X"CD",X"A0",X"8D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"00",X"42",X"7E",X"BE",X"28",X"FD",X"C3",X"18",X"03",X"7C",X"FE",X"C7",X"D8",X"FE",X"D8",
		X"3F",X"C9",X"2B",X"2B",X"36",X"9F",X"2B",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"CE",X"13",X"3E",X"00",X"32",X"01",
		X"70",X"76",X"0F",X"FE",X"0A",X"38",X"01",X"3C",X"32",X"E0",X"49",X"78",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"FE",X"0A",X"38",X"01",X"3C",X"32",X"00",X"4A",X"76",X"00",X"00",X"00",X"00",X"00",
		X"60",X"04",X"19",X"47",X"80",X"03",X"03",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"81",
		X"01",X"03",X"81",X"01",X"89",X"00",X"0F",X"00",X"00",X"02",X"05",X"04",X"75",X"81",X"86",X"00",
		X"00",X"0B",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"18",X"B1",X"00",X"35",X"B2",X"0F",X"B0",X"00",X"00",X"11",X"B3",
		X"29",X"00",X"04",X"28",X"44",X"28",X"04",X"00",X"04",X"00",X"04",X"28",X"04",X"28",X"19",X"A7",
		X"38",X"28",X"78",X"28",X"38",X"08",X"38",X"08",X"38",X"28",X"F8",X"28",X"11",X"00",X"44",X"28",
		X"04",X"10",X"04",X"10",X"04",X"28",X"11",X"00",X"19",X"AE",X"40",X"2F",X"00",X"1F",X"00",X"1F",
		X"00",X"2F",X"11",X"00",X"04",X"28",X"44",X"28",X"04",X"20",X"04",X"20",X"04",X"28",X"84",X"28",
		X"11",X"00",X"54",X"29",X"14",X"01",X"14",X"01",X"14",X"29",X"19",X"BD",X"50",X"2A",X"10",X"0A",
		X"10",X"0A",X"10",X"2A",X"29",X"11",X"99",X"B5",X"44",X"2E",X"04",X"26",X"04",X"26",X"04",X"2E",
		X"19",X"BD",X"10",X"6A",X"50",X"6A",X"10",X"5A",X"10",X"5A",X"10",X"6A",X"10",X"6A",X"11",X"00",
		X"14",X"29",X"54",X"29",X"14",X"11",X"14",X"11",X"14",X"29",X"14",X"29",X"11",X"00",X"11",X"00",
		X"71",X"28",X"31",X"08",X"31",X"08",X"31",X"28",X"11",X"00",X"67",X"AB",X"15",X"E7",X"15",X"E7",
		X"27",X"2B",X"29",X"22",X"58",X"2C",X"38",X"18",X"38",X"18",X"D8",X"2C",X"11",X"00",X"21",X"00",
		X"21",X"01",X"21",X"02",X"21",X"03",X"21",X"04",X"21",X"05",X"6D",X"EC",X"2D",X"0C",X"2D",X"0C",
		X"2D",X"EC",X"11",X"00",X"43",X"2C",X"C5",X"02",X"05",X"02",X"03",X"2C",X"11",X"00",X"00",X"2C",
		X"43",X"31",X"03",X"01",X"03",X"01",X"03",X"31",X"00",X"2C",X"11",X"00",X"04",X"2B",X"44",X"2B",
		X"38",X"08",X"38",X"08",X"04",X"2B",X"C4",X"2B",X"11",X"00",X"44",X"30",X"04",X"20",X"04",X"20",
		X"04",X"30",X"29",X"33",X"11",X"00",X"5C",X"28",X"00",X"1F",X"00",X"1F",X"1C",X"28",X"11",X"00",
		X"20",X"28",X"4B",X"30",X"0B",X"10",X"0B",X"10",X"0B",X"30",X"A0",X"28",X"11",X"00",X"44",X"33",
		X"1C",X"20",X"1C",X"20",X"04",X"33",X"11",X"00",X"40",X"2C",X"00",X"1C",X"00",X"1C",X"00",X"2C",
		X"11",X"00",X"11",X"00",X"5C",X"33",X"1C",X"03",X"1C",X"43",X"1C",X"73",X"29",X"44",X"04",X"30",
		X"44",X"30",X"00",X"24",X"00",X"24",X"04",X"30",X"04",X"30",X"11",X"00",X"1C",X"28",X"78",X"28",
		X"38",X"08",X"38",X"08",X"38",X"28",X"1C",X"28",X"11",X"00",X"11",X"00",X"47",X"33",X"07",X"03",
		X"07",X"03",X"07",X"33",X"11",X"00",X"41",X"28",X"09",X"08",X"09",X"08",X"01",X"28",X"11",X"00",
		X"47",X"28",X"38",X"18",X"38",X"18",X"C7",X"28",X"29",X"55",X"21",X"00",X"21",X"01",X"21",X"02",
		X"21",X"03",X"21",X"04",X"21",X"05",X"7F",X"30",X"07",X"27",X"07",X"27",X"3F",X"30",X"11",X"00",
		X"58",X"2C",X"18",X"0C",X"18",X"0C",X"18",X"2C",X"11",X"00",X"8C",X"86",X"87",X"88",X"89",X"8A",
		X"8B",X"15",X"07",X"00",X"07",X"00",X"07",X"05",X"07",X"8D",X"00",X"8C",X"15",X"15",X"01",X"15",
		X"01",X"15",X"05",X"15",X"8C",X"8C",X"80",X"81",X"82",X"83",X"84",X"85",X"8C",X"90",X"15",X"25",
		X"02",X"25",X"02",X"25",X"05",X"25",X"8C",X"15",X"02",X"04",X"02",X"04",X"02",X"05",X"02",X"8C",
		X"15",X"05",X"00",X"35",X"00",X"35",X"05",X"05",X"8D",X"11",X"15",X"07",X"02",X"67",X"02",X"67",
		X"05",X"07",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"15",X"17",X"01",X"17",X"01",X"17",X"05",
		X"17",X"8C",X"15",X"26",X"03",X"26",X"03",X"26",X"05",X"26",X"8C",X"86",X"87",X"88",X"89",X"8A",
		X"8B",X"05",X"27",X"01",X"27",X"01",X"27",X"05",X"27",X"8D",X"22",X"8C",X"15",X"15",X"02",X"05",
		X"02",X"05",X"05",X"15",X"8C",X"8C",X"80",X"81",X"82",X"83",X"84",X"85",X"8C",X"8C",X"15",X"15",
		X"00",X"15",X"00",X"15",X"05",X"15",X"8C",X"15",X"02",X"03",X"02",X"03",X"02",X"05",X"02",X"8C",
		X"05",X"25",X"01",X"15",X"01",X"15",X"05",X"25",X"8C",X"15",X"17",X"00",X"07",X"00",X"07",X"05",
		X"17",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"15",X"27",X"02",X"27",X"02",X"27",X"05",X"27",
		X"8C",X"05",X"17",X"00",X"17",X"00",X"17",X"05",X"17",X"8C",X"CE",X"CC",X"CF",X"79",X"52",X"48",
		X"62",X"E9",X"52",X"48",X"62",X"49",X"52",X"48",X"62",X"CD",X"33",X"CE",X"CC",X"CE",X"D0",X"45",
		X"14",X"41",X"14",X"41",X"14",X"45",X"14",X"CC",X"CC",X"CC",X"CF",X"69",X"04",X"F8",X"14",X"49",
		X"04",X"48",X"04",X"49",X"14",X"48",X"04",X"CC",X"CE",X"CC",X"CE",X"CC",X"49",X"32",X"58",X"42",
		X"49",X"32",X"48",X"42",X"79",X"32",X"48",X"42",X"8C",X"8E",X"8D",X"44",X"8C",X"8C",X"8E",X"8C",
		X"8C",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8C",X"8E",X"8C",X"59",X"62",X"68",X"52",X"49",
		X"32",X"48",X"42",X"8C",X"8E",X"11",X"1F",X"13",X"09",X"00",X"0B",X"0B",X"0B",X"0B",X"11",X"11",
		X"41",X"0B",X"B1",X"00",X"20",X"0B",X"11",X"11",X"65",X"87",X"11",X"13",X"0A",X"00",X"0B",X"12",
		X"0B",X"11",X"0C",X"00",X"0B",X"0B",X"21",X"11",X"65",X"87",X"11",X"31",X"0A",X"00",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"21",X"11",X"80",X"81",X"A0",X"85",X"21",X"22",X"92",X"00",X"12",X"12",
		X"12",X"32",X"B1",X"80",X"B0",X"89",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"81",X"20",
		X"21",X"22",X"92",X"84",X"12",X"32",X"31",X"B0",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"80",X"81",X"20",X"21",X"A2",X"86",X"23",X"93",X"00",X"13",X"13",X"13",X"24",X"25",X"26",
		X"96",X"84",X"16",X"75",X"73",X"71",X"60",X"00",X"80",X"17",X"80",X"8A",X"00",X"00",X"00",X"40",
		X"51",X"53",X"55",X"96",X"84",X"16",X"57",X"18",X"98",X"14",X"18",X"18",X"18",X"77",X"B6",X"80",
		X"35",X"34",X"33",X"92",X"00",X"12",X"12",X"12",X"71",X"60",X"00",X"00",X"80",X"10",X"00",X"00",
		X"00",X"00",X"40",X"51",X"53",X"55",X"96",X"02",X"16",X"16",X"16",X"27",X"28",X"29",X"2A",X"2B",
		X"9B",X"00",X"1B",X"1B",X"1B",X"2C",X"2D",X"2E",X"9E",X"10",X"1E",X"1E",X"1E",X"7D",X"7B",X"F9",
		X"80",X"77",X"96",X"01",X"16",X"16",X"16",X"36",X"35",X"B4",X"80",X"33",X"32",X"31",X"30",X"00",
		X"80",X"8A",X"80",X"17",X"00",X"00",X"00",X"00",X"00",X"40",X"51",X"53",X"55",X"57",X"98",X"02",
		X"18",X"18",X"18",X"29",X"2A",X"2B",X"1B",X"9B",X"84",X"1B",X"2C",X"2D",X"2E",X"9E",X"17",X"1E",
		X"1E",X"1E",X"7D",X"7B",X"79",X"F7",X"80",X"75",X"73",X"71",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"87",X"52",X"93",X"80",X"13",X"13",X"13",X"72",X"70",X"00",X"00",X"00",
		X"3E",X"FF",X"32",X"00",X"78",X"C3",X"E9",X"A6",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"37",X"81",
		X"E0",X"80",X"0B",X"83",X"E0",X"82",X"2F",X"8B",X"8B",X"8B",X"01",X"83",X"E0",X"E0",X"0D",X"E0",
		X"E0",X"82",X"0D",X"84",X"84",X"84",X"0C",X"84",X"84",X"85",X"15",X"86",X"84",X"85",X"0A",X"86",
		X"84",X"84",X"13",X"87",X"87",X"87",X"02",X"88",X"88",X"88",X"04",X"8A",X"8A",X"8A",X"07",X"8B",
		X"8B",X"8B",X"01",X"3A",X"15",X"41",X"FE",X"14",X"CA",X"1E",X"1B",X"CD",X"55",X"0F",X"CD",X"00",
		X"0D",X"C3",X"CB",X"17",X"05",X"3A",X"34",X"50",X"B8",X"D9",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7C",X"0F",X"0F",X"0F",X"E6",X"1F",X"5F",X"16",X"48",X"87",X"4F",X"06",
		X"50",X"0A",X"95",X"D6",X"0F",X"47",X"07",X"07",X"E6",X"E0",X"4F",X"78",X"07",X"07",X"E6",X"03",
		X"47",X"EB",X"09",X"C9",X"8E",X"2B",X"8E",X"2B",X"57",X"19",X"8E",X"2B",X"8E",X"2B",X"AC",X"33",
		X"B0",X"36",X"00",X"00",X"3A",X"0C",X"41",X"07",X"C6",X"84",X"6F",X"26",X"08",X"5E",X"23",X"56",
		X"EB",X"E9",X"3A",X"0D",X"41",X"A7",X"20",X"53",X"2A",X"02",X"41",X"3A",X"0B",X"41",X"47",X"3A",
		X"00",X"42",X"E6",X"03",X"B8",X"30",X"01",X"2C",X"CD",X"A2",X"01",X"7C",X"FE",X"CD",X"30",X"53",
		X"7D",X"FE",X"E0",X"38",X"03",X"2E",X"E0",X"7D",X"32",X"40",X"50",X"D6",X"10",X"32",X"44",X"50",
		X"7C",X"32",X"43",X"50",X"32",X"47",X"50",X"22",X"02",X"41",X"2A",X"09",X"41",X"CD",X"D3",X"01",
		X"7D",X"FE",X"E0",X"38",X"03",X"2E",X"E0",X"7D",X"FE",X"22",X"30",X"03",X"2E",X"22",X"7D",X"32",
		X"4C",X"50",X"32",X"09",X"41",X"D6",X"0F",X"32",X"48",X"50",X"C9",X"00",X"00",X"00",X"21",X"0D",
		X"41",X"35",X"20",X"D6",X"21",X"07",X"41",X"CB",X"46",X"20",X"04",X"CB",X"CE",X"18",X"15",X"CB",
		X"D6",X"18",X"11",X"3A",X"09",X"41",X"95",X"C6",X"0C",X"FE",X"18",X"38",X"07",X"3E",X"08",X"32",
		X"0D",X"41",X"18",X"B6",X"2A",X"09",X"41",X"22",X"02",X"41",X"3E",X"00",X"32",X"4C",X"50",X"3E",
		X"07",X"32",X"4A",X"50",X"3E",X"73",X"32",X"04",X"41",X"3E",X"0F",X"32",X"08",X"41",X"21",X"03",
		X"05",X"22",X"4D",X"50",X"3E",X"01",X"32",X"0C",X"41",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"A6",X"69",X"9A",X"66",X"66",X"59",X"56",X"56",X"55",X"55",X"54",X"14",X"45",
		X"44",X"10",X"04",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"41",X"10",X"44",X"44",X"51",
		X"54",X"54",X"55",X"56",X"96",X"65",X"66",X"9A",X"A6",X"69",X"AA",X"AA",X"AA",X"06",X"03",X"21",
		X"50",X"50",X"7E",X"A7",X"28",X"2F",X"35",X"23",X"23",X"23",X"7D",X"00",X"E6",X"0C",X"0F",X"C6",
		X"0E",X"5F",X"16",X"41",X"1A",X"07",X"07",X"4F",X"12",X"30",X"33",X"13",X"1A",X"3C",X"FE",X"8D",
		X"20",X"02",X"3E",X"60",X"12",X"5F",X"16",X"09",X"1A",X"A1",X"28",X"26",X"E6",X"AA",X"28",X"01",
		X"35",X"23",X"10",X"CE",X"C9",X"3A",X"00",X"42",X"E6",X"3F",X"20",X"0C",X"CD",X"FA",X"18",X"00",
		X"00",X"00",X"30",X"04",X"C6",X"50",X"36",X"F1",X"23",X"23",X"23",X"77",X"18",X"E3",X"13",X"1A",
		X"18",X"D3",X"34",X"18",X"DC",X"A0",X"4B",X"68",X"66",X"60",X"6C",X"63",X"69",X"5E",X"01",X"5E",
		X"5E",X"64",X"65",X"5E",X"6A",X"61",X"67",X"69",X"63",X"5E",X"5E",X"68",X"66",X"60",X"6C",X"63",
		X"69",X"5E",X"02",X"FF",X"3F",X"49",X"61",X"69",X"63",X"62",X"65",X"6B",X"FF",X"BF",X"4B",X"65",
		X"74",X"64",X"6B",X"FF",X"21",X"E5",X"09",X"3E",X"02",X"18",X"02",X"3E",X"01",X"08",X"01",X"1F",
		X"00",X"5E",X"23",X"56",X"23",X"7E",X"FE",X"FF",X"28",X"07",X"12",X"EB",X"ED",X"42",X"EB",X"18",
		X"F3",X"23",X"08",X"3D",X"20",X"E7",X"C9",X"3E",X"14",X"18",X"02",X"3E",X"01",X"08",X"3A",X"01",
		X"40",X"3C",X"FE",X"14",X"20",X"01",X"AF",X"32",X"01",X"40",X"C6",X"02",X"5F",X"16",X"42",X"D6",
		X"14",X"30",X"0F",X"C6",X"06",X"38",X"10",X"C6",X"06",X"38",X"11",X"C6",X"06",X"21",X"E1",X"4A",
		X"18",X"0D",X"21",X"5F",X"48",X"18",X"08",X"21",X"61",X"48",X"18",X"03",X"21",X"A1",X"49",X"0F",
		X"0F",X"0F",X"4F",X"06",X"00",X"09",X"1A",X"77",X"08",X"3D",X"20",X"C1",X"C9",X"80",X"81",X"82",
		X"80",X"82",X"81",X"80",X"81",X"80",X"81",X"82",X"80",X"A9",X"A7",X"A9",X"A7",X"AB",X"A7",X"AB",
		X"AD",X"A9",X"A7",X"A9",X"AB",X"AF",X"AF",X"AB",X"A7",X"A9",X"AB",X"A9",X"A7",X"A9",X"AB",X"A7",
		X"AB",X"A7",X"A9",X"AD",X"B1",X"AF",X"A9",X"4E",X"4E",X"66",X"63",X"6B",X"67",X"64",X"4E",X"4E",
		X"4E",X"63",X"6F",X"60",X"61",X"4E",X"63",X"69",X"67",X"6B",X"6A",X"4E",X"4E",X"63",X"6F",X"60",
		X"61",X"4E",X"4E",X"4E",X"4E",X"19",X"67",X"18",X"63",X"69",X"5E",X"0A",X"07",X"07",X"E6",X"E0",
		X"5F",X"0A",X"07",X"07",X"E6",X"03",X"57",X"19",X"C9",X"A7",X"ED",X"52",X"BC",X"C0",X"26",X"4B",
		X"C9",X"CD",X"EF",X"13",X"36",X"07",X"23",X"23",X"36",X"07",X"11",X"20",X"00",X"21",X"1B",X"48",
		X"0E",X"03",X"E5",X"06",X"20",X"36",X"9D",X"19",X"10",X"FB",X"E1",X"23",X"0D",X"20",X"F3",X"C9",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"04",X"04",X"07",X"04",X"04",X"07",X"06",X"07",
		X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"04",X"04",X"07",X"06",
		X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"04",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"02",X"02",X"07",X"07",X"07",
		X"07",X"06",X"02",X"02",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",
		X"02",X"07",X"01",X"04",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"04",X"04",X"2A",X"00",X"41",X"54",X"5D",X"01",X"34",X"50",X"0A",X"E6",
		X"07",X"C0",X"7D",X"FE",X"1A",X"28",X"10",X"FE",X"D8",X"20",X"05",X"7C",X"FE",X"05",X"28",X"1C",
		X"23",X"23",X"22",X"00",X"41",X"18",X"38",X"3A",X"15",X"41",X"FE",X"01",X"00",X"00",X"21",X"14",
		X"41",X"36",X"89",X"21",X"1A",X"05",X"3C",X"32",X"15",X"41",X"18",X"E4",X"3A",X"15",X"41",X"FE",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"DA",X"05",X"22",X"00",X"41",X"21",X"B3",
		X"02",X"22",X"14",X"41",X"C9",X"21",X"14",X"41",X"36",X"98",X"21",X"1A",X"05",X"18",X"D7",X"21",
		X"3A",X"48",X"D5",X"CD",X"CB",X"0A",X"D1",X"1A",X"E6",X"07",X"3D",X"20",X"4A",X"1A",X"E6",X"3F",
		X"FE",X"09",X"20",X"0B",X"36",X"84",X"06",X"0E",X"2B",X"36",X"81",X"10",X"FB",X"18",X"34",X"30",
		X"15",X"01",X"06",X"04",X"36",X"88",X"2B",X"36",X"80",X"2B",X"36",X"82",X"10",X"F8",X"41",X"2B",
		X"36",X"82",X"10",X"FB",X"18",X"1D",X"FE",X"19",X"28",X"54",X"D8",X"FE",X"29",X"38",X"77",X"28",
		X"63",X"13",X"1A",X"E6",X"38",X"0F",X"0F",X"0F",X"C6",X"83",X"77",X"06",X"0A",X"2B",X"36",X"81",
		X"10",X"FB",X"1B",X"2B",X"C3",X"AF",X"0C",X"13",X"1A",X"E6",X"38",X"0F",X"0F",X"0F",X"C6",X"83",
		X"77",X"2B",X"1A",X"E6",X"C0",X"07",X"07",X"4F",X"07",X"81",X"C6",X"7D",X"4F",X"06",X"0A",X"1B",
		X"1A",X"E6",X"07",X"28",X"08",X"08",X"0A",X"77",X"2B",X"08",X"3D",X"20",X"F8",X"03",X"1A",X"E6",
		X"38",X"28",X"5C",X"08",X"0A",X"77",X"2B",X"08",X"D6",X"08",X"20",X"F7",X"18",X"51",X"1A",X"07",
		X"30",X"04",X"2B",X"2B",X"2B",X"2B",X"13",X"1A",X"5F",X"16",X"0A",X"06",X"08",X"1A",X"77",X"2B",
		X"13",X"10",X"FA",X"C9",X"13",X"1A",X"16",X"0B",X"5F",X"21",X"35",X"50",X"06",X"11",X"1A",X"77",
		X"2B",X"2B",X"13",X"10",X"F9",X"C9",X"13",X"1A",X"A7",X"28",X"0F",X"FE",X"05",X"28",X"0B",X"CD",
		X"72",X"03",X"36",X"88",X"2B",X"36",X"88",X"2B",X"18",X"07",X"06",X"05",X"36",X"88",X"2B",X"10",
		X"FB",X"C6",X"C5",X"4F",X"06",X"0A",X"0A",X"77",X"FE",X"18",X"C0",X"22",X"02",X"40",X"C9",X"03",
		X"13",X"1A",X"E6",X"07",X"28",X"08",X"08",X"0A",X"77",X"2B",X"08",X"3D",X"20",X"F8",X"1B",X"1A",
		X"06",X"0A",X"E6",X"C0",X"C8",X"D5",X"11",X"20",X"00",X"07",X"30",X"1C",X"06",X"A2",X"07",X"30",
		X"02",X"06",X"A5",X"7D",X"E6",X"E0",X"C6",X"0D",X"6F",X"70",X"3E",X"47",X"CD",X"D9",X"0A",X"05",
		X"70",X"CD",X"D9",X"0A",X"05",X"70",X"D1",X"C9",X"3A",X"14",X"41",X"4F",X"3C",X"CD",X"46",X"87",
		X"3E",X"47",X"36",X"7F",X"2B",X"36",X"7E",X"CD",X"D9",X"0A",X"36",X"7C",X"23",X"36",X"7D",X"CD",
		X"D9",X"0A",X"0A",X"77",X"3E",X"47",X"CD",X"D9",X"0A",X"0A",X"3D",X"77",X"D1",X"C9",X"00",X"00",
		X"21",X"DA",X"4B",X"01",X"34",X"50",X"0A",X"E6",X"07",X"3D",X"20",X"0A",X"CD",X"CB",X"0A",X"06",
		X"11",X"36",X"5E",X"2B",X"10",X"FB",X"21",X"3A",X"50",X"06",X"14",X"35",X"2D",X"2D",X"10",X"FB",
		X"C9",X"FF",X"CE",X"4B",X"6D",X"67",X"4E",X"8D",X"FF",X"F1",X"4B",X"69",X"63",X"60",X"62",X"6C",
		X"FF",X"2F",X"48",X"66",X"6E",X"6E",X"63",X"FF",X"32",X"4B",X"6B",X"74",X"62",X"6A",X"FF",X"21",
		X"02",X"48",X"01",X"1C",X"20",X"11",X"20",X"00",X"78",X"E5",X"47",X"36",X"5E",X"19",X"10",X"FB",
		X"E1",X"23",X"0D",X"20",X"F4",X"C9",X"CD",X"67",X"36",X"7E",X"BE",X"28",X"FD",X"10",X"F7",X"C9",
		X"CD",X"38",X"83",X"CD",X"33",X"87",X"06",X"D0",X"C5",X"CD",X"66",X"0B",X"CD",X"00",X"0D",X"C1",
		X"10",X"F6",X"06",X"07",X"21",X"AB",X"4B",X"11",X"20",X"00",X"36",X"8A",X"19",X"10",X"FB",X"21",
		X"AC",X"4B",X"36",X"9B",X"06",X"03",X"19",X"36",X"9C",X"19",X"36",X"9B",X"10",X"F8",X"21",X"29",
		X"0D",X"CD",X"D0",X"9C",X"11",X"03",X"20",X"0E",X"0A",X"06",X"02",X"3A",X"02",X"41",X"3C",X"32",
		X"02",X"41",X"32",X"40",X"50",X"D6",X"10",X"32",X"44",X"50",X"CD",X"56",X"0D",X"15",X"28",X"3A",
		X"0D",X"20",X"E6",X"7B",X"1D",X"FE",X"03",X"28",X"13",X"FE",X"02",X"28",X"21",X"D5",X"3E",X"5E",
		X"32",X"AF",X"4B",X"21",X"22",X"0D",X"CD",X"1B",X"0A",X"D1",X"18",X"CB",X"D5",X"21",X"71",X"4B",
		X"01",X"01",X"05",X"CD",X"45",X"0D",X"3E",X"9E",X"32",X"B0",X"4B",X"D1",X"18",X"B9",X"3E",X"5E",
		X"32",X"B0",X"4B",X"3E",X"9E",X"32",X"AF",X"4B",X"18",X"AD",X"06",X"40",X"CD",X"56",X"0D",X"21",
		X"6E",X"4B",X"01",X"01",X"04",X"CD",X"45",X"0D",X"3E",X"40",X"32",X"16",X"42",X"C3",X"18",X"03",
		X"E5",X"21",X"03",X"42",X"3A",X"07",X"41",X"0F",X"30",X"02",X"2E",X"0F",X"E5",X"06",X"05",X"79",
		X"0D",X"D6",X"05",X"38",X"0D",X"4F",X"05",X"7E",X"C6",X"05",X"FE",X"0A",X"38",X"0E",X"D6",X"0A",
		X"77",X"23",X"7E",X"3C",X"FE",X"0A",X"20",X"04",X"AF",X"77",X"10",X"F5",X"77",X"E1",X"79",X"A7",
		X"20",X"DA",X"E1",X"C9",X"4F",X"C3",X"6C",X"2C",X"00",X"00",X"00",X"00",X"A7",X"ED",X"52",X"7C",
		X"FE",X"47",X"C0",X"26",X"4B",X"C9",X"3A",X"02",X"41",X"D6",X"18",X"32",X"48",X"50",X"3A",X"03",
		X"41",X"32",X"4B",X"50",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"05",X"6F",X"26",X"41",X"7E",X"07",
		X"07",X"07",X"47",X"3A",X"00",X"42",X"E6",X"7C",X"0E",X"17",X"B8",X"30",X"11",X"0D",X"FE",X"14",
		X"28",X"0C",X"0D",X"FE",X"0C",X"28",X"07",X"0D",X"FE",X"04",X"28",X"02",X"0E",X"17",X"79",X"32",
		X"49",X"50",X"C9",X"00",X"00",X"19",X"10",X"04",X"47",X"09",X"11",X"04",X"47",X"D1",X"17",X"07",
		X"47",X"F1",X"03",X"07",X"A7",X"F1",X"0C",X"07",X"C7",X"F1",X"0A",X"07",X"C7",X"F1",X"08",X"07",
		X"97",X"F1",X"2F",X"06",X"A7",X"80",X"80",X"81",X"81",X"82",X"82",X"80",X"81",X"81",X"80",X"80",
		X"82",X"82",X"80",X"B7",X"AD",X"AB",X"B5",X"A9",X"B7",X"B7",X"B7",X"AD",X"A7",X"B7",X"B7",X"B7",
		X"A9",X"B5",X"B7",X"AB",X"B7",X"B7",X"B7",X"B5",X"B3",X"B5",X"B7",X"B1",X"B1",X"A9",X"AB",X"B1",
		X"AD",X"AF",X"4E",X"67",X"6E",X"65",X"6A",X"60",X"61",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"04",
		X"04",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"04",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"06",X"04",X"06",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"3A",X"15",X"41",X"FE",X"02",X"DA",X"68",X"26",X"FE",X"0A",X"D2",
		X"EB",X"12",X"2A",X"00",X"41",X"54",X"5D",X"01",X"34",X"50",X"0A",X"E6",X"07",X"C0",X"21",X"3A",
		X"48",X"D5",X"CD",X"CB",X"0A",X"D1",X"1A",X"CB",X"77",X"28",X"08",X"E5",X"23",X"36",X"DE",X"CD",
		X"F7",X"13",X"E1",X"FE",X"80",X"38",X"04",X"FE",X"E0",X"38",X"59",X"E6",X"0F",X"C6",X"83",X"77",
		X"2B",X"D5",X"13",X"1A",X"E6",X"0F",X"47",X"1A",X"E6",X"F0",X"0F",X"0F",X"0F",X"C6",X"A5",X"5F",
		X"16",X"0E",X"1A",X"77",X"2B",X"13",X"1A",X"77",X"2B",X"1B",X"10",X"F6",X"D1",X"1A",X"E6",X"F0",
		X"FE",X"E0",X"28",X"48",X"FE",X"F0",X"28",X"49",X"CB",X"6F",X"28",X"0C",X"7D",X"E6",X"E0",X"C6",
		X"0D",X"32",X"04",X"40",X"7C",X"32",X"05",X"40",X"1A",X"07",X"07",X"06",X"0E",X"CD",X"B2",X"0C",
		X"EB",X"23",X"7D",X"FE",X"39",X"28",X"2F",X"FE",X"99",X"28",X"3B",X"FE",X"F4",X"28",X"4C",X"23",
		X"22",X"00",X"41",X"C9",X"D5",X"E6",X"BF",X"FE",X"90",X"20",X"63",X"11",X"A8",X"0A",X"2B",X"2B",
		X"06",X"07",X"1A",X"77",X"2B",X"13",X"10",X"FA",X"D1",X"EB",X"18",X"D6",X"22",X"0A",X"40",X"18",
		X"CF",X"CD",X"AA",X"11",X"18",X"CA",X"3A",X"15",X"41",X"FE",X"05",X"18",X"03",X"21",X"D9",X"05",
		X"3C",X"32",X"15",X"41",X"18",X"C9",X"3A",X"15",X"41",X"FE",X"07",X"00",X"00",X"3E",X"04",X"CD",
		X"FE",X"13",X"3E",X"03",X"18",X"EA",X"21",X"39",X"06",X"18",X"E5",X"7C",X"FE",X"06",X"20",X"AF",
		X"3A",X"15",X"41",X"FE",X"06",X"18",X"05",X"21",X"99",X"06",X"18",X"D4",X"3E",X"01",X"32",X"0C",
		X"41",X"21",X"F5",X"06",X"22",X"00",X"41",X"21",X"B3",X"0B",X"22",X"14",X"41",X"C9",X"FE",X"8E",
		X"20",X"04",X"36",X"DF",X"18",X"A2",X"38",X"05",X"11",X"D3",X"0E",X"18",X"93",X"FE",X"8C",X"28",
		X"F3",X"38",X"09",X"13",X"1A",X"16",X"0F",X"C3",X"CD",X"10",X"00",X"00",X"FE",X"82",X"20",X"11",
		X"F5",X"3E",X"8F",X"32",X"5B",X"50",X"3E",X"F1",X"32",X"58",X"50",X"3E",X"01",X"32",X"0E",X"40",
		X"F1",X"01",X"03",X"08",X"D6",X"86",X"38",X"15",X"28",X"2E",X"FE",X"05",X"28",X"2A",X"2B",X"2B",
		X"36",X"9F",X"2B",X"36",X"89",X"2B",X"0D",X"28",X"24",X"36",X"88",X"18",X"F5",X"01",X"06",X"0F",
		X"C6",X"06",X"28",X"14",X"FE",X"05",X"28",X"10",X"2B",X"2B",X"36",X"9F",X"2B",X"36",X"88",X"2B",
		X"36",X"89",X"0D",X"20",X"F7",X"2B",X"18",X"0C",X"36",X"88",X"2B",X"10",X"FB",X"FE",X"02",X"20",
		X"03",X"22",X"02",X"40",X"C6",X"C5",X"4F",X"06",X"0A",X"0A",X"77",X"18",X"87",X"CD",X"68",X"0C",
		X"D1",X"C3",X"D0",X"0F",X"2A",X"00",X"42",X"C3",X"08",X"14",X"00",X"01",X"34",X"50",X"0A",X"E6",
		X"07",X"FE",X"01",X"C0",X"2A",X"02",X"40",X"CD",X"13",X"11",X"20",X"05",X"AF",X"32",X"03",X"40",
		X"C9",X"2A",X"02",X"40",X"7C",X"A7",X"C8",X"0A",X"0E",X"23",X"E6",X"20",X"20",X"02",X"0E",X"27",
		X"2B",X"71",X"2B",X"0D",X"71",X"CD",X"52",X"96",X"A7",X"CD",X"6E",X"11",X"0D",X"0D",X"71",X"23",
		X"0C",X"71",X"C9",X"7D",X"E6",X"E0",X"C6",X"1A",X"6F",X"E5",X"21",X"BA",X"4B",X"CD",X"CB",X"0A",
		X"D1",X"A7",X"ED",X"52",X"C8",X"11",X"00",X"04",X"A7",X"ED",X"52",X"C9",X"CD",X"C4",X"8D",X"A7",
		X"C8",X"4F",X"21",X"5B",X"50",X"7E",X"0D",X"20",X"07",X"FE",X"47",X"28",X"0E",X"35",X"18",X"10",
		X"FE",X"C7",X"28",X"03",X"34",X"18",X"09",X"3E",X"01",X"18",X"02",X"3E",X"02",X"32",X"0E",X"40",
		X"2E",X"58",X"35",X"20",X"05",X"AF",X"32",X"0E",X"40",X"C9",X"3A",X"00",X"42",X"E6",X"3F",X"28",
		X"09",X"FE",X"20",X"C0",X"3E",X"08",X"32",X"59",X"50",X"C9",X"3E",X"09",X"18",X"F8",X"3E",X"47",
		X"C3",X"D9",X"0A",X"B1",X"01",X"34",X"50",X"0A",X"E6",X"07",X"FE",X"02",X"C0",X"2A",X"0A",X"40",
		X"CD",X"13",X"11",X"20",X"05",X"AF",X"32",X"0B",X"40",X"C9",X"2A",X"0A",X"40",X"7C",X"A7",X"C8",
		X"0A",X"0E",X"23",X"E6",X"40",X"28",X"0A",X"01",X"73",X"11",X"11",X"20",X"00",X"D5",X"C3",X"E0",
		X"0C",X"CD",X"01",X"11",X"CD",X"6E",X"11",X"C3",X"CE",X"14",X"D5",X"CD",X"97",X"11",X"D1",X"22",
		X"0C",X"40",X"C9",X"01",X"34",X"50",X"0A",X"E6",X"07",X"FE",X"02",X"C0",X"2A",X"0C",X"40",X"CD",
		X"13",X"11",X"20",X"05",X"AF",X"32",X"0D",X"40",X"C9",X"2A",X"0C",X"40",X"7C",X"A7",X"C8",X"11",
		X"20",X"00",X"0A",X"E6",X"18",X"C0",X"0A",X"E6",X"60",X"0F",X"0F",X"0F",X"00",X"C6",X"A8",X"77",
		X"19",X"3C",X"77",X"C9",X"3A",X"00",X"42",X"0F",X"38",X"0B",X"21",X"12",X"50",X"06",X"07",X"35",
		X"2B",X"2B",X"10",X"FB",X"00",X"01",X"12",X"50",X"0A",X"E6",X"07",X"FE",X"02",X"C0",X"21",X"C9",
		X"4B",X"CD",X"CB",X"0A",X"06",X"07",X"36",X"5E",X"2B",X"10",X"FB",X"01",X"12",X"50",X"0A",X"CD",
		X"01",X"18",X"00",X"C0",X"ED",X"5F",X"FE",X"40",X"D0",X"21",X"29",X"48",X"CD",X"CB",X"0A",X"0E",
		X"A2",X"3A",X"12",X"50",X"07",X"30",X"0A",X"2B",X"2B",X"2B",X"0E",X"A5",X"22",X"08",X"40",X"18",
		X"03",X"22",X"06",X"40",X"CD",X"A1",X"93",X"71",X"CD",X"6E",X"11",X"0D",X"71",X"CD",X"D9",X"0A",
		X"0D",X"71",X"C9",X"21",X"54",X"50",X"3A",X"00",X"42",X"47",X"0E",X"0A",X"E6",X"3F",X"FE",X"38",
		X"28",X"05",X"FE",X"18",X"20",X"0A",X"0C",X"79",X"32",X"55",X"50",X"3C",X"3C",X"32",X"51",X"50",
		X"3A",X"0F",X"40",X"A7",X"20",X"0F",X"78",X"FE",X"40",X"D2",X"C2",X"9F",X"3A",X"00",X"68",X"E6",
		X"40",X"28",X"01",X"35",X"35",X"35",X"7E",X"2E",X"50",X"77",X"11",X"0F",X"40",X"1A",X"A7",X"28",
		X"16",X"2E",X"53",X"FE",X"50",X"38",X"07",X"FE",X"9F",X"20",X"07",X"AF",X"12",X"C9",X"35",X"35",
		X"18",X"02",X"34",X"34",X"3C",X"12",X"C9",X"CD",X"A1",X"87",X"96",X"FE",X"80",X"C0",X"CB",X"50",
		X"C0",X"3E",X"01",X"12",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",
		X"00",X"42",X"06",X"10",X"CB",X"67",X"28",X"08",X"06",X"0E",X"CB",X"6F",X"28",X"02",X"06",X"12",
		X"78",X"32",X"41",X"50",X"3C",X"32",X"45",X"50",X"C9",X"00",X"00",X"FE",X"0D",X"D2",X"BE",X"15",
		X"01",X"34",X"50",X"0A",X"E6",X"07",X"C0",X"21",X"3A",X"48",X"CD",X"CB",X"0A",X"E5",X"2A",X"00",
		X"41",X"4E",X"EB",X"21",X"16",X"41",X"06",X"0F",X"7E",X"FE",X"0F",X"79",X"20",X"2A",X"F5",X"13",
		X"C3",X"ED",X"3D",X"20",X"1C",X"11",X"F5",X"06",X"3A",X"15",X"41",X"3C",X"32",X"15",X"41",X"FE",
		X"0D",X"20",X"0E",X"F1",X"E1",X"3E",X"04",X"00",X"00",X"00",X"21",X"26",X"07",X"C3",X"00",X"8A",
		X"C9",X"F1",X"06",X"F0",X"0F",X"0F",X"0F",X"0F",X"70",X"EB",X"22",X"00",X"41",X"11",X"20",X"00",
		X"E1",X"E6",X"0F",X"C8",X"E5",X"3D",X"28",X"44",X"3D",X"28",X"22",X"3D",X"28",X"2A",X"3D",X"28",
		X"13",X"E1",X"FE",X"05",X"30",X"3A",X"3D",X"47",X"07",X"80",X"C6",X"94",X"77",X"2B",X"3C",X"77",
		X"2B",X"3C",X"77",X"C9",X"7D",X"D6",X"0E",X"6F",X"22",X"08",X"40",X"18",X"07",X"7D",X"D6",X"07",
		X"6F",X"22",X"04",X"40",X"0E",X"A2",X"18",X"09",X"7D",X"D6",X"0A",X"6F",X"22",X"06",X"40",X"0E",
		X"A5",X"71",X"CD",X"6E",X"11",X"0D",X"71",X"CD",X"D9",X"0A",X"0D",X"71",X"E1",X"36",X"DF",X"C9",
		X"01",X"89",X"0A",X"D6",X"05",X"28",X"05",X"3D",X"20",X"07",X"0E",X"8D",X"D5",X"CD",X"E0",X"0C",
		X"C9",X"0E",X"AD",X"3D",X"28",X"05",X"3D",X"20",X"19",X"0E",X"AF",X"2C",X"22",X"02",X"40",X"C9",
		X"CD",X"6E",X"11",X"36",X"F4",X"23",X"36",X"F5",X"CD",X"D9",X"0A",X"71",X"CD",X"6E",X"11",X"0D",
		X"71",X"C9",X"06",X"19",X"21",X"35",X"50",X"36",X"04",X"2B",X"2B",X"10",X"FA",X"C9",X"F5",X"C5",
		X"47",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"56",X"32",X"E0",X"49",X"78",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"56",X"32",X"00",X"4A",X"C1",X"F1",X"C9",X"21",
		X"37",X"50",X"36",X"07",X"23",X"23",X"C9",X"23",X"36",X"DE",X"23",X"36",X"DE",X"C9",X"32",X"37",
		X"50",X"32",X"39",X"50",X"32",X"3B",X"50",X"C9",X"7D",X"4D",X"44",X"00",X"E6",X"0F",X"FE",X"08",
		X"C0",X"21",X"06",X"40",X"CB",X"48",X"28",X"08",X"2E",X"04",X"CB",X"50",X"28",X"02",X"2E",X"08",
		X"06",X"03",X"C5",X"5E",X"23",X"56",X"E5",X"1A",X"FE",X"A5",X"28",X"04",X"FE",X"8F",X"20",X"11",
		X"EB",X"78",X"FE",X"03",X"18",X"07",X"0E",X"5F",X"CD",X"00",X"11",X"18",X"04",X"79",X"CD",X"F8",
		X"10",X"E1",X"23",X"7D",X"FE",X"0A",X"20",X"02",X"2E",X"04",X"C1",X"10",X"D5",X"C9",X"FE",X"00",
		X"28",X"28",X"4F",X"C5",X"E5",X"2A",X"0C",X"40",X"2B",X"19",X"19",X"C1",X"A7",X"ED",X"42",X"20",
		X"06",X"AF",X"32",X"0D",X"40",X"18",X"0F",X"2A",X"0A",X"40",X"CD",X"6E",X"11",X"2B",X"AF",X"ED",
		X"42",X"20",X"03",X"32",X"0B",X"40",X"C1",X"C3",X"6C",X"2C",X"E5",X"2A",X"11",X"40",X"EB",X"2A",
		X"00",X"41",X"ED",X"52",X"11",X"24",X"00",X"ED",X"52",X"1E",X"20",X"30",X"14",X"3A",X"13",X"40",
		X"C6",X"02",X"FE",X"0A",X"38",X"02",X"3E",X"09",X"47",X"07",X"4F",X"07",X"07",X"81",X"4F",X"18",
		X"13",X"01",X"1E",X"03",X"ED",X"5F",X"E6",X"03",X"28",X"0A",X"01",X"28",X"04",X"FE",X"01",X"28",
		X"03",X"01",X"32",X"05",X"E1",X"23",X"70",X"CD",X"6E",X"11",X"36",X"00",X"CD",X"D9",X"0A",X"36",
		X"00",X"78",X"32",X"13",X"40",X"2A",X"00",X"41",X"22",X"11",X"40",X"C3",X"6C",X"2C",X"36",X"5E",
		X"CD",X"D9",X"0A",X"36",X"5E",X"C9",X"7C",X"FE",X"C7",X"38",X"0E",X"FE",X"D8",X"30",X"0A",X"3A",
		X"0C",X"41",X"A7",X"C8",X"FE",X"05",X"D0",X"18",X"03",X"37",X"C9",X"00",X"E5",X"11",X"EA",X"08",
		X"19",X"11",X"0A",X"00",X"06",X"03",X"E5",X"D5",X"C5",X"CD",X"64",X"08",X"7E",X"C1",X"D1",X"FE",
		X"94",X"38",X"05",X"FE",X"A0",X"DA",X"1F",X"15",X"CD",X"77",X"93",X"CA",X"16",X"15",X"E1",X"19",
		X"10",X"E4",X"E1",X"A7",X"C9",X"00",X"F1",X"C1",X"F1",X"C5",X"16",X"00",X"C3",X"74",X"02",X"3A",
		X"07",X"41",X"47",X"E6",X"01",X"3C",X"07",X"A0",X"00",X"00",X"3E",X"01",X"32",X"14",X"40",X"E1",
		X"E1",X"A7",X"C9",X"3E",X"02",X"32",X"0C",X"41",X"2A",X"02",X"41",X"22",X"09",X"41",X"7D",X"32",
		X"4C",X"50",X"3E",X"2F",X"32",X"49",X"50",X"3D",X"32",X"4D",X"50",X"3E",X"04",X"CD",X"2E",X"18",
		X"ED",X"5F",X"E6",X"03",X"32",X"0B",X"41",X"3E",X"3E",X"32",X"41",X"50",X"3C",X"32",X"45",X"50",
		X"3E",X"C7",X"32",X"4F",X"50",X"CD",X"5D",X"19",X"E1",X"E1",X"A7",X"C9",X"3A",X"0C",X"41",X"FE",
		X"02",X"C8",X"C3",X"46",X"0E",X"61",X"67",X"6E",X"6D",X"69",X"60",X"6B",X"1A",X"66",X"60",X"6B",
		X"65",X"67",X"6E",X"6A",X"5E",X"01",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7E",X"D6",X"A6",X"D8",X"FE",X"12",X"3F",X"C9",X"A7",X"A9",X"AB",
		X"AD",X"AF",X"B1",X"B3",X"B5",X"B7",X"CB",X"67",X"20",X"0B",X"E6",X"0F",X"C6",X"9D",X"4F",X"06",
		X"15",X"D5",X"C3",X"E0",X"0C",X"E6",X"0F",X"07",X"C6",X"A7",X"4F",X"C3",X"AC",X"9C",X"FE",X"14",
		X"D2",X"00",X"00",X"01",X"34",X"50",X"0A",X"E6",X"07",X"C0",X"21",X"3A",X"48",X"CD",X"CB",X"0A",
		X"E5",X"CD",X"40",X"2E",X"4E",X"7D",X"FE",X"50",X"28",X"1F",X"FE",X"F2",X"28",X"27",X"FE",X"0E",
		X"20",X"31",X"7C",X"FE",X"20",X"20",X"2C",X"3E",X"14",X"32",X"15",X"41",X"E1",X"3E",X"03",X"32",
		X"0C",X"41",X"21",X"01",X"20",X"C3",X"C5",X"87",X"00",X"3A",X"15",X"41",X"FE",X"0E",X"28",X"0F",
		X"21",X"25",X"07",X"18",X"0A",X"3A",X"15",X"41",X"FE",X"12",X"18",X"03",X"21",X"50",X"07",X"3C",
		X"32",X"15",X"41",X"23",X"CB",X"79",X"28",X"02",X"56",X"23",X"7C",X"FE",X"08",X"20",X"03",X"21",
		X"00",X"20",X"22",X"00",X"41",X"79",X"E1",X"E6",X"0F",X"28",X"06",X"47",X"36",X"C0",X"2B",X"10",
		X"FB",X"79",X"E6",X"70",X"28",X"13",X"0F",X"0F",X"0F",X"0F",X"C6",X"C0",X"77",X"FE",X"C5",X"28",
		X"04",X"FE",X"C7",X"20",X"03",X"3D",X"2B",X"77",X"2B",X"CB",X"79",X"C8",X"7A",X"11",X"20",X"00",
		X"CB",X"7F",X"20",X"04",X"CD",X"A6",X"15",X"C9",X"FE",X"8F",X"20",X"03",X"2B",X"18",X"09",X"FE",
		X"81",X"30",X"03",X"23",X"18",X"02",X"20",X"04",X"22",X"02",X"40",X"C9",X"FE",X"83",X"30",X"04",
		X"22",X"0A",X"40",X"C9",X"20",X"04",X"22",X"15",X"40",X"C9",X"FE",X"85",X"30",X"04",X"C3",X"EE",
		X"17",X"00",X"D6",X"88",X"38",X"07",X"01",X"FF",X"4B",X"C5",X"C3",X"48",X"13",X"01",X"0E",X"03",
		X"FE",X"FD",X"28",X"0A",X"01",X"00",X"11",X"FE",X"FE",X"28",X"03",X"01",X"02",X"0F",X"21",X"35",
		X"50",X"36",X"01",X"2B",X"2B",X"10",X"FA",X"79",X"A7",X"C8",X"36",X"07",X"2B",X"2B",X"3D",X"18",
		X"F7",X"01",X"34",X"50",X"0A",X"E6",X"07",X"FE",X"03",X"C0",X"2A",X"15",X"40",X"CD",X"13",X"11",
		X"20",X"05",X"AF",X"32",X"16",X"40",X"C9",X"2A",X"15",X"40",X"7C",X"A7",X"C8",X"0A",X"0E",X"23",
		X"E6",X"40",X"28",X"0E",X"CD",X"01",X"11",X"CD",X"6E",X"11",X"36",X"5E",X"CD",X"D9",X"0A",X"36",
		X"5E",X"C9",X"0E",X"B5",X"11",X"20",X"00",X"CD",X"AB",X"13",X"C9",X"2B",X"2B",X"CD",X"6E",X"11",
		X"00",X"00",X"00",X"C3",X"D9",X"0A",X"CD",X"EB",X"16",X"01",X"5E",X"05",X"71",X"2B",X"71",X"23",
		X"19",X"10",X"F9",X"C9",X"21",X"19",X"40",X"D9",X"2A",X"17",X"40",X"7C",X"A7",X"C8",X"01",X"34",
		X"50",X"E5",X"CD",X"13",X"11",X"E1",X"20",X"05",X"D9",X"2B",X"36",X"00",X"C9",X"3A",X"00",X"42",
		X"E6",X"03",X"FE",X"03",X"C0",X"11",X"20",X"00",X"D9",X"7E",X"34",X"D9",X"47",X"FE",X"0C",X"30",
		X"40",X"E6",X"03",X"28",X"1C",X"3D",X"28",X"11",X"3D",X"20",X"28",X"36",X"E3",X"00",X"00",X"00",
		X"CD",X"6E",X"11",X"36",X"E3",X"00",X"00",X"00",X"C9",X"36",X"E1",X"CD",X"6E",X"11",X"36",X"E1",
		X"C9",X"06",X"02",X"C3",X"10",X"2C",X"71",X"2B",X"10",X"FC",X"CD",X"6E",X"11",X"C1",X"23",X"71",
		X"10",X"FC",X"C9",X"36",X"E2",X"2B",X"36",X"E3",X"CD",X"6E",X"11",X"36",X"E3",X"23",X"36",X"E2",
		X"C9",X"3A",X"15",X"41",X"FE",X"0D",X"28",X"04",X"FE",X"10",X"20",X"13",X"78",X"FE",X"0D",X"38",
		X"0B",X"28",X"08",X"06",X"04",X"D9",X"36",X"00",X"D9",X"18",X"C8",X"2B",X"C3",X"EB",X"97",X"FE",
		X"0E",X"28",X"18",X"FE",X"11",X"28",X"14",X"78",X"FE",X"0D",X"38",X"F0",X"28",X"ED",X"FE",X"0E",
		X"28",X"17",X"E5",X"2B",X"2B",X"CD",X"2F",X"2C",X"E1",X"18",X"D8",X"78",X"FE",X"0D",X"38",X"0B",
		X"E5",X"CD",X"2F",X"2C",X"E1",X"06",X"02",X"18",X"CC",X"2B",X"2B",X"CD",X"EB",X"16",X"CD",X"E2",
		X"97",X"71",X"2B",X"00",X"71",X"23",X"0C",X"19",X"10",X"F7",X"C9",X"3A",X"15",X"41",X"FE",X"0E",
		X"38",X"0F",X"FE",X"15",X"30",X"0B",X"3A",X"12",X"50",X"47",X"CD",X"54",X"08",X"00",X"CA",X"EA",
		X"11",X"C3",X"E4",X"11",X"21",X"1C",X"40",X"D9",X"2A",X"1A",X"40",X"C3",X"0B",X"17",X"3A",X"18",
		X"40",X"A7",X"20",X"04",X"22",X"17",X"40",X"C9",X"22",X"1A",X"40",X"C9",X"00",X"00",X"00",X"00",
		X"11",X"D9",X"B8",X"20",X"03",X"F6",X"01",X"C9",X"D9",X"E6",X"7F",X"FE",X"02",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"4A",
		X"50",X"32",X"4E",X"50",X"C9",X"00",X"39",X"07",X"40",X"00",X"39",X"07",X"40",X"00",X"39",X"07",
		X"54",X"01",X"20",X"04",X"44",X"F1",X"21",X"04",X"44",X"01",X"22",X"04",X"54",X"F1",X"23",X"04",
		X"54",X"3A",X"55",X"50",X"D6",X"0A",X"FE",X"02",X"D0",X"3A",X"15",X"41",X"FE",X"0A",X"30",X"06",
		X"CD",X"2C",X"11",X"C3",X"43",X"12",X"2A",X"00",X"41",X"11",X"06",X"07",X"ED",X"52",X"38",X"F0",
		X"3A",X"54",X"50",X"FE",X"F1",X"38",X"F6",X"3E",X"01",X"32",X"04",X"60",X"32",X"18",X"41",X"21",
		X"35",X"18",X"01",X"0C",X"00",X"11",X"50",X"50",X"ED",X"B0",X"32",X"17",X"41",X"C9",X"DA",X"8D",
		X"09",X"FE",X"2C",X"30",X"0A",X"3E",X"2C",X"01",X"10",X"00",X"21",X"41",X"18",X"18",X"E4",X"FE",
		X"2E",X"38",X"03",X"C9",X"00",X"00",X"21",X"50",X"50",X"7E",X"06",X"04",X"FE",X"FF",X"20",X"09",
		X"21",X"17",X"41",X"34",X"21",X"5C",X"50",X"18",X"39",X"3A",X"00",X"42",X"0F",X"D0",X"34",X"23",
		X"23",X"23",X"23",X"10",X"F9",X"2B",X"11",X"0E",X"41",X"1A",X"07",X"07",X"4F",X"12",X"30",X"0C",
		X"13",X"1A",X"3C",X"FE",X"8D",X"20",X"02",X"3E",X"60",X"12",X"18",X"02",X"13",X"1A",X"5F",X"16",
		X"09",X"06",X"04",X"1A",X"A1",X"28",X"0B",X"E6",X"AA",X"C8",X"35",X"2B",X"2B",X"2B",X"2B",X"10",
		X"F9",X"C9",X"34",X"2B",X"2B",X"2B",X"2B",X"10",X"F9",X"C9",X"3A",X"17",X"41",X"3C",X"32",X"17",
		X"41",X"FE",X"20",X"D0",X"ED",X"5F",X"0F",X"0F",X"FE",X"40",X"C9",X"21",X"02",X"60",X"AF",X"06",
		X"05",X"77",X"23",X"10",X"FC",X"C3",X"E1",X"0A",X"3A",X"15",X"41",X"FE",X"0D",X"DA",X"27",X"02",
		X"7E",X"FE",X"C1",X"C8",X"37",X"C9",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"0F",X"14",X"19",
		X"1E",X"28",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"56",X"0D",X"AF",X"32",X"40",X"40",X"32",X"00",X"40",X"3E",X"F2",X"32",X"24",X"41",X"C9",
		X"3E",X"F2",X"32",X"4C",X"50",X"18",X"E9",X"CD",X"43",X"19",X"C3",X"A2",X"08",X"32",X"4B",X"50",
		X"C3",X"43",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"3F",X"97",X"06",X"1B",
		X"35",X"2B",X"2B",X"10",X"FB",X"01",X"3A",X"50",X"0A",X"E6",X"07",X"FE",X"07",X"C0",X"21",X"3D",
		X"48",X"CD",X"CB",X"0A",X"06",X"1B",X"36",X"5E",X"2B",X"10",X"FB",X"21",X"00",X"41",X"34",X"7E",
		X"C6",X"1D",X"32",X"1F",X"40",X"21",X"23",X"48",X"22",X"1D",X"40",X"21",X"0B",X"08",X"D9",X"21",
		X"11",X"20",X"D9",X"46",X"23",X"56",X"23",X"4E",X"23",X"7D",X"FE",X"1E",X"28",X"54",X"7E",X"23",
		X"D9",X"47",X"3A",X"01",X"41",X"4F",X"79",X"37",X"9E",X"30",X"04",X"C6",X"1B",X"38",X"07",X"23",
		X"23",X"23",X"10",X"F2",X"18",X"DC",X"08",X"2B",X"3A",X"1F",X"40",X"96",X"23",X"23",X"28",X"25",
		X"38",X"EE",X"3C",X"BE",X"28",X"06",X"30",X"E8",X"D9",X"5A",X"18",X"02",X"D9",X"59",X"D9",X"C5",
		X"E5",X"01",X"3A",X"50",X"2A",X"1D",X"40",X"CD",X"CB",X"0A",X"08",X"85",X"6F",X"D9",X"7B",X"D9",
		X"77",X"E1",X"C1",X"18",X"CB",X"7E",X"D9",X"3D",X"20",X"05",X"79",X"FE",X"85",X"28",X"DE",X"58",
		X"18",X"DC",X"3A",X"1D",X"40",X"C6",X"1A",X"32",X"1D",X"40",X"D9",X"2B",X"06",X"20",X"3A",X"1F",
		X"40",X"BE",X"28",X"06",X"23",X"23",X"23",X"10",X"F8",X"C9",X"23",X"3A",X"01",X"41",X"96",X"23",
		X"38",X"25",X"96",X"30",X"1D",X"2F",X"FE",X"1B",X"38",X"02",X"3E",X"1A",X"3C",X"08",X"E5",X"2A",
		X"1D",X"40",X"C5",X"01",X"3A",X"50",X"CD",X"CB",X"0A",X"08",X"47",X"36",X"E0",X"2B",X"10",X"FB",
		X"C1",X"E1",X"3A",X"1F",X"40",X"18",X"CF",X"2F",X"FE",X"1A",X"30",X"F6",X"3C",X"5F",X"3E",X"1B",
		X"93",X"BE",X"38",X"01",X"7E",X"08",X"E5",X"2A",X"1D",X"40",X"7D",X"93",X"6F",X"18",X"D3",X"00",
		X"CD",X"43",X"97",X"06",X"1B",X"34",X"2B",X"2B",X"10",X"FB",X"01",X"3A",X"50",X"0A",X"E6",X"07",
		X"C0",X"21",X"DD",X"4B",X"CD",X"CB",X"0A",X"06",X"1B",X"36",X"5E",X"2B",X"10",X"FB",X"21",X"00",
		X"41",X"35",X"7E",X"32",X"1F",X"40",X"21",X"C3",X"4B",X"22",X"1D",X"40",X"C3",X"9B",X"19",X"CD",
		X"31",X"1F",X"3E",X"01",X"32",X"02",X"60",X"21",X"07",X"50",X"06",X"1B",X"36",X"04",X"23",X"23",
		X"10",X"FA",X"C9",X"3A",X"21",X"40",X"A7",X"C8",X"AF",X"32",X"21",X"40",X"3A",X"07",X"41",X"0F",
		X"3A",X"00",X"68",X"D8",X"3A",X"00",X"60",X"C9",X"3A",X"00",X"41",X"FE",X"3C",X"30",X"0B",X"3A",
		X"20",X"40",X"D6",X"03",X"28",X"04",X"AF",X"32",X"20",X"40",X"3A",X"22",X"40",X"A7",X"28",X"06",
		X"CD",X"60",X"29",X"C3",X"00",X"28",X"3A",X"03",X"41",X"FE",X"2F",X"38",X"14",X"FE",X"CF",X"38",
		X"1C",X"47",X"3A",X"01",X"41",X"A7",X"28",X"15",X"3E",X"C8",X"32",X"03",X"41",X"3E",X"01",X"18",
		X"07",X"C6",X"08",X"32",X"03",X"41",X"3E",X"80",X"32",X"22",X"40",X"18",X"D3",X"21",X"20",X"40",
		X"7E",X"A7",X"28",X"13",X"3D",X"28",X"27",X"CD",X"A3",X"1A",X"CB",X"57",X"18",X"03",X"CB",X"5F",
		X"C8",X"3E",X"02",X"32",X"20",X"40",X"C9",X"3A",X"00",X"41",X"FE",X"91",X"38",X"03",X"36",X"02",
		X"C9",X"CD",X"6B",X"19",X"CD",X"D2",X"1B",X"CD",X"A3",X"1A",X"3E",X"02",X"18",X"E5",X"3A",X"00",
		X"41",X"FE",X"3D",X"30",X"03",X"36",X"02",X"C9",X"CD",X"60",X"1A",X"CD",X"F5",X"29",X"CD",X"A3",
		X"1A",X"E6",X"08",X"18",X"E5",X"3A",X"22",X"40",X"A7",X"C0",X"3A",X"19",X"41",X"26",X"44",X"FE",
		X"42",X"20",X"02",X"3E",X"00",X"3C",X"3C",X"6F",X"32",X"19",X"41",X"7E",X"A7",X"C8",X"34",X"FE",
		X"02",X"28",X"10",X"FE",X"18",X"D8",X"36",X"00",X"06",X"7F",X"7D",X"FE",X"87",X"18",X"06",X"06",
		X"F7",X"18",X"02",X"06",X"BB",X"26",X"22",X"5E",X"23",X"56",X"2A",X"00",X"41",X"EB",X"CD",X"26",
		X"9B",X"24",X"05",X"CD",X"26",X"9B",X"2C",X"05",X"05",X"CD",X"26",X"9B",X"25",X"04",X"CD",X"26",
		X"9B",X"2C",X"06",X"5E",X"CD",X"26",X"9B",X"C9",X"06",X"80",X"C5",X"CD",X"3A",X"31",X"2A",X"02",
		X"41",X"2D",X"CD",X"B1",X"02",X"06",X"01",X"CD",X"56",X"0D",X"C1",X"10",X"ED",X"CD",X"28",X"87",
		X"06",X"30",X"CD",X"56",X"0D",X"C3",X"18",X"03",X"CD",X"56",X"0D",X"C3",X"E5",X"2A",X"3A",X"1A",
		X"41",X"FE",X"4F",X"DA",X"96",X"2B",X"C3",X"57",X"8C",X"35",X"55",X"6B",X"8F",X"AA",X"D6",X"FE",
		X"00",X"00",X"01",X"3A",X"50",X"0A",X"E6",X"07",X"FE",X"01",X"C0",X"3A",X"00",X"41",X"C6",X"1D",
		X"32",X"1F",X"40",X"21",X"3D",X"48",X"22",X"1D",X"40",X"01",X"F5",X"F4",X"11",X"F7",X"F6",X"D9",
		X"21",X"D0",X"21",X"06",X"08",X"3A",X"1F",X"40",X"4F",X"79",X"96",X"28",X"27",X"3D",X"CA",X"78",
		X"1C",X"23",X"23",X"10",X"F4",X"D9",X"78",X"FE",X"F4",X"20",X"0B",X"01",X"AD",X"AC",X"11",X"AF",
		X"AE",X"D9",X"06",X"11",X"18",X"E3",X"FE",X"AC",X"C0",X"01",X"7D",X"7C",X"11",X"7F",X"7E",X"D9",
		X"06",X"21",X"18",X"D5",X"23",X"3A",X"01",X"41",X"37",X"9E",X"38",X"1D",X"20",X"D4",X"C5",X"E5",
		X"26",X"44",X"2B",X"7E",X"A7",X"20",X"0B",X"CD",X"0D",X"2A",X"D9",X"7A",X"D9",X"77",X"E1",X"C1",
		X"18",X"C0",X"CD",X"0D",X"2A",X"36",X"BA",X"18",X"F5",X"FE",X"E5",X"38",X"B5",X"C5",X"E5",X"47",
		X"26",X"44",X"2B",X"7E",X"A7",X"78",X"20",X"11",X"CD",X"16",X"2A",X"D9",X"7B",X"D9",X"77",X"2B",
		X"7D",X"E6",X"1F",X"FE",X"02",X"20",X"D3",X"18",X"D5",X"CD",X"16",X"2A",X"36",X"BB",X"2B",X"7D",
		X"E6",X"1F",X"FE",X"02",X"20",X"CF",X"18",X"C6",X"23",X"3A",X"01",X"41",X"37",X"9E",X"38",X"19",
		X"20",X"BE",X"C5",X"E5",X"26",X"44",X"2B",X"7E",X"A7",X"20",X"07",X"CD",X"0D",X"2A",X"D9",X"78",
		X"18",X"AA",X"CD",X"0D",X"2A",X"36",X"B8",X"18",X"DD",X"FE",X"E5",X"38",X"A3",X"C5",X"E5",X"47",
		X"26",X"44",X"2B",X"7E",X"A7",X"78",X"20",X"11",X"CD",X"16",X"2A",X"D9",X"79",X"D9",X"77",X"2B",
		X"7D",X"E6",X"1F",X"FE",X"02",X"20",X"D7",X"18",X"BD",X"CD",X"16",X"2A",X"36",X"B9",X"2B",X"7D",
		X"E6",X"1F",X"FE",X"02",X"20",X"CF",X"18",X"AE",X"3A",X"01",X"41",X"32",X"1F",X"40",X"21",X"DD",
		X"4B",X"18",X"0B",X"3A",X"01",X"41",X"C6",X"1A",X"32",X"1F",X"40",X"21",X"C3",X"4B",X"22",X"1D",
		X"40",X"01",X"F5",X"F4",X"11",X"F7",X"F6",X"D9",X"21",X"D1",X"21",X"06",X"08",X"3A",X"1F",X"40",
		X"4F",X"79",X"96",X"28",X"27",X"3D",X"CA",X"76",X"1D",X"23",X"23",X"10",X"F4",X"D9",X"78",X"FE",
		X"F4",X"20",X"0B",X"01",X"AD",X"AC",X"11",X"AF",X"AE",X"D9",X"06",X"11",X"18",X"E3",X"FE",X"AC",
		X"C0",X"01",X"7D",X"7C",X"11",X"7F",X"7E",X"D9",X"06",X"21",X"18",X"D5",X"2B",X"3A",X"00",X"41",
		X"37",X"9E",X"23",X"38",X"1D",X"20",X"D2",X"C5",X"E5",X"26",X"44",X"2B",X"7E",X"A7",X"20",X"0B",
		X"CD",X"0D",X"2A",X"D9",X"79",X"D9",X"77",X"E1",X"C1",X"18",X"BE",X"CD",X"0D",X"2A",X"36",X"B9",
		X"18",X"F5",X"FE",X"E2",X"38",X"B3",X"C5",X"E5",X"F5",X"26",X"44",X"2B",X"7E",X"A7",X"28",X"13",
		X"F1",X"F5",X"CD",X"CB",X"2A",X"D9",X"36",X"BB",X"F1",X"28",X"DC",X"11",X"20",X"00",X"CD",X"D9",
		X"0A",X"18",X"DB",X"F1",X"F5",X"CD",X"CB",X"2A",X"7B",X"D9",X"77",X"F1",X"28",X"C9",X"11",X"20",
		X"00",X"CD",X"D9",X"0A",X"18",X"BD",X"2B",X"3A",X"00",X"41",X"37",X"9E",X"23",X"38",X"19",X"20",
		X"B8",X"C5",X"E5",X"26",X"44",X"2B",X"7E",X"A7",X"20",X"07",X"CD",X"0D",X"2A",X"D9",X"78",X"18",
		X"A4",X"CD",X"0D",X"2A",X"36",X"B8",X"18",X"9F",X"FE",X"E2",X"38",X"9D",X"C5",X"E5",X"F5",X"26",
		X"44",X"2B",X"7E",X"A7",X"28",X"13",X"F1",X"F5",X"CD",X"CB",X"2A",X"D9",X"36",X"BA",X"F1",X"28",
		X"86",X"11",X"20",X"00",X"CD",X"D9",X"0A",X"18",X"DB",X"F1",X"F5",X"CD",X"CB",X"2A",X"7A",X"D9",
		X"77",X"F1",X"28",X"D2",X"11",X"20",X"00",X"CD",X"D9",X"0A",X"18",X"C1",X"DD",X"7E",X"00",X"FE",
		X"F8",X"D2",X"47",X"1E",X"6F",X"DD",X"7E",X"03",X"FE",X"E7",X"38",X"05",X"DD",X"36",X"00",X"FF",
		X"C9",X"67",X"E5",X"11",X"F8",X"06",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"E0",X"FD",X"7E",X"02",
		X"20",X"03",X"07",X"07",X"07",X"E1",X"4F",X"E6",X"E0",X"28",X"02",X"2C",X"2C",X"79",X"E6",X"0E",
		X"28",X"02",X"2D",X"2D",X"79",X"E6",X"83",X"28",X"02",X"24",X"24",X"79",X"E6",X"38",X"28",X"02",
		X"25",X"25",X"FD",X"7E",X"01",X"5F",X"16",X"2A",X"1A",X"57",X"FD",X"7E",X"00",X"47",X"07",X"07",
		X"FD",X"77",X"00",X"30",X"08",X"1C",X"7B",X"FE",X"93",X"20",X"02",X"1E",X"81",X"78",X"A2",X"28",
		X"09",X"E6",X"AA",X"79",X"20",X"02",X"0F",X"0F",X"07",X"4F",X"DD",X"74",X"03",X"DD",X"75",X"00",
		X"FD",X"73",X"01",X"FD",X"71",X"02",X"C9",X"21",X"9D",X"40",X"3A",X"00",X"42",X"E6",X"06",X"C0",
		X"7E",X"3C",X"28",X"01",X"77",X"06",X"03",X"FE",X"31",X"38",X"06",X"06",X"01",X"FE",X"61",X"30",
		X"02",X"A0",X"C0",X"3A",X"54",X"41",X"3C",X"3C",X"20",X"02",X"3E",X"E0",X"32",X"54",X"41",X"6F",
		X"26",X"21",X"5E",X"23",X"56",X"2A",X"00",X"41",X"7A",X"94",X"FE",X"1A",X"D0",X"4F",X"7B",X"95",
		X"FE",X"1D",X"D0",X"07",X"07",X"07",X"C6",X"0F",X"DD",X"77",X"00",X"3E",X"1A",X"91",X"07",X"07",
		X"07",X"C6",X"0F",X"DD",X"77",X"03",X"3E",X"60",X"32",X"6A",X"40",X"C9",X"00",X"00",X"00",X"00",
		X"21",X"58",X"50",X"11",X"A0",X"40",X"3A",X"00",X"42",X"4F",X"A7",X"08",X"1A",X"FE",X"09",X"30",
		X"1E",X"7E",X"FE",X"F8",X"30",X"2E",X"34",X"CB",X"71",X"20",X"02",X"35",X"35",X"2E",X"5B",X"79",
		X"E6",X"03",X"20",X"01",X"35",X"7E",X"FE",X"E7",X"D8",X"3E",X"FF",X"32",X"58",X"50",X"C9",X"7E",
		X"FE",X"F8",X"30",X"2E",X"CB",X"69",X"20",X"04",X"35",X"35",X"18",X"02",X"34",X"34",X"2E",X"5B",
		X"CB",X"41",X"18",X"DE",X"08",X"20",X"18",X"3A",X"01",X"42",X"E6",X"03",X"C0",X"1A",X"3C",X"12",
		X"3A",X"40",X"50",X"C6",X"18",X"77",X"3E",X"E6",X"32",X"5B",X"50",X"32",X"43",X"40",X"C9",X"AF",
		X"18",X"F9",X"08",X"20",X"FA",X"3A",X"01",X"42",X"0F",X"D8",X"18",X"E4",X"CD",X"3C",X"0E",X"05",
		X"C2",X"D2",X"8C",X"C3",X"E0",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"02",X"44",X"06",X"42",X"36",X"00",X"23",X"10",X"FB",X"C9",X"00",
		X"00",X"22",X"00",X"41",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"50",X"6F",X"26",X"41",X"7E",X"D6",
		X"01",X"D8",X"3E",X"05",X"32",X"A0",X"40",X"3E",X"80",X"32",X"9D",X"40",X"C9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"04",X"C5",X"3A",X"1E",
		X"41",X"FE",X"A1",X"20",X"02",X"3E",X"85",X"3C",X"32",X"1E",X"41",X"6F",X"26",X"2D",X"5E",X"16",
		X"03",X"2A",X"00",X"41",X"EB",X"3A",X"00",X"42",X"E6",X"06",X"07",X"C6",X"A2",X"4F",X"06",X"2D",
		X"C5",X"DD",X"E1",X"0E",X"03",X"DD",X"46",X"00",X"C5",X"CD",X"98",X"1B",X"C1",X"DD",X"23",X"24",
		X"0D",X"20",X"F2",X"C1",X"10",X"C7",X"C9",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"50",X"6F",X"26",
		X"41",X"7E",X"06",X"E0",X"A7",X"28",X"07",X"06",X"60",X"3D",X"28",X"02",X"06",X"20",X"3A",X"00",
		X"42",X"A0",X"C0",X"C3",X"BE",X"3F",X"CD",X"3B",X"0A",X"3E",X"08",X"32",X"07",X"41",X"3E",X"FF",
		X"32",X"00",X"78",X"AF",X"32",X"03",X"68",X"32",X"00",X"60",X"C3",X"58",X"9C",X"00",X"A7",X"C2",
		X"91",X"80",X"3A",X"15",X"41",X"FE",X"14",X"C2",X"B0",X"3B",X"C3",X"21",X"3C",X"32",X"A1",X"40",
		X"0E",X"5A",X"CD",X"00",X"0E",X"AF",X"32",X"62",X"40",X"C3",X"58",X"99",X"00",X"00",X"00",X"00",
		X"00",X"ED",X"A8",X"04",X"AF",X"FD",X"28",X"04",X"AF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"52",X"54",X"56",X"58",X"5A",X"5C",X"7C",X"7A",X"78",X"76",X"74",X"72",X"70",X"98",X"00",
		X"1F",X"22",X"21",X"1F",X"21",X"25",X"1F",X"20",X"21",X"43",X"1D",X"05",X"47",X"19",X"05",X"4B",
		X"15",X"09",X"53",X"11",X"09",X"5B",X"0D",X"09",X"63",X"07",X"0A",X"3D",X"02",X"71",X"3D",X"01",
		X"71",X"3D",X"00",X"71",X"26",X"2B",X"26",X"27",X"2A",X"2E",X"28",X"29",X"18",X"54",X"22",X"09",
		X"5C",X"1E",X"09",X"64",X"1A",X"09",X"73",X"1A",X"08",X"7A",X"16",X"09",X"82",X"12",X"08",X"7C",
		X"0D",X"04",X"8A",X"0A",X"06",X"90",X"0F",X"04",X"98",X"0B",X"04",X"A0",X"0A",X"04",X"98",X"13",
		X"08",X"A6",X"0F",X"05",X"8C",X"1B",X"08",X"84",X"22",X"08",X"8C",X"2A",X"08",X"7C",X"2A",X"08",
		X"84",X"32",X"08",X"7C",X"39",X"08",X"54",X"32",X"04",X"58",X"39",X"04",X"60",X"39",X"04",X"68",
		X"3E",X"05",X"5C",X"40",X"04",X"62",X"45",X"04",X"68",X"4A",X"05",X"74",X"4A",X"04",X"68",X"26",
		X"05",X"68",X"35",X"05",X"64",X"31",X"05",X"5C",X"2D",X"09",X"5C",X"2A",X"0D",X"73",X"26",X"09",
		X"73",X"41",X"09",X"94",X"22",X"09",X"9C",X"1E",X"09",X"A4",X"1A",X"07",X"4B",X"3E",X"09",X"53",
		X"46",X"0A",X"A7",X"22",X"07",X"63",X"51",X"05",X"62",X"50",X"05",X"61",X"4F",X"05",X"60",X"4E",
		X"05",X"5F",X"4D",X"05",X"5E",X"4C",X"05",X"5D",X"4B",X"05",X"5C",X"4A",X"05",X"5B",X"49",X"05",
		X"5A",X"48",X"05",X"59",X"47",X"05",X"78",X"51",X"05",X"79",X"50",X"05",X"7A",X"4F",X"05",X"7B",
		X"4E",X"05",X"7C",X"4D",X"05",X"7D",X"4C",X"05",X"7E",X"4B",X"05",X"7F",X"4A",X"05",X"80",X"49",
		X"05",X"81",X"48",X"05",X"82",X"47",X"05",X"83",X"46",X"05",X"84",X"45",X"05",X"85",X"44",X"05",
		X"86",X"43",X"05",X"87",X"42",X"05",X"88",X"41",X"05",X"89",X"40",X"05",X"8A",X"3F",X"05",X"8B",
		X"3E",X"05",X"8C",X"3D",X"05",X"8D",X"3C",X"05",X"8E",X"3B",X"05",X"8F",X"3A",X"05",X"90",X"39",
		X"05",X"91",X"38",X"05",X"92",X"37",X"05",X"93",X"36",X"05",X"94",X"35",X"05",X"95",X"34",X"05",
		X"96",X"33",X"05",X"97",X"32",X"05",X"98",X"31",X"05",X"99",X"30",X"05",X"9A",X"2F",X"05",X"9B",
		X"2E",X"05",X"9C",X"2D",X"05",X"9D",X"2C",X"05",X"9E",X"2B",X"05",X"9F",X"2A",X"05",X"A0",X"29",
		X"05",X"A1",X"28",X"05",X"A2",X"27",X"05",X"A3",X"26",X"05",X"A4",X"25",X"05",X"A5",X"24",X"05",
		X"A6",X"23",X"05",X"6D",X"02",X"06",X"26",X"2C",X"20",X"3D",X"03",X"1D",X"3E",X"03",X"1D",X"3F",
		X"03",X"1D",X"AB",X"03",X"1F",X"AC",X"03",X"1F",X"AD",X"03",X"1F",X"43",X"1E",X"03",X"47",X"1A",
		X"03",X"4B",X"16",X"03",X"53",X"12",X"03",X"5B",X"0E",X"03",X"63",X"08",X"05",X"6C",X"03",X"04",
		X"54",X"23",X"07",X"5C",X"1F",X"03",X"64",X"1B",X"03",X"7A",X"17",X"03",X"82",X"13",X"03",X"5C",
		X"2B",X"02",X"64",X"2E",X"03",X"68",X"32",X"03",X"68",X"27",X"03",X"6C",X"27",X"0E",X"73",X"27",
		X"1A",X"7B",X"27",X"1A",X"94",X"23",X"13",X"9C",X"1F",X"03",X"A4",X"1B",X"03",X"53",X"3F",X"07",
		X"4B",X"2C",X"12",X"27",X"2C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"52",X"6A",X"52",X"6C",X"52",X"6E",X"52",X"70",X"52",X"72",X"52",X"74",X"52",X"76",X"52",
		X"59",X"20",X"6B",X"18",X"80",X"12",X"98",X"11",X"87",X"20",X"73",X"24",X"5A",X"2C",X"7C",X"34",
		X"92",X"34",X"5C",X"3E",X"6B",X"48",X"73",X"42",X"84",X"42",X"48",X"28",X"9C",X"1B",X"A9",X"03",
		X"40",X"28",X"32",X"23",X"3C",X"23",X"42",X"22",X"46",X"1E",X"4A",X"1A",X"50",X"16",X"58",X"12",
		X"66",X"08",X"6A",X"08",X"76",X"03",X"84",X"03",X"94",X"03",X"9B",X"03",X"A4",X"03",X"7C",X"0E",
		X"8E",X"0B",X"91",X"10",X"98",X"0C",X"A6",X"10",X"9C",X"14",X"87",X"13",X"80",X"17",X"59",X"23",
		X"51",X"2B",X"60",X"2E",X"54",X"33",X"68",X"36",X"86",X"33",X"78",X"42",X"64",X"46",X"69",X"4B",
		X"75",X"4B",X"81",X"2B",X"54",X"1F",X"06",X"54",X"29",X"06",X"7E",X"29",X"07",X"95",X"29",X"05",
		X"4F",X"32",X"06",X"87",X"32",X"0A",X"56",X"3A",X"06",X"80",X"3A",X"06",X"78",X"4A",X"0A",X"A4",
		X"26",X"04",X"A4",X"26",X"04",X"A4",X"27",X"03",X"A4",X"28",X"02",X"A4",X"29",X"01",X"9B",X"2F",
		X"04",X"9B",X"30",X"03",X"9B",X"31",X"02",X"9B",X"32",X"01",X"90",X"3A",X"04",X"90",X"3B",X"03",
		X"90",X"3C",X"02",X"90",X"3D",X"01",X"87",X"43",X"04",X"87",X"44",X"03",X"87",X"45",X"02",X"87",
		X"46",X"01",X"7C",X"4E",X"04",X"7C",X"4F",X"03",X"7C",X"50",X"02",X"7C",X"51",X"01",X"A6",X"23",
		X"05",X"A5",X"24",X"05",X"A4",X"25",X"05",X"9B",X"2E",X"05",X"92",X"37",X"05",X"91",X"38",X"05",
		X"90",X"39",X"05",X"87",X"42",X"05",X"7D",X"4C",X"05",X"7C",X"4D",X"05",X"AA",X"1F",X"01",X"A9",
		X"20",X"02",X"A8",X"21",X"03",X"A7",X"22",X"04",X"9F",X"2A",X"01",X"9E",X"2B",X"02",X"9D",X"2C",
		X"03",X"9C",X"2D",X"04",X"96",X"33",X"01",X"95",X"34",X"02",X"94",X"35",X"03",X"93",X"36",X"04",
		X"8B",X"3E",X"01",X"8A",X"3F",X"02",X"89",X"40",X"03",X"88",X"41",X"04",X"81",X"48",X"01",X"80",
		X"49",X"02",X"7E",X"4B",X"04",X"7E",X"33",X"03",X"65",X"3B",X"03",X"64",X"39",X"03",X"73",X"39",
		X"0D",X"61",X"42",X"0C",X"75",X"42",X"0F",X"48",X"02",X"04",X"54",X"02",X"04",X"60",X"02",X"04",
		X"78",X"02",X"04",X"84",X"02",X"04",X"90",X"02",X"04",X"9C",X"02",X"04",X"6D",X"02",X"06",X"21",
		X"23",X"0B",X"26",X"2C",X"02",X"5D",X"0D",X"02",X"8C",X"0D",X"02",X"5F",X"16",X"02",X"6C",X"16",
		X"03",X"73",X"16",X"03",X"8C",X"16",X"02",X"5F",X"20",X"03",X"6C",X"22",X"04",X"73",X"22",X"04",
		X"8C",X"20",X"03",X"61",X"2A",X"03",X"8C",X"2A",X"03",X"7B",X"33",X"02",X"62",X"3B",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"32",X"23",X"3C",X"23",X"4B",X"0D",X"58",X"0D",X"A3",X"0B",X"48",
		X"16",X"50",X"16",X"7D",X"16",X"A4",X"17",X"9A",X"1B",X"4E",X"20",X"5A",X"20",X"88",X"20",X"4C",
		X"2A",X"5B",X"2A",X"5D",X"33",X"5C",X"3B",X"7C",X"3B",X"64",X"44",X"66",X"4B",X"73",X"4B",X"A0",
		X"2E",X"97",X"37",X"8C",X"42",X"83",X"4C",X"4F",X"03",X"59",X"03",X"67",X"03",X"7E",X"03",X"8A",
		X"03",X"96",X"03",X"A2",X"03",X"65",X"0B",X"78",X"0C",X"84",X"10",X"90",X"0D",X"9C",X"11",X"69",
		X"1D",X"75",X"1D",X"91",X"16",X"98",X"24",X"63",X"2A",X"76",X"2A",X"6A",X"33",X"74",X"33",X"85",
		X"33",X"6B",X"3B",X"71",X"53",X"6D",X"53",X"6E",X"55",X"6F",X"53",X"70",X"55",X"20",X"2F",X"26",
		X"2F",X"5D",X"10",X"8B",X"10",X"8D",X"0D",X"5D",X"16",X"8D",X"16",X"8D",X"20",X"5F",X"2A",X"6B",
		X"44",X"73",X"44",X"6B",X"4B",X"2A",X"2C",X"2E",X"2C",X"32",X"2C",X"36",X"2C",X"3A",X"2C",X"3E",
		X"2E",X"41",X"31",X"1F",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9E",X"0D",X"1E",X"1E",X"1E",X"16",X"96",X"04",X"16",X"16",X"75",X"F3",X"04",X"71",X"60",X"80",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F3",X"E1",X"80",X"F0",X"E2",X"80",X"F0",X"E3",
		X"80",X"F0",X"E4",X"80",X"F2",X"E5",X"80",X"F3",X"56",X"80",X"F0",X"40",X"00",X"00",X"80",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F2",X"30",X"80",X"F0",X"21",X"80",X"F1",X"E2",X"80",X"F0",
		X"E3",X"80",X"F0",X"77",X"80",X"F0",X"68",X"80",X"F0",X"E9",X"80",X"03",X"00",X"00",X"80",X"0A",
		X"00",X"00",X"00",X"80",X"02",X"80",X"03",X"00",X"00",X"80",X"03",X"00",X"00",X"80",X"0A",X"00",
		X"00",X"00",X"00",X"80",X"F3",X"90",X"80",X"F2",X"70",X"80",X"F1",X"50",X"80",X"F2",X"4A",X"80",
		X"F3",X"6B",X"80",X"F0",X"EC",X"80",X"F0",X"ED",X"80",X"F2",X"E4",X"A0",X"F5",X"35",X"A1",X"F0",
		X"20",X"22",X"92",X"01",X"92",X"0B",X"12",X"12",X"12",X"92",X"02",X"32",X"31",X"B0",X"04",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"F2",X"10",X"80",X"F2",X"02",X"80",
		X"F3",X"E3",X"A0",X"F5",X"54",X"A1",X"F0",X"35",X"A2",X"F0",X"20",X"A3",X"F0",X"40",X"93",X"FC",
		X"60",X"13",X"13",X"13",X"24",X"25",X"26",X"96",X"07",X"16",X"75",X"73",X"F1",X"04",X"60",X"80",
		X"01",X"80",X"01",X"80",X"0B",X"00",X"00",X"00",X"80",X"02",X"80",X"06",X"50",X"D2",X"06",X"54",
		X"56",X"97",X"0D",X"17",X"17",X"17",X"76",X"74",X"13",X"93",X"08",X"13",X"13",X"72",X"70",X"80",
		X"02",X"80",X"F3",X"E1",X"80",X"F2",X"E2",X"80",X"F3",X"E3",X"80",X"F2",X"E4",X"D0",X"F0",X"35",
		X"D2",X"F0",X"20",X"54",X"95",X"0C",X"15",X"15",X"15",X"74",X"F2",X"04",X"70",X"00",X"50",X"91",
		X"01",X"91",X"01",X"91",X"01",X"91",X"01",X"91",X"01",X"52",X"13",X"93",X"04",X"13",X"13",X"54",
		X"56",X"97",X"0B",X"17",X"17",X"17",X"97",X"01",X"97",X"01",X"76",X"95",X"09",X"15",X"56",X"58",
		X"99",X"0D",X"19",X"19",X"19",X"78",X"76",X"F4",X"04",X"72",X"91",X"12",X"91",X"21",X"91",X"32",
		X"91",X"41",X"91",X"52",X"91",X"61",X"91",X"72",X"91",X"81",X"D2",X"90",X"93",X"A0",X"93",X"B9",
		X"93",X"C0",X"54",X"56",X"58",X"99",X"0C",X"19",X"19",X"19",X"92",X"0A",X"12",X"12",X"12",X"71",
		X"E0",X"F0",X"E1",X"80",X"F4",X"EE",X"80",X"F0",X"EF",X"80",X"F2",X"E3",X"80",X"F3",X"E4",X"80",
		X"F2",X"35",X"80",X"F3",X"20",X"80",X"02",X"00",X"00",X"00",X"80",X"F3",X"E1",X"80",X"F0",X"E2",
		X"80",X"F0",X"E3",X"80",X"F0",X"E4",X"80",X"F2",X"E5",X"80",X"F3",X"56",X"80",X"F0",X"40",X"00",
		X"00",X"80",X"0A",X"00",X"00",X"00",X"00",X"00",X"80",X"F2",X"30",X"80",X"F0",X"21",X"80",X"F1",
		X"E2",X"80",X"F0",X"E3",X"80",X"F0",X"77",X"80",X"F0",X"68",X"80",X"F0",X"E9",X"80",X"03",X"00",
		X"00",X"80",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"01",X"00",X"90",X"02",X"12",X"14",X"31",X"B1",X"03",X"31",X"04",
		X"04",X"04",X"04",X"06",X"06",X"06",X"06",X"06",X"06",X"02",X"02",X"02",X"02",X"02",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"05",X"05",X"05",X"05",X"05",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"06",X"06",X"06",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"05",X"05",X"06",X"06",X"06",X"00",X"50",X"51",X"B2",X"04",X"32",X"32",
		X"32",X"32",X"33",X"33",X"33",X"33",X"32",X"B2",X"06",X"32",X"32",X"32",X"14",X"16",X"37",X"B7",
		X"05",X"37",X"37",X"37",X"76",X"74",X"33",X"33",X"33",X"33",X"33",X"00",X"80",X"07",X"00",X"00",
		X"00",X"10",X"12",X"35",X"35",X"35",X"35",X"56",X"57",X"18",X"B9",X"07",X"39",X"39",X"39",X"80",
		X"08",X"80",X"09",X"80",X"0A",X"80",X"0B",X"80",X"0C",X"80",X"0D",X"80",X"0E",X"00",X"37",X"B7",
		X"01",X"37",X"37",X"00",X"80",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"5E",X"41",X"7E",X"7E",X"2A",X"55",X"41",X"7E",X"7E",X"C9",X"D3",X"C2",X"E0",X"13",X"2E",
		X"14",X"7E",X"FE",X"4F",X"C8",X"C3",X"E0",X"13",X"3A",X"34",X"50",X"E6",X"07",X"CA",X"66",X"0B",
		X"C3",X"31",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"1D",X"1D",X"2E",X"2E",X"40",X"53",X"AC",X"1D",X"2E",X"2E",X"40",X"53",X"AC",X"1D",X"2E",
		X"2E",X"40",X"53",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3B",X"02",X"3B",X"02",X"3B",X"02",X"FC",X"01",X"FC",X"01",X"01",X"00",X"3B",X"02",X"3B",X"02",
		X"01",X"00",X"FC",X"01",X"FC",X"01",X"01",X"00",X"3B",X"02",X"3B",X"02",X"01",X"00",X"FC",X"01",
		X"FC",X"01",X"01",X"00",X"3B",X"02",X"3B",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"F5",X"0F",X"E6",X"1F",X"C6",X"80",X"4F",X"06",X"26",X"21",X"00",X"58",X"11",X"00",
		X"59",X"AF",X"12",X"0A",X"77",X"3E",X"01",X"12",X"36",X"01",X"3E",X"08",X"12",X"36",X"0F",X"F1",
		X"4F",X"FE",X"BF",X"30",X"0C",X"AF",X"32",X"01",X"60",X"79",X"E6",X"3E",X"C6",X"A0",X"4F",X"18",
		X"10",X"79",X"E6",X"3E",X"C6",X"A0",X"4F",X"0A",X"D6",X"FC",X"28",X"02",X"3E",X"FF",X"3C",X"32",
		X"01",X"60",X"3E",X"02",X"12",X"0A",X"77",X"3E",X"03",X"12",X"03",X"0A",X"77",X"3E",X"0A",X"12",
		X"36",X"00",X"3E",X"09",X"C3",X"3A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"22",X"40",X"0F",X"30",X"3A",X"01",X"3A",X"50",X"21",X"24",X"48",X"CD",X"CB",X"0A",X"3E",
		X"1E",X"06",X"00",X"E5",X"54",X"5D",X"1D",X"0E",X"1A",X"ED",X"B0",X"E1",X"11",X"20",X"00",X"19",
		X"3D",X"20",X"F0",X"01",X"3A",X"50",X"21",X"3D",X"48",X"CD",X"CB",X"0A",X"11",X"20",X"00",X"06",
		X"1E",X"36",X"5E",X"19",X"10",X"FB",X"21",X"01",X"41",X"35",X"3E",X"02",X"C3",X"93",X"2A",X"00",
		X"0F",X"D0",X"AF",X"32",X"22",X"40",X"CD",X"C8",X"1C",X"3A",X"01",X"41",X"32",X"1F",X"40",X"21",
		X"DD",X"4B",X"22",X"1D",X"40",X"21",X"0B",X"08",X"D9",X"21",X"11",X"20",X"D9",X"46",X"23",X"56",
		X"23",X"4E",X"23",X"7D",X"FE",X"1E",X"CA",X"1E",X"29",X"7E",X"23",X"D9",X"47",X"3A",X"1F",X"40",
		X"BE",X"28",X"07",X"23",X"23",X"23",X"10",X"F8",X"18",X"E2",X"2B",X"5E",X"23",X"23",X"4E",X"0D",
		X"08",X"3A",X"00",X"41",X"57",X"7B",X"92",X"38",X"08",X"28",X"43",X"FE",X"1E",X"30",X"05",X"18",
		X"6A",X"81",X"38",X"05",X"3A",X"1F",X"40",X"18",X"DB",X"C5",X"E5",X"28",X"22",X"4F",X"C5",X"2A",
		X"1D",X"40",X"01",X"3A",X"50",X"CD",X"CB",X"0A",X"C1",X"0C",X"06",X"1E",X"11",X"20",X"00",X"0D",
		X"28",X"16",X"D9",X"7A",X"D9",X"77",X"CD",X"3C",X"0E",X"10",X"F4",X"E1",X"C1",X"18",X"D5",X"2A",
		X"1D",X"40",X"01",X"3A",X"50",X"CD",X"CB",X"0A",X"D9",X"79",X"D9",X"77",X"18",X"ED",X"C5",X"E5",
		X"06",X"1E",X"C5",X"2A",X"1D",X"40",X"01",X"3A",X"50",X"CD",X"CB",X"0A",X"D9",X"08",X"20",X"0C",
		X"79",X"FE",X"85",X"78",X"20",X"01",X"79",X"D9",X"77",X"C1",X"18",X"CF",X"78",X"D9",X"77",X"11",
		X"20",X"00",X"CD",X"3C",X"0E",X"C1",X"05",X"28",X"C2",X"18",X"B1",X"C5",X"E5",X"57",X"0F",X"0F",
		X"0F",X"E6",X"E0",X"5F",X"3E",X"1E",X"92",X"47",X"7A",X"0F",X"0F",X"0F",X"E6",X"03",X"57",X"2A",
		X"1D",X"40",X"A7",X"ED",X"52",X"C5",X"01",X"3A",X"50",X"CD",X"CB",X"0A",X"18",X"BE",X"D9",X"2B",
		X"06",X"20",X"3A",X"00",X"41",X"57",X"7E",X"92",X"FE",X"1E",X"30",X"30",X"57",X"23",X"3A",X"1F",
		X"40",X"96",X"38",X"29",X"23",X"BE",X"30",X"20",X"E5",X"C5",X"7A",X"0F",X"0F",X"0F",X"E6",X"E0",
		X"5F",X"7A",X"0F",X"0F",X"0F",X"E6",X"03",X"57",X"2A",X"1D",X"40",X"A7",X"ED",X"52",X"01",X"3A",
		X"50",X"CD",X"CB",X"0A",X"36",X"E0",X"C1",X"E1",X"23",X"10",X"C7",X"C9",X"23",X"23",X"18",X"F8",
		X"3A",X"22",X"40",X"07",X"30",X"3A",X"01",X"3A",X"50",X"21",X"1C",X"48",X"CD",X"CB",X"0A",X"3E",
		X"20",X"06",X"00",X"E5",X"54",X"5D",X"1C",X"0E",X"1A",X"ED",X"B8",X"E1",X"11",X"20",X"00",X"19",
		X"3D",X"20",X"F0",X"01",X"3A",X"50",X"21",X"23",X"48",X"CD",X"CB",X"0A",X"11",X"20",X"00",X"06",
		X"1E",X"36",X"5E",X"19",X"10",X"FB",X"21",X"01",X"41",X"34",X"3E",X"40",X"C3",X"97",X"2A",X"00",
		X"07",X"D0",X"AF",X"32",X"22",X"40",X"CD",X"D3",X"1C",X"3A",X"01",X"41",X"C6",X"1A",X"32",X"1F",
		X"40",X"21",X"C3",X"4B",X"22",X"1D",X"40",X"C3",X"55",X"28",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"3A",X"50",X"0A",X"E6",X"07",X"FE",X"02",X"C0",X"3A",X"00",
		X"41",X"32",X"1F",X"40",X"21",X"DD",X"4B",X"22",X"1D",X"40",X"C3",X"E9",X"1B",X"01",X"3A",X"50",
		X"2A",X"1D",X"40",X"C3",X"CB",X"0A",X"2A",X"1D",X"40",X"85",X"3C",X"6F",X"01",X"3A",X"50",X"CD",
		X"CB",X"0A",X"C9",X"00",X"66",X"2E",X"6D",X"06",X"5E",X"CD",X"26",X"9B",X"2E",X"72",X"CD",X"26",
		X"9B",X"24",X"C9",X"01",X"06",X"5E",X"C5",X"CD",X"26",X"9B",X"2D",X"C1",X"0D",X"20",X"F7",X"2E",
		X"72",X"C9",X"3A",X"00",X"42",X"E6",X"7F",X"FE",X"05",X"38",X"0E",X"21",X"1F",X"2D",X"01",X"05",
		X"00",X"ED",X"B9",X"C0",X"79",X"06",X"23",X"18",X"02",X"06",X"7F",X"87",X"C6",X"11",X"6F",X"26",
		X"2D",X"5E",X"23",X"56",X"2A",X"00",X"41",X"EB",X"CD",X"98",X"1B",X"24",X"05",X"CD",X"98",X"1B",
		X"2C",X"05",X"05",X"CD",X"98",X"1B",X"25",X"04",X"CD",X"98",X"1B",X"06",X"5E",X"2C",X"C3",X"98",
		X"1B",X"90",X"99",X"64",X"00",X"01",X"04",X"90",X"61",X"66",X"66",X"66",X"98",X"00",X"02",X"08",
		X"60",X"92",X"99",X"0E",X"FC",X"18",X"02",X"0E",X"04",X"32",X"22",X"40",X"3A",X"15",X"41",X"FE",
		X"14",X"C0",X"06",X"03",X"21",X"53",X"50",X"79",X"86",X"77",X"23",X"23",X"23",X"23",X"10",X"F7",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"1D",X"40",X"2F",X"0F",
		X"0F",X"0F",X"47",X"E6",X"E0",X"4F",X"78",X"E6",X"03",X"47",X"A7",X"ED",X"42",X"01",X"3A",X"50",
		X"CD",X"CB",X"0A",X"D9",X"C9",X"2A",X"00",X"41",X"EB",X"21",X"1A",X"41",X"7E",X"E6",X"7F",X"23",
		X"BE",X"28",X"2A",X"38",X"35",X"34",X"66",X"2E",X"71",X"01",X"02",X"8D",X"CB",X"44",X"28",X"02",
		X"06",X"8F",X"E5",X"C5",X"CD",X"26",X"9B",X"2D",X"05",X"CD",X"26",X"9B",X"2D",X"C1",X"0D",X"20",
		X"F2",X"E1",X"24",X"78",X"FE",X"95",X"28",X"41",X"01",X"02",X"95",X"18",X"E5",X"CD",X"F4",X"97",
		X"66",X"24",X"2E",X"72",X"DD",X"21",X"B1",X"2C",X"18",X"45",X"2B",X"35",X"7E",X"FE",X"83",X"20",
		X"0F",X"21",X"72",X"03",X"CD",X"33",X"2A",X"24",X"CD",X"33",X"2A",X"24",X"CD",X"33",X"2A",X"C9",
		X"30",X"09",X"FE",X"08",X"D0",X"C3",X"78",X"99",X"00",X"00",X"00",X"E6",X"7F",X"67",X"2E",X"72",
		X"24",X"24",X"CD",X"33",X"2A",X"25",X"25",X"18",X"12",X"3A",X"00",X"42",X"E6",X"03",X"C0",X"21",
		X"1A",X"41",X"7E",X"FE",X"4F",X"30",X"21",X"34",X"CD",X"24",X"2A",X"DD",X"21",X"A5",X"2C",X"01",
		X"02",X"06",X"C5",X"DD",X"46",X"00",X"CD",X"26",X"9B",X"2D",X"C1",X"DD",X"23",X"10",X"F3",X"06",
		X"06",X"2E",X"72",X"24",X"0D",X"20",X"EB",X"C9",X"36",X"D0",X"23",X"36",X"D1",X"C9",X"CD",X"F2",
		X"9C",X"C3",X"54",X"02",X"00",X"00",X"F1",X"E1",X"F1",X"7C",X"E6",X"F8",X"3D",X"67",X"22",X"02",
		X"41",X"21",X"48",X"50",X"06",X"05",X"36",X"F8",X"23",X"23",X"23",X"23",X"10",X"F8",X"3A",X"1A",
		X"41",X"F5",X"CD",X"E5",X"2A",X"3A",X"1A",X"41",X"47",X"F1",X"B8",X"30",X"1C",X"3A",X"22",X"40",
		X"A7",X"28",X"08",X"CD",X"60",X"29",X"CD",X"00",X"28",X"18",X"F2",X"3E",X"80",X"32",X"22",X"40",
		X"06",X"02",X"C5",X"CD",X"60",X"29",X"C1",X"10",X"F9",X"3A",X"1A",X"41",X"FE",X"D0",X"28",X"07",
		X"06",X"01",X"CD",X"56",X"0D",X"18",X"C7",X"3E",X"73",X"32",X"04",X"41",X"C3",X"E0",X"2C",X"00",
		X"3A",X"20",X"41",X"A7",X"28",X"02",X"AF",X"C9",X"3A",X"15",X"41",X"C9",X"00",X"00",X"00",X"00",
		X"FF",X"2D",X"05",X"A0",X"FF",X"2D",X"05",X"A0",X"FF",X"2C",X"03",X"A0",X"A9",X"2A",X"01",X"47",
		X"3A",X"20",X"41",X"A7",X"20",X"06",X"0E",X"5E",X"C5",X"C3",X"56",X"17",X"0E",X"02",X"C5",X"E5",
		X"CD",X"20",X"2E",X"2B",X"10",X"FA",X"E1",X"CD",X"6E",X"11",X"C1",X"0D",X"20",X"F0",X"C9",X"3A",
		X"20",X"41",X"A7",X"CA",X"F6",X"16",X"CD",X"EB",X"16",X"06",X"05",X"CD",X"20",X"2E",X"2B",X"CD",
		X"20",X"2E",X"23",X"19",X"10",X"F5",X"C9",X"7D",X"A7",X"28",X"02",X"2E",X"01",X"22",X"1F",X"41",
		X"C9",X"3A",X"00",X"60",X"E6",X"20",X"C8",X"3A",X"07",X"41",X"C9",X"22",X"24",X"41",X"3E",X"20",
		X"32",X"62",X"40",X"C9",X"3E",X"05",X"32",X"63",X"40",X"C3",X"00",X"0E",X"3E",X"01",X"32",X"66",
		X"40",X"C3",X"38",X"9A",X"3E",X"01",X"32",X"67",X"40",X"C3",X"5A",X"8B",X"32",X"02",X"60",X"32",
		X"06",X"60",X"C9",X"00",X"00",X"26",X"50",X"7E",X"32",X"6B",X"40",X"1A",X"C9",X"77",X"3E",X"30",
		X"32",X"6C",X"40",X"C3",X"E4",X"38",X"32",X"5A",X"50",X"3E",X"30",X"32",X"6C",X"40",X"C9",X"32",
		X"5E",X"50",X"18",X"F5",X"00",X"9D",X"8D",X"8C",X"8D",X"8C",X"93",X"9C",X"9B",X"9A",X"90",X"91",
		X"92",X"A1",X"8D",X"8C",X"8D",X"8C",X"99",X"A0",X"9F",X"9E",X"96",X"97",X"98",X"00",X"00",X"00",
		X"00",X"3A",X"15",X"41",X"FE",X"14",X"C0",X"3A",X"00",X"41",X"FE",X"20",X"D8",X"11",X"50",X"50",
		X"21",X"00",X"2C",X"01",X"10",X"00",X"ED",X"B0",X"F1",X"C3",X"E0",X"2C",X"00",X"00",X"00",X"00",
		X"CD",X"00",X"8C",X"CD",X"B8",X"1A",X"CD",X"A0",X"3C",X"CD",X"3B",X"0A",X"CD",X"45",X"1B",X"CD",
		X"E5",X"2A",X"CD",X"9B",X"A0",X"CD",X"9C",X"37",X"CD",X"B5",X"37",X"CD",X"B2",X"2D",X"CD",X"DA",
		X"2D",X"CD",X"A9",X"3A",X"CD",X"70",X"84",X"21",X"00",X"42",X"7E",X"BE",X"28",X"FD",X"C3",X"E0",
		X"2C",X"A6",X"1F",X"9C",X"2A",X"92",X"33",X"87",X"3B",X"7D",X"44",X"10",X"20",X"30",X"50",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"15",
		X"41",X"FE",X"14",X"C2",X"67",X"8A",X"E1",X"E5",X"11",X"F3",X"10",X"19",X"CD",X"64",X"08",X"7E",
		X"FE",X"E0",X"20",X"05",X"16",X"00",X"C3",X"73",X"02",X"2B",X"7E",X"FE",X"E0",X"CA",X"81",X"36",
		X"E1",X"E5",X"11",X"00",X"0D",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"E0",X"C2",X"D3",X"02",X"C3",
		X"89",X"36",X"7D",X"CD",X"EC",X"8C",X"E5",X"CD",X"60",X"29",X"CD",X"00",X"28",X"E1",X"3A",X"01",
		X"41",X"A7",X"C8",X"7C",X"FE",X"CF",X"D8",X"D6",X"08",X"67",X"32",X"03",X"41",X"E5",X"CD",X"06",
		X"28",X"CD",X"42",X"28",X"E1",X"C9",X"48",X"54",X"60",X"78",X"84",X"90",X"9C",X"4A",X"56",X"62",
		X"7A",X"86",X"92",X"9E",X"49",X"55",X"61",X"79",X"85",X"91",X"9D",X"4B",X"57",X"63",X"7B",X"87",
		X"93",X"9F",X"A2",X"A2",X"A3",X"5E",X"A2",X"A3",X"5E",X"5E",X"A3",X"5E",X"5E",X"5E",X"5E",X"5E",
		X"5E",X"5E",X"3A",X"00",X"42",X"E6",X"10",X"3E",X"2A",X"20",X"02",X"3E",X"17",X"32",X"5D",X"50",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"00",X"41",X"FE",X"91",X"C0",
		X"3A",X"02",X"41",X"FE",X"DC",X"D8",X"3A",X"04",X"41",X"FE",X"75",X"D0",X"3A",X"01",X"41",X"FE",
		X"20",X"28",X"0D",X"CD",X"60",X"29",X"CD",X"00",X"28",X"CD",X"66",X"29",X"CD",X"A2",X"29",X"C9",
		X"21",X"36",X"07",X"22",X"00",X"41",X"3E",X"0E",X"32",X"15",X"41",X"3E",X"01",X"32",X"1F",X"41",
		X"3E",X"F8",X"00",X"32",X"54",X"50",X"32",X"58",X"50",X"CD",X"78",X"89",X"F1",X"C3",X"98",X"1B",
		X"7D",X"E6",X"1F",X"C6",X"A2",X"FE",X"AE",X"38",X"04",X"FE",X"B7",X"38",X"02",X"3E",X"5E",X"77",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"1F",X"41",X"A7",X"28",X"13",X"06",X"03",X"23",X"36",X"DE",X"10",X"FB",X"FE",X"04",X"38",
		X"0C",X"FE",X"1D",X"30",X"13",X"3C",X"32",X"1F",X"41",X"2A",X"00",X"41",X"C9",X"06",X"18",X"2B",
		X"2B",X"2B",X"36",X"5E",X"10",X"FB",X"18",X"ED",X"47",X"28",X"12",X"CD",X"F0",X"2B",X"FE",X"10",
		X"38",X"E7",X"78",X"FE",X"2F",X"20",X"DE",X"F1",X"F1",X"C3",X"AA",X"30",X"00",X"AF",X"CD",X"7C",
		X"2C",X"78",X"18",X"D1",X"95",X"5E",X"5E",X"5E",X"96",X"92",X"5E",X"5E",X"96",X"93",X"7F",X"7E",
		X"96",X"93",X"7D",X"7C",X"96",X"93",X"AD",X"5E",X"96",X"93",X"AC",X"5E",X"96",X"93",X"5E",X"5E",
		X"96",X"93",X"5E",X"5E",X"5E",X"8E",X"7F",X"7E",X"96",X"93",X"5E",X"5E",X"5E",X"8F",X"7D",X"7C",
		X"96",X"93",X"91",X"91",X"91",X"8F",X"AD",X"5E",X"96",X"94",X"5E",X"5E",X"5E",X"90",X"AC",X"5E",
		X"97",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"3E",X"01",X"32",X"04",X"60",X"00",X"00",X"00",
		X"C3",X"AA",X"30",X"06",X"06",X"06",X"06",X"06",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",
		X"02",X"02",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"04",X"04",X"04",X"04",X"04",X"06",X"06",
		X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"02",X"41",X"0F",X"0F",X"0F",X"E6",X"1F",X"47",X"3A",
		X"00",X"41",X"C6",X"10",X"80",X"FE",X"34",X"38",X"05",X"3E",X"02",X"32",X"20",X"41",X"01",X"34",
		X"50",X"0A",X"E6",X"07",X"C0",X"21",X"3A",X"48",X"CD",X"CB",X"0A",X"EB",X"2A",X"00",X"41",X"4E",
		X"79",X"EB",X"E6",X"0F",X"28",X"06",X"47",X"36",X"C0",X"2B",X"10",X"FB",X"79",X"E6",X"70",X"28",
		X"13",X"0F",X"0F",X"0F",X"0F",X"C6",X"C0",X"77",X"FE",X"C5",X"28",X"04",X"FE",X"C7",X"20",X"03",
		X"3D",X"2B",X"77",X"2B",X"CB",X"79",X"CA",X"5C",X"30",X"13",X"1A",X"4F",X"E6",X"0F",X"28",X"51",
		X"FE",X"03",X"28",X"09",X"30",X"0E",X"3D",X"28",X"07",X"36",X"8D",X"18",X"44",X"36",X"8D",X"2B",
		X"36",X"8C",X"18",X"3D",X"FE",X"06",X"28",X"0C",X"30",X"0D",X"FE",X"05",X"28",X"01",X"23",X"22",
		X"02",X"40",X"18",X"2D",X"2B",X"18",X"F8",X"FE",X"09",X"28",X"0A",X"30",X"16",X"FE",X"08",X"28",
		X"08",X"3E",X"0D",X"18",X"06",X"3E",X"0F",X"18",X"02",X"3E",X"0E",X"32",X"15",X"41",X"22",X"17",
		X"40",X"18",X"0E",X"D5",X"C5",X"E5",X"C6",X"93",X"11",X"20",X"00",X"CD",X"AE",X"15",X"E1",X"C1",
		X"D1",X"79",X"E6",X"F0",X"28",X"29",X"FE",X"F0",X"28",X"27",X"D6",X"10",X"0F",X"FE",X"38",X"30",
		X"07",X"0F",X"C6",X"84",X"06",X"04",X"18",X"06",X"D6",X"38",X"C6",X"A0",X"06",X"08",X"D5",X"5F",
		X"16",X"2E",X"7D",X"E6",X"E0",X"C6",X"0B",X"6F",X"1A",X"77",X"13",X"2B",X"10",X"FA",X"D1",X"18",
		X"4B",X"13",X"1A",X"D5",X"4F",X"E6",X"0F",X"28",X"17",X"07",X"47",X"07",X"80",X"C6",X"0A",X"5F",
		X"16",X"31",X"7D",X"E6",X"E0",X"C6",X"0C",X"CD",X"EE",X"93",X"1A",X"77",X"13",X"23",X"10",X"FA",
		X"79",X"FE",X"E0",X"30",X"1D",X"E6",X"E0",X"07",X"07",X"07",X"CD",X"20",X"33",X"00",X"6F",X"11",
		X"25",X"40",X"CB",X"61",X"28",X"02",X"1E",X"2F",X"06",X"05",X"1A",X"A7",X"28",X"07",X"13",X"13",
		X"10",X"F8",X"D1",X"18",X"07",X"7C",X"12",X"1B",X"7D",X"12",X"18",X"F6",X"EB",X"3A",X"20",X"41",
		X"4F",X"7D",X"FE",X"B9",X"28",X"0B",X"FE",X"56",X"28",X"16",X"FE",X"95",X"20",X"23",X"C3",X"5E",
		X"89",X"79",X"FE",X"02",X"00",X"00",X"21",X"BA",X"24",X"79",X"3C",X"32",X"20",X"41",X"18",X"12",
		X"7C",X"FE",X"25",X"20",X"0C",X"23",X"18",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"E8",X"23",X"22",X"00",X"41",X"EB",X"7D",X"E6",X"E0",X"C6",X"0C",X"6F",X"01",X"AE",X"09",X"7E",
		X"FE",X"5E",X"20",X"01",X"71",X"23",X"0C",X"10",X"F6",X"C9",X"06",X"0F",X"21",X"35",X"50",X"36",
		X"03",X"2B",X"2B",X"10",X"FA",X"06",X"09",X"36",X"01",X"2B",X"2B",X"10",X"FA",X"3E",X"01",X"32",
		X"20",X"41",X"32",X"03",X"60",X"AF",X"32",X"02",X"60",X"21",X"F0",X"23",X"22",X"00",X"41",X"3E",
		X"05",X"32",X"0C",X"41",X"C3",X"CC",X"87",X"2B",X"2B",X"35",X"35",X"C3",X"DA",X"37",X"34",X"26",
		X"50",X"1A",X"86",X"CD",X"B9",X"97",X"2B",X"18",X"F1",X"3A",X"07",X"41",X"E6",X"08",X"C0",X"C3",
		X"D3",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7D",X"E6",X"E0",X"C6",X"0C",X"6F",X"7E",X"FE",X"C0",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5E",X"5E",X"5E",X"87",X"5E",X"5E",X"80",X"5E",X"87",X"5E",X"5E",X"5E",X"81",X"85",X"5E",X"5E",
		X"5E",X"5E",X"82",X"5E",X"86",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"86",X"5E",X"5E",X"5E",X"5E",
		X"5E",X"5E",X"86",X"5E",X"81",X"83",X"86",X"87",X"5E",X"5E",X"82",X"5E",X"86",X"5E",X"5E",X"87",
		X"5E",X"5E",X"5E",X"86",X"87",X"5E",X"5E",X"5E",X"5E",X"5E",X"87",X"5E",X"80",X"5E",X"5E",X"87",
		X"5E",X"5E",X"81",X"84",X"85",X"5E",X"5E",X"5E",X"81",X"85",X"5E",X"86",X"87",X"5E",X"80",X"5E",
		X"87",X"86",X"5E",X"5E",X"81",X"84",X"5E",X"5E",X"86",X"5E",X"3A",X"20",X"41",X"A7",X"20",X"11",
		X"3A",X"15",X"41",X"FE",X"14",X"CA",X"21",X"1B",X"CD",X"55",X"0F",X"CD",X"00",X"0D",X"C3",X"16",
		X"88",X"FE",X"12",X"D2",X"80",X"35",X"3D",X"28",X"0F",X"FE",X"04",X"D2",X"A7",X"31",X"3A",X"00",
		X"42",X"0F",X"D8",X"CD",X"4E",X"2F",X"18",X"03",X"CD",X"36",X"2F",X"CD",X"00",X"0D",X"3A",X"34",
		X"50",X"47",X"D9",X"CD",X"EA",X"11",X"C9",X"3A",X"00",X"42",X"0F",X"D8",X"01",X"34",X"50",X"0A",
		X"E6",X"07",X"C2",X"9B",X"31",X"21",X"3A",X"48",X"CD",X"CB",X"0A",X"EB",X"2A",X"00",X"41",X"4E",
		X"EB",X"79",X"E6",X"7F",X"28",X"2F",X"CB",X"61",X"28",X"75",X"79",X"E6",X"0F",X"28",X"06",X"47",
		X"36",X"C0",X"2B",X"10",X"FB",X"79",X"E6",X"60",X"28",X"0D",X"FE",X"40",X"38",X"10",X"28",X"12",
		X"36",X"C7",X"2B",X"36",X"C6",X"18",X"0D",X"36",X"C5",X"2B",X"36",X"C4",X"18",X"06",X"36",X"C1",
		X"18",X"02",X"36",X"C2",X"2B",X"CB",X"79",X"28",X"44",X"13",X"1A",X"FE",X"03",X"28",X"08",X"30",
		X"0F",X"3D",X"28",X"07",X"2B",X"18",X"04",X"7D",X"D6",X"08",X"6F",X"22",X"02",X"40",X"18",X"2D",
		X"FE",X"08",X"30",X"0E",X"C6",X"99",X"D5",X"E5",X"11",X"20",X"00",X"CD",X"AE",X"15",X"E1",X"D1",
		X"18",X"1B",X"FE",X"0D",X"30",X"7C",X"2B",X"2B",X"36",X"B7",X"FE",X"09",X"20",X"0F",X"D5",X"E5",
		X"11",X"58",X"50",X"21",X"F1",X"1F",X"01",X"08",X"00",X"ED",X"B0",X"E1",X"D1",X"18",X"14",X"00",
		X"00",X"00",X"00",X"00",X"7D",X"E6",X"E0",X"C6",X"0C",X"6F",X"79",X"E6",X"0F",X"47",X"36",X"C0",
		X"23",X"10",X"FB",X"CD",X"96",X"30",X"EB",X"3A",X"20",X"41",X"4F",X"7D",X"FE",X"D8",X"28",X"10",
		X"FE",X"F8",X"28",X"1D",X"FE",X"1B",X"28",X"2C",X"FE",X"46",X"20",X"2F",X"3E",X"08",X"18",X"09",
		X"79",X"FE",X"05",X"28",X"09",X"FE",X"0D",X"00",X"00",X"21",X"F9",X"25",X"18",X"10",X"23",X"18",
		X"0D",X"79",X"FE",X"07",X"28",X"05",X"21",X"D9",X"25",X"18",X"03",X"21",X"B9",X"25",X"3C",X"32",
		X"20",X"41",X"18",X"08",X"79",X"FE",X"0A",X"20",X"E0",X"18",X"E3",X"23",X"22",X"00",X"41",X"C3",
		X"9B",X"31",X"06",X"0A",X"36",X"B7",X"2B",X"10",X"FB",X"18",X"92",X"3A",X"20",X"41",X"A7",X"C8",
		X"FE",X"12",X"D0",X"01",X"34",X"50",X"0A",X"E6",X"07",X"FE",X"02",X"20",X"44",X"21",X"25",X"40",
		X"7E",X"A7",X"20",X"09",X"23",X"23",X"7D",X"FE",X"39",X"20",X"F5",X"18",X"34",X"56",X"2B",X"5E",
		X"23",X"E5",X"EB",X"E5",X"CD",X"13",X"11",X"20",X"06",X"E1",X"E1",X"36",X"00",X"18",X"E5",X"E1",
		X"D1",X"D5",X"3A",X"34",X"50",X"E6",X"08",X"20",X"09",X"7B",X"FE",X"2E",X"30",X"0D",X"C3",X"2C",
		X"97",X"00",X"7B",X"FE",X"2E",X"38",X"04",X"C3",X"36",X"97",X"00",X"CD",X"20",X"2E",X"E1",X"18",
		X"C3",X"3A",X"59",X"50",X"FE",X"A8",X"C0",X"3A",X"00",X"42",X"0F",X"D8",X"3A",X"58",X"50",X"FE",
		X"F0",X"C3",X"BB",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"47",X"7D",X"E6",X"E0",X"C6",X"0F",X"80",X"C9",X"3A",X"07",X"41",X"47",X"E6",X"01",X"3C",X"07",
		X"A0",X"28",X"18",X"3E",X"17",X"32",X"49",X"50",X"7C",X"FE",X"C7",X"D0",X"24",X"24",X"7D",X"CD",
		X"3A",X"02",X"E5",X"06",X"01",X"CD",X"50",X"19",X"E1",X"18",X"ED",X"11",X"4F",X"50",X"7C",X"12",
		X"32",X"4B",X"50",X"7D",X"32",X"4C",X"50",X"D6",X"0F",X"32",X"48",X"50",X"3E",X"3E",X"32",X"41",
		X"50",X"3C",X"32",X"45",X"50",X"3E",X"05",X"32",X"49",X"50",X"3D",X"32",X"4D",X"50",X"3E",X"04",
		X"32",X"4E",X"50",X"32",X"4A",X"50",X"1A",X"FE",X"C7",X"30",X"06",X"3C",X"3C",X"12",X"32",X"4B",
		X"50",X"7C",X"FE",X"C7",X"30",X"0E",X"24",X"7D",X"CD",X"3A",X"02",X"E5",X"06",X"01",X"CD",X"40",
		X"19",X"E1",X"18",X"E2",X"3E",X"F1",X"32",X"4C",X"50",X"3E",X"05",X"32",X"4E",X"50",X"3E",X"07",
		X"32",X"4A",X"50",X"3E",X"03",X"32",X"4D",X"50",X"C9",X"00",X"00",X"00",X"3A",X"00",X"42",X"0F",
		X"D8",X"CD",X"FF",X"9C",X"FE",X"2F",X"20",X"13",X"06",X"04",X"3A",X"00",X"42",X"E6",X"20",X"20",
		X"02",X"06",X"06",X"78",X"32",X"41",X"50",X"3C",X"32",X"45",X"50",X"2A",X"02",X"41",X"CD",X"A2",
		X"01",X"CD",X"D3",X"01",X"3A",X"03",X"41",X"BC",X"D2",X"63",X"34",X"E5",X"11",X"F3",X"10",X"19",
		X"CD",X"64",X"08",X"11",X"20",X"00",X"7E",X"FE",X"C1",X"28",X"0B",X"FE",X"93",X"28",X"07",X"FE",
		X"8F",X"20",X"4E",X"00",X"00",X"00",X"2B",X"1E",X"A0",X"CD",X"3C",X"0E",X"0E",X"08",X"1E",X"20",
		X"19",X"0D",X"28",X"2A",X"7E",X"D6",X"A6",X"38",X"F7",X"FE",X"08",X"30",X"F3",X"0F",X"38",X"F0",
		X"C6",X"2B",X"4F",X"06",X"03",X"CD",X"20",X"2E",X"19",X"CD",X"20",X"2E",X"10",X"FA",X"2B",X"CD",
		X"20",X"2E",X"CD",X"3C",X"0E",X"CD",X"20",X"2E",X"06",X"19",X"0A",X"CD",X"34",X"0E",X"E1",X"7C",
		X"3C",X"E6",X"F8",X"67",X"3E",X"73",X"32",X"04",X"41",X"3E",X"0F",X"32",X"08",X"41",X"C3",X"B1",
		X"02",X"C3",X"5B",X"34",X"00",X"7E",X"FE",X"C1",X"20",X"09",X"E1",X"E1",X"CD",X"3B",X"8B",X"3E",
		X"98",X"18",X"E3",X"19",X"19",X"7E",X"FE",X"C1",X"28",X"F0",X"E1",X"7D",X"E6",X"1F",X"FE",X"1B",
		X"30",X"94",X"E1",X"E5",X"11",X"F3",X"05",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"C0",X"20",X"06",
		X"CD",X"00",X"31",X"00",X"28",X"D5",X"E1",X"7C",X"FE",X"4D",X"38",X"10",X"FE",X"54",X"30",X"0C",
		X"3E",X"2E",X"32",X"41",X"50",X"3C",X"CD",X"0E",X"97",X"C3",X"B1",X"02",X"3A",X"5C",X"50",X"95",
		X"FE",X"04",X"30",X"F5",X"3A",X"59",X"50",X"FE",X"A8",X"20",X"EE",X"3A",X"43",X"50",X"FE",X"9F",
		X"CA",X"E2",X"3D",X"30",X"03",X"3C",X"18",X"01",X"3D",X"32",X"43",X"50",X"32",X"47",X"50",X"06",
		X"01",X"CD",X"56",X"0D",X"18",X"E5",X"00",X"00",X"00",X"3A",X"20",X"41",X"3D",X"FE",X"2F",X"D0",
		X"2A",X"21",X"41",X"CD",X"17",X"97",X"19",X"7C",X"FE",X"4C",X"20",X"02",X"26",X"48",X"22",X"21",
		X"41",X"7E",X"FE",X"A4",X"28",X"07",X"FE",X"A5",X"28",X"03",X"FE",X"5E",X"C0",X"23",X"7E",X"FE",
		X"C0",X"28",X"0A",X"FE",X"AE",X"28",X"06",X"FE",X"80",X"D8",X"FE",X"83",X"D0",X"2B",X"ED",X"5F",
		X"E6",X"02",X"20",X"03",X"36",X"A4",X"C9",X"36",X"A5",X"C9",X"AF",X"32",X"48",X"50",X"CD",X"C7",
		X"97",X"06",X"60",X"CD",X"62",X"93",X"01",X"10",X"06",X"21",X"43",X"50",X"35",X"2E",X"47",X"35",
		X"2E",X"5B",X"35",X"2E",X"5F",X"35",X"C5",X"06",X"02",X"CD",X"56",X"0D",X"C1",X"10",X"EA",X"06",
		X"06",X"C5",X"CD",X"66",X"29",X"C1",X"0D",X"20",X"E0",X"06",X"98",X"21",X"5B",X"50",X"34",X"2E",
		X"5F",X"34",X"C5",X"06",X"02",X"CD",X"56",X"0D",X"C1",X"10",X"F0",X"3E",X"00",X"32",X"58",X"50",
		X"32",X"5C",X"50",X"3E",X"12",X"32",X"20",X"41",X"3A",X"43",X"50",X"32",X"03",X"41",X"3E",X"03",
		X"32",X"3B",X"50",X"32",X"39",X"50",X"3E",X"01",X"32",X"37",X"50",X"21",X"35",X"50",X"06",X"18",
		X"36",X"07",X"2B",X"2B",X"10",X"FA",X"21",X"1B",X"48",X"11",X"20",X"00",X"06",X"20",X"36",X"A5",
		X"23",X"36",X"AE",X"23",X"36",X"AF",X"2B",X"2B",X"19",X"10",X"F3",X"CD",X"90",X"36",X"C9",X"00",
		X"01",X"34",X"50",X"0A",X"E6",X"07",X"C2",X"97",X"3A",X"21",X"23",X"41",X"35",X"20",X"05",X"36",
		X"10",X"2E",X"20",X"34",X"21",X"28",X"48",X"CD",X"CB",X"0A",X"11",X"20",X"00",X"3A",X"20",X"41",
		X"FE",X"30",X"30",X"42",X"0A",X"E6",X"18",X"FE",X"18",X"20",X"3B",X"ED",X"5F",X"E6",X"10",X"20",
		X"35",X"E5",X"ED",X"5F",X"E6",X"0F",X"85",X"6F",X"0E",X"A8",X"E6",X"02",X"20",X"02",X"0E",X"AB",
		X"71",X"CD",X"3C",X"0E",X"0D",X"71",X"CD",X"3C",X"0E",X"0D",X"71",X"19",X"19",X"7D",X"E6",X"07",
		X"20",X"05",X"22",X"02",X"40",X"18",X"0E",X"2B",X"36",X"7F",X"2B",X"36",X"7E",X"CD",X"3C",X"0E",
		X"36",X"7C",X"23",X"36",X"7D",X"E1",X"3A",X"20",X"41",X"FE",X"2C",X"DA",X"97",X"3A",X"7D",X"E6",
		X"E0",X"C6",X"1D",X"6F",X"06",X"05",X"36",X"AD",X"2B",X"10",X"FB",X"3A",X"23",X"41",X"E6",X"03",
		X"C2",X"97",X"3A",X"36",X"AC",X"C3",X"97",X"3A",X"CD",X"C0",X"83",X"CD",X"24",X"1F",X"21",X"4D",
		X"9D",X"3A",X"07",X"41",X"47",X"E6",X"01",X"3C",X"07",X"A0",X"28",X"02",X"2E",X"3B",X"CD",X"17",
		X"0A",X"11",X"20",X"00",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"52",X"4F",X"06",X"41",X"0A",X"21",
		X"DE",X"4A",X"06",X"0C",X"A7",X"28",X"09",X"D6",X"02",X"30",X"09",X"AF",X"36",X"1E",X"18",X"06",
		X"36",X"1D",X"18",X"02",X"36",X"1F",X"F5",X"CD",X"3C",X"0E",X"F1",X"10",X"E7",X"CB",X"45",X"C0",
		X"21",X"DF",X"4A",X"18",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"07",X"41",X"E6",X"08",X"28",X"07",X"2A",X"14",
		X"42",X"7C",X"B5",X"20",X"04",X"21",X"00",X"42",X"C9",X"F1",X"C9",X"3E",X"01",X"32",X"5A",X"50",
		X"C9",X"3E",X"9D",X"32",X"04",X"41",X"C3",X"D3",X"02",X"E1",X"26",X"BF",X"C3",X"D4",X"02",X"00",
		X"CD",X"BC",X"87",X"C6",X"10",X"32",X"21",X"41",X"3E",X"41",X"32",X"23",X"41",X"32",X"02",X"60",
		X"3E",X"04",X"32",X"42",X"50",X"3E",X"06",X"32",X"0C",X"41",X"C3",X"D9",X"3A",X"00",X"00",X"00",
		X"3A",X"3B",X"40",X"A7",X"28",X"06",X"3D",X"32",X"3B",X"40",X"18",X"03",X"32",X"3C",X"40",X"CD",
		X"FF",X"9C",X"2A",X"02",X"41",X"7C",X"FE",X"D3",X"38",X"09",X"3E",X"20",X"32",X"41",X"50",X"3C",
		X"32",X"45",X"50",X"CD",X"A2",X"01",X"CD",X"D3",X"01",X"E5",X"11",X"F3",X"10",X"19",X"CD",X"64",
		X"08",X"7E",X"FE",X"AD",X"28",X"60",X"FE",X"A6",X"38",X"48",X"FE",X"AC",X"30",X"44",X"11",X"20",
		X"00",X"2B",X"7E",X"FE",X"7F",X"28",X"0D",X"FE",X"7D",X"28",X"0C",X"19",X"7E",X"FE",X"7D",X"28",
		X"06",X"E1",X"18",X"3A",X"CD",X"3C",X"0E",X"CD",X"3C",X"0E",X"36",X"00",X"19",X"36",X"00",X"2B",
		X"36",X"5E",X"19",X"36",X"5E",X"23",X"3A",X"3C",X"40",X"3C",X"FE",X"09",X"28",X"03",X"32",X"3C",
		X"40",X"77",X"07",X"47",X"07",X"07",X"80",X"CD",X"34",X"0E",X"3E",X"60",X"32",X"3B",X"40",X"E1",
		X"18",X"0C",X"E1",X"7C",X"FE",X"D7",X"38",X"0B",X"FE",X"F0",X"30",X"07",X"26",X"D7",X"3E",X"73",
		X"32",X"04",X"41",X"C3",X"B1",X"02",X"E1",X"3E",X"B8",X"32",X"43",X"50",X"32",X"47",X"50",X"CD",
		X"77",X"37",X"F1",X"00",X"00",X"CD",X"E2",X"9A",X"C3",X"AE",X"89",X"C2",X"8E",X"38",X"2B",X"2B",
		X"7E",X"D6",X"06",X"77",X"C3",X"DA",X"37",X"3A",X"15",X"41",X"FE",X"0A",X"DA",X"93",X"8A",X"3E",
		X"07",X"32",X"72",X"40",X"C3",X"90",X"8A",X"CD",X"47",X"93",X"3E",X"10",X"32",X"41",X"50",X"3C",
		X"32",X"45",X"50",X"C9",X"CD",X"CF",X"12",X"CD",X"70",X"9F",X"06",X"B0",X"CD",X"56",X"0D",X"C9",
		X"CD",X"84",X"37",X"C3",X"18",X"03",X"CD",X"84",X"37",X"C3",X"E0",X"2C",X"DD",X"21",X"50",X"50",
		X"FD",X"21",X"0E",X"41",X"CD",X"8B",X"A7",X"DD",X"21",X"54",X"50",X"FD",X"21",X"11",X"41",X"CD",
		X"B2",X"9F",X"C3",X"A0",X"1E",X"3A",X"00",X"42",X"07",X"07",X"07",X"07",X"32",X"06",X"60",X"C9",
		X"00",X"00",X"00",X"3A",X"20",X"41",X"FE",X"12",X"DA",X"6C",X"15",X"C3",X"66",X"9C",X"0F",X"D8",
		X"21",X"50",X"50",X"06",X"04",X"7E",X"FE",X"F8",X"38",X"09",X"23",X"23",X"23",X"23",X"10",X"F5",
		X"C3",X"D1",X"38",X"23",X"23",X"7E",X"FE",X"04",X"20",X"13",X"CD",X"92",X"97",X"00",X"E6",X"08",
		X"3E",X"2C",X"20",X"01",X"3C",X"77",X"2B",X"7E",X"D6",X"04",X"77",X"18",X"DD",X"26",X"40",X"7E",
		X"A7",X"20",X"04",X"26",X"50",X"18",X"D5",X"3D",X"28",X"1E",X"3D",X"28",X"51",X"3D",X"20",X"5E",
		X"23",X"7E",X"FE",X"3A",X"28",X"2B",X"5E",X"16",X"8B",X"1A",X"4F",X"35",X"CA",X"C0",X"97",X"00",
		X"26",X"50",X"7E",X"91",X"C3",X"E3",X"30",X"00",X"23",X"5E",X"23",X"56",X"13",X"7B",X"FE",X"23",
		X"20",X"03",X"11",X"D3",X"2E",X"72",X"2B",X"73",X"CD",X"85",X"2C",X"86",X"77",X"2B",X"C3",X"D7",
		X"30",X"3A",X"02",X"41",X"26",X"50",X"2B",X"2B",X"2B",X"96",X"FE",X"D0",X"38",X"A9",X"26",X"40",
		X"23",X"23",X"23",X"ED",X"5F",X"E6",X"07",X"C6",X"30",X"77",X"26",X"50",X"18",X"DF",X"26",X"50",
		X"23",X"7E",X"FE",X"DA",X"30",X"D7",X"26",X"40",X"5E",X"16",X"8B",X"C3",X"DE",X"30",X"3D",X"28",
		X"10",X"3D",X"28",X"28",X"3D",X"28",X"36",X"3D",X"28",X"42",X"26",X"50",X"3D",X"C3",X"5B",X"37",
		X"00",X"26",X"50",X"2B",X"3A",X"00",X"42",X"E6",X"02",X"0F",X"C6",X"2E",X"77",X"23",X"23",X"CD",
		X"A6",X"A7",X"30",X"A8",X"2B",X"2B",X"2B",X"36",X"FF",X"C3",X"DA",X"37",X"26",X"50",X"23",X"3A",
		X"53",X"50",X"77",X"2B",X"2B",X"2B",X"3A",X"50",X"50",X"D6",X"04",X"18",X"1D",X"26",X"50",X"23",
		X"3A",X"57",X"50",X"77",X"2B",X"2B",X"2B",X"3A",X"54",X"50",X"18",X"ED",X"3A",X"3F",X"40",X"4F",
		X"3A",X"34",X"50",X"91",X"C6",X"F5",X"26",X"50",X"2B",X"2B",X"77",X"23",X"36",X"2E",X"C3",X"DB",
		X"37",X"3A",X"20",X"41",X"FE",X"18",X"30",X"2F",X"2E",X"50",X"06",X"04",X"7E",X"FE",X"F8",X"30",
		X"07",X"23",X"23",X"23",X"23",X"10",X"F5",X"C9",X"ED",X"5F",X"E6",X"0F",X"20",X"F3",X"ED",X"5F",
		X"4F",X"3A",X"00",X"42",X"00",X"00",X"E6",X"70",X"81",X"D6",X"C0",X"30",X"E4",X"36",X"F1",X"C6",
		X"E0",X"23",X"23",X"23",X"C3",X"8D",X"2C",X"4F",X"FE",X"1A",X"D8",X"20",X"1E",X"3A",X"23",X"41",
		X"FE",X"10",X"20",X"17",X"3E",X"02",X"32",X"52",X"50",X"32",X"56",X"50",X"CD",X"7B",X"36",X"32",
		X"5E",X"50",X"3E",X"27",X"32",X"51",X"50",X"32",X"55",X"50",X"C9",X"3A",X"00",X"42",X"E6",X"1F",
		X"FE",X"0E",X"28",X"06",X"21",X"58",X"50",X"C3",X"F6",X"39",X"2E",X"50",X"06",X"02",X"7E",X"FE",
		X"F8",X"30",X"09",X"23",X"23",X"23",X"23",X"10",X"F5",X"C3",X"F6",X"39",X"36",X"F1",X"23",X"23",
		X"23",X"79",X"FE",X"2C",X"30",X"0A",X"ED",X"5F",X"E6",X"30",X"28",X"59",X"FE",X"20",X"20",X"16",
		X"ED",X"5F",X"E6",X"0F",X"07",X"07",X"C6",X"6F",X"77",X"26",X"40",X"36",X"D3",X"23",X"36",X"2E",
		X"2B",X"2B",X"36",X"01",X"18",X"48",X"FE",X"30",X"28",X"51",X"79",X"FE",X"20",X"38",X"4C",X"C5",
		X"E5",X"2B",X"2B",X"2B",X"36",X"F9",X"21",X"3B",X"48",X"01",X"36",X"50",X"CD",X"CB",X"0A",X"22",
		X"3D",X"40",X"3A",X"34",X"50",X"32",X"3F",X"40",X"36",X"93",X"11",X"20",X"00",X"CD",X"3C",X"0E",
		X"36",X"92",X"CD",X"3C",X"0E",X"36",X"91",X"E1",X"C1",X"7D",X"C6",X"05",X"6F",X"7E",X"FE",X"F8",
		X"30",X"36",X"C3",X"34",X"39",X"36",X"E2",X"26",X"40",X"36",X"3A",X"2B",X"36",X"03",X"26",X"50",
		X"7D",X"C6",X"06",X"6F",X"7E",X"FE",X"F8",X"38",X"E9",X"18",X"10",X"ED",X"5F",X"E6",X"0F",X"C6",
		X"20",X"77",X"26",X"40",X"36",X"00",X"2B",X"36",X"02",X"18",X"E3",X"36",X"F1",X"3E",X"07",X"90",
		X"26",X"40",X"23",X"23",X"77",X"C3",X"34",X"39",X"36",X"F1",X"23",X"23",X"23",X"36",X"CF",X"26",
		X"40",X"2B",X"36",X"07",X"18",X"EF",X"06",X"02",X"7E",X"FE",X"F8",X"30",X"31",X"26",X"40",X"23",
		X"23",X"7E",X"26",X"50",X"FE",X"04",X"28",X"28",X"FE",X"08",X"28",X"24",X"FE",X"09",X"28",X"20",
		X"2B",X"2B",X"CD",X"90",X"93",X"96",X"FE",X"F0",X"38",X"14",X"23",X"23",X"23",X"3A",X"03",X"41",
		X"96",X"00",X"00",X"30",X"0C",X"26",X"40",X"2B",X"36",X"04",X"C3",X"78",X"96",X"00",X"23",X"23",
		X"23",X"23",X"10",X"C4",X"2A",X"3D",X"40",X"7E",X"FE",X"93",X"C0",X"3A",X"34",X"50",X"4F",X"3A",
		X"3F",X"40",X"91",X"D6",X"F1",X"4F",X"3A",X"02",X"41",X"81",X"FE",X"80",X"D8",X"06",X"25",X"3A",
		X"03",X"41",X"FE",X"B7",X"30",X"01",X"04",X"3A",X"58",X"50",X"FE",X"F8",X"30",X"1C",X"3A",X"5C",
		X"50",X"FE",X"F8",X"D8",X"78",X"32",X"5D",X"50",X"D6",X"1D",X"32",X"5E",X"40",X"79",X"2F",X"D6",
		X"04",X"32",X"5C",X"50",X"3E",X"C7",X"C3",X"82",X"96",X"00",X"78",X"32",X"59",X"50",X"D6",X"1D",
		X"32",X"5A",X"40",X"79",X"2F",X"D6",X"04",X"32",X"58",X"50",X"3E",X"C7",X"C3",X"87",X"96",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"DB",X"4B",X"01",X"34",X"50",X"3D",X"C2",X"9B",
		X"31",X"CD",X"CB",X"0A",X"36",X"5E",X"C3",X"9B",X"31",X"2A",X"24",X"41",X"7D",X"FE",X"F2",X"38",
		X"13",X"C3",X"B5",X"A7",X"E6",X"01",X"3C",X"47",X"3A",X"00",X"40",X"A0",X"C8",X"2A",X"02",X"41",
		X"C3",X"5B",X"2C",X"00",X"C6",X"08",X"6F",X"22",X"24",X"41",X"32",X"4C",X"50",X"7C",X"32",X"4F",
		X"50",X"CD",X"F0",X"3A",X"AF",X"32",X"00",X"40",X"C9",X"3E",X"04",X"32",X"52",X"50",X"32",X"56",
		X"50",X"32",X"5A",X"50",X"32",X"5E",X"50",X"C9",X"3A",X"20",X"41",X"A7",X"C0",X"C3",X"D4",X"10",
		X"7D",X"FE",X"D9",X"D0",X"E5",X"11",X"00",X"0C",X"19",X"CD",X"5C",X"97",X"7E",X"FE",X"20",X"38",
		X"04",X"FE",X"28",X"38",X"5E",X"FE",X"86",X"28",X"22",X"FE",X"87",X"28",X"2D",X"FE",X"93",X"C2",
		X"A7",X"3B",X"3A",X"20",X"41",X"FE",X"12",X"DA",X"A7",X"3B",X"36",X"A4",X"11",X"20",X"00",X"CD",
		X"3C",X"0E",X"36",X"A4",X"CD",X"3C",X"0E",X"36",X"A4",X"18",X"75",X"3A",X"20",X"41",X"A7",X"28",
		X"76",X"FE",X"12",X"30",X"72",X"01",X"24",X"40",X"18",X"0D",X"3A",X"20",X"41",X"A7",X"28",X"67",
		X"FE",X"12",X"30",X"63",X"01",X"2E",X"40",X"CD",X"20",X"2E",X"EB",X"3E",X"05",X"08",X"0A",X"6F",
		X"03",X"0A",X"67",X"A7",X"ED",X"52",X"28",X"07",X"03",X"08",X"3D",X"20",X"F0",X"18",X"41",X"AF",
		X"02",X"18",X"3D",X"11",X"20",X"00",X"D6",X"24",X"30",X"02",X"C6",X"04",X"28",X"0C",X"3D",X"28",
		X"0A",X"3D",X"20",X"01",X"23",X"CD",X"3C",X"0E",X"18",X"01",X"23",X"3E",X"5E",X"77",X"2B",X"77",
		X"19",X"77",X"CD",X"3A",X"97",X"06",X"05",X"DD",X"21",X"02",X"40",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"A7",X"ED",X"52",X"20",X"04",X"DD",X"36",X"01",X"00",X"DD",X"23",X"DD",X"23",X"10",X"EB",
		X"E1",X"3E",X"60",X"32",X"40",X"40",X"C9",X"E1",X"EB",X"3A",X"20",X"41",X"C3",X"CE",X"1F",X"00",
		X"3A",X"51",X"50",X"D6",X"0C",X"28",X"03",X"3D",X"20",X"1D",X"3A",X"50",X"50",X"93",X"FE",X"0C",
		X"30",X"15",X"3A",X"53",X"50",X"D6",X"01",X"92",X"FE",X"0C",X"30",X"0B",X"C3",X"F3",X"3B",X"00",
		X"3E",X"C7",X"32",X"53",X"50",X"18",X"CA",X"3A",X"55",X"50",X"D6",X"0B",X"28",X"03",X"3D",X"20",
		X"1C",X"3A",X"54",X"50",X"93",X"FE",X"0C",X"30",X"14",X"3A",X"57",X"50",X"C6",X"05",X"92",X"FE",
		X"0B",X"30",X"0A",X"3E",X"F1",X"32",X"50",X"50",X"32",X"54",X"50",X"18",X"A4",X"3A",X"59",X"50",
		X"D6",X"08",X"28",X"02",X"3D",X"C0",X"3A",X"58",X"50",X"93",X"FE",X"0C",X"D0",X"3A",X"5B",X"50",
		X"C6",X"05",X"92",X"FE",X"12",X"D0",X"3E",X"01",X"32",X"58",X"50",X"18",X"84",X"FE",X"14",X"20",
		X"38",X"06",X"03",X"21",X"50",X"50",X"7E",X"C6",X"0A",X"93",X"FE",X"13",X"38",X"07",X"23",X"23",
		X"23",X"23",X"10",X"F2",X"C9",X"23",X"23",X"23",X"7E",X"C6",X"03",X"92",X"FE",X"10",X"30",X"F1",
		X"2B",X"2B",X"00",X"00",X"00",X"2B",X"36",X"FF",X"3E",X"60",X"32",X"40",X"40",X"18",X"DF",X"23",
		X"23",X"77",X"3E",X"60",X"32",X"40",X"40",X"18",X"D6",X"3A",X"20",X"41",X"C3",X"91",X"80",X"06",
		X"04",X"21",X"50",X"50",X"7E",X"93",X"FE",X"0C",X"38",X"07",X"23",X"23",X"23",X"23",X"10",X"F4",
		X"C9",X"23",X"23",X"23",X"7E",X"C6",X"05",X"92",X"FE",X"12",X"30",X"F1",X"2B",X"2B",X"3E",X"60",
		X"32",X"40",X"40",X"2B",X"36",X"F9",X"18",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"40",X"40",X"7E",X"A7",X"CA",X"C3",X"37",X"FE",X"60",X"28",X"18",X"FE",X"50",X"28",X"10",
		X"FE",X"40",X"28",X"31",X"FE",X"30",X"28",X"08",X"FE",X"20",X"20",X"31",X"3E",X"1E",X"18",X"27",
		X"3E",X"1D",X"18",X"23",X"3A",X"4C",X"50",X"C6",X"09",X"32",X"48",X"50",X"CD",X"5F",X"8A",X"3A",
		X"4F",X"50",X"C6",X"04",X"32",X"4B",X"50",X"0F",X"0F",X"E6",X"3E",X"32",X"42",X"40",X"4F",X"06",
		X"50",X"0A",X"32",X"41",X"40",X"3E",X"1C",X"32",X"49",X"50",X"35",X"18",X"07",X"3D",X"20",X"FA",
		X"3E",X"17",X"18",X"F3",X"3A",X"42",X"40",X"4F",X"06",X"50",X"0A",X"47",X"3A",X"41",X"40",X"90",
		X"47",X"3A",X"49",X"40",X"90",X"32",X"48",X"50",X"3A",X"20",X"41",X"FE",X"12",X"D8",X"C3",X"CB",
		X"37",X"E5",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"5E",X"20",X"03",X"E1",X"A7",X"C9",X"FE",X"AE",
		X"38",X"04",X"FE",X"B7",X"38",X"F5",X"E1",X"37",X"C9",X"67",X"2D",X"11",X"F0",X"0C",X"CD",X"11",
		X"3D",X"30",X"01",X"2C",X"C3",X"D5",X"3D",X"D6",X"08",X"BC",X"38",X"0C",X"24",X"11",X"F8",X"0E",
		X"CD",X"11",X"3D",X"30",X"0D",X"25",X"18",X"0A",X"25",X"11",X"F8",X"08",X"CD",X"11",X"3D",X"30",
		X"01",X"24",X"7D",X"FE",X"F8",X"C9",X"7E",X"D6",X"80",X"28",X"02",X"AF",X"C9",X"CD",X"70",X"3D",
		X"3E",X"01",X"37",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7D",X"E6",X"1F",X"07",X"07",X"07",X"4F",X"7D",X"E6",X"E0",X"6F",X"EB",X"21",X"00",X"4C",X"A7",
		X"ED",X"52",X"7D",X"84",X"0F",X"0F",X"47",X"3A",X"34",X"50",X"80",X"6F",X"61",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"27",X"32",X"59",X"50",X"32",X"5D",X"50",
		X"21",X"22",X"02",X"22",X"51",X"50",X"22",X"55",X"50",X"C3",X"4E",X"2F",X"3A",X"59",X"50",X"FE",
		X"A8",X"20",X"04",X"3A",X"5C",X"50",X"C9",X"F1",X"C3",X"B1",X"02",X"28",X"0A",X"3D",X"32",X"58",
		X"50",X"C6",X"10",X"32",X"5C",X"50",X"C9",X"3E",X"27",X"32",X"59",X"50",X"32",X"5D",X"50",X"3E",
		X"F8",X"32",X"5C",X"50",X"C9",X"3A",X"00",X"42",X"0F",X"D2",X"52",X"3D",X"3A",X"03",X"41",X"C3",
		X"37",X"3D",X"3E",X"F8",X"32",X"50",X"50",X"32",X"54",X"50",X"C3",X"FA",X"34",X"7B",X"FE",X"07",
		X"28",X"05",X"FE",X"26",X"C3",X"13",X"13",X"3E",X"01",X"32",X"04",X"60",X"C3",X"31",X"13",X"00",
		X"00",X"44",X"44",X"44",X"46",X"44",X"46",X"64",X"64",X"66",X"26",X"26",X"22",X"22",X"26",X"22",
		X"22",X"26",X"62",X"62",X"62",X"62",X"66",X"66",X"46",X"46",X"64",X"44",X"44",X"54",X"54",X"45",
		X"44",X"54",X"44",X"45",X"44",X"44",X"46",X"54",X"64",X"66",X"66",X"62",X"62",X"62",X"22",X"26",
		X"22",X"45",X"22",X"26",X"26",X"66",X"46",X"46",X"46",X"44",X"44",X"45",X"55",X"55",X"11",X"15",
		X"15",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"20",X"41",X"A7",X"C8",X"FE",X"12",X"D0",X"C3",X"96",X"A7",X"A7",X"28",X"5F",X"6F",X"26",
		X"3E",X"3A",X"44",X"40",X"FE",X"F0",X"28",X"0C",X"3E",X"F0",X"32",X"44",X"40",X"A6",X"0F",X"0F",
		X"0F",X"0F",X"18",X"11",X"7D",X"FE",X"7A",X"20",X"01",X"AF",X"3C",X"6F",X"32",X"43",X"40",X"3E",
		X"0F",X"32",X"44",X"40",X"A6",X"4F",X"CB",X"51",X"28",X"07",X"3A",X"53",X"50",X"3C",X"32",X"53",
		X"50",X"CB",X"49",X"20",X"09",X"CB",X"41",X"20",X"0D",X"3A",X"50",X"50",X"18",X"04",X"3A",X"50",
		X"50",X"3D",X"3D",X"32",X"50",X"50",X"3A",X"50",X"50",X"FE",X"F8",X"30",X"0C",X"3A",X"53",X"50",
		X"FE",X"C7",X"38",X"09",X"3E",X"F8",X"32",X"50",X"50",X"AF",X"32",X"43",X"40",X"3A",X"45",X"40",
		X"A7",X"28",X"63",X"6F",X"26",X"3E",X"3A",X"46",X"40",X"FE",X"F0",X"28",X"0C",X"3E",X"F0",X"32",
		X"46",X"40",X"A6",X"0F",X"0F",X"0F",X"0F",X"18",X"11",X"7D",X"FE",X"7A",X"20",X"01",X"AF",X"3C",
		X"6F",X"32",X"45",X"40",X"3E",X"0F",X"32",X"46",X"40",X"A6",X"4F",X"CB",X"51",X"28",X"07",X"3A",
		X"57",X"50",X"3C",X"32",X"57",X"50",X"CB",X"41",X"20",X"0A",X"CB",X"49",X"28",X"0D",X"3A",X"54",
		X"50",X"3C",X"18",X"04",X"3A",X"54",X"50",X"3D",X"32",X"54",X"50",X"3A",X"54",X"50",X"FE",X"F8",
		X"38",X"06",X"AF",X"32",X"45",X"40",X"18",X"0E",X"3A",X"57",X"50",X"FE",X"C7",X"38",X"07",X"3E",
		X"F8",X"32",X"54",X"50",X"18",X"EC",X"3A",X"47",X"40",X"A7",X"28",X"18",X"3A",X"50",X"50",X"6F",
		X"3A",X"53",X"50",X"CD",X"29",X"3D",X"38",X"04",X"AF",X"32",X"47",X"40",X"7D",X"32",X"50",X"50",
		X"7C",X"32",X"53",X"50",X"3A",X"48",X"40",X"A7",X"28",X"18",X"3A",X"54",X"50",X"6F",X"3A",X"57",
		X"50",X"CD",X"29",X"3D",X"38",X"04",X"AF",X"32",X"48",X"40",X"7D",X"32",X"54",X"50",X"7C",X"32",
		X"57",X"50",X"3A",X"59",X"50",X"FE",X"27",X"20",X"0F",X"3A",X"58",X"50",X"FE",X"F8",X"30",X"08",
		X"D6",X"04",X"CD",X"59",X"A0",X"32",X"58",X"50",X"3A",X"5D",X"50",X"FE",X"27",X"20",X"0C",X"3A",
		X"5C",X"50",X"FE",X"F8",X"30",X"05",X"D6",X"04",X"CD",X"65",X"A0",X"C3",X"97",X"1F",X"3A",X"20",
		X"41",X"FE",X"05",X"D2",X"0C",X"80",X"3A",X"43",X"40",X"A7",X"20",X"1A",X"3A",X"34",X"50",X"E6",
		X"08",X"28",X"13",X"2A",X"95",X"40",X"CD",X"56",X"3D",X"30",X"0B",X"32",X"43",X"40",X"7D",X"32",
		X"50",X"50",X"7C",X"32",X"53",X"50",X"3A",X"45",X"40",X"A7",X"C0",X"3A",X"34",X"50",X"E6",X"08",
		X"C0",X"2A",X"95",X"40",X"CD",X"56",X"3D",X"D0",X"C3",X"00",X"80",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
