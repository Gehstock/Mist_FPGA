-- Sixteen level by Three voice YM2149 volume_table[C][B][A]
-- Data measured by Paulo Simoes. Copyright 2012 Paulo Simoes.
-- original 16 bit data reduced to 10 bit

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity vol_table is
  port (
    CLK         : in    std_logic;
    ADDR_A      : in    std_logic_vector(11 downto 0);
    DATA_A      : out   std_logic_vector(9 downto 0);
    ADDR_B      : in    std_logic_vector(11 downto 0);
    DATA_B      : out   std_logic_vector(9 downto 0)
    );
end;

architecture RTL of vol_table is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(9 downto 0);
  constant voltable : ROM_ARRAY := (
	"00"&x"00","00"&x"01","00"&x"03","00"&x"06","00"&x"09","00"&x"0d","00"&x"13","00"&x"1a","00"&x"27","00"&x"36","00"&x"50","00"&x"6e","00"&x"a1","00"&x"e4","01"&x"66","10"&x"1a",
	"00"&x"01","00"&x"04","00"&x"06","00"&x"08","00"&x"0c","00"&x"0f","00"&x"16","00"&x"1d","00"&x"2a","00"&x"38","00"&x"52","00"&x"70","00"&x"a4","00"&x"e6","01"&x"67","10"&x"1a",
	"00"&x"03","00"&x"06","00"&x"08","00"&x"0a","00"&x"0e","00"&x"11","00"&x"18","00"&x"1f","00"&x"2c","00"&x"3a","00"&x"54","00"&x"72","00"&x"a5","00"&x"e8","01"&x"68","10"&x"1a",
	"00"&x"06","00"&x"08","00"&x"0a","00"&x"0c","00"&x"10","00"&x"14","00"&x"1a","00"&x"21","00"&x"2e","00"&x"3d","00"&x"56","00"&x"74","00"&x"a7","00"&x"e9","01"&x"69","10"&x"1b",
	"00"&x"09","00"&x"0c","00"&x"0e","00"&x"10","00"&x"13","00"&x"17","00"&x"1e","00"&x"25","00"&x"31","00"&x"40","00"&x"5a","00"&x"77","00"&x"aa","00"&x"ec","01"&x"6b","10"&x"1b",
	"00"&x"0d","00"&x"0f","00"&x"11","00"&x"14","00"&x"17","00"&x"1b","00"&x"21","00"&x"29","00"&x"35","00"&x"43","00"&x"5d","00"&x"7a","00"&x"ad","00"&x"ef","01"&x"6d","10"&x"1c",
	"00"&x"13","00"&x"16","00"&x"18","00"&x"1a","00"&x"1e","00"&x"21","00"&x"28","00"&x"2f","00"&x"3b","00"&x"4a","00"&x"63","00"&x"80","00"&x"b3","00"&x"f4","01"&x"71","10"&x"1d",
	"00"&x"1a","00"&x"1d","00"&x"1f","00"&x"21","00"&x"25","00"&x"29","00"&x"2f","00"&x"36","00"&x"42","00"&x"50","00"&x"6a","00"&x"85","00"&x"b9","00"&x"f9","01"&x"75","10"&x"1f",
	"00"&x"27","00"&x"2a","00"&x"2c","00"&x"2e","00"&x"31","00"&x"35","00"&x"3b","00"&x"42","00"&x"4e","00"&x"5c","00"&x"75","00"&x"90","00"&x"c3","01"&x"03","01"&x"7d","10"&x"22",
	"00"&x"36","00"&x"38","00"&x"3a","00"&x"3d","00"&x"40","00"&x"43","00"&x"4a","00"&x"50","00"&x"5c","00"&x"6a","00"&x"82","00"&x"9d","00"&x"d0","01"&x"0e","01"&x"87","10"&x"28",
	"00"&x"50","00"&x"52","00"&x"54","00"&x"56","00"&x"5a","00"&x"5d","00"&x"63","00"&x"6a","00"&x"75","00"&x"82","00"&x"98","00"&x"b4","00"&x"e6","01"&x"22","01"&x"99","10"&x"34",
	"00"&x"6e","00"&x"70","00"&x"72","00"&x"74","00"&x"77","00"&x"7a","00"&x"80","00"&x"85","00"&x"90","00"&x"9d","00"&x"b4","00"&x"cf","01"&x"01","01"&x"3b","01"&x"af","10"&x"44",
	"00"&x"a1","00"&x"a4","00"&x"a5","00"&x"a7","00"&x"aa","00"&x"ad","00"&x"b3","00"&x"b9","00"&x"c3","00"&x"d0","00"&x"e6","01"&x"01","01"&x"2f","01"&x"6a","01"&x"dc","10"&x"69",
	"00"&x"e4","00"&x"e6","00"&x"e8","00"&x"e9","00"&x"ec","00"&x"ef","00"&x"f4","00"&x"f9","01"&x"03","01"&x"0e","01"&x"22","01"&x"3b","01"&x"6a","01"&x"a3","10"&x"14","10"&x"9a",
	"01"&x"66","01"&x"67","01"&x"68","01"&x"69","01"&x"6b","01"&x"6d","01"&x"71","01"&x"75","01"&x"7d","01"&x"87","01"&x"99","01"&x"af","01"&x"dc","10"&x"14","10"&x"79","10"&x"f3",
	"10"&x"1a","10"&x"1a","10"&x"1a","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1d","10"&x"1f","10"&x"22","10"&x"28","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"01","00"&x"04","00"&x"06","00"&x"08","00"&x"0c","00"&x"0f","00"&x"16","00"&x"1d","00"&x"2a","00"&x"38","00"&x"52","00"&x"70","00"&x"a4","00"&x"e6","01"&x"67","10"&x"1a",
	"00"&x"04","00"&x"07","00"&x"09","00"&x"0b","00"&x"0e","00"&x"12","00"&x"19","00"&x"20","00"&x"2c","00"&x"3b","00"&x"55","00"&x"72","00"&x"a6","00"&x"e8","01"&x"68","10"&x"1b",
	"00"&x"06","00"&x"09","00"&x"0b","00"&x"0d","00"&x"10","00"&x"14","00"&x"1b","00"&x"22","00"&x"2e","00"&x"3d","00"&x"57","00"&x"74","00"&x"a8","00"&x"ea","01"&x"6a","10"&x"1b",
	"00"&x"08","00"&x"0b","00"&x"0d","00"&x"0f","00"&x"12","00"&x"16","00"&x"1d","00"&x"24","00"&x"30","00"&x"3f","00"&x"59","00"&x"76","00"&x"a9","00"&x"eb","01"&x"6b","10"&x"1b",
	"00"&x"0c","00"&x"0e","00"&x"10","00"&x"12","00"&x"16","00"&x"1a","00"&x"20","00"&x"27","00"&x"34","00"&x"42","00"&x"5c","00"&x"79","00"&x"ac","00"&x"ee","01"&x"6c","10"&x"1b",
	"00"&x"0f","00"&x"12","00"&x"14","00"&x"16","00"&x"1a","00"&x"1d","00"&x"24","00"&x"2b","00"&x"37","00"&x"46","00"&x"5f","00"&x"7c","00"&x"af","00"&x"f1","01"&x"6e","10"&x"1c",
	"00"&x"16","00"&x"19","00"&x"1b","00"&x"1d","00"&x"20","00"&x"24","00"&x"2a","00"&x"31","00"&x"3e","00"&x"4c","00"&x"65","00"&x"81","00"&x"b5","00"&x"f5","01"&x"72","10"&x"1d",
	"00"&x"1d","00"&x"20","00"&x"22","00"&x"24","00"&x"27","00"&x"2b","00"&x"31","00"&x"39","00"&x"45","00"&x"53","00"&x"6c","00"&x"87","00"&x"bb","00"&x"fb","01"&x"77","10"&x"1f",
	"00"&x"2a","00"&x"2c","00"&x"2e","00"&x"30","00"&x"34","00"&x"37","00"&x"3e","00"&x"45","00"&x"51","00"&x"5f","00"&x"78","00"&x"92","00"&x"c5","01"&x"05","01"&x"7f","10"&x"22",
	"00"&x"38","00"&x"3b","00"&x"3d","00"&x"3f","00"&x"42","00"&x"46","00"&x"4c","00"&x"53","00"&x"5f","00"&x"6d","00"&x"84","00"&x"9f","00"&x"d2","01"&x"0f","01"&x"88","10"&x"28",
	"00"&x"52","00"&x"55","00"&x"57","00"&x"59","00"&x"5c","00"&x"5f","00"&x"65","00"&x"6c","00"&x"78","00"&x"84","00"&x"9a","00"&x"b6","00"&x"e8","01"&x"24","01"&x"9a","10"&x"34",
	"00"&x"70","00"&x"72","00"&x"74","00"&x"76","00"&x"79","00"&x"7c","00"&x"81","00"&x"87","00"&x"92","00"&x"9f","00"&x"b6","00"&x"d1","01"&x"02","01"&x"3d","01"&x"b0","10"&x"44",
	"00"&x"a4","00"&x"a6","00"&x"a8","00"&x"a9","00"&x"ac","00"&x"af","00"&x"b5","00"&x"bb","00"&x"c5","00"&x"d2","00"&x"e8","01"&x"02","01"&x"31","01"&x"6c","01"&x"dc","10"&x"69",
	"00"&x"e6","00"&x"e8","00"&x"ea","00"&x"eb","00"&x"ee","00"&x"f1","00"&x"f5","00"&x"fb","01"&x"05","01"&x"0f","01"&x"24","01"&x"3d","01"&x"6c","01"&x"a4","10"&x"14","10"&x"9a",
	"01"&x"67","01"&x"68","01"&x"6a","01"&x"6b","01"&x"6c","01"&x"6e","01"&x"72","01"&x"77","01"&x"7f","01"&x"88","01"&x"9a","01"&x"b0","01"&x"dc","10"&x"14","10"&x"79","10"&x"f3",
	"10"&x"1a","10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1d","10"&x"1f","10"&x"22","10"&x"28","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"03","00"&x"06","00"&x"08","00"&x"0a","00"&x"0e","00"&x"11","00"&x"18","00"&x"1f","00"&x"2c","00"&x"3a","00"&x"54","00"&x"72","00"&x"a5","00"&x"e8","01"&x"68","10"&x"1a",
	"00"&x"06","00"&x"09","00"&x"0b","00"&x"0d","00"&x"10","00"&x"14","00"&x"1b","00"&x"22","00"&x"2e","00"&x"3d","00"&x"57","00"&x"74","00"&x"a8","00"&x"ea","01"&x"6a","10"&x"1b",
	"00"&x"08","00"&x"0b","00"&x"0d","00"&x"0f","00"&x"12","00"&x"16","00"&x"1d","00"&x"24","00"&x"30","00"&x"3f","00"&x"59","00"&x"76","00"&x"a9","00"&x"eb","01"&x"6b","10"&x"1b",
	"00"&x"0a","00"&x"0d","00"&x"0f","00"&x"11","00"&x"15","00"&x"18","00"&x"1f","00"&x"26","00"&x"33","00"&x"41","00"&x"5b","00"&x"78","00"&x"ab","00"&x"ed","01"&x"6c","10"&x"1b",
	"00"&x"0e","00"&x"10","00"&x"12","00"&x"15","00"&x"18","00"&x"1c","00"&x"22","00"&x"2a","00"&x"36","00"&x"44","00"&x"5e","00"&x"7b","00"&x"ae","00"&x"ef","01"&x"6e","10"&x"1c",
	"00"&x"11","00"&x"14","00"&x"16","00"&x"18","00"&x"1c","00"&x"20","00"&x"26","00"&x"2d","00"&x"3a","00"&x"48","00"&x"61","00"&x"7e","00"&x"b1","00"&x"f2","01"&x"70","10"&x"1c",
	"00"&x"18","00"&x"1b","00"&x"1d","00"&x"1f","00"&x"22","00"&x"26","00"&x"2c","00"&x"33","00"&x"40","00"&x"4e","00"&x"67","00"&x"83","00"&x"b6","00"&x"f7","01"&x"73","10"&x"1d",
	"00"&x"1f","00"&x"22","00"&x"24","00"&x"26","00"&x"2a","00"&x"2d","00"&x"33","00"&x"3b","00"&x"47","00"&x"55","00"&x"6e","00"&x"89","00"&x"bd","00"&x"fc","01"&x"78","10"&x"1f",
	"00"&x"2c","00"&x"2e","00"&x"30","00"&x"33","00"&x"36","00"&x"3a","00"&x"40","00"&x"47","00"&x"53","00"&x"61","00"&x"79","00"&x"94","00"&x"c7","01"&x"06","01"&x"7f","10"&x"23",
	"00"&x"3a","00"&x"3d","00"&x"3f","00"&x"41","00"&x"44","00"&x"48","00"&x"4e","00"&x"55","00"&x"61","00"&x"6f","00"&x"85","00"&x"a1","00"&x"d4","01"&x"10","01"&x"89","10"&x"28",
	"00"&x"54","00"&x"57","00"&x"59","00"&x"5b","00"&x"5e","00"&x"61","00"&x"67","00"&x"6e","00"&x"79","00"&x"85","00"&x"9c","00"&x"b8","00"&x"ea","01"&x"25","01"&x"9b","10"&x"34",
	"00"&x"72","00"&x"74","00"&x"76","00"&x"78","00"&x"7b","00"&x"7e","00"&x"83","00"&x"89","00"&x"94","00"&x"a1","00"&x"b8","00"&x"d3","01"&x"04","01"&x"3e","01"&x"b1","10"&x"44",
	"00"&x"a5","00"&x"a8","00"&x"a9","00"&x"ab","00"&x"ae","00"&x"b1","00"&x"b6","00"&x"bd","00"&x"c7","00"&x"d4","00"&x"ea","01"&x"04","01"&x"32","01"&x"6c","01"&x"dd","10"&x"69",
	"00"&x"e8","00"&x"ea","00"&x"eb","00"&x"ed","00"&x"ef","00"&x"f2","00"&x"f7","00"&x"fc","01"&x"06","01"&x"10","01"&x"25","01"&x"3e","01"&x"6c","01"&x"a5","10"&x"15","10"&x"9a",
	"01"&x"68","01"&x"6a","01"&x"6b","01"&x"6c","01"&x"6e","01"&x"70","01"&x"73","01"&x"78","01"&x"7f","01"&x"89","01"&x"9b","01"&x"b1","01"&x"dd","10"&x"15","10"&x"79","10"&x"f3",
	"10"&x"1a","10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1c","10"&x"1d","10"&x"1f","10"&x"23","10"&x"28","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"06","00"&x"08","00"&x"0a","00"&x"0c","00"&x"10","00"&x"14","00"&x"1a","00"&x"21","00"&x"2e","00"&x"3d","00"&x"56","00"&x"74","00"&x"a7","00"&x"e9","01"&x"69","10"&x"1b",
	"00"&x"08","00"&x"0b","00"&x"0d","00"&x"0f","00"&x"12","00"&x"16","00"&x"1d","00"&x"24","00"&x"30","00"&x"3f","00"&x"59","00"&x"76","00"&x"a9","00"&x"eb","01"&x"6b","10"&x"1b",
	"00"&x"0a","00"&x"0d","00"&x"0f","00"&x"11","00"&x"15","00"&x"18","00"&x"1f","00"&x"26","00"&x"33","00"&x"41","00"&x"5b","00"&x"78","00"&x"ab","00"&x"ed","01"&x"6c","10"&x"1b",
	"00"&x"0c","00"&x"0f","00"&x"11","00"&x"13","00"&x"17","00"&x"1b","00"&x"21","00"&x"28","00"&x"35","00"&x"43","00"&x"5d","00"&x"7a","00"&x"ad","00"&x"ee","01"&x"6d","10"&x"1c",
	"00"&x"10","00"&x"12","00"&x"15","00"&x"17","00"&x"1a","00"&x"1e","00"&x"24","00"&x"2c","00"&x"38","00"&x"46","00"&x"60","00"&x"7d","00"&x"b0","00"&x"f1","01"&x"6f","10"&x"1c",
	"00"&x"14","00"&x"16","00"&x"18","00"&x"1b","00"&x"1e","00"&x"22","00"&x"28","00"&x"2f","00"&x"3c","00"&x"4a","00"&x"63","00"&x"80","00"&x"b3","00"&x"f4","01"&x"71","10"&x"1c",
	"00"&x"1a","00"&x"1d","00"&x"1f","00"&x"21","00"&x"24","00"&x"28","00"&x"2e","00"&x"35","00"&x"42","00"&x"50","00"&x"69","00"&x"84","00"&x"b8","00"&x"f8","01"&x"74","10"&x"1e",
	"00"&x"21","00"&x"24","00"&x"26","00"&x"28","00"&x"2c","00"&x"2f","00"&x"35","00"&x"3d","00"&x"49","00"&x"57","00"&x"70","00"&x"8a","00"&x"be","00"&x"fe","01"&x"79","10"&x"1f",
	"00"&x"2e","00"&x"30","00"&x"33","00"&x"35","00"&x"38","00"&x"3c","00"&x"42","00"&x"49","00"&x"55","00"&x"63","00"&x"7b","00"&x"95","00"&x"c9","01"&x"08","01"&x"80","10"&x"23",
	"00"&x"3d","00"&x"3f","00"&x"41","00"&x"43","00"&x"46","00"&x"4a","00"&x"50","00"&x"57","00"&x"63","00"&x"71","00"&x"87","00"&x"a3","00"&x"d5","01"&x"12","01"&x"8a","10"&x"29",
	"00"&x"56","00"&x"59","00"&x"5b","00"&x"5d","00"&x"60","00"&x"63","00"&x"69","00"&x"70","00"&x"7b","00"&x"87","00"&x"9e","00"&x"b9","00"&x"eb","01"&x"26","01"&x"9c","10"&x"34",
	"00"&x"74","00"&x"76","00"&x"78","00"&x"7a","00"&x"7d","00"&x"80","00"&x"84","00"&x"8a","00"&x"95","00"&x"a3","00"&x"b9","00"&x"d4","01"&x"05","01"&x"3f","01"&x"b1","10"&x"44",
	"00"&x"a7","00"&x"a9","00"&x"ab","00"&x"ad","00"&x"b0","00"&x"b3","00"&x"b8","00"&x"be","00"&x"c9","00"&x"d5","00"&x"eb","01"&x"05","01"&x"33","01"&x"6d","01"&x"dd","10"&x"69",
	"00"&x"e9","00"&x"eb","00"&x"ed","00"&x"ee","00"&x"f1","00"&x"f4","00"&x"f8","00"&x"fe","01"&x"08","01"&x"12","01"&x"26","01"&x"3f","01"&x"6d","01"&x"a5","10"&x"15","10"&x"9a",
	"01"&x"69","01"&x"6b","01"&x"6c","01"&x"6d","01"&x"6f","01"&x"71","01"&x"74","01"&x"79","01"&x"80","01"&x"8a","01"&x"9c","01"&x"b1","01"&x"dd","10"&x"15","10"&x"79","10"&x"f3",
	"10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1e","10"&x"1f","10"&x"23","10"&x"29","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"09","00"&x"0c","00"&x"0e","00"&x"10","00"&x"13","00"&x"17","00"&x"1e","00"&x"25","00"&x"31","00"&x"40","00"&x"5a","00"&x"77","00"&x"aa","00"&x"ec","01"&x"6b","10"&x"1b",
	"00"&x"0c","00"&x"0e","00"&x"10","00"&x"12","00"&x"16","00"&x"1a","00"&x"20","00"&x"27","00"&x"34","00"&x"42","00"&x"5c","00"&x"79","00"&x"ac","00"&x"ee","01"&x"6c","10"&x"1b",
	"00"&x"0e","00"&x"10","00"&x"12","00"&x"15","00"&x"18","00"&x"1c","00"&x"22","00"&x"2a","00"&x"36","00"&x"44","00"&x"5e","00"&x"7b","00"&x"ae","00"&x"ef","01"&x"6e","10"&x"1c",
	"00"&x"10","00"&x"12","00"&x"15","00"&x"17","00"&x"1a","00"&x"1e","00"&x"24","00"&x"2c","00"&x"38","00"&x"46","00"&x"60","00"&x"7d","00"&x"b0","00"&x"f1","01"&x"6f","10"&x"1c",
	"00"&x"13","00"&x"16","00"&x"18","00"&x"1a","00"&x"1d","00"&x"21","00"&x"28","00"&x"2f","00"&x"3b","00"&x"4a","00"&x"63","00"&x"80","00"&x"b2","00"&x"f3","01"&x"70","10"&x"1c",
	"00"&x"17","00"&x"1a","00"&x"1c","00"&x"1e","00"&x"21","00"&x"25","00"&x"2c","00"&x"32","00"&x"3f","00"&x"4d","00"&x"66","00"&x"82","00"&x"b6","00"&x"f6","01"&x"72","10"&x"1d",
	"00"&x"1e","00"&x"20","00"&x"22","00"&x"24","00"&x"28","00"&x"2c","00"&x"32","00"&x"39","00"&x"45","00"&x"53","00"&x"6c","00"&x"87","00"&x"bb","00"&x"fb","01"&x"76","10"&x"1e",
	"00"&x"25","00"&x"27","00"&x"2a","00"&x"2c","00"&x"2f","00"&x"32","00"&x"39","00"&x"40","00"&x"4c","00"&x"5a","00"&x"73","00"&x"8d","00"&x"c1","01"&x"00","01"&x"7a","10"&x"20",
	"00"&x"31","00"&x"34","00"&x"36","00"&x"38","00"&x"3b","00"&x"3f","00"&x"45","00"&x"4c","00"&x"58","00"&x"66","00"&x"7e","00"&x"98","00"&x"cb","01"&x"0a","01"&x"82","10"&x"23",
	"00"&x"40","00"&x"42","00"&x"44","00"&x"46","00"&x"4a","00"&x"4d","00"&x"53","00"&x"5a","00"&x"66","00"&x"74","00"&x"8a","00"&x"a5","00"&x"d8","01"&x"14","01"&x"8c","10"&x"29",
	"00"&x"5a","00"&x"5c","00"&x"5e","00"&x"60","00"&x"63","00"&x"66","00"&x"6c","00"&x"73","00"&x"7e","00"&x"8a","00"&x"a1","00"&x"bc","00"&x"ed","01"&x"28","01"&x"9d","10"&x"34",
	"00"&x"77","00"&x"79","00"&x"7b","00"&x"7d","00"&x"80","00"&x"82","00"&x"87","00"&x"8d","00"&x"98","00"&x"a5","00"&x"bc","00"&x"d7","01"&x"07","01"&x"41","01"&x"b2","10"&x"44",
	"00"&x"aa","00"&x"ac","00"&x"ae","00"&x"b0","00"&x"b2","00"&x"b6","00"&x"bb","00"&x"c1","00"&x"cb","00"&x"d8","00"&x"ed","01"&x"07","01"&x"35","01"&x"6f","01"&x"de","10"&x"69",
	"00"&x"ec","00"&x"ee","00"&x"ef","00"&x"f1","00"&x"f3","00"&x"f6","00"&x"fb","01"&x"00","01"&x"0a","01"&x"14","01"&x"28","01"&x"41","01"&x"6f","01"&x"a6","10"&x"15","10"&x"9a",
	"01"&x"6b","01"&x"6c","01"&x"6e","01"&x"6f","01"&x"70","01"&x"72","01"&x"76","01"&x"7a","01"&x"82","01"&x"8c","01"&x"9d","01"&x"b2","01"&x"de","10"&x"15","10"&x"79","10"&x"f3",
	"10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1d","10"&x"1e","10"&x"20","10"&x"23","10"&x"29","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"0d","00"&x"0f","00"&x"11","00"&x"14","00"&x"17","00"&x"1b","00"&x"21","00"&x"29","00"&x"35","00"&x"43","00"&x"5d","00"&x"7a","00"&x"ad","00"&x"ef","01"&x"6d","10"&x"1c",
	"00"&x"0f","00"&x"12","00"&x"14","00"&x"16","00"&x"1a","00"&x"1d","00"&x"24","00"&x"2b","00"&x"37","00"&x"46","00"&x"5f","00"&x"7c","00"&x"af","00"&x"f1","01"&x"6e","10"&x"1c",
	"00"&x"11","00"&x"14","00"&x"16","00"&x"18","00"&x"1c","00"&x"20","00"&x"26","00"&x"2d","00"&x"3a","00"&x"48","00"&x"61","00"&x"7e","00"&x"b1","00"&x"f2","01"&x"70","10"&x"1c",
	"00"&x"14","00"&x"16","00"&x"18","00"&x"1b","00"&x"1e","00"&x"22","00"&x"28","00"&x"2f","00"&x"3c","00"&x"4a","00"&x"63","00"&x"80","00"&x"b3","00"&x"f4","01"&x"71","10"&x"1c",
	"00"&x"17","00"&x"1a","00"&x"1c","00"&x"1e","00"&x"21","00"&x"25","00"&x"2c","00"&x"32","00"&x"3f","00"&x"4d","00"&x"66","00"&x"82","00"&x"b6","00"&x"f6","01"&x"72","10"&x"1d",
	"00"&x"1b","00"&x"1d","00"&x"20","00"&x"22","00"&x"25","00"&x"29","00"&x"2f","00"&x"36","00"&x"42","00"&x"51","00"&x"6a","00"&x"85","00"&x"b9","00"&x"f9","01"&x"74","10"&x"1e",
	"00"&x"21","00"&x"24","00"&x"26","00"&x"28","00"&x"2c","00"&x"2f","00"&x"35","00"&x"3c","00"&x"48","00"&x"57","00"&x"70","00"&x"8a","00"&x"be","00"&x"fe","01"&x"78","10"&x"1f",
	"00"&x"29","00"&x"2b","00"&x"2d","00"&x"2f","00"&x"32","00"&x"36","00"&x"3c","00"&x"43","00"&x"4f","00"&x"5d","00"&x"76","00"&x"90","00"&x"c4","01"&x"03","01"&x"7c","10"&x"20",
	"00"&x"35","00"&x"37","00"&x"3a","00"&x"3c","00"&x"3f","00"&x"42","00"&x"48","00"&x"4f","00"&x"5b","00"&x"69","00"&x"81","00"&x"9b","00"&x"ce","01"&x"0c","01"&x"84","10"&x"24",
	"00"&x"43","00"&x"46","00"&x"48","00"&x"4a","00"&x"4d","00"&x"51","00"&x"57","00"&x"5d","00"&x"69","00"&x"77","00"&x"8d","00"&x"a8","00"&x"db","01"&x"16","01"&x"8e","10"&x"29",
	"00"&x"5d","00"&x"5f","00"&x"61","00"&x"63","00"&x"66","00"&x"6a","00"&x"70","00"&x"76","00"&x"81","00"&x"8d","00"&x"a4","00"&x"bf","00"&x"f0","01"&x"2a","01"&x"9f","10"&x"35",
	"00"&x"7a","00"&x"7c","00"&x"7e","00"&x"80","00"&x"82","00"&x"85","00"&x"8a","00"&x"90","00"&x"9b","00"&x"a8","00"&x"bf","00"&x"da","01"&x"09","01"&x"43","01"&x"b4","10"&x"44",
	"00"&x"ad","00"&x"af","00"&x"b1","00"&x"b3","00"&x"b6","00"&x"b9","00"&x"be","00"&x"c4","00"&x"ce","00"&x"db","00"&x"f0","01"&x"09","01"&x"37","01"&x"71","01"&x"df","10"&x"69",
	"00"&x"ef","00"&x"f1","00"&x"f2","00"&x"f4","00"&x"f6","00"&x"f9","00"&x"fe","01"&x"03","01"&x"0c","01"&x"16","01"&x"2a","01"&x"43","01"&x"71","01"&x"a8","10"&x"16","10"&x"9a",
	"01"&x"6d","01"&x"6e","01"&x"70","01"&x"71","01"&x"72","01"&x"74","01"&x"78","01"&x"7c","01"&x"84","01"&x"8e","01"&x"9f","01"&x"b4","01"&x"df","10"&x"16","10"&x"79","10"&x"f3",
	"10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1d","10"&x"1e","10"&x"1f","10"&x"20","10"&x"24","10"&x"29","10"&x"35","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"13","00"&x"16","00"&x"18","00"&x"1a","00"&x"1e","00"&x"21","00"&x"28","00"&x"2f","00"&x"3b","00"&x"4a","00"&x"63","00"&x"80","00"&x"b3","00"&x"f4","01"&x"71","10"&x"1d",
	"00"&x"16","00"&x"19","00"&x"1b","00"&x"1d","00"&x"20","00"&x"24","00"&x"2a","00"&x"31","00"&x"3e","00"&x"4c","00"&x"65","00"&x"81","00"&x"b5","00"&x"f5","01"&x"72","10"&x"1d",
	"00"&x"18","00"&x"1b","00"&x"1d","00"&x"1f","00"&x"22","00"&x"26","00"&x"2c","00"&x"33","00"&x"40","00"&x"4e","00"&x"67","00"&x"83","00"&x"b6","00"&x"f7","01"&x"73","10"&x"1d",
	"00"&x"1a","00"&x"1d","00"&x"1f","00"&x"21","00"&x"24","00"&x"28","00"&x"2e","00"&x"35","00"&x"42","00"&x"50","00"&x"69","00"&x"84","00"&x"b8","00"&x"f8","01"&x"74","10"&x"1e",
	"00"&x"1e","00"&x"20","00"&x"22","00"&x"24","00"&x"28","00"&x"2c","00"&x"32","00"&x"39","00"&x"45","00"&x"53","00"&x"6c","00"&x"87","00"&x"bb","00"&x"fb","01"&x"76","10"&x"1e",
	"00"&x"21","00"&x"24","00"&x"26","00"&x"28","00"&x"2c","00"&x"2f","00"&x"35","00"&x"3c","00"&x"48","00"&x"57","00"&x"70","00"&x"8a","00"&x"be","00"&x"fe","01"&x"78","10"&x"1f",
	"00"&x"28","00"&x"2a","00"&x"2c","00"&x"2e","00"&x"32","00"&x"35","00"&x"3c","00"&x"43","00"&x"4f","00"&x"5d","00"&x"75","00"&x"90","00"&x"c3","01"&x"02","01"&x"7c","10"&x"20",
	"00"&x"2f","00"&x"31","00"&x"33","00"&x"35","00"&x"39","00"&x"3c","00"&x"43","00"&x"4a","00"&x"55","00"&x"63","00"&x"7c","00"&x"96","00"&x"c9","01"&x"08","01"&x"80","10"&x"21",
	"00"&x"3b","00"&x"3e","00"&x"40","00"&x"42","00"&x"45","00"&x"48","00"&x"4f","00"&x"55","00"&x"61","00"&x"6f","00"&x"85","00"&x"a1","00"&x"d3","01"&x"10","01"&x"87","10"&x"25",
	"00"&x"4a","00"&x"4c","00"&x"4e","00"&x"50","00"&x"53","00"&x"57","00"&x"5d","00"&x"63","00"&x"6f","00"&x"7d","00"&x"92","00"&x"ae","00"&x"e0","01"&x"1b","01"&x"91","10"&x"2a",
	"00"&x"63","00"&x"65","00"&x"67","00"&x"69","00"&x"6c","00"&x"70","00"&x"75","00"&x"7c","00"&x"85","00"&x"92","00"&x"a9","00"&x"c4","00"&x"f5","01"&x"2f","01"&x"a1","10"&x"35",
	"00"&x"80","00"&x"81","00"&x"83","00"&x"84","00"&x"87","00"&x"8a","00"&x"90","00"&x"96","00"&x"a1","00"&x"ae","00"&x"c4","00"&x"df","01"&x"0d","01"&x"47","01"&x"b6","10"&x"45",
	"00"&x"b3","00"&x"b5","00"&x"b6","00"&x"b8","00"&x"bb","00"&x"be","00"&x"c3","00"&x"c9","00"&x"d3","00"&x"e0","00"&x"f5","01"&x"0d","01"&x"3b","01"&x"74","01"&x"e0","10"&x"69",
	"00"&x"f4","00"&x"f5","00"&x"f7","00"&x"f8","00"&x"fb","00"&x"fe","01"&x"02","01"&x"08","01"&x"10","01"&x"1b","01"&x"2f","01"&x"47","01"&x"74","01"&x"aa","10"&x"17","10"&x"9a",
	"01"&x"71","01"&x"72","01"&x"73","01"&x"74","01"&x"76","01"&x"78","01"&x"7c","01"&x"80","01"&x"87","01"&x"91","01"&x"a1","01"&x"b6","01"&x"e0","10"&x"17","10"&x"79","10"&x"f3",
	"10"&x"1d","10"&x"1d","10"&x"1d","10"&x"1e","10"&x"1e","10"&x"1f","10"&x"20","10"&x"21","10"&x"25","10"&x"2a","10"&x"35","10"&x"45","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"1a","00"&x"1d","00"&x"1f","00"&x"21","00"&x"25","00"&x"29","00"&x"2f","00"&x"36","00"&x"42","00"&x"50","00"&x"6a","00"&x"85","00"&x"b9","00"&x"f9","01"&x"75","10"&x"1f",
	"00"&x"1d","00"&x"20","00"&x"22","00"&x"24","00"&x"27","00"&x"2b","00"&x"31","00"&x"39","00"&x"45","00"&x"53","00"&x"6c","00"&x"87","00"&x"bb","00"&x"fb","01"&x"77","10"&x"1f",
	"00"&x"1f","00"&x"22","00"&x"24","00"&x"26","00"&x"2a","00"&x"2d","00"&x"33","00"&x"3b","00"&x"47","00"&x"55","00"&x"6e","00"&x"89","00"&x"bd","00"&x"fc","01"&x"78","10"&x"1f",
	"00"&x"21","00"&x"24","00"&x"26","00"&x"28","00"&x"2c","00"&x"2f","00"&x"35","00"&x"3d","00"&x"49","00"&x"57","00"&x"70","00"&x"8a","00"&x"be","00"&x"fe","01"&x"79","10"&x"1f",
	"00"&x"25","00"&x"27","00"&x"2a","00"&x"2c","00"&x"2f","00"&x"32","00"&x"39","00"&x"40","00"&x"4c","00"&x"5a","00"&x"73","00"&x"8d","00"&x"c1","01"&x"00","01"&x"7a","10"&x"20",
	"00"&x"29","00"&x"2b","00"&x"2d","00"&x"2f","00"&x"32","00"&x"36","00"&x"3c","00"&x"43","00"&x"4f","00"&x"5d","00"&x"76","00"&x"90","00"&x"c4","01"&x"03","01"&x"7c","10"&x"20",
	"00"&x"2f","00"&x"31","00"&x"33","00"&x"35","00"&x"39","00"&x"3c","00"&x"43","00"&x"4a","00"&x"55","00"&x"63","00"&x"7c","00"&x"96","00"&x"c9","01"&x"08","01"&x"80","10"&x"21",
	"00"&x"36","00"&x"39","00"&x"3b","00"&x"3d","00"&x"40","00"&x"43","00"&x"4a","00"&x"50","00"&x"5c","00"&x"6a","00"&x"82","00"&x"9c","00"&x"cf","01"&x"0c","01"&x"84","10"&x"23",
	"00"&x"42","00"&x"45","00"&x"47","00"&x"49","00"&x"4c","00"&x"4f","00"&x"55","00"&x"5c","00"&x"68","00"&x"76","00"&x"8c","00"&x"a7","00"&x"d9","01"&x"15","01"&x"8b","10"&x"26",
	"00"&x"50","00"&x"53","00"&x"55","00"&x"57","00"&x"5a","00"&x"5d","00"&x"63","00"&x"6a","00"&x"76","00"&x"82","00"&x"99","00"&x"b4","00"&x"e5","01"&x"20","01"&x"94","10"&x"2c",
	"00"&x"6a","00"&x"6c","00"&x"6e","00"&x"70","00"&x"73","00"&x"76","00"&x"7c","00"&x"82","00"&x"8c","00"&x"99","00"&x"af","00"&x"ca","00"&x"fa","01"&x"33","01"&x"a4","10"&x"36",
	"00"&x"85","00"&x"87","00"&x"89","00"&x"8a","00"&x"8d","00"&x"90","00"&x"96","00"&x"9c","00"&x"a7","00"&x"b4","00"&x"ca","00"&x"e4","01"&x"11","01"&x"4b","01"&x"b9","10"&x"46",
	"00"&x"b9","00"&x"bb","00"&x"bd","00"&x"be","00"&x"c1","00"&x"c4","00"&x"c9","00"&x"cf","00"&x"d9","00"&x"e5","00"&x"fa","01"&x"11","01"&x"3f","01"&x"78","01"&x"e3","10"&x"6a",
	"00"&x"f9","00"&x"fb","00"&x"fc","00"&x"fe","01"&x"00","01"&x"03","01"&x"08","01"&x"0c","01"&x"15","01"&x"20","01"&x"33","01"&x"4b","01"&x"78","01"&x"ad","10"&x"18","10"&x"9a",
	"01"&x"75","01"&x"77","01"&x"78","01"&x"79","01"&x"7a","01"&x"7c","01"&x"80","01"&x"84","01"&x"8b","01"&x"94","01"&x"a4","01"&x"b9","01"&x"e3","10"&x"18","10"&x"79","10"&x"f3",
	"10"&x"1f","10"&x"1f","10"&x"1f","10"&x"1f","10"&x"20","10"&x"20","10"&x"21","10"&x"23","10"&x"26","10"&x"2c","10"&x"36","10"&x"46","10"&x"6a","10"&x"9a","10"&x"f3","11"&x"61",
	"00"&x"27","00"&x"2a","00"&x"2c","00"&x"2e","00"&x"31","00"&x"35","00"&x"3b","00"&x"42","00"&x"4e","00"&x"5c","00"&x"75","00"&x"90","00"&x"c3","01"&x"03","01"&x"7d","10"&x"22",
	"00"&x"2a","00"&x"2c","00"&x"2e","00"&x"30","00"&x"34","00"&x"37","00"&x"3e","00"&x"45","00"&x"51","00"&x"5f","00"&x"78","00"&x"92","00"&x"c5","01"&x"05","01"&x"7f","10"&x"22",
	"00"&x"2c","00"&x"2e","00"&x"30","00"&x"33","00"&x"36","00"&x"3a","00"&x"40","00"&x"47","00"&x"53","00"&x"61","00"&x"79","00"&x"94","00"&x"c7","01"&x"06","01"&x"7f","10"&x"23",
	"00"&x"2e","00"&x"30","00"&x"33","00"&x"35","00"&x"38","00"&x"3c","00"&x"42","00"&x"49","00"&x"55","00"&x"63","00"&x"7b","00"&x"95","00"&x"c9","01"&x"08","01"&x"80","10"&x"23",
	"00"&x"31","00"&x"34","00"&x"36","00"&x"38","00"&x"3b","00"&x"3f","00"&x"45","00"&x"4c","00"&x"58","00"&x"66","00"&x"7e","00"&x"98","00"&x"cb","01"&x"0a","01"&x"82","10"&x"23",
	"00"&x"35","00"&x"37","00"&x"3a","00"&x"3c","00"&x"3f","00"&x"42","00"&x"48","00"&x"4f","00"&x"5b","00"&x"69","00"&x"81","00"&x"9b","00"&x"ce","01"&x"0c","01"&x"84","10"&x"24",
	"00"&x"3b","00"&x"3e","00"&x"40","00"&x"42","00"&x"45","00"&x"48","00"&x"4f","00"&x"55","00"&x"61","00"&x"6f","00"&x"85","00"&x"a1","00"&x"d3","01"&x"10","01"&x"87","10"&x"25",
	"00"&x"42","00"&x"45","00"&x"47","00"&x"49","00"&x"4c","00"&x"4f","00"&x"55","00"&x"5c","00"&x"68","00"&x"76","00"&x"8c","00"&x"a7","00"&x"d9","01"&x"15","01"&x"8b","10"&x"26",
	"00"&x"4e","00"&x"51","00"&x"53","00"&x"55","00"&x"58","00"&x"5b","00"&x"61","00"&x"68","00"&x"74","00"&x"81","00"&x"97","00"&x"b2","00"&x"e3","01"&x"1e","01"&x"92","10"&x"2a",
	"00"&x"5c","00"&x"5f","00"&x"61","00"&x"63","00"&x"66","00"&x"69","00"&x"6f","00"&x"76","00"&x"81","00"&x"8c","00"&x"a3","00"&x"be","00"&x"ef","01"&x"29","01"&x"9b","10"&x"2f",
	"00"&x"75","00"&x"78","00"&x"79","00"&x"7b","00"&x"7e","00"&x"81","00"&x"85","00"&x"8c","00"&x"97","00"&x"a3","00"&x"ba","00"&x"d4","01"&x"03","01"&x"3c","01"&x"aa","10"&x"39",
	"00"&x"90","00"&x"92","00"&x"94","00"&x"95","00"&x"98","00"&x"9b","00"&x"a1","00"&x"a7","00"&x"b2","00"&x"be","00"&x"d4","00"&x"ee","01"&x"1a","01"&x"53","01"&x"bf","10"&x"48",
	"00"&x"c3","00"&x"c5","00"&x"c7","00"&x"c9","00"&x"cb","00"&x"ce","00"&x"d3","00"&x"d9","00"&x"e3","00"&x"ef","01"&x"03","01"&x"1a","01"&x"47","01"&x"7f","01"&x"e7","10"&x"6b",
	"01"&x"03","01"&x"05","01"&x"06","01"&x"08","01"&x"0a","01"&x"0c","01"&x"10","01"&x"15","01"&x"1e","01"&x"29","01"&x"3c","01"&x"53","01"&x"7f","01"&x"b3","10"&x"1b","10"&x"9b",
	"01"&x"7d","01"&x"7f","01"&x"7f","01"&x"80","01"&x"82","01"&x"84","01"&x"87","01"&x"8b","01"&x"92","01"&x"9b","01"&x"aa","01"&x"bf","01"&x"e7","10"&x"1b","10"&x"7a","10"&x"f3",
	"10"&x"22","10"&x"22","10"&x"23","10"&x"23","10"&x"23","10"&x"24","10"&x"25","10"&x"26","10"&x"2a","10"&x"2f","10"&x"39","10"&x"48","10"&x"6b","10"&x"9b","10"&x"f3","11"&x"61",
	"00"&x"36","00"&x"38","00"&x"3a","00"&x"3d","00"&x"40","00"&x"43","00"&x"4a","00"&x"50","00"&x"5c","00"&x"6a","00"&x"82","00"&x"9d","00"&x"d0","01"&x"0e","01"&x"87","10"&x"28",
	"00"&x"38","00"&x"3b","00"&x"3d","00"&x"3f","00"&x"42","00"&x"46","00"&x"4c","00"&x"53","00"&x"5f","00"&x"6d","00"&x"84","00"&x"9f","00"&x"d2","01"&x"0f","01"&x"88","10"&x"28",
	"00"&x"3a","00"&x"3d","00"&x"3f","00"&x"41","00"&x"44","00"&x"48","00"&x"4e","00"&x"55","00"&x"61","00"&x"6f","00"&x"85","00"&x"a1","00"&x"d4","01"&x"10","01"&x"89","10"&x"28",
	"00"&x"3d","00"&x"3f","00"&x"41","00"&x"43","00"&x"46","00"&x"4a","00"&x"50","00"&x"57","00"&x"63","00"&x"71","00"&x"87","00"&x"a3","00"&x"d5","01"&x"12","01"&x"8a","10"&x"29",
	"00"&x"40","00"&x"42","00"&x"44","00"&x"46","00"&x"4a","00"&x"4d","00"&x"53","00"&x"5a","00"&x"66","00"&x"74","00"&x"8a","00"&x"a5","00"&x"d8","01"&x"14","01"&x"8c","10"&x"29",
	"00"&x"43","00"&x"46","00"&x"48","00"&x"4a","00"&x"4d","00"&x"51","00"&x"57","00"&x"5d","00"&x"69","00"&x"77","00"&x"8d","00"&x"a8","00"&x"db","01"&x"16","01"&x"8e","10"&x"29",
	"00"&x"4a","00"&x"4c","00"&x"4e","00"&x"50","00"&x"53","00"&x"57","00"&x"5d","00"&x"63","00"&x"6f","00"&x"7d","00"&x"92","00"&x"ae","00"&x"e0","01"&x"1b","01"&x"91","10"&x"2a",
	"00"&x"50","00"&x"53","00"&x"55","00"&x"57","00"&x"5a","00"&x"5d","00"&x"63","00"&x"6a","00"&x"76","00"&x"82","00"&x"99","00"&x"b4","00"&x"e5","01"&x"20","01"&x"94","10"&x"2c",
	"00"&x"5c","00"&x"5f","00"&x"61","00"&x"63","00"&x"66","00"&x"69","00"&x"6f","00"&x"76","00"&x"81","00"&x"8c","00"&x"a3","00"&x"be","00"&x"ef","01"&x"29","01"&x"9b","10"&x"2f",
	"00"&x"6a","00"&x"6d","00"&x"6f","00"&x"71","00"&x"74","00"&x"77","00"&x"7d","00"&x"82","00"&x"8c","00"&x"99","00"&x"b0","00"&x"cb","00"&x"fb","01"&x"33","01"&x"a2","10"&x"34",
	"00"&x"82","00"&x"84","00"&x"85","00"&x"87","00"&x"8a","00"&x"8d","00"&x"92","00"&x"99","00"&x"a3","00"&x"b0","00"&x"c6","00"&x"e0","01"&x"0d","01"&x"46","01"&x"b2","10"&x"3d",
	"00"&x"9d","00"&x"9f","00"&x"a1","00"&x"a3","00"&x"a5","00"&x"a8","00"&x"ae","00"&x"b4","00"&x"be","00"&x"cb","00"&x"e0","00"&x"f9","01"&x"25","01"&x"5d","01"&x"c6","10"&x"4c",
	"00"&x"d0","00"&x"d2","00"&x"d4","00"&x"d5","00"&x"d8","00"&x"db","00"&x"e0","00"&x"e5","00"&x"ef","00"&x"fb","01"&x"0d","01"&x"25","01"&x"51","01"&x"87","01"&x"ed","10"&x"6e",
	"01"&x"0e","01"&x"0f","01"&x"10","01"&x"12","01"&x"14","01"&x"16","01"&x"1b","01"&x"20","01"&x"29","01"&x"33","01"&x"46","01"&x"5d","01"&x"87","01"&x"ba","10"&x"20","10"&x"9c",
	"01"&x"87","01"&x"88","01"&x"89","01"&x"8a","01"&x"8c","01"&x"8e","01"&x"91","01"&x"94","01"&x"9b","01"&x"a2","01"&x"b2","01"&x"c6","01"&x"ed","10"&x"20","10"&x"7c","10"&x"f3",
	"10"&x"28","10"&x"28","10"&x"28","10"&x"29","10"&x"29","10"&x"29","10"&x"2a","10"&x"2c","10"&x"2f","10"&x"34","10"&x"3d","10"&x"4c","10"&x"6e","10"&x"9c","10"&x"f3","11"&x"61",
	"00"&x"50","00"&x"52","00"&x"54","00"&x"56","00"&x"5a","00"&x"5d","00"&x"63","00"&x"6a","00"&x"75","00"&x"82","00"&x"98","00"&x"b4","00"&x"e6","01"&x"22","01"&x"99","10"&x"34",
	"00"&x"52","00"&x"55","00"&x"57","00"&x"59","00"&x"5c","00"&x"5f","00"&x"65","00"&x"6c","00"&x"78","00"&x"84","00"&x"9a","00"&x"b6","00"&x"e8","01"&x"24","01"&x"9a","10"&x"34",
	"00"&x"54","00"&x"57","00"&x"59","00"&x"5b","00"&x"5e","00"&x"61","00"&x"67","00"&x"6e","00"&x"79","00"&x"85","00"&x"9c","00"&x"b8","00"&x"ea","01"&x"25","01"&x"9b","10"&x"34",
	"00"&x"56","00"&x"59","00"&x"5b","00"&x"5d","00"&x"60","00"&x"63","00"&x"69","00"&x"70","00"&x"7b","00"&x"87","00"&x"9e","00"&x"b9","00"&x"eb","01"&x"26","01"&x"9c","10"&x"34",
	"00"&x"5a","00"&x"5c","00"&x"5e","00"&x"60","00"&x"63","00"&x"66","00"&x"6c","00"&x"73","00"&x"7e","00"&x"8a","00"&x"a1","00"&x"bc","00"&x"ed","01"&x"28","01"&x"9d","10"&x"34",
	"00"&x"5d","00"&x"5f","00"&x"61","00"&x"63","00"&x"66","00"&x"6a","00"&x"70","00"&x"76","00"&x"81","00"&x"8d","00"&x"a4","00"&x"bf","00"&x"f0","01"&x"2a","01"&x"9f","10"&x"35",
	"00"&x"63","00"&x"65","00"&x"67","00"&x"69","00"&x"6c","00"&x"70","00"&x"75","00"&x"7c","00"&x"85","00"&x"92","00"&x"a9","00"&x"c4","00"&x"f5","01"&x"2f","01"&x"a1","10"&x"35",
	"00"&x"6a","00"&x"6c","00"&x"6e","00"&x"70","00"&x"73","00"&x"76","00"&x"7c","00"&x"82","00"&x"8c","00"&x"99","00"&x"af","00"&x"ca","00"&x"fa","01"&x"33","01"&x"a4","10"&x"36",
	"00"&x"75","00"&x"78","00"&x"79","00"&x"7b","00"&x"7e","00"&x"81","00"&x"85","00"&x"8c","00"&x"97","00"&x"a3","00"&x"ba","00"&x"d4","01"&x"03","01"&x"3c","01"&x"aa","10"&x"39",
	"00"&x"82","00"&x"84","00"&x"85","00"&x"87","00"&x"8a","00"&x"8d","00"&x"92","00"&x"99","00"&x"a3","00"&x"b0","00"&x"c6","00"&x"e0","01"&x"0d","01"&x"46","01"&x"b2","10"&x"3d",
	"00"&x"98","00"&x"9a","00"&x"9c","00"&x"9e","00"&x"a1","00"&x"a4","00"&x"a9","00"&x"af","00"&x"ba","00"&x"c6","00"&x"dc","00"&x"f5","01"&x"21","01"&x"58","01"&x"c2","10"&x"47",
	"00"&x"b4","00"&x"b6","00"&x"b8","00"&x"b9","00"&x"bc","00"&x"bf","00"&x"c4","00"&x"ca","00"&x"d4","00"&x"e0","00"&x"f5","01"&x"0c","01"&x"38","01"&x"6e","01"&x"d5","10"&x"55",
	"00"&x"e6","00"&x"e8","00"&x"ea","00"&x"eb","00"&x"ed","00"&x"f0","00"&x"f5","00"&x"fa","01"&x"03","01"&x"0d","01"&x"21","01"&x"38","01"&x"63","01"&x"97","01"&x"fa","10"&x"75",
	"01"&x"22","01"&x"24","01"&x"25","01"&x"26","01"&x"28","01"&x"2a","01"&x"2f","01"&x"33","01"&x"3c","01"&x"46","01"&x"58","01"&x"6e","01"&x"97","01"&x"c8","10"&x"2a","10"&x"a0",
	"01"&x"99","01"&x"9a","01"&x"9b","01"&x"9c","01"&x"9d","01"&x"9f","01"&x"a1","01"&x"a4","01"&x"aa","01"&x"b2","01"&x"c2","01"&x"d5","01"&x"fa","10"&x"2a","10"&x"82","10"&x"f5",
	"10"&x"34","10"&x"34","10"&x"34","10"&x"34","10"&x"34","10"&x"35","10"&x"35","10"&x"36","10"&x"39","10"&x"3d","10"&x"47","10"&x"55","10"&x"75","10"&x"a0","10"&x"f5","11"&x"61",
	"00"&x"6e","00"&x"70","00"&x"72","00"&x"74","00"&x"77","00"&x"7a","00"&x"80","00"&x"85","00"&x"90","00"&x"9d","00"&x"b4","00"&x"cf","01"&x"01","01"&x"3b","01"&x"af","10"&x"44",
	"00"&x"70","00"&x"72","00"&x"74","00"&x"76","00"&x"79","00"&x"7c","00"&x"81","00"&x"87","00"&x"92","00"&x"9f","00"&x"b6","00"&x"d1","01"&x"02","01"&x"3d","01"&x"b0","10"&x"44",
	"00"&x"72","00"&x"74","00"&x"76","00"&x"78","00"&x"7b","00"&x"7e","00"&x"83","00"&x"89","00"&x"94","00"&x"a1","00"&x"b8","00"&x"d3","01"&x"04","01"&x"3e","01"&x"b1","10"&x"44",
	"00"&x"74","00"&x"76","00"&x"78","00"&x"7a","00"&x"7d","00"&x"80","00"&x"84","00"&x"8a","00"&x"95","00"&x"a3","00"&x"b9","00"&x"d4","01"&x"05","01"&x"3f","01"&x"b1","10"&x"44",
	"00"&x"77","00"&x"79","00"&x"7b","00"&x"7d","00"&x"80","00"&x"82","00"&x"87","00"&x"8d","00"&x"98","00"&x"a5","00"&x"bc","00"&x"d7","01"&x"07","01"&x"41","01"&x"b2","10"&x"44",
	"00"&x"7a","00"&x"7c","00"&x"7e","00"&x"80","00"&x"82","00"&x"85","00"&x"8a","00"&x"90","00"&x"9b","00"&x"a8","00"&x"bf","00"&x"da","01"&x"09","01"&x"43","01"&x"b4","10"&x"44",
	"00"&x"80","00"&x"81","00"&x"83","00"&x"84","00"&x"87","00"&x"8a","00"&x"90","00"&x"96","00"&x"a1","00"&x"ae","00"&x"c4","00"&x"df","01"&x"0d","01"&x"47","01"&x"b6","10"&x"45",
	"00"&x"85","00"&x"87","00"&x"89","00"&x"8a","00"&x"8d","00"&x"90","00"&x"96","00"&x"9c","00"&x"a7","00"&x"b4","00"&x"ca","00"&x"e4","01"&x"11","01"&x"4b","01"&x"b9","10"&x"46",
	"00"&x"90","00"&x"92","00"&x"94","00"&x"95","00"&x"98","00"&x"9b","00"&x"a1","00"&x"a7","00"&x"b2","00"&x"be","00"&x"d4","00"&x"ee","01"&x"1a","01"&x"53","01"&x"bf","10"&x"48",
	"00"&x"9d","00"&x"9f","00"&x"a1","00"&x"a3","00"&x"a5","00"&x"a8","00"&x"ae","00"&x"b4","00"&x"be","00"&x"cb","00"&x"e0","00"&x"f9","01"&x"25","01"&x"5d","01"&x"c6","10"&x"4c",
	"00"&x"b4","00"&x"b6","00"&x"b8","00"&x"b9","00"&x"bc","00"&x"bf","00"&x"c4","00"&x"ca","00"&x"d4","00"&x"e0","00"&x"f5","01"&x"0c","01"&x"38","01"&x"6e","01"&x"d5","10"&x"55",
	"00"&x"cf","00"&x"d1","00"&x"d3","00"&x"d4","00"&x"d7","00"&x"da","00"&x"df","00"&x"e4","00"&x"ee","00"&x"f9","01"&x"0c","01"&x"23","01"&x"4e","01"&x"84","01"&x"e7","10"&x"63",
	"01"&x"01","01"&x"02","01"&x"04","01"&x"05","01"&x"07","01"&x"09","01"&x"0d","01"&x"11","01"&x"1a","01"&x"25","01"&x"38","01"&x"4e","01"&x"78","01"&x"a9","10"&x"0b","10"&x"80",
	"01"&x"3b","01"&x"3d","01"&x"3e","01"&x"3f","01"&x"41","01"&x"43","01"&x"47","01"&x"4b","01"&x"53","01"&x"5d","01"&x"6e","01"&x"84","01"&x"a9","01"&x"da","10"&x"37","10"&x"a9",
	"01"&x"af","01"&x"b0","01"&x"b1","01"&x"b1","01"&x"b2","01"&x"b4","01"&x"b6","01"&x"b9","01"&x"bf","01"&x"c6","01"&x"d5","01"&x"e7","10"&x"0b","10"&x"37","10"&x"8c","10"&x"f9",
	"10"&x"44","10"&x"44","10"&x"44","10"&x"44","10"&x"44","10"&x"44","10"&x"45","10"&x"46","10"&x"48","10"&x"4c","10"&x"55","10"&x"63","10"&x"80","10"&x"a9","10"&x"f9","11"&x"61",
	"00"&x"a1","00"&x"a4","00"&x"a5","00"&x"a7","00"&x"aa","00"&x"ad","00"&x"b3","00"&x"b9","00"&x"c3","00"&x"d0","00"&x"e6","01"&x"01","01"&x"2f","01"&x"6a","01"&x"dc","10"&x"69",
	"00"&x"a4","00"&x"a6","00"&x"a8","00"&x"a9","00"&x"ac","00"&x"af","00"&x"b5","00"&x"bb","00"&x"c5","00"&x"d2","00"&x"e8","01"&x"02","01"&x"31","01"&x"6c","01"&x"dc","10"&x"69",
	"00"&x"a5","00"&x"a8","00"&x"a9","00"&x"ab","00"&x"ae","00"&x"b1","00"&x"b6","00"&x"bd","00"&x"c7","00"&x"d4","00"&x"ea","01"&x"04","01"&x"32","01"&x"6c","01"&x"dd","10"&x"69",
	"00"&x"a7","00"&x"a9","00"&x"ab","00"&x"ad","00"&x"b0","00"&x"b3","00"&x"b8","00"&x"be","00"&x"c9","00"&x"d5","00"&x"eb","01"&x"05","01"&x"33","01"&x"6d","01"&x"dd","10"&x"69",
	"00"&x"aa","00"&x"ac","00"&x"ae","00"&x"b0","00"&x"b2","00"&x"b6","00"&x"bb","00"&x"c1","00"&x"cb","00"&x"d8","00"&x"ed","01"&x"07","01"&x"35","01"&x"6f","01"&x"de","10"&x"69",
	"00"&x"ad","00"&x"af","00"&x"b1","00"&x"b3","00"&x"b6","00"&x"b9","00"&x"be","00"&x"c4","00"&x"ce","00"&x"db","00"&x"f0","01"&x"09","01"&x"37","01"&x"71","01"&x"df","10"&x"69",
	"00"&x"b3","00"&x"b5","00"&x"b6","00"&x"b8","00"&x"bb","00"&x"be","00"&x"c3","00"&x"c9","00"&x"d3","00"&x"e0","00"&x"f5","01"&x"0d","01"&x"3b","01"&x"74","01"&x"e0","10"&x"69",
	"00"&x"b9","00"&x"bb","00"&x"bd","00"&x"be","00"&x"c1","00"&x"c4","00"&x"c9","00"&x"cf","00"&x"d9","00"&x"e5","00"&x"fa","01"&x"11","01"&x"3f","01"&x"78","01"&x"e3","10"&x"6a",
	"00"&x"c3","00"&x"c5","00"&x"c7","00"&x"c9","00"&x"cb","00"&x"ce","00"&x"d3","00"&x"d9","00"&x"e3","00"&x"ef","01"&x"03","01"&x"1a","01"&x"47","01"&x"7f","01"&x"e7","10"&x"6b",
	"00"&x"d0","00"&x"d2","00"&x"d4","00"&x"d5","00"&x"d8","00"&x"db","00"&x"e0","00"&x"e5","00"&x"ef","00"&x"fb","01"&x"0d","01"&x"25","01"&x"51","01"&x"87","01"&x"ed","10"&x"6e",
	"00"&x"e6","00"&x"e8","00"&x"ea","00"&x"eb","00"&x"ed","00"&x"f0","00"&x"f5","00"&x"fa","01"&x"03","01"&x"0d","01"&x"21","01"&x"38","01"&x"63","01"&x"97","01"&x"fa","10"&x"75",
	"01"&x"01","01"&x"02","01"&x"04","01"&x"05","01"&x"07","01"&x"09","01"&x"0d","01"&x"11","01"&x"1a","01"&x"25","01"&x"38","01"&x"4e","01"&x"78","01"&x"a9","10"&x"0b","10"&x"80",
	"01"&x"2f","01"&x"31","01"&x"32","01"&x"33","01"&x"35","01"&x"37","01"&x"3b","01"&x"3f","01"&x"47","01"&x"51","01"&x"63","01"&x"78","01"&x"9e","01"&x"ce","10"&x"2c","10"&x"9b",
	"01"&x"6a","01"&x"6c","01"&x"6c","01"&x"6d","01"&x"6f","01"&x"71","01"&x"74","01"&x"78","01"&x"7f","01"&x"87","01"&x"97","01"&x"a9","01"&x"ce","01"&x"fd","10"&x"54","10"&x"c0",
	"01"&x"dc","01"&x"dc","01"&x"dd","01"&x"dd","01"&x"de","01"&x"df","01"&x"e0","01"&x"e3","01"&x"e7","01"&x"ed","01"&x"fa","10"&x"0b","10"&x"2c","10"&x"54","10"&x"a4","11"&x"09",
	"10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"6a","10"&x"6b","10"&x"6e","10"&x"75","10"&x"80","10"&x"9b","10"&x"c0","11"&x"09","11"&x"67",
	"00"&x"e4","00"&x"e6","00"&x"e8","00"&x"e9","00"&x"ec","00"&x"ef","00"&x"f4","00"&x"f9","01"&x"03","01"&x"0e","01"&x"22","01"&x"3b","01"&x"6a","01"&x"a3","10"&x"14","10"&x"9a",
	"00"&x"e6","00"&x"e8","00"&x"ea","00"&x"eb","00"&x"ee","00"&x"f1","00"&x"f5","00"&x"fb","01"&x"05","01"&x"0f","01"&x"24","01"&x"3d","01"&x"6c","01"&x"a4","10"&x"14","10"&x"9a",
	"00"&x"e8","00"&x"ea","00"&x"eb","00"&x"ed","00"&x"ef","00"&x"f2","00"&x"f7","00"&x"fc","01"&x"06","01"&x"10","01"&x"25","01"&x"3e","01"&x"6c","01"&x"a5","10"&x"15","10"&x"9a",
	"00"&x"e9","00"&x"eb","00"&x"ed","00"&x"ee","00"&x"f1","00"&x"f4","00"&x"f8","00"&x"fe","01"&x"08","01"&x"12","01"&x"26","01"&x"3f","01"&x"6d","01"&x"a5","10"&x"15","10"&x"9a",
	"00"&x"ec","00"&x"ee","00"&x"ef","00"&x"f1","00"&x"f3","00"&x"f6","00"&x"fb","01"&x"00","01"&x"0a","01"&x"14","01"&x"28","01"&x"41","01"&x"6f","01"&x"a6","10"&x"15","10"&x"9a",
	"00"&x"ef","00"&x"f1","00"&x"f2","00"&x"f4","00"&x"f6","00"&x"f9","00"&x"fe","01"&x"03","01"&x"0c","01"&x"16","01"&x"2a","01"&x"43","01"&x"71","01"&x"a8","10"&x"16","10"&x"9a",
	"00"&x"f4","00"&x"f5","00"&x"f7","00"&x"f8","00"&x"fb","00"&x"fe","01"&x"02","01"&x"08","01"&x"10","01"&x"1b","01"&x"2f","01"&x"47","01"&x"74","01"&x"aa","10"&x"17","10"&x"9a",
	"00"&x"f9","00"&x"fb","00"&x"fc","00"&x"fe","01"&x"00","01"&x"03","01"&x"08","01"&x"0c","01"&x"15","01"&x"20","01"&x"33","01"&x"4b","01"&x"78","01"&x"ad","10"&x"18","10"&x"9a",
	"01"&x"03","01"&x"05","01"&x"06","01"&x"08","01"&x"0a","01"&x"0c","01"&x"10","01"&x"15","01"&x"1e","01"&x"29","01"&x"3c","01"&x"53","01"&x"7f","01"&x"b3","10"&x"1b","10"&x"9b",
	"01"&x"0e","01"&x"0f","01"&x"10","01"&x"12","01"&x"14","01"&x"16","01"&x"1b","01"&x"20","01"&x"29","01"&x"33","01"&x"46","01"&x"5d","01"&x"87","01"&x"ba","10"&x"20","10"&x"9c",
	"01"&x"22","01"&x"24","01"&x"25","01"&x"26","01"&x"28","01"&x"2a","01"&x"2f","01"&x"33","01"&x"3c","01"&x"46","01"&x"58","01"&x"6e","01"&x"97","01"&x"c8","10"&x"2a","10"&x"a0",
	"01"&x"3b","01"&x"3d","01"&x"3e","01"&x"3f","01"&x"41","01"&x"43","01"&x"47","01"&x"4b","01"&x"53","01"&x"5d","01"&x"6e","01"&x"84","01"&x"a9","01"&x"da","10"&x"37","10"&x"a9",
	"01"&x"6a","01"&x"6c","01"&x"6c","01"&x"6d","01"&x"6f","01"&x"71","01"&x"74","01"&x"78","01"&x"7f","01"&x"87","01"&x"97","01"&x"a9","01"&x"ce","01"&x"fd","10"&x"54","10"&x"c0",
	"01"&x"a3","01"&x"a4","01"&x"a5","01"&x"a5","01"&x"a6","01"&x"a8","01"&x"aa","01"&x"ad","01"&x"b3","01"&x"ba","01"&x"c8","01"&x"da","01"&x"fd","10"&x"29","10"&x"7b","10"&x"e0",
	"10"&x"14","10"&x"14","10"&x"15","10"&x"15","10"&x"15","10"&x"16","10"&x"17","10"&x"18","10"&x"1b","10"&x"20","10"&x"2a","10"&x"37","10"&x"54","10"&x"7b","10"&x"c6","11"&x"25",
	"10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9b","10"&x"9c","10"&x"a0","10"&x"a9","10"&x"c0","10"&x"e0","11"&x"25","11"&x"7a",
	"01"&x"66","01"&x"67","01"&x"68","01"&x"69","01"&x"6b","01"&x"6d","01"&x"71","01"&x"75","01"&x"7d","01"&x"87","01"&x"99","01"&x"af","01"&x"dc","10"&x"14","10"&x"79","10"&x"f3",
	"01"&x"67","01"&x"68","01"&x"6a","01"&x"6b","01"&x"6c","01"&x"6e","01"&x"72","01"&x"77","01"&x"7f","01"&x"88","01"&x"9a","01"&x"b0","01"&x"dc","10"&x"14","10"&x"79","10"&x"f3",
	"01"&x"68","01"&x"6a","01"&x"6b","01"&x"6c","01"&x"6e","01"&x"70","01"&x"73","01"&x"78","01"&x"7f","01"&x"89","01"&x"9b","01"&x"b1","01"&x"dd","10"&x"15","10"&x"79","10"&x"f3",
	"01"&x"69","01"&x"6b","01"&x"6c","01"&x"6d","01"&x"6f","01"&x"71","01"&x"74","01"&x"79","01"&x"80","01"&x"8a","01"&x"9c","01"&x"b1","01"&x"dd","10"&x"15","10"&x"79","10"&x"f3",
	"01"&x"6b","01"&x"6c","01"&x"6e","01"&x"6f","01"&x"70","01"&x"72","01"&x"76","01"&x"7a","01"&x"82","01"&x"8c","01"&x"9d","01"&x"b2","01"&x"de","10"&x"15","10"&x"79","10"&x"f3",
	"01"&x"6d","01"&x"6e","01"&x"70","01"&x"71","01"&x"72","01"&x"74","01"&x"78","01"&x"7c","01"&x"84","01"&x"8e","01"&x"9f","01"&x"b4","01"&x"df","10"&x"16","10"&x"79","10"&x"f3",
	"01"&x"71","01"&x"72","01"&x"73","01"&x"74","01"&x"76","01"&x"78","01"&x"7c","01"&x"80","01"&x"87","01"&x"91","01"&x"a1","01"&x"b6","01"&x"e0","10"&x"17","10"&x"79","10"&x"f3",
	"01"&x"75","01"&x"77","01"&x"78","01"&x"79","01"&x"7a","01"&x"7c","01"&x"80","01"&x"84","01"&x"8b","01"&x"94","01"&x"a4","01"&x"b9","01"&x"e3","10"&x"18","10"&x"79","10"&x"f3",
	"01"&x"7d","01"&x"7f","01"&x"7f","01"&x"80","01"&x"82","01"&x"84","01"&x"87","01"&x"8b","01"&x"92","01"&x"9b","01"&x"aa","01"&x"bf","01"&x"e7","10"&x"1b","10"&x"7a","10"&x"f3",
	"01"&x"87","01"&x"88","01"&x"89","01"&x"8a","01"&x"8c","01"&x"8e","01"&x"91","01"&x"94","01"&x"9b","01"&x"a2","01"&x"b2","01"&x"c6","01"&x"ed","10"&x"20","10"&x"7c","10"&x"f3",
	"01"&x"99","01"&x"9a","01"&x"9b","01"&x"9c","01"&x"9d","01"&x"9f","01"&x"a1","01"&x"a4","01"&x"aa","01"&x"b2","01"&x"c2","01"&x"d5","01"&x"fa","10"&x"2a","10"&x"82","10"&x"f5",
	"01"&x"af","01"&x"b0","01"&x"b1","01"&x"b1","01"&x"b2","01"&x"b4","01"&x"b6","01"&x"b9","01"&x"bf","01"&x"c6","01"&x"d5","01"&x"e7","10"&x"0b","10"&x"37","10"&x"8c","10"&x"f9",
	"01"&x"dc","01"&x"dc","01"&x"dd","01"&x"dd","01"&x"de","01"&x"df","01"&x"e0","01"&x"e3","01"&x"e7","01"&x"ed","01"&x"fa","10"&x"0b","10"&x"2c","10"&x"54","10"&x"a4","11"&x"09",
	"10"&x"14","10"&x"14","10"&x"15","10"&x"15","10"&x"15","10"&x"16","10"&x"17","10"&x"18","10"&x"1b","10"&x"20","10"&x"2a","10"&x"37","10"&x"54","10"&x"7b","10"&x"c6","11"&x"25",
	"10"&x"79","10"&x"79","10"&x"79","10"&x"79","10"&x"79","10"&x"79","10"&x"79","10"&x"79","10"&x"7a","10"&x"7c","10"&x"82","10"&x"8c","10"&x"a4","10"&x"c6","11"&x"0c","11"&x"62",
	"10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f5","10"&x"f9","11"&x"09","11"&x"25","11"&x"62","11"&x"b1",
	"10"&x"1a","10"&x"1a","10"&x"1a","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1d","10"&x"1f","10"&x"22","10"&x"28","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1a","10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1d","10"&x"1f","10"&x"22","10"&x"28","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1a","10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1c","10"&x"1d","10"&x"1f","10"&x"23","10"&x"28","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1b","10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1e","10"&x"1f","10"&x"23","10"&x"29","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1b","10"&x"1b","10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1d","10"&x"1e","10"&x"20","10"&x"23","10"&x"29","10"&x"34","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1c","10"&x"1d","10"&x"1e","10"&x"1f","10"&x"20","10"&x"24","10"&x"29","10"&x"35","10"&x"44","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1d","10"&x"1d","10"&x"1d","10"&x"1e","10"&x"1e","10"&x"1f","10"&x"20","10"&x"21","10"&x"25","10"&x"2a","10"&x"35","10"&x"45","10"&x"69","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"1f","10"&x"1f","10"&x"1f","10"&x"1f","10"&x"20","10"&x"20","10"&x"21","10"&x"23","10"&x"26","10"&x"2c","10"&x"36","10"&x"46","10"&x"6a","10"&x"9a","10"&x"f3","11"&x"61",
	"10"&x"22","10"&x"22","10"&x"23","10"&x"23","10"&x"23","10"&x"24","10"&x"25","10"&x"26","10"&x"2a","10"&x"2f","10"&x"39","10"&x"48","10"&x"6b","10"&x"9b","10"&x"f3","11"&x"61",
	"10"&x"28","10"&x"28","10"&x"28","10"&x"29","10"&x"29","10"&x"29","10"&x"2a","10"&x"2c","10"&x"2f","10"&x"34","10"&x"3d","10"&x"4c","10"&x"6e","10"&x"9c","10"&x"f3","11"&x"61",
	"10"&x"34","10"&x"34","10"&x"34","10"&x"34","10"&x"34","10"&x"35","10"&x"35","10"&x"36","10"&x"39","10"&x"3d","10"&x"47","10"&x"55","10"&x"75","10"&x"a0","10"&x"f5","11"&x"61",
	"10"&x"44","10"&x"44","10"&x"44","10"&x"44","10"&x"44","10"&x"44","10"&x"45","10"&x"46","10"&x"48","10"&x"4c","10"&x"55","10"&x"63","10"&x"80","10"&x"a9","10"&x"f9","11"&x"61",
	"10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"69","10"&x"6a","10"&x"6b","10"&x"6e","10"&x"75","10"&x"80","10"&x"9b","10"&x"c0","11"&x"09","11"&x"67",
	"10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9a","10"&x"9b","10"&x"9c","10"&x"a0","10"&x"a9","10"&x"c0","10"&x"e0","11"&x"25","11"&x"7a",
	"10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f3","10"&x"f5","10"&x"f9","11"&x"09","11"&x"25","11"&x"62","11"&x"b1",
	"11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"61","11"&x"67","11"&x"7a","11"&x"b1","11"&x"f9"
);

signal ROM : ROM_ARRAY := voltable;

begin

process(CLK)
begin
	if rising_edge(CLK) then
		DATA_A <= ROM(to_integer(unsigned(ADDR_A)));
		DATA_B <= ROM(to_integer(unsigned(ADDR_B)));
	end if;
end process;
end RTL;
