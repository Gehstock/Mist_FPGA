library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg4_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg4_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"CD",X"EE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"DD",X"EE",X"EE",X"FC",X"CF",X"FC",X"C0",X"FE",X"E0",X"FE",X"E0",
		X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",
		X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"00",X"CC",X"FF",X"EC",X"CC",X"FC",X"CC",X"EC",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"00",
		X"EC",X"FF",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"CC",X"FF",X"EC",X"CC",X"EC",X"CC",X"EC",X"EE",X"EC",X"FF",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",
		X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",X"FF",X"F0",X"FC",X"C0",X"FD",X"D0",X"FE",X"E0",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EF",X"FE",X"FF",X"FE",X"11",X"11",X"44",X"44",
		X"DD",X"EE",X"FC",X"CC",X"EC",X"DD",X"EC",X"FF",X"EC",X"FF",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"33",X"32",X"33",X"23",X"23",X"33",X"32",X"33",X"32",X"33",X"23",X"33",X"33",X"23",X"33",X"32",
		X"CC",X"FF",X"DC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"11",X"11",X"77",X"77",X"99",X"99",X"11",X"11",X"66",X"66",X"AB",X"A6",X"BA",X"B6",X"AB",X"A8",
		X"11",X"11",X"77",X"77",X"99",X"99",X"11",X"11",X"66",X"61",X"AB",X"61",X"B3",X"61",X"AB",X"61",
		X"DD",X"DD",X"CC",X"CC",X"FD",X"FF",X"DC",X"69",X"DC",X"B9",X"DC",X"A8",X"DC",X"B8",X"CE",X"F8",
		X"DD",X"DD",X"CC",X"CC",X"FD",X"FF",X"DC",X"91",X"DC",X"91",X"DC",X"81",X"DC",X"81",X"CE",X"F1",
		X"08",X"88",X"08",X"88",X"08",X"88",X"08",X"88",X"08",X"88",X"08",X"88",X"08",X"88",X"18",X"88",
		X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",
		X"88",X"88",X"99",X"99",X"74",X"74",X"88",X"88",X"77",X"77",X"88",X"88",X"99",X"90",X"88",X"88",
		X"88",X"88",X"99",X"90",X"74",X"00",X"88",X"00",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"8F",X"77",X"FC",X"78",X"CC",X"8F",X"CE",X"FC",X"FC",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"88",X"88",X"77",X"77",X"99",X"99",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CD",X"CC",X"DD",X"CD",X"FF",
		X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1E",X"DD",X"11",X"FF",X"11",X"11",X"DD",X"DD",X"DC",X"CC",
		X"DD",X"11",X"FF",X"1D",X"11",X"1D",X"DD",X"D1",X"11",X"D1",X"C1",X"F1",X"CC",X"11",X"CC",X"CD",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"11",X"11",X"BB",X"BB",X"22",X"22",X"03",X"1B",X"11",X"11",X"BB",X"BB",X"22",X"22",X"03",X"1B",
		X"11",X"11",X"BB",X"BB",X"22",X"22",X"80",X"78",X"11",X"11",X"BB",X"BB",X"22",X"22",X"80",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",X"33",X"00",X"77",X"77",
		X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",X"77",X"77",X"99",X"97",X"11",X"17",
		X"11",X"17",X"11",X"17",X"11",X"17",X"11",X"17",X"11",X"17",X"11",X"17",X"99",X"97",X"77",X"77",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"F0",X"CC",X"CF",X"EC",X"CC",X"EC",X"EC",X"EC",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"FF",X"CC",X"CC",
		X"CF",X"00",X"CC",X"FF",X"EC",X"CC",X"EC",X"CC",X"EF",X"EE",X"FF",X"FF",X"11",X"11",X"88",X"88",
		X"00",X"00",X"FE",X"00",X"CC",X"00",X"CE",X"00",X"EC",X"00",X"EE",X"C0",X"11",X"E0",X"88",X"00",
		X"77",X"77",X"18",X"19",X"77",X"77",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"70",X"91",X"00",X"77",X"00",X"18",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"77",X"FF",X"77",X"CC",X"77",X"CC",X"F7",X"EE",X"FF",X"EF",X"CC",X"FE",X"CC",X"EC",X"FE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"F7",X"77",X"FF",X"77",
		X"FD",X"1F",X"8F",X"1E",X"18",X"EC",X"11",X"FD",X"F1",X"8F",X"EF",X"88",X"EE",X"11",X"EE",X"FF",
		X"CC",X"77",X"CC",X"F7",X"FE",X"FF",X"1F",X"CC",X"1E",X"CC",X"EC",X"FE",X"FD",X"1F",X"8F",X"1C",
		X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",
		X"77",X"71",X"77",X"77",X"77",X"77",X"17",X"77",X"91",X"77",X"99",X"77",X"91",X"17",X"91",X"91",
		X"99",X"99",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",X"8C",X"98",X"EC",X"F8",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"77",X"CC",X"77",X"CC",X"77",
		X"FE",X"FF",X"FF",X"CC",X"1E",X"CC",X"EC",X"FE",X"FD",X"FF",X"8F",X"1E",X"78",X"EC",X"11",X"FD",
		X"FF",X"FF",X"CC",X"CC",X"DC",X"DD",X"FF",X"EE",X"CC",X"FF",X"CC",X"FE",X"FE",X"FF",X"FF",X"CC",
		X"77",X"8F",X"77",X"78",X"77",X"11",X"77",X"77",X"77",X"77",X"11",X"77",X"1C",X"77",X"EC",X"F7",
		X"1E",X"CC",X"EC",X"FE",X"FD",X"FE",X"8F",X"EC",X"78",X"FD",X"11",X"7F",X"1C",X"88",X"EC",X"F8",
		X"FF",X"FF",X"CC",X"CC",X"DC",X"DD",X"EC",X"EE",X"EC",X"FF",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"FF",X"FF",X"CC",X"CC",X"DC",X"DD",X"EC",X"EE",X"EC",X"FF",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"FC",X"FE",X"CF",X"FE",X"CC",X"FE",X"EC",X"FE",X"FE",X"CF",X"1F",X"CC",X"7D",X"EC",X"ED",X"FE",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"FC",X"FE",X"CF",X"FE",X"CC",X"FF",
		X"CC",X"C1",X"CC",X"D1",X"CC",X"D1",X"CC",X"D1",X"CC",X"1D",X"CC",X"1D",X"CC",X"1E",X"CD",X"11",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"DE",X"D1",X"E1",X"DD",X"1C",X"CD",X"DC",X"CD",X"DC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"DC",X"CD",X"DC",X"DD",X"DD",X"FF",X"EF",X"11",X"11",X"DD",X"1D",X"DC",X"1D",X"CC",X"1D",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1E",X"DC",X"11",X"FD",
		X"DD",X"DD",X"FF",X"FF",X"11",X"11",X"DD",X"D1",X"CC",X"D1",X"CC",X"D1",X"CC",X"D1",X"CC",X"D1",
		X"DD",X"1F",X"DD",X"D1",X"CC",X"DD",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"1C",X"CC",X"CC",X"CC",X"CC",X"CC",X"1C",X"DD",X"1D",X"DE",X"1D",X"EE",X"1E",X"11",X"11",
		X"CC",X"11",X"CC",X"1C",X"CC",X"CC",X"CD",X"CC",X"DD",X"CD",X"DD",X"DD",X"EE",X"EE",X"11",X"11",
		X"EC",X"FE",X"EC",X"FE",X"FF",X"FE",X"CC",X"FE",X"CC",X"CF",X"EC",X"CC",X"EC",X"EC",X"EC",X"EE",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"FF",X"FE",X"CC",X"FF",X"CC",X"CC",
		X"9D",X"77",X"89",X"77",X"88",X"77",X"88",X"97",X"11",X"89",X"91",X"18",X"91",X"11",X"91",X"91",
		X"19",X"EC",X"71",X"FD",X"77",X"8F",X"77",X"99",X"77",X"11",X"77",X"77",X"17",X"77",X"91",X"D7",
		X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"9C",X"91",X"EC",X"F8",
		X"99",X"77",X"91",X"77",X"91",X"11",X"91",X"91",X"99",X"98",X"91",X"91",X"9C",X"91",X"EC",X"F9",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"11",X"77",X"1A",X"77",X"AA",X"77",X"1A",
		X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"17",X"11",X"87",X"1A",X"87",X"BB",X"87",X"1B",X"87",
		X"77",X"1A",X"77",X"1A",X"77",X"AA",X"77",X"1B",X"77",X"1B",X"77",X"22",X"77",X"22",X"77",X"77",
		X"1B",X"87",X"1B",X"87",X"BB",X"87",X"1B",X"87",X"1B",X"87",X"22",X"87",X"22",X"87",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",
		X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"18",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"22",X"77",X"22",X"77",X"77",
		X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"28",X"77",X"77",X"77",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EF",X"FE",X"FF",X"FE",X"11",X"11",X"88",X"88",
		X"EC",X"FF",X"EC",X"CC",X"EC",X"CC",X"EC",X"FE",X"EF",X"FE",X"FF",X"FE",X"11",X"11",X"88",X"88",
		X"00",X"C0",X"FF",X"E0",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"3B",X"00",X"3B",X"00",X"33",X"00",X"33",X"00",X"FF",X"00",X"EE",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"8F",X"66",X"FC",X"44",X"CC",X"7F",X"CE",X"FC",X"FC",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"66",X"FF",X"44",X"CC",X"77",X"CC",X"11",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"CC",X"CD",X"CC",X"DD",X"CC",X"D1",X"CC",X"D1",X"CC",X"1D",X"CC",X"1D",X"CD",X"1E",X"DD",X"11",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"DD",X"11",X"CD",X"DD",X"DD",X"CC",X"FF",X"CC",X"11",X"CC",X"C1",X"CC",X"CC",X"CC",X"CC",
		X"DC",X"CC",X"ED",X"DD",X"1E",X"FF",X"11",X"11",X"11",X"DD",X"D1",X"CC",X"1D",X"CC",X"1D",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",
		X"EE",X"CC",X"11",X"CC",X"D1",X"CC",X"DD",X"DC",X"DC",X"ED",X"DC",X"EF",X"ED",X"11",X"1F",X"1D",
		X"CC",X"DD",X"DD",X"DE",X"FF",X"F1",X"11",X"11",X"DD",X"DD",X"CC",X"DD",X"CC",X"CD",X"CC",X"CD",
		X"11",X"DD",X"DD",X"DC",X"DC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"FF",X"CC",
		X"00",X"00",X"00",X"FF",X"00",X"CC",X"FF",X"CD",X"CC",X"EE",X"CC",X"FF",X"EC",X"FE",X"EC",X"FE",
		X"CC",X"EE",X"CC",X"FE",X"DC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"33",X"11",X"33",X"11",X"11",X"55",X"55",X"66",X"66",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"11",X"55",X"55",X"66",X"66",
		X"77",X"77",X"18",X"18",X"77",X"77",X"81",X"81",X"81",X"81",X"99",X"99",X"99",X"99",X"88",X"88",
		X"99",X"99",X"99",X"99",X"91",X"99",X"91",X"99",X"81",X"88",X"81",X"88",X"71",X"77",X"79",X"77",
		X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"CD",X"FE",X"FF",X"FE",X"FF",X"FE",X"11",X"11",X"88",X"88",
		X"CD",X"FF",X"CD",X"FF",X"CD",X"FF",X"CD",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"11",X"88",X"88",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FF",X"EC",X"FC",X"EF",X"CC",X"FC",X"CE",
		X"EC",X"FC",X"EC",X"CC",X"FF",X"CE",X"CC",X"EF",X"CC",X"F1",X"CD",X"18",X"CC",X"88",X"EC",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"CC",X"FC",X"CC",X"CC",X"EE",
		X"00",X"00",X"00",X"FF",X"00",X"CC",X"FF",X"CC",X"CC",X"FE",X"CC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FE",X"EC",X"FF",X"EF",X"CC",X"FC",X"CC",X"CC",X"EE",
		X"EC",X"FE",X"EC",X"FF",X"EC",X"CC",X"FF",X"CC",X"CC",X"DE",X"CC",X"FE",X"EC",X"FE",X"EC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"99",X"02",X"AA",X"08",X"00",X"08",X"00",X"00",X"02",
		X"27",X"00",X"89",X"90",X"9A",X"00",X"9A",X"00",X"89",X"00",X"98",X"90",X"78",X"00",X"97",X"A0",
		X"00",X"00",X"00",X"89",X"29",X"99",X"9A",X"7A",X"99",X"99",X"00",X"09",X"70",X"AA",X"99",X"99",
		X"A9",X"A0",X"98",X"A0",X"88",X"A0",X"AA",X"A0",X"2A",X"00",X"8A",X"00",X"8A",X"20",X"AA",X"82",
		X"77",X"77",X"18",X"17",X"77",X"71",X"44",X"87",X"88",X"88",X"11",X"88",X"11",X"11",X"11",X"11",
		X"1F",X"FE",X"81",X"FE",X"48",X"FE",X"77",X"FE",X"17",X"1E",X"71",X"81",X"87",X"48",X"88",X"77",
		X"99",X"11",X"99",X"99",X"99",X"99",X"99",X"99",X"88",X"89",X"88",X"88",X"77",X"88",X"77",X"77",
		X"18",X"17",X"11",X"71",X"91",X"87",X"99",X"88",X"99",X"88",X"89",X"99",X"88",X"89",X"88",X"88",
		X"44",X"44",X"77",X"77",X"11",X"11",X"19",X"99",X"19",X"66",X"19",X"67",X"19",X"77",X"19",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"66",X"66",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"66",X"66",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"44",X"44",X"77",X"74",X"11",X"74",X"99",X"74",X"97",X"74",X"99",X"74",X"66",X"74",X"76",X"74",
		X"11",X"11",X"11",X"18",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"22",X"88",X"22",X"28",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"CE",X"F0",
		X"DD",X"D0",X"CC",X"DF",X"FF",X"F0",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"CE",X"F0",
		X"44",X"44",X"77",X"77",X"11",X"11",X"18",X"88",X"18",X"88",X"18",X"99",X"18",X"77",X"18",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"77",X"99",X"79",X"88",X"98",X"88",X"88",X"88",
		X"CC",X"CD",X"CC",X"DD",X"CC",X"D1",X"CC",X"D1",X"DD",X"1D",X"FF",X"1E",X"11",X"1E",X"DD",X"11",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"D1",X"CC",X"DD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"DC",X"DD",X"DD",X"FF",X"EF",X"11",X"11",X"DD",X"11",X"DC",X"D1",X"CC",X"D1",X"CC",
		X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"DD",X"DD",X"FF",X"FF",X"11",X"11",X"DD",X"D1",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"DC",X"CC",
		X"CC",X"DD",X"CC",X"CD",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"ED",X"CC",X"ED",X"DD",X"1E",X"FF",X"11",X"11",X"D1",X"DD",X"D1",X"DC",X"D1",X"CC",X"D1",X"CC",
		X"18",X"77",X"19",X"77",X"17",X"79",X"17",X"77",X"17",X"77",X"17",X"79",X"19",X"77",X"18",X"77",
		X"88",X"88",X"98",X"88",X"79",X"88",X"77",X"88",X"77",X"88",X"79",X"88",X"98",X"88",X"88",X"88",
		X"18",X"77",X"18",X"77",X"18",X"99",X"18",X"88",X"18",X"88",X"14",X"44",X"77",X"77",X"11",X"11",
		X"88",X"88",X"98",X"88",X"79",X"88",X"77",X"99",X"77",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"88",X"89",X"88",X"99",X"88",X"77",X"89",X"77",X"89",X"77",X"88",X"77",X"88",X"99",X"88",X"89",
		X"98",X"71",X"79",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"79",X"71",X"98",X"71",
		X"88",X"97",X"88",X"77",X"89",X"79",X"97",X"98",X"77",X"98",X"44",X"44",X"77",X"77",X"11",X"11",
		X"98",X"71",X"98",X"71",X"79",X"71",X"98",X"61",X"88",X"71",X"44",X"71",X"76",X"71",X"11",X"11",
		X"EE",X"EE",X"CC",X"CC",X"FF",X"FF",X"EC",X"88",X"EC",X"88",X"EC",X"88",X"EC",X"88",X"CD",X"F8",
		X"EE",X"EE",X"CC",X"CC",X"FF",X"FF",X"EC",X"71",X"EC",X"71",X"EC",X"71",X"EC",X"71",X"CD",X"F1",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"98",X"97",X"98",X"89",X"79",X"88",X"77",X"88",X"97",
		X"44",X"41",X"77",X"71",X"11",X"71",X"88",X"71",X"88",X"71",X"78",X"71",X"98",X"71",X"98",X"71",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"87",X"DC",X"87",X"DC",X"87",X"DC",X"87",X"CE",X"F7",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"CE",X"F0",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"88",X"DC",X"88",X"DC",X"88",X"DC",X"88",X"CE",X"F8",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"CE",X"F0",
		X"F7",X"77",X"FF",X"77",X"CC",X"77",X"CC",X"F7",X"EE",X"FF",X"FF",X"CC",X"11",X"CC",X"77",X"EE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"F7",X"77",X"FF",X"77",
		X"77",X"FF",X"88",X"11",X"77",X"77",X"17",X"77",X"F1",X"88",X"EF",X"77",X"EE",X"11",X"EE",X"FF",
		X"CC",X"77",X"CC",X"F7",X"EE",X"FF",X"FF",X"CC",X"11",X"CC",X"77",X"EE",X"77",X"FF",X"88",X"11",
		X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",
		X"77",X"71",X"77",X"77",X"77",X"77",X"17",X"77",X"91",X"77",X"99",X"77",X"91",X"17",X"91",X"91",
		X"99",X"99",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",X"91",X"91",X"8C",X"99",X"EC",X"F9",
		X"77",X"77",X"77",X"77",X"77",X"77",X"99",X"77",X"99",X"77",X"FF",X"DD",X"CC",X"EE",X"CC",X"DD",
		X"44",X"44",X"88",X"81",X"77",X"77",X"99",X"99",X"94",X"84",X"94",X"84",X"98",X"48",X"98",X"48",
		X"44",X"44",X"88",X"81",X"77",X"71",X"99",X"71",X"84",X"71",X"84",X"71",X"48",X"71",X"48",X"71",
		X"78",X"87",X"78",X"87",X"78",X"87",X"78",X"87",X"78",X"87",X"78",X"87",X"78",X"87",X"78",X"87",
		X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",
		X"44",X"44",X"77",X"77",X"99",X"92",X"92",X"77",X"99",X"77",X"97",X"77",X"97",X"77",X"27",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"77",X"99",X"77",X"77",X"99",X"99",X"97",X"99",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"77",X"77",X"99",X"77",X"77",X"77",X"87",X"77",
		X"44",X"44",X"77",X"71",X"99",X"71",X"79",X"71",X"79",X"71",X"77",X"71",X"77",X"71",X"77",X"71",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",
		X"77",X"99",X"78",X"99",X"88",X"79",X"88",X"89",X"99",X"99",X"99",X"78",X"79",X"88",X"77",X"88",
		X"27",X"77",X"97",X"77",X"97",X"77",X"99",X"77",X"92",X"77",X"99",X"92",X"77",X"77",X"11",X"11",
		X"97",X"88",X"99",X"88",X"77",X"77",X"77",X"99",X"77",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"87",X"97",X"79",X"97",X"99",X"79",X"99",X"79",X"88",X"79",X"88",X"79",X"78",X"97",X"97",X"97",
		X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",
		X"97",X"77",X"77",X"77",X"99",X"77",X"77",X"77",X"77",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"77",X"71",X"77",X"71",X"77",X"71",X"79",X"71",X"79",X"71",X"99",X"71",X"77",X"71",X"11",X"11",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"CE",X"F0",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"CE",X"F0",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"77",X"77",X"99",X"77",X"77",X"77",X"87",X"77",
		X"44",X"41",X"77",X"71",X"11",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",
		X"27",X"00",X"0A",X"70",X"00",X"80",X"0A",X"98",X"2A",X"AA",X"92",X"9A",X"A7",X"22",X"9A",X"99",
		X"00",X"00",X"00",X"00",X"20",X"00",X"97",X"00",X"A9",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"99",X"A0",X"99",X"AA",X"99",X"92",X"99",X"78",X"AA",X"89",X"77",X"99",X"8A",X"99",X"70",X"88",
		X"00",X"00",X"22",X"00",X"99",X"00",X"17",X"82",X"99",X"99",X"00",X"01",X"70",X"00",X"99",X"90",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"DD",X"EE",X"ED",X"CC",X"FD",X"CC",X"ED",X"EE",X"ED",X"EE",X"ED",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"DD",X"DE",X"EE",X"DE",X"FF",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",
		X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",
		X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",
		X"77",X"77",X"11",X"29",X"82",X"82",X"27",X"98",X"79",X"99",X"29",X"88",X"82",X"82",X"98",X"27",
		X"77",X"77",X"11",X"71",X"82",X"87",X"27",X"98",X"79",X"99",X"29",X"88",X"82",X"82",X"98",X"27",
		X"99",X"79",X"88",X"29",X"82",X"82",X"27",X"98",X"79",X"99",X"79",X"88",X"77",X"87",X"99",X"99",
		X"99",X"79",X"88",X"79",X"82",X"87",X"27",X"98",X"79",X"99",X"79",X"88",X"77",X"87",X"99",X"99",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"66",X"44",X"44",X"77",X"77",X"11",X"11",
		X"76",X"71",X"66",X"71",X"99",X"71",X"97",X"71",X"99",X"71",X"44",X"71",X"77",X"71",X"11",X"11",
		X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",
		X"FD",X"EF",X"FD",X"EF",X"FD",X"EF",X"FD",X"EF",X"FD",X"EF",X"FD",X"EF",X"FD",X"EF",X"FD",X"EF",
		X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",
		X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",
		X"FF",X"ED",X"CC",X"ED",X"DD",X"ED",X"EE",X"ED",X"FF",X"ED",X"CC",X"ED",X"DD",X"FF",X"EE",X"FF",
		X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"DE",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"FF",X"00",X"EC",X"0F",X"0E",X"FC",X"00",X"CC",X"0E",X"CE",X"CC",X"EF",X"E1",X"11",X"00",X"88",
		X"FF",X"CC",X"CC",X"CC",X"CC",X"EE",X"ED",X"FE",X"FF",X"FE",X"FF",X"FE",X"11",X"11",X"88",X"88",
		X"22",X"22",X"11",X"11",X"22",X"77",X"08",X"88",X"00",X"88",X"00",X"11",X"00",X"00",X"00",X"00",
		X"77",X"77",X"18",X"18",X"77",X"77",X"81",X"81",X"81",X"81",X"11",X"11",X"11",X"11",X"11",X"11",
		X"EF",X"18",X"FF",X"47",X"F1",X"71",X"18",X"17",X"87",X"78",X"47",X"88",X"71",X"88",X"17",X"11",
		X"77",X"77",X"81",X"81",X"77",X"77",X"44",X"47",X"88",X"87",X"81",X"11",X"11",X"11",X"11",X"11",
		X"78",X"11",X"88",X"19",X"81",X"99",X"19",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"77",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"77",X"77",X"77",X"77",
		X"88",X"88",X"99",X"99",X"07",X"47",X"88",X"88",X"77",X"77",X"00",X"88",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"70",X"77",X"00",X"77",X"0F",X"70",X"FC",X"DD",X"CD",X"EF",X"CE",X"FC",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CC",X"CF",X"DC",X"FC",X"ED",X"CC",X"EF",X"CE",X"FC",X"CD",X"CC",X"CC",X"CE",X"FC",
		X"CC",X"CC",X"CE",X"FC",X"CD",X"9F",X"CC",X"99",X"FC",X"87",X"9F",X"71",X"99",X"17",X"87",X"77",
		X"CD",X"9F",X"CC",X"99",X"FC",X"87",X"9F",X"71",X"99",X"17",X"87",X"77",X"7C",X"77",X"EC",X"F7",
		X"71",X"77",X"17",X"77",X"77",X"77",X"77",X"71",X"D7",X"17",X"77",X"97",X"7C",X"97",X"EC",X"F7",
		X"78",X"17",X"89",X"77",X"91",X"77",X"17",X"77",X"77",X"77",X"77",X"79",X"77",X"11",X"77",X"71",
		X"EE",X"88",X"ED",X"88",X"D9",X"88",X"88",X"88",X"88",X"88",X"11",X"18",X"71",X"71",X"71",X"71",
		X"71",X"78",X"19",X"79",X"71",X"71",X"71",X"71",X"78",X"78",X"79",X"79",X"7C",X"71",X"EC",X"F8",
		X"78",X"78",X"79",X"79",X"71",X"71",X"71",X"71",X"78",X"78",X"79",X"71",X"7C",X"71",X"EC",X"F8",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"7F",X"77",X"FF",X"77",X"FC",X"7F",X"CC",
		X"77",X"FF",X"7F",X"CC",X"FF",X"CC",X"FC",X"EE",X"CC",X"FF",X"CE",X"11",X"EF",X"77",X"F1",X"77",
		X"FF",X"CE",X"FC",X"EF",X"CC",X"F1",X"CE",X"17",X"EF",X"77",X"F1",X"78",X"17",X"87",X"77",X"71",
		X"17",X"88",X"77",X"77",X"78",X"11",X"87",X"FF",X"71",X"EE",X"11",X"EE",X"FF",X"EE",X"EE",X"EE",
		X"88",X"88",X"77",X"77",X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",
		X"88",X"88",X"77",X"79",X"99",X"79",X"91",X"79",X"91",X"79",X"91",X"79",X"99",X"79",X"91",X"79",
		X"88",X"88",X"77",X"77",X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"99",X"99",X"91",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"91",X"91",X"91",X"91",X"98",X"98",X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"91",
		X"91",X"91",X"91",X"91",X"98",X"98",X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"91",
		X"98",X"98",X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"98",X"98",X"77",X"77",X"99",X"99",
		X"98",X"98",X"99",X"99",X"91",X"91",X"91",X"91",X"91",X"91",X"98",X"98",X"77",X"77",X"99",X"99",
		X"91",X"79",X"91",X"79",X"98",X"79",X"99",X"79",X"91",X"79",X"91",X"79",X"91",X"79",X"91",X"79",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"79",X"99",X"79",X"91",X"79",X"91",X"79",X"91",X"79",X"98",X"79",X"77",X"79",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"77",X"16",X"77",X"16",X"77",X"16",X"77",X"16",X"77",X"16",X"77",X"16",X"77",X"16",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"19",X"77",X"19",X"77",X"19",X"67",X"19",X"66",X"19",X"99",X"44",X"44",X"77",X"77",X"11",X"11",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"66",X"44",X"44",X"77",X"77",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"EE",X"EE",X"CC",X"CC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"A7",X"66",X"7E",X"EE",X"7E",X"CC",X"8E",X"BB",X"8E",X"BB",X"8E",X"BB",X"8B",X"BB",X"8B",X"BB",
		X"68",X"22",X"88",X"72",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"BE",X"DD",X"EE",X"DD",X"EE",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"D7",X"DD",X"DD",X"DD",X"BB",X"DB",X"BB",X"DB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"BB",X"DD",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"88",X"BB",X"88",
		X"DD",X"8B",X"DD",X"88",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",
		X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",
		X"69",X"78",X"EE",X"77",X"DD",X"98",X"BB",X"98",X"BB",X"99",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",
		X"66",X"66",X"EE",X"EE",X"ED",X"DD",X"DB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"9D",X"DD",X"9D",X"DB",X"9D",X"DB",X"9D",X"BB",X"9D",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"8B",X"B7",X"8B",X"B7",X"8B",X"B7",X"8B",X"B7",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",
		X"97",X"70",X"97",X"70",X"97",X"70",X"97",X"70",X"97",X"70",X"97",X"70",X"97",X"70",X"97",X"70",
		X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",
		X"97",X"70",X"C7",X"77",X"B9",X"77",X"B9",X"77",X"B9",X"77",X"B9",X"77",X"B9",X"77",X"B9",X"77",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"EE",
		X"98",X"77",X"98",X"77",X"98",X"77",X"98",X"77",X"98",X"77",X"98",X"77",X"98",X"77",X"BB",X"77",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"88",X"BB",X"BB",
		X"B9",X"77",X"B9",X"77",X"B9",X"77",X"B9",X"77",X"B8",X"77",X"B8",X"77",X"77",X"77",X"98",X"77",
		X"BD",X"DD",X"DD",X"DD",X"DD",X"BB",X"DB",X"BD",X"DB",X"DB",X"DB",X"BB",X"DB",X"BD",X"DB",X"BD",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"AA",X"DD",X"8A",X"BB",X"8A",X"BB",X"8A",X"DB",X"8A",X"B9",X"8A",X"B9",X"88",X"B9",X"88",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",
		X"BE",X"DE",X"EE",X"ED",X"EE",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BE",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"8D",X"DD",X"D8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",
		X"DD",X"AA",X"DD",X"8A",X"BB",X"8A",X"BB",X"8A",X"BB",X"8A",X"8B",X"8A",X"8B",X"88",X"8B",X"88",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"8B",X"88",X"8B",X"88",X"B8",X"88",X"B8",X"88",X"B8",X"88",X"B8",X"88",X"B9",X"88",X"B9",X"88",
		X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",
		X"BE",X"ED",X"EE",X"DD",X"EE",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BE",
		X"DD",X"D9",X"DE",X"D9",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",
		X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",
		X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",
		X"DD",X"ED",X"DD",X"ED",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",
		X"DD",X"BB",X"DD",X"8B",X"9B",X"8B",X"9B",X"8B",X"9B",X"8B",X"9B",X"8B",X"9B",X"88",X"B9",X"88",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",X"B9",X"88",
		X"66",X"66",X"EE",X"EE",X"EE",X"DD",X"EE",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",
		X"66",X"66",X"EE",X"EE",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"EE",X"BB",X"ED",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"27",X"66",X"7E",X"EE",X"7E",X"CC",X"8E",X"BB",X"8E",X"BB",X"8E",X"BB",X"8B",X"BB",X"8B",X"BB",
		X"68",X"22",X"88",X"72",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",
		X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",
		X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",
		X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",
		X"66",X"66",X"EE",X"EE",X"EE",X"DD",X"EE",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",
		X"99",X"77",X"B9",X"77",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"66",X"8B",X"E8",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"66",X"BB",X"EE",X"86",X"DD",X"EE",X"BB",X"DE",X"BB",X"ED",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",
		X"BB",X"BB",X"66",X"66",X"EE",X"EE",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"66",X"66",X"8E",X"EE",X"89",X"DD",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"B8",X"BB",X"B8",
		X"66",X"00",X"EE",X"90",X"DD",X"87",X"BA",X"87",X"BA",X"87",X"BA",X"87",X"BA",X"87",X"BA",X"87",
		X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"BB",
		X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"66",X"66",X"EE",X"EE",X"EE",X"DD",X"EE",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",
		X"99",X"77",X"B9",X"77",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"66",X"8D",X"E8",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"E9",X"7D",X"EE",X"77",X"DD",X"98",X"BB",X"98",X"BB",X"99",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",
		X"EE",X"EE",X"EE",X"EE",X"ED",X"DD",X"DB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"DD",X"EE",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",
		X"99",X"77",X"B9",X"77",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"EE",X"8B",X"E8",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"BE",X"EE",X"EE",X"EE",X"EE",X"DD",X"EE",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",
		X"EE",X"EE",X"EE",X"EE",X"CC",X"CC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"B7",X"EE",X"7E",X"EE",X"7E",X"CC",X"8E",X"BB",X"8E",X"BB",X"8E",X"BB",X"8B",X"BB",X"8B",X"BB",
		X"EE",X"8B",X"E8",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"DD",X"EE",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",X"ED",X"BB",
		X"99",X"77",X"B9",X"77",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"EE",X"8D",X"E8",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",X"88",X"77",
		X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",X"B8",X"87",
		X"69",X"72",X"EE",X"77",X"DD",X"98",X"BB",X"98",X"BB",X"99",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",
		X"66",X"66",X"EE",X"EE",X"ED",X"DD",X"DB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"E7",X"60",X"7E",X"E0",X"7E",X"C0",X"8E",X"B0",X"8E",X"B0",X"8E",X"B0",X"8B",X"B0",X"8B",X"B0",
		X"BB",X"BB",X"DD",X"7B",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",
		X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",
		X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"2E",X"E2",X"2E",X"66",X"E6",X"6C",X"66",X"CE",X"66",X"EE",X"CC",X"EE",X"CE",X"EE",X"CE",X"EE",
		X"EE",X"EE",X"66",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"DE",X"EE",X"ED",X"EE",
		X"CC",X"EE",X"2B",X"EE",X"BC",X"EE",X"BC",X"EE",X"BC",X"CC",X"2B",X"CC",X"22",X"BB",X"22",X"22",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",X"ED",X"CB",X"CC",X"BB",X"BB",X"22",X"22",X"22",X"22",X"22",
		X"66",X"22",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6D",X"D6",X"DD",X"D6",
		X"66",X"66",X"66",X"66",X"66",X"66",X"EC",X"66",X"EC",X"66",X"EC",X"DD",X"6E",X"DD",X"6E",X"CD",
		X"66",X"66",X"DD",X"66",X"ED",X"DE",X"EE",X"EE",X"CC",X"EC",X"BB",X"CB",X"22",X"BB",X"22",X"22",
		X"6E",X"CC",X"EE",X"CC",X"CC",X"EE",X"BB",X"CC",X"22",X"BB",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"66",X"66",X"EE",X"66",X"66",X"6E",X"66",X"6E",X"66",X"ED",X"66",X"ED",X"EE",X"E6",X"DD",
		X"22",X"66",X"66",X"66",X"E6",X"66",X"6E",X"66",X"66",X"66",X"66",X"66",X"ED",X"66",X"D6",X"66",
		X"66",X"66",X"E6",X"66",X"EE",X"66",X"DD",X"EE",X"CC",X"DD",X"BB",X"CD",X"22",X"BC",X"22",X"2B",
		X"66",X"66",X"66",X"EE",X"66",X"ED",X"6E",X"DC",X"ED",X"CB",X"DC",X"B2",X"CB",X"22",X"B2",X"22",
		X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"60",X"00",X"66",X"00",X"06",X"00",
		X"60",X"00",X"06",X"00",X"00",X"60",X"00",X"66",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"60",
		X"06",X"00",X"06",X"00",X"06",X"00",X"00",X"00",X"00",X"66",X"66",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"60",X"00",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"24",X"22",X"20",X"12",X"14",X"14",X"10",X"11",X"21",X"1D",X"14",X"41",X"D0",X"10",X"41",X"2A",
		X"41",X"1D",X"41",X"11",X"01",X"4D",X"D0",X"11",X"4D",X"1D",X"01",X"4D",X"4D",X"02",X"41",X"4D",
		X"0D",X"04",X"4A",X"A0",X"0E",X"CA",X"AA",X"CD",X"A4",X"0D",X"0A",X"EE",X"EA",X"EA",X"EE",X"EE",
		X"0A",X"0A",X"04",X"DE",X"A0",X"00",X"00",X"AA",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"ED",
		X"14",X"C4",X"C2",X"C1",X"1C",X"2C",X"C2",X"04",X"1C",X"4C",X"0C",X"CC",X"4C",X"4B",X"02",X"0C",
		X"14",X"40",X"C2",X"11",X"4C",X"02",X"0C",X"20",X"24",X"4C",X"2C",X"04",X"0C",X"2B",X"B4",X"4B",
		X"B0",X"B4",X"4B",X"B0",X"0B",X"B4",X"BB",X"1B",X"42",X"4B",X"B0",X"0B",X"B4",X"BB",X"B0",X"BB",
		X"C0",X"0B",X"1B",X"1C",X"BB",X"0B",X"B4",X"BB",X"B0",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"F4",X"0B",X"20",X"1C",X"CF",X"C4",X"10",X"C1",X"2C",X"1F",X"F4",X"41",X"C0",X"B0",X"4B",X"2B",
		X"4C",X"F0",X"4C",X"B1",X"0F",X"4C",X"C0",X"C1",X"4C",X"1B",X"01",X"4F",X"4C",X"02",X"4C",X"4B",
		X"0C",X"BF",X"4B",X"B0",X"FC",X"BB",X"0B",X"CB",X"B4",X"BB",X"B0",X"BB",X"BF",X"BB",X"B0",X"BB",
		X"0C",X"FB",X"FB",X"0B",X"04",X"BB",X"B0",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"14",X"A4",X"A2",X"A1",X"1A",X"2A",X"F2",X"04",X"1A",X"4A",X"0A",X"BF",X"4E",X"4B",X"02",X"0B",
		X"14",X"40",X"A2",X"11",X"4B",X"F2",X"FA",X"20",X"24",X"4A",X"2A",X"04",X"0A",X"AA",X"A4",X"4A",
		X"B0",X"B4",X"FE",X"E0",X"0B",X"EF",X"BB",X"1B",X"42",X"FE",X"E0",X"0E",X"EF",X"EE",X"EE",X"E0",
		X"A0",X"0E",X"EA",X"FE",X"BD",X"0E",X"B4",X"EE",X"E0",X"EE",X"EB",X"00",X"0B",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"1A",
		X"28",X"22",X"22",X"82",X"21",X"21",X"12",X"12",X"21",X"21",X"11",X"11",X"01",X"01",X"00",X"00",
		X"28",X"22",X"22",X"82",X"21",X"22",X"12",X"12",X"21",X"21",X"11",X"11",X"01",X"01",X"00",X"00",
		X"A0",X"A0",X"AA",X"AA",X"BA",X"BA",X"BB",X"DB",X"BC",X"DB",X"CC",X"DB",X"AA",X"CB",X"AA",X"CC",
		X"A0",X"A0",X"AA",X"AA",X"BA",X"BA",X"BB",X"CB",X"CE",X"CC",X"BE",X"CC",X"B0",X"CE",X"BA",X"CA",
		X"62",X"21",X"12",X"26",X"10",X"21",X"12",X"21",X"11",X"11",X"31",X"11",X"11",X"00",X"00",X"00",
		X"21",X"16",X"21",X"21",X"26",X"22",X"21",X"11",X"11",X"11",X"31",X"31",X"11",X"00",X"00",X"00",
		X"00",X"AA",X"AA",X"AA",X"CC",X"AB",X"BC",X"AA",X"CD",X"BA",X"CD",X"BA",X"CD",X"BB",X"CD",X"BB",
		X"00",X"AA",X"AA",X"AA",X"AA",X"BB",X"BB",X"BB",X"BB",X"BC",X"BB",X"BC",X"BD",X"BD",X"BD",X"BB",
		X"50",X"05",X"01",X"50",X"81",X"81",X"05",X"05",X"20",X"80",X"22",X"02",X"52",X"25",X"00",X"00",
		X"18",X"05",X"50",X"80",X"51",X"01",X"08",X"11",X"20",X"25",X"25",X"20",X"50",X"5C",X"0C",X"0C",
		X"CC",X"CC",X"CC",X"BB",X"BB",X"CC",X"CC",X"CC",X"CC",X"BB",X"CC",X"CC",X"CB",X"CC",X"CC",X"CC",
		X"BB",X"CC",X"CC",X"BC",X"BB",X"CB",X"CC",X"CC",X"CC",X"CB",X"CC",X"BB",X"BC",X"CC",X"CC",X"CC",
		X"12",X"12",X"23",X"21",X"21",X"11",X"11",X"10",X"11",X"00",X"11",X"0A",X"01",X"AA",X"C1",X"CB",
		X"21",X"22",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"10",X"10",X"10",X"1A",X"0A",
		X"C1",X"CD",X"C0",X"CE",X"C0",X"DE",X"CA",X"EE",X"CA",X"EE",X"EB",X"EE",X"EB",X"EE",X"ED",X"EE",
		X"1A",X"0A",X"1A",X"AA",X"1B",X"AA",X"0B",X"AA",X"0B",X"AD",X"AB",X"AD",X"AB",X"AD",X"BB",X"DD",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"C0",X"CC",X"0C",X"C0",X"CC",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"0C",X"CC",X"CC",X"CC",
		X"BB",X"BB",X"CC",X"BC",X"BB",X"BC",X"BB",X"BB",X"BB",X"CA",X"CA",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"AB",X"BB",X"BA",X"BB",X"BA",X"BB",X"BC",X"BB",X"CB",X"AB",X"CB",X"AB",X"BB",X"CB",X"AB",X"BA",
		X"CB",X"BC",X"BA",X"BC",X"BA",X"AB",X"BC",X"BA",X"CC",X"BA",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BA",X"BA",X"BA",X"BB",X"BB",X"BB",X"CC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"14",X"14",X"22",X"11",X"11",X"21",X"72",X"04",X"11",X"4E",X"0D",X"D7",X"42",X"4E",X"02",X"01",
		X"14",X"40",X"11",X"11",X"41",X"72",X"72",X"20",X"24",X"4B",X"2D",X"04",X"0A",X"2B",X"A4",X"4B",
		X"E0",X"E4",X"7D",X"E0",X"0E",X"E7",X"EE",X"1E",X"42",X"7E",X"E0",X"0E",X"E7",X"EE",X"E0",X"EE",
		X"A0",X"0D",X"1A",X"7D",X"AA",X"0D",X"B4",X"BD",X"B0",X"AD",X"BB",X"BD",X"BB",X"BD",X"BB",X"DD",
		X"DE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",
		X"CE",X"DD",X"CE",X"DD",X"CE",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",
		X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",
		X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"DC",X"DD",X"DC",X"DD",X"DC",X"DD",
		X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",
		X"DC",X"DD",X"DD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",
		X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"1E",X"DD",X"1E",X"D1",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DC",X"EE",X"D1",X"EE",X"D1",X"EE",X"16",X"22",
		X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"AD",X"BB",X"AD",X"BB",X"AD",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",
		X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",
		X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"AA",X"BB",X"AA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AD",X"BA",X"AD",X"BA",X"AD",X"BA",X"AD",
		X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"22",X"BB",
		X"BB",X"AD",X"BB",X"AD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"82",X"21",X"22",
		X"ED",X"EE",X"EE",X"EE",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"DD",X"EB",X"DE",X"DA",X"DE",X"EB",
		X"AB",X"DD",X"AB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"AA",X"DD",X"BB",X"DE",X"BB",X"DD",
		X"DE",X"EB",X"DE",X"EE",X"DE",X"EE",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"DE",X"DD",X"ED",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"BD",X"BD",X"DD",X"BD",X"DD",X"AD",X"DD",X"BD",X"BD",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"CE",
		X"BD",X"DD",X"BD",X"DE",X"BD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DD",X"DD",X"DD",X"DD",X"EB",
		X"DD",X"EE",X"DD",X"EC",X"DD",X"EE",X"DD",X"EE",X"DD",X"DE",X"EB",X"2E",X"12",X"21",X"22",X"22",
		X"DD",X"EB",X"DD",X"EB",X"DD",X"DB",X"DD",X"DD",X"DD",X"DD",X"11",X"11",X"22",X"21",X"22",X"22",
		X"BD",X"EE",X"BD",X"EE",X"AD",X"EE",X"0D",X"EE",X"AD",X"EE",X"0D",X"EE",X"CD",X"EB",X"DD",X"BB",
		X"CC",X"BB",X"B0",X"AE",X"B0",X"EE",X"BA",X"EE",X"AA",X"DE",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",
		X"DD",X"BB",X"DD",X"CC",X"CD",X"AA",X"DD",X"DA",X"DD",X"DA",X"DE",X"DD",X"DE",X"ED",X"22",X"ED",
		X"BB",X"AA",X"BB",X"AC",X"CB",X"CC",X"EA",X"0C",X"EE",X"0C",X"EE",X"A0",X"EE",X"A1",X"EE",X"11",
		X"BD",X"EE",X"BD",X"EE",X"AD",X"EE",X"0D",X"EE",X"AD",X"EE",X"0D",X"EE",X"CD",X"EB",X"DD",X"BB",
		X"CC",X"BB",X"B0",X"AE",X"B0",X"EE",X"BA",X"EE",X"AA",X"DE",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",
		X"DD",X"BB",X"DD",X"CC",X"CD",X"AA",X"DD",X"DA",X"DD",X"DA",X"DE",X"DD",X"DE",X"ED",X"DE",X"ED",
		X"BB",X"AA",X"BB",X"AC",X"CB",X"CC",X"EA",X"0C",X"EE",X"0C",X"EE",X"A0",X"EE",X"A0",X"EE",X"A0",
		X"CB",X"DE",X"CC",X"DE",X"CC",X"EE",X"CC",X"EE",X"EE",X"CA",X"EE",X"CB",X"EE",X"AC",X"EE",X"AC",
		X"0B",X"C0",X"A0",X"CD",X"AB",X"CD",X"0B",X"DD",X"BB",X"DD",X"BB",X"BA",X"CB",X"BB",X"CE",X"BB",
		X"DB",X"BC",X"D0",X"BC",X"BB",X"BD",X"BB",X"CD",X"BB",X"CD",X"BB",X"CE",X"BC",X"EE",X"BC",X"EE",
		X"EE",X"CC",X"EE",X"AC",X"EE",X"A0",X"DE",X"A0",X"DD",X"CC",X"BD",X"CC",X"CC",X"CC",X"AC",X"CC",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"CE",
		X"BD",X"DD",X"BD",X"DE",X"BD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DD",X"DD",X"DD",X"DD",X"EB",
		X"DD",X"EE",X"DD",X"EC",X"DD",X"EE",X"DD",X"EE",X"DD",X"DE",X"EB",X"1E",X"11",X"11",X"21",X"21",
		X"DD",X"EB",X"DD",X"EB",X"DD",X"DB",X"DD",X"DD",X"DD",X"DD",X"11",X"11",X"11",X"11",X"22",X"11",
		X"DB",X"DB",X"BD",X"BD",X"DB",X"DC",X"CC",X"CD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"CD",X"CC",
		X"DB",X"DB",X"BD",X"CC",X"CC",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DC",X"CC",X"CC",X"DE",
		X"CC",X"CD",X"DE",X"DE",X"ED",X"ED",X"DE",X"DE",X"ED",X"ED",X"DE",X"DC",X"DC",X"CB",X"BD",X"BD",
		X"ED",X"ED",X"DE",X"DE",X"ED",X"ED",X"DE",X"DE",X"ED",X"CC",X"CD",X"BD",X"DB",X"DB",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"60",X"60",X"00",X"06",X"00",X"06",X"00",X"60",X"00",X"00",X"60",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
