library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"66",X"33",X"33",X"33",X"22",X"CC",X"00",X"11",X"22",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"00",
		X"EE",X"33",X"77",X"EE",X"88",X"00",X"FF",X"00",X"33",X"66",X"00",X"11",X"33",X"66",X"77",X"00",
		X"FF",X"66",X"CC",X"EE",X"33",X"33",X"EE",X"00",X"77",X"00",X"00",X"11",X"00",X"44",X"33",X"00",
		X"EE",X"66",X"66",X"66",X"FF",X"66",X"66",X"00",X"00",X"11",X"22",X"44",X"77",X"00",X"00",X"00",
		X"FF",X"00",X"EE",X"33",X"33",X"33",X"EE",X"00",X"77",X"66",X"77",X"00",X"00",X"44",X"33",X"00",
		X"EE",X"00",X"00",X"EE",X"33",X"33",X"EE",X"00",X"11",X"22",X"66",X"77",X"66",X"66",X"33",X"00",
		X"FF",X"33",X"66",X"CC",X"88",X"88",X"88",X"00",X"77",X"44",X"00",X"00",X"11",X"11",X"11",X"00",
		X"EE",X"33",X"33",X"CC",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"11",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"FF",X"33",X"22",X"CC",X"00",X"33",X"66",X"66",X"33",X"00",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"44",X"00",X"00",X"00",
		X"CC",X"AA",X"DD",X"AA",X"99",X"AA",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",
		X"CC",X"22",X"99",X"11",X"11",X"99",X"22",X"CC",X"33",X"44",X"99",X"AA",X"AA",X"99",X"44",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"33",X"33",X"FF",X"33",X"33",X"00",X"11",X"22",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"EE",X"33",X"33",X"EE",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"77",X"00",
		X"EE",X"33",X"00",X"00",X"00",X"33",X"EE",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"CC",X"66",X"33",X"33",X"33",X"66",X"CC",X"00",X"77",X"66",X"66",X"66",X"66",X"66",X"77",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"EE",X"33",X"00",X"77",X"33",X"33",X"FF",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"33",X"33",X"33",X"FF",X"33",X"33",X"33",X"00",X"66",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"EE",X"88",X"88",X"88",X"88",X"88",X"EE",X"00",X"77",X"11",X"11",X"11",X"11",X"11",X"77",X"00",
		X"FF",X"66",X"66",X"66",X"66",X"66",X"CC",X"00",X"11",X"00",X"00",X"00",X"66",X"66",X"33",X"00",
		X"33",X"66",X"CC",X"88",X"CC",X"66",X"33",X"00",X"66",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"33",X"33",X"33",X"33",X"33",X"77",X"00",
		X"33",X"77",X"FF",X"BB",X"33",X"33",X"33",X"00",X"66",X"77",X"77",X"66",X"66",X"66",X"66",X"00",
		X"33",X"33",X"BB",X"FF",X"77",X"33",X"33",X"00",X"66",X"77",X"77",X"66",X"66",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"33",X"EE",X"00",X"00",X"00",X"77",X"66",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"33",X"FF",X"22",X"DD",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"EE",X"CC",X"66",X"33",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"EE",X"33",X"00",X"EE",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"33",X"00",X"66",X"33",X"00",
		X"EE",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"77",X"11",X"11",X"11",X"11",X"11",X"11",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"33",X"33",X"33",X"33",X"66",X"CC",X"88",X"00",X"66",X"66",X"66",X"66",X"33",X"11",X"00",X"00",
		X"33",X"33",X"33",X"BB",X"FF",X"77",X"22",X"00",X"66",X"66",X"66",X"66",X"77",X"77",X"22",X"00",
		X"33",X"66",X"CC",X"CC",X"EE",X"77",X"33",X"00",X"66",X"77",X"33",X"11",X"33",X"66",X"44",X"00",
		X"66",X"66",X"66",X"CC",X"88",X"88",X"88",X"00",X"66",X"66",X"66",X"33",X"11",X"11",X"11",X"00",
		X"FF",X"77",X"EE",X"CC",X"88",X"00",X"FF",X"00",X"77",X"00",X"00",X"11",X"33",X"77",X"77",X"00",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"0E",X"0C",X"00",X"11",X"11",X"11",X"11",X"33",X"0F",X"07",
		X"00",X"00",X"00",X"88",X"CC",X"0E",X"0C",X"0E",X"00",X"00",X"03",X"07",X"03",X"07",X"CF",X"EF",
		X"00",X"80",X"50",X"8A",X"0A",X"0C",X"08",X"08",X"00",X"00",X"77",X"FF",X"7F",X"0F",X"0F",X"0F",
		X"00",X"70",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"10",X"10",X"10",X"10",
		X"00",X"88",X"FF",X"11",X"11",X"33",X"EE",X"EE",X"FF",X"11",X"FF",X"EE",X"EE",X"FF",X"FF",X"FF",
		X"CC",X"00",X"33",X"FF",X"FF",X"EE",X"CC",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"88",X"FF",X"77",X"77",X"FF",X"FF",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"77",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"00",X"CC",X"FF",X"FF",X"77",X"33",X"00",
		X"66",X"9F",X"9F",X"66",X"00",X"00",X"00",X"00",X"66",X"9F",X"9F",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"03",X"0F",X"03",X"01",X"03",X"0F",X"03",X"08",X"0C",X"0F",X"0C",X"08",X"0C",X"0F",X"0C",
		X"01",X"03",X"0F",X"03",X"01",X"03",X"0F",X"01",X"08",X"0C",X"0F",X"0C",X"08",X"0C",X"0F",X"08",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"EE",X"CC",X"CC",X"CC",X"EE",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"02",X"04",X"08",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"04",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"0C",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"0A",X"02",X"02",X"09",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"02",X"0A",X"0A",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"04",
		X"02",X"0A",X"0A",X"01",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"02",X"01",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"0E",X"01",X"01",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"20",X"40",X"C0",X"B0",X"E0",X"00",X"00",X"10",X"10",X"30",X"20",X"78",X"3C",X"1E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"4F",X"2F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"4F",X"2F",X"9F",X"0F",X"0F",X"0E",X"08",X"00",X"03",X"13",X"07",X"47",X"2F",X"0F",X"0F",X"0E",
		X"03",X"03",X"05",X"09",X"01",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"03",X"0C",X"00",X"00",
		X"CE",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"33",X"75",X"FB",X"FB",X"FF",X"FF",X"77",X"33",
		X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"74",X"FD",X"FD",X"FF",
		X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"0C",X"4E",X"0F",X"8F",
		X"8C",X"0C",X"80",X"00",X"00",X"00",X"00",X"00",X"2F",X"FC",X"FC",X"CC",X"CC",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2F",X"3C",X"70",X"00",X"11",X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",
		X"00",X"08",X"0C",X"8C",X"8C",X"0C",X"08",X"00",X"E0",X"D2",X"C3",X"87",X"0F",X"1F",X"0F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"D2",X"1E",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"01",X"03",X"03",X"03",X"03",X"01",X"00",
		X"0E",X"0F",X"0B",X"0F",X"0E",X"06",X"0C",X"0C",X"00",X"03",X"07",X"0A",X"0F",X"05",X"0F",X"0A",
		X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"0F",X"0D",X"0E",X"78",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"83",X"C3",X"83",X"C2",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",
		X"83",X"82",X"83",X"83",X"B0",X"70",X"F0",X"E0",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"F0",
		X"A0",X"B0",X"80",X"F0",X"00",X"F0",X"88",X"88",X"20",X"20",X"20",X"A8",X"6C",X"7C",X"FF",X"4F",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"4F",X"FF",X"4F",X"4F",X"FF",X"4E",X"4C",X"00",
		X"00",X"00",X"00",X"77",X"2F",X"2F",X"FF",X"2F",X"00",X"00",X"00",X"00",X"11",X"13",X"33",X"17",
		X"2F",X"FF",X"2F",X"2F",X"FF",X"2F",X"2F",X"FF",X"17",X"FF",X"9F",X"9F",X"FF",X"17",X"13",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0A",
		X"1E",X"3C",X"3C",X"68",X"E0",X"C0",X"C0",X"00",X"0F",X"0A",X"0F",X"0B",X"1E",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"86",
		X"0F",X"0A",X"0F",X"0E",X"87",X"F0",X"F0",X"F0",X"87",X"C3",X"C3",X"61",X"70",X"30",X"30",X"00",
		X"10",X"20",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"00",X"F0",X"76",X"FC",X"F9",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"EE",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"77",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"67",X"DF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"8E",X"4E",X"FF",X"88",X"0C",X"0F",X"AF",X"3F",X"2F",X"6F",
		X"8E",X"0E",X"4E",X"8C",X"0C",X"08",X"00",X"00",X"AF",X"3F",X"6F",X"AF",X"3F",X"2F",X"6F",X"0E",
		X"33",X"00",X"13",X"0F",X"4F",X"9F",X"9F",X"BF",X"00",X"00",X"00",X"00",X"01",X"03",X"27",X"17",
		X"9F",X"DF",X"BF",X"9F",X"DF",X"3F",X"1F",X"03",X"27",X"17",X"07",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"88",X"CC",
		X"00",X"88",X"CC",X"CC",X"CC",X"4C",X"08",X"00",X"FF",X"FF",X"FF",X"FF",X"0F",X"0A",X"0F",X"0A",
		X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"0E",X"0B",X"0E",X"05",X"00",X"11",X"33",X"33",X"33",X"23",X"01",X"00",
		X"20",X"20",X"24",X"0E",X"0E",X"0B",X"07",X"07",X"00",X"00",X"00",X"00",X"03",X"0E",X"0D",X"03",
		X"0D",X"0D",X"0B",X"0A",X"06",X"0C",X"08",X"00",X"0E",X"0E",X"01",X"07",X"0F",X"0E",X"01",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",
		X"08",X"0F",X"00",X"00",X"01",X"0F",X"0E",X"0F",X"07",X"01",X"00",X"00",X"00",X"07",X"03",X"01",
		X"00",X"C0",X"80",X"0E",X"0F",X"2F",X"0F",X"8F",X"60",X"F0",X"B4",X"87",X"87",X"1F",X"0F",X"8F",
		X"0F",X"0E",X"8E",X"0C",X"0C",X"08",X"00",X"00",X"0F",X"2F",X"0F",X"8F",X"2F",X"0F",X"0F",X"0C",
		X"30",X"F0",X"D2",X"3C",X"3C",X"9E",X"0F",X"0F",X"00",X"00",X"30",X"01",X"03",X"07",X"07",X"17",
		X"2F",X"0F",X"4F",X"0F",X"0F",X"07",X"01",X"00",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"00",X"00",X"6E",X"BF",X"DF",X"CF",X"AF",X"6F",
		X"7F",X"7F",X"7F",X"FF",X"EE",X"CC",X"88",X"00",X"FF",X"0F",X"FF",X"6F",X"AF",X"DF",X"BF",X"6E",
		X"00",X"00",X"07",X"5F",X"DF",X"DF",X"DF",X"5F",X"00",X"00",X"00",X"00",X"01",X"13",X"27",X"37",
		X"8F",X"0F",X"8F",X"5F",X"DF",X"DF",X"DF",X"0F",X"7F",X"0F",X"7F",X"37",X"27",X"13",X"01",X"00",
		X"0C",X"0F",X"0C",X"0F",X"0F",X"0F",X"09",X"09",X"00",X"00",X"09",X"09",X"0B",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"EE",X"EE",X"FF",X"FF",X"EE",X"CC",X"88",
		X"04",X"0F",X"0F",X"0F",X"03",X"88",X"EE",X"FF",X"00",X"03",X"03",X"00",X"00",X"11",X"33",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"FF",
		X"80",X"80",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"10",X"B0",X"B0",X"E1",X"86",X"01",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0E",X"0E",X"0C",X"08",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"07",X"0D",X"0E",X"CF",X"8F",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"17",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"17",X"17",X"03",X"03",X"01",X"01",X"00",X"00",
		X"E0",X"C0",X"E0",X"70",X"F0",X"F0",X"10",X"00",X"70",X"90",X"E0",X"F0",X"F0",X"E8",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"EE",X"44",X"44",X"CC",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"77",X"BF",X"FF",X"FF",X"DD",X"00",X"00",X"00",X"00",X"00",X"11",X"23",X"33",
		X"DD",X"BB",X"FF",X"44",X"77",X"EE",X"EE",X"88",X"11",X"77",X"BF",X"FF",X"66",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"CC",X"CC",X"44",X"66",X"EE",X"FF",
		X"66",X"AA",X"AA",X"FF",X"FF",X"33",X"FF",X"EE",X"FF",X"FF",X"BB",X"DD",X"EE",X"77",X"DD",X"FF",
		X"88",X"FF",X"FF",X"EE",X"FF",X"FF",X"77",X"DD",X"33",X"33",X"66",X"CC",X"DD",X"DD",X"CC",X"77",
		X"EE",X"66",X"55",X"55",X"44",X"66",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"0C",X"07",X"00",X"F0",X"F0",X"F0",X"F8",X"FC",X"0F",X"0E",X"0C",
		X"00",X"00",X"10",X"70",X"F0",X"F0",X"F0",X"F1",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"F2",X"F2",X"F3",X"F1",X"F1",X"0F",X"00",X"03",X"30",X"30",X"30",X"10",X"00",X"01",X"00",X"00",
		X"01",X"02",X"0C",X"0C",X"0C",X"84",X"84",X"80",X"00",X"00",X"01",X"0F",X"01",X"07",X"30",X"70",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"73",X"F3",X"F0",X"F8",X"E8",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"71",X"F1",X"FC",X"FC",X"E0",X"00",X"00",X"00",X"00",X"10",X"F0",X"30",X"10",
		X"00",X"88",X"CC",X"EE",X"EE",X"2E",X"0F",X"8D",X"22",X"77",X"FF",X"FF",X"FF",X"AF",X"0F",X"0F",
		X"8D",X"0D",X"8D",X"0D",X"0F",X"0C",X"0C",X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"22",X"33",X"77",X"FF",X"FF",X"DF",X"DF",X"CF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"8F",X"8F",X"8F",X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"02",X"0C",X"0E",X"C3",X"E5",X"C3",X"0E",X"0F",
		X"78",X"68",X"68",X"68",X"C0",X"00",X"00",X"00",X"EF",X"CF",X"0F",X"EF",X"EF",X"0E",X"01",X"01",
		X"08",X"07",X"1E",X"78",X"F4",X"78",X"1F",X"0F",X"00",X"00",X"00",X"01",X"01",X"01",X"08",X"09",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"07",X"13",X"13",X"13",X"01",X"00",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"88",X"FF",X"11",X"11",X"33",X"EE",X"EE",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"77",
		X"FF",X"88",X"FF",X"77",X"70",X"FF",X"FF",X"F8",X"FF",X"11",X"FF",X"EE",X"E0",X"FF",X"FF",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"00",
		X"F3",X"F3",X"FF",X"FE",X"FE",X"FF",X"FE",X"FF",X"FC",X"FC",X"F9",X"F7",X"F7",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"02",X"04",X"08",X"0E",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"0C",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"00",X"00",X"00",X"00",
		X"0A",X"02",X"02",X"09",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"01",X"00",X"04",X"03",X"00",X"00",X"00",X"00",
		X"02",X"0A",X"0A",X"01",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",
		X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"07",X"00",X"00",X"00",X"00",
		X"02",X"0A",X"0A",X"01",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"0F",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"02",X"01",X"09",X"06",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"0E",X"01",X"01",X"0E",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"00",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"01",X"07",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"11",X"00",X"01",
		X"EF",X"EF",X"CF",X"AF",X"EF",X"CF",X"08",X"00",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"08",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"00",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"06",X"00",X"11",X"33",X"33",X"33",X"11",X"00",X"00",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",X"05",X"05",X"0E",X"0E",X"0E",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"03",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"0C",X"0E",X"E1",X"F2",X"F0",X"0F",X"0E",
		X"00",X"88",X"CC",X"CC",X"CC",X"88",X"00",X"08",X"08",X"0E",X"0F",X"07",X"03",X"00",X"00",X"00",
		X"07",X"07",X"07",X"0F",X"0F",X"0F",X"01",X"02",X"7F",X"7F",X"3F",X"5F",X"7F",X"3F",X"01",X"00",
		X"00",X"00",X"00",X"00",X"08",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"03",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"0C",X"0E",X"E1",X"F2",X"F0",X"0F",X"0E",
		X"00",X"88",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"06",
		X"07",X"07",X"07",X"0F",X"0F",X"07",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"0A",X"0A",
		X"00",X"00",X"00",X"00",X"06",X"06",X"04",X"0C",X"00",X"00",X"00",X"01",X"01",X"04",X"0E",X"06",
		X"08",X"07",X"0F",X"0F",X"0F",X"1F",X"27",X"2F",X"02",X"0C",X"0E",X"0F",X"0F",X"0E",X"8C",X"8E",
		X"0C",X"08",X"00",X"00",X"06",X"0C",X"08",X"00",X"03",X"01",X"01",X"01",X"00",X"00",X"01",X"03",
		X"4F",X"8F",X"8F",X"8F",X"5F",X"0F",X"08",X"00",X"4F",X"4F",X"8F",X"8F",X"0E",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0C",X"00",X"00",X"00",X"01",X"05",X"0C",X"0C",X"06",
		X"08",X"07",X"0F",X"0F",X"0F",X"1F",X"27",X"2F",X"02",X"0C",X"0E",X"0F",X"0F",X"0E",X"8C",X"4F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"07",X"03",X"01",X"01",X"0C",X"07",X"07",X"00",
		X"2F",X"2F",X"4F",X"4F",X"2F",X"0F",X"00",X"00",X"4F",X"2F",X"2F",X"4E",X"8E",X"0F",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"01",X"01",X"01",X"08",X"09",
		X"08",X"07",X"1E",X"78",X"F4",X"78",X"1F",X"0F",X"02",X"0C",X"0E",X"C3",X"E5",X"C3",X"0E",X"0F",
		X"68",X"68",X"68",X"68",X"C0",X"00",X"00",X"00",X"07",X"13",X"13",X"13",X"01",X"00",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"EF",X"CF",X"0F",X"EF",X"EF",X"0E",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"06",X"00",X"00",X"00",X"01",X"01",X"04",X"0C",X"0D",
		X"08",X"07",X"0F",X"0F",X"0F",X"1F",X"27",X"2F",X"02",X"0C",X"0E",X"0F",X"0F",X"0E",X"8C",X"8F",
		X"0C",X"08",X"08",X"08",X"00",X"00",X"00",X"08",X"07",X"03",X"03",X"03",X"01",X"00",X"01",X"03",
		X"4F",X"8F",X"8F",X"8F",X"5F",X"0F",X"08",X"00",X"4F",X"4F",X"8F",X"8F",X"0F",X"0E",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"02",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"01",X"07",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"01",X"11",X"33",X"33",X"33",X"11",X"00",X"00",
		X"EF",X"6F",X"8F",X"EF",X"EF",X"CF",X"04",X"03",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"04",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"00",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"06",X"00",X"11",X"33",X"07",X"33",X"11",X"00",X"03",
		X"EF",X"8F",X"6F",X"EF",X"EF",X"CF",X"04",X"09",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"04",X"08",
		X"00",X"08",X"0C",X"0F",X"86",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"77",
		X"00",X"11",X"09",X"05",X"8F",X"BF",X"DF",X"EF",X"00",X"0F",X"E5",X"F0",X"78",X"0F",X"0F",X"0F",
		X"00",X"00",X"06",X"0E",X"0C",X"0C",X"08",X"00",X"77",X"33",X"03",X"02",X"02",X"00",X"00",X"00",
		X"CF",X"8F",X"0F",X"07",X"0F",X"09",X"08",X"00",X"0E",X"0E",X"0C",X"0D",X"0F",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"00",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"06",X"00",X"11",X"33",X"33",X"33",X"11",X"00",X"00",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",X"05",X"05",X"0E",X"0E",X"0E",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0E",X"0C",X"01",X"01",X"03",X"07",X"16",X"34",X"36",X"34",
		X"00",X"0E",X"0F",X"87",X"87",X"87",X"87",X"0F",X"00",X"03",X"03",X"01",X"01",X"0C",X"0E",X"0F",
		X"0C",X"08",X"08",X"0E",X"00",X"08",X"00",X"00",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6F",X"EF",X"DF",X"BF",X"FF",X"77",X"33",X"00",X"0F",X"0F",X"8F",X"CE",X"CE",X"CF",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"02",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"01",X"07",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"01",X"11",X"33",X"33",X"33",X"11",X"00",X"00",
		X"EF",X"6F",X"8F",X"EF",X"EF",X"CF",X"04",X"03",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"04",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"00",X"00",
		X"00",X"03",X"07",X"78",X"F4",X"F0",X"0F",X"07",X"02",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"06",X"00",X"11",X"33",X"07",X"33",X"11",X"00",X"03",
		X"EF",X"8F",X"6F",X"EF",X"EF",X"CF",X"04",X"09",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"04",X"08",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"67",X"57",X"33",X"00",X"00",X"00",X"00",X"EE",X"BF",X"5F",X"EE",X"00",
		X"00",X"00",X"88",X"4C",X"4C",X"88",X"00",X"00",X"00",X"00",X"11",X"11",X"04",X"00",X"00",X"00",
		X"77",X"AF",X"2F",X"5F",X"8F",X"DF",X"33",X"00",X"EE",X"5F",X"2F",X"2F",X"EF",X"1F",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"67",X"57",X"33",X"00",X"00",X"00",X"00",X"EE",X"BF",X"5F",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"88",X"4C",X"4C",X"88",X"00",X"00",X"00",X"00",X"11",X"11",X"04",X"00",X"00",X"00",
		X"77",X"AF",X"2F",X"5F",X"8F",X"DF",X"33",X"00",X"EE",X"5F",X"2F",X"2F",X"EF",X"1F",X"CC",X"00",
		X"00",X"00",X"00",X"02",X"0C",X"03",X"84",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"76",
		X"00",X"00",X"02",X"05",X"0A",X"0F",X"CF",X"EF",X"00",X"00",X"08",X"04",X"08",X"03",X"0F",X"4B",
		X"0C",X"87",X"0C",X"0F",X"84",X"8A",X"89",X"00",X"FF",X"77",X"11",X"00",X"00",X"00",X"11",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"88",X"00",X"2D",X"8F",X"ED",X"CF",X"FF",X"33",X"11",X"00",
		X"00",X"00",X"02",X"04",X"08",X"03",X"0C",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"76",
		X"00",X"00",X"05",X"05",X"0A",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"04",X"08",X"03",X"0F",X"CB",
		X"0F",X"84",X"0F",X"0C",X"0A",X"89",X"CC",X"00",X"FF",X"77",X"11",X"00",X"11",X"11",X"33",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"00",X"00",X"ED",X"CF",X"ED",X"FF",X"FF",X"33",X"00",X"00",
		X"CC",X"CC",X"0E",X"00",X"00",X"06",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"02",X"05",
		X"02",X"02",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"01",X"03",
		X"00",X"01",X"07",X"0F",X"3C",X"E0",X"00",X"00",X"06",X"0C",X"08",X"87",X"01",X"02",X"04",X"06",
		X"0E",X"08",X"66",X"6E",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"00",X"03",X"03",X"0E",X"0A",X"02",X"0A",X"07",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"01",X"07",X"0F",X"02",X"06",
		X"00",X"01",X"07",X"0F",X"3C",X"E0",X"00",X"00",X"04",X"08",X"08",X"87",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"02",X"07",X"0E",X"0E",X"08",X"00",X"00",X"00",X"00",X"0C",X"0E",X"06",X"01",
		X"00",X"00",X"00",X"00",X"60",X"02",X"02",X"07",X"00",X"00",X"00",X"00",X"60",X"04",X"04",X"0E",
		X"00",X"0C",X"00",X"0C",X"00",X"08",X"04",X"08",X"00",X"07",X"08",X"03",X"04",X"09",X"02",X"04",
		X"2F",X"1F",X"1F",X"1F",X"2F",X"03",X"00",X"00",X"4F",X"8F",X"8F",X"8F",X"4F",X"0C",X"00",X"00",
		X"00",X"02",X"06",X"0C",X"09",X"0B",X"0E",X"08",X"00",X"00",X"08",X"04",X"02",X"0E",X"06",X"01",
		X"00",X"00",X"00",X"00",X"60",X"02",X"02",X"07",X"00",X"00",X"00",X"00",X"60",X"04",X"04",X"0E",
		X"00",X"0E",X"01",X"0C",X"02",X"09",X"04",X"02",X"00",X"03",X"00",X"03",X"00",X"01",X"02",X"01",
		X"2F",X"1F",X"1F",X"1F",X"2F",X"03",X"00",X"00",X"4F",X"8F",X"8F",X"8F",X"4F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"0C",X"03",X"11",
		X"00",X"FF",X"FF",X"FF",X"F9",X"FD",X"FF",X"FF",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",
		X"00",X"00",X"00",X"88",X"BB",X"CC",X"CC",X"00",X"33",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"CC",X"00",X"CC",X"00",X"00",X"99",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"03",X"1D",
		X"00",X"FF",X"FF",X"FF",X"F9",X"FD",X"FF",X"FF",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",
		X"00",X"00",X"00",X"22",X"AA",X"CC",X"00",X"00",X"33",X"11",X"00",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"66",X"EE",X"FF",X"FF",X"33",X"00",X"CC",X"00",X"00",X"66",X"FF",X"FF",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"71",X"31",X"10",X"00",
		X"00",X"80",X"D0",X"D0",X"FD",X"F5",X"D2",X"0F",X"00",X"C0",X"E0",X"F0",X"FC",X"E4",X"C1",X"0E",
		X"00",X"00",X"20",X"42",X"42",X"48",X"08",X"00",X"03",X"00",X"01",X"02",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"F0",X"07",X"70",X"07",X"30",X"00",X"8F",X"0C",X"E0",X"0C",X"C2",X"1E",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"30",X"70",X"71",X"31",X"14",X"03",
		X"00",X"80",X"D0",X"D0",X"FD",X"F5",X"D2",X"0F",X"00",X"C0",X"E0",X"F0",X"FC",X"E4",X"C0",X"0F",
		X"00",X"08",X"00",X"00",X"48",X"4A",X"08",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"07",X"70",X"07",X"70",X"03",X"00",X"8E",X"0D",X"0E",X"C0",X"0E",X"D2",X"18",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
