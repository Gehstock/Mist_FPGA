LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
PACKAGE rom_pack IS

  TYPE arr8  IS ARRAY(natural RANGE<>) OF unsigned(7 DOWNTO 0);

  CONSTANT INIT_SL31253 : arr8 := (
    x"70",x"0B",x"70",x"5C",x"0A",x"1F",x"25",x"40",x"94",x"F8",x"67",x"6B",x"20",x"28",x"5C",x"2A",
    x"08",x"00",x"16",x"25",x"55",x"94",x"04",x"29",x"08",x"02",x"20",x"D6",x"53",x"28",x"00",x"D0",
    x"20",x"4A",x"50",x"28",x"00",x"99",x"63",x"6C",x"74",x"5C",x"44",x"6F",x"5C",x"25",x"03",x"91",
    x"F0",x"28",x"01",x"35",x"28",x"02",x"24",x"28",x"00",x"88",x"28",x"02",x"DA",x"28",x"00",x"88",
    x"28",x"02",x"E8",x"28",x"00",x"88",x"21",x"04",x"84",x"07",x"28",x"03",x"8C",x"28",x"03",x"99",
    x"28",x"06",x"58",x"28",x"04",x"67",x"28",x"03",x"D3",x"63",x"6F",x"4C",x"25",x"02",x"94",x"04",
    x"28",x"04",x"47",x"64",x"6F",x"4C",x"1F",x"5C",x"70",x"B0",x"A0",x"21",x"04",x"94",x"04",x"28",
    x"02",x"24",x"63",x"6C",x"2A",x"00",x"83",x"4C",x"12",x"8E",x"16",x"55",x"28",x"00",x"8F",x"70",
    x"B5",x"90",x"B5",x"22",x"13",x"07",x"03",x"03",x"64",x"6E",x"4E",x"51",x"4C",x"50",x"1C",x"20",
    x"FF",x"56",x"36",x"94",x"FE",x"35",x"94",x"F8",x"1C",x"08",x"28",x"01",x"07",x"20",x"33",x"51",
    x"20",x"13",x"52",x"28",x"06",x"79",x"20",x"8B",x"50",x"28",x"06",x"79",x"28",x"00",x"C1",x"20",
    x"33",x"51",x"20",x"13",x"52",x"7D",x"50",x"28",x"06",x"79",x"28",x"06",x"79",x"28",x"01",x"1E",
    x"0C",x"A0",x"18",x"21",x"0F",x"84",x"FB",x"54",x"20",x"FF",x"55",x"35",x"94",x"FE",x"90",x"C0",
    x"08",x"28",x"01",x"07",x"70",x"52",x"20",x"7E",x"51",x"43",x"22",x"10",x"50",x"28",x"06",x"79",
    x"75",x"51",x"7D",x"50",x"28",x"06",x"79",x"31",x"41",x"25",x"70",x"81",x"F6",x"42",x"24",x"05",
    x"52",x"63",x"6F",x"73",x"FC",x"84",x"08",x"42",x"25",x"30",x"81",x"DB",x"70",x"53",x"42",x"25",
    x"40",x"81",x"D4",x"28",x"01",x"1E",x"0C",x"0A",x"57",x"67",x"6B",x"4C",x"0B",x"00",x"5C",x"0A",
    x"1F",x"0B",x"01",x"5C",x"0A",x"1F",x"0B",x"0A",x"67",x"6B",x"5C",x"47",x"0B",x"1C",x"0A",x"57",
    x"67",x"6B",x"4C",x"24",x"FF",x"0B",x"4C",x"05",x"0A",x"24",x"FF",x"0B",x"4C",x"04",x"0A",x"67",
    x"6B",x"5C",x"47",x"0B",x"1C",x"08",x"28",x"01",x"07",x"63",x"6F",x"4C",x"64",x"6D",x"25",x"01",
    x"84",x"0E",x"20",x"53",x"5D",x"7C",x"5E",x"20",x"D0",x"53",x"28",x"00",x"D0",x"90",x"2F",x"20",
    x"17",x"5D",x"20",x"FF",x"5C",x"20",x"D6",x"53",x"28",x"00",x"D0",x"20",x"11",x"51",x"78",x"52",
    x"28",x"01",x"F6",x"20",x"11",x"51",x"20",x"25",x"52",x"28",x"01",x"F6",x"20",x"5C",x"51",x"78",
    x"52",x"28",x"01",x"F6",x"20",x"5C",x"51",x"20",x"25",x"52",x"28",x"01",x"F6",x"20",x"14",x"51",
    x"76",x"52",x"28",x"02",x"0E",x"20",x"14",x"51",x"20",x"2E",x"52",x"28",x"02",x"0E",x"20",x"99",
    x"62",x"6E",x"5D",x"5C",x"28",x"02",x"AC",x"28",x"02",x"B5",x"64",x"6A",x"72",x"5C",x"90",x"05",
    x"08",x"28",x"01",x"07",x"62",x"68",x"20",x"17",x"5C",x"6B",x"5C",x"20",x"1C",x"51",x"20",x"1A",
    x"52",x"20",x"B0",x"50",x"28",x"06",x"79",x"20",x"38",x"51",x"20",x"1B",x"52",x"20",x"55",x"50",
    x"28",x"06",x"79",x"20",x"52",x"51",x"20",x"1A",x"52",x"20",x"71",x"50",x"28",x"06",x"79",x"64",
    x"6D",x"4C",x"13",x"81",x"06",x"28",x"04",x"47",x"90",x"19",x"20",x"11",x"51",x"20",x"1A",x"52",
    x"20",x"B2",x"50",x"28",x"06",x"79",x"20",x"5E",x"51",x"20",x"1A",x"52",x"20",x"73",x"50",x"28",
    x"06",x"79",x"28",x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",x"78",x"53",x"20",x"81",x"50",x"28",
    x"06",x"79",x"41",x"24",x"FA",x"51",x"42",x"1F",x"52",x"33",x"94",x"F1",x"90",x"E5",x"08",x"28",
    x"01",x"07",x"20",x"46",x"53",x"20",x"92",x"50",x"28",x"06",x"79",x"41",x"24",x"FB",x"51",x"33",
    x"94",x"F4",x"90",x"CF",x"08",x"28",x"01",x"07",x"20",x"85",x"50",x"28",x"00",x"99",x"44",x"25",
    x"08",x"94",x"05",x"28",x"01",x"1E",x"0C",x"25",x"02",x"94",x"0D",x"20",x"8E",x"50",x"28",x"00",
    x"99",x"63",x"6C",x"44",x"5C",x"90",x"E2",x"25",x"01",x"94",x"DE",x"20",x"8C",x"50",x"28",x"00",
    x"99",x"2A",x"02",x"6C",x"44",x"12",x"8E",x"16",x"67",x"69",x"5D",x"70",x"5C",x"66",x"6F",x"7F",
    x"5C",x"28",x"02",x"71",x"64",x"6D",x"4C",x"22",x"20",x"5C",x"90",x"BD",x"02",x"05",x"10",x"10",
    x"20",x"08",x"28",x"01",x"07",x"67",x"6A",x"4E",x"54",x"4C",x"53",x"14",x"22",x"80",x"50",x"20",
    x"2A",x"51",x"20",x"33",x"52",x"28",x"06",x"79",x"43",x"21",x"0F",x"22",x"80",x"50",x"28",x"06",
    x"79",x"20",x"91",x"50",x"28",x"06",x"79",x"44",x"14",x"22",x"80",x"50",x"28",x"06",x"79",x"44",
    x"21",x"0F",x"22",x"80",x"50",x"28",x"06",x"79",x"28",x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",
    x"6E",x"20",x"17",x"90",x"08",x"08",x"28",x"01",x"07",x"6F",x"20",x"50",x"62",x"51",x"20",x"33",
    x"52",x"71",x"24",x"66",x"DC",x"5C",x"14",x"22",x"40",x"50",x"28",x"06",x"79",x"4C",x"21",x"0F",
    x"22",x"40",x"50",x"28",x"06",x"79",x"28",x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",x"20",x"B0",
    x"54",x"62",x"69",x"70",x"B4",x"A4",x"90",x"0D",x"08",x"28",x"01",x"07",x"20",x"71",x"54",x"62",
    x"6C",x"70",x"B1",x"A1",x"18",x"F1",x"50",x"4D",x"51",x"4C",x"52",x"71",x"F0",x"84",x"05",x"41",
    x"24",x"02",x"51",x"72",x"F0",x"84",x"05",x"41",x"24",x"FE",x"51",x"74",x"F0",x"84",x"05",x"42",
    x"24",x"02",x"52",x"78",x"F0",x"84",x"05",x"42",x"24",x"FE",x"52",x"63",x"6F",x"4C",x"25",x"02",
    x"91",x"36",x"94",x"17",x"71",x"F4",x"94",x"0B",x"41",x"25",x"2D",x"81",x"04",x"20",x"2D",x"51",
    x"90",x"09",x"41",x"25",x"3D",x"91",x"04",x"20",x"3D",x"51",x"41",x"25",x"52",x"81",x"04",x"20",
    x"52",x"51",x"25",x"1A",x"91",x"04",x"20",x"1A",x"51",x"42",x"25",x"2B",x"81",x"04",x"20",x"2B",
    x"52",x"25",x"09",x"91",x"03",x"79",x"52",x"64",x"6F",x"4C",x"21",x"03",x"25",x"03",x"94",x"24",
    x"62",x"68",x"71",x"F4",x"84",x"02",x"6B",x"20",x"10",x"F0",x"84",x"02",x"3C",x"20",x"20",x"F0",
    x"84",x"04",x"4C",x"1F",x"5C",x"4C",x"25",x"16",x"94",x"03",x"20",x"1D",x"25",x"1E",x"94",x"03",
    x"20",x"17",x"5C",x"44",x"50",x"28",x"06",x"79",x"28",x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",
    x"68",x"20",x"B2",x"53",x"70",x"B4",x"A4",x"90",x"0C",x"08",x"28",x"01",x"07",x"6A",x"20",x"73",
    x"53",x"70",x"B1",x"A1",x"18",x"50",x"63",x"4D",x"51",x"4C",x"52",x"40",x"21",x"80",x"84",x"05",
    x"42",x"24",x"02",x"52",x"40",x"21",x"40",x"84",x"03",x"32",x"32",x"42",x"25",x"14",x"91",x"04",
    x"20",x"14",x"52",x"25",x"20",x"81",x"04",x"20",x"20",x"52",x"43",x"50",x"28",x"06",x"79",x"28",
    x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",x"64",x"68",x"4D",x"51",x"4D",x"52",x"4D",x"53",x"4D",
    x"54",x"4C",x"25",x"00",x"84",x"0D",x"70",x"5C",x"43",x"13",x"C3",x"C3",x"53",x"44",x"13",x"C4",
    x"C4",x"54",x"41",x"C3",x"51",x"42",x"C4",x"52",x"64",x"6D",x"20",x"44",x"FC",x"84",x"3D",x"28");

  CONSTANT INIT_SL31254 : arr8 := (
    x"04",x"9C",x"64",x"6A",x"41",x"50",x"25",x"5C",x"81",x"07",x"28",x"04",x"3F",x"20",x"5C",x"51",
    x"41",x"50",x"25",x"14",x"91",x"07",x"28",x"04",x"3F",x"20",x"14",x"51",x"6B",x"42",x"50",x"25",
    x"08",x"91",x"07",x"28",x"04",x"3F",x"20",x"09",x"52",x"42",x"50",x"25",x"2E",x"81",x"07",x"28",
    x"04",x"3F",x"20",x"2E",x"52",x"20",x"55",x"50",x"28",x"06",x"79",x"28",x"01",x"1E",x"0C",x"4C",
    x"18",x"1F",x"5C",x"20",x"40",x"B5",x"1C",x"08",x"28",x"01",x"07",x"20",x"36",x"51",x"7A",x"52",
    x"75",x"54",x"20",x"81",x"50",x"28",x"06",x"79",x"41",x"24",x"FA",x"51",x"42",x"24",x"08",x"52",
    x"34",x"94",x"F0",x"28",x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",x"67",x"68",x"4C",x"22",x"00",
    x"84",x"27",x"70",x"5C",x"6A",x"71",x"50",x"18",x"DC",x"24",x"66",x"D0",x"5C",x"25",x"99",x"94",
    x"15",x"20",x"59",x"5E",x"71",x"50",x"18",x"DC",x"24",x"66",x"D0",x"25",x"99",x"94",x"06",x"28",
    x"02",x"24",x"90",x"05",x"5C",x"28",x"02",x"71",x"28",x"01",x"1E",x"0C",x"08",x"28",x"01",x"07",
    x"64",x"6F",x"71",x"FC",x"84",x"13",x"62",x"6C",x"28",x"05",x"FC",x"30",x"84",x"3B",x"62",x"69",
    x"28",x"05",x"FC",x"30",x"84",x"30",x"90",x"11",x"62",x"69",x"28",x"05",x"FC",x"30",x"84",x"26",
    x"62",x"6C",x"28",x"05",x"FC",x"30",x"84",x"21",x"64",x"6D",x"4C",x"21",x"04",x"94",x"04",x"29",
    x"05",x"9D",x"63",x"68",x"28",x"05",x"FC",x"30",x"84",x"7C",x"63",x"6A",x"28",x"05",x"FC",x"30",
    x"84",x"78",x"29",x"05",x"88",x"68",x"90",x"02",x"6B",x"62",x"4D",x"54",x"4D",x"4C",x"57",x"64",
    x"6D",x"4C",x"13",x"44",x"81",x"21",x"2A",x"05",x"0E",x"77",x"54",x"37",x"37",x"44",x"C7",x"53",
    x"42",x"18",x"1F",x"C3",x"84",x"04",x"34",x"81",x"F5",x"44",x"8E",x"16",x"90",x"0B",x"04",x"04",
    x"05",x"06",x"00",x"01",x"02",x"03",x"24",x"E9",x"2A",x"05",x"47",x"13",x"8E",x"16",x"55",x"16",
    x"56",x"64",x"6A",x"4C",x"22",x"00",x"91",x"13",x"45",x"18",x"1F",x"55",x"6D",x"4C",x"13",x"6A",
    x"91",x"05",x"46",x"18",x"1F",x"56",x"41",x"24",x"02",x"51",x"45",x"5D",x"46",x"5D",x"72",x"5C",
    x"20",x"80",x"B5",x"28",x"01",x"1E",x"0C",x"02",x"00",x"02",x"01",x"02",x"02",x"01",x"02",x"01",
    x"FE",x"02",x"FE",x"02",x"FF",x"71",x"53",x"90",x"03",x"72",x"53",x"64",x"6A",x"4C",x"33",x"84",
    x"07",x"22",x"00",x"81",x"07",x"90",x"08",x"22",x"00",x"81",x"04",x"18",x"1F",x"5C",x"20",x"80",
    x"B5",x"6B",x"4C",x"22",x"00",x"94",x"10",x"62",x"69",x"4C",x"21",x"01",x"84",x"04",x"72",x"90",
    x"03",x"20",x"FE",x"64",x"6B",x"5C",x"90",x"6C",x"42",x"25",x"14",x"81",x"0E",x"25",x"24",x"91",
    x"0A",x"41",x"25",x"14",x"81",x"14",x"25",x"5C",x"91",x"10",x"29",x"05",x"43",x"41",x"25",x"14",
    x"81",x"08",x"25",x"5C",x"91",x"04",x"29",x"05",x"43",x"64",x"6A",x"4D",x"13",x"91",x"05",x"24",
    x"02",x"90",x"03",x"24",x"FE",x"C1",x"51",x"6B",x"4C",x"C2",x"52",x"20",x"55",x"50",x"28",x"06",
    x"79",x"64",x"6B",x"70",x"5C",x"64",x"68",x"4C",x"25",x"30",x"91",x"06",x"28",x"02",x"B5",x"90",
    x"04",x"28",x"02",x"AC",x"20",x"FF",x"55",x"28",x"00",x"8F",x"63",x"6F",x"4C",x"25",x"02",x"94",
    x"10",x"62",x"6E",x"4D",x"25",x"15",x"84",x"06",x"4C",x"25",x"15",x"94",x"04",x"28",x"02",x"24",
    x"28",x"01",x"A0",x"28",x"01",x"1E",x"28",x"01",x"1E",x"29",x"00",x"37",x"08",x"28",x"01",x"07",
    x"4C",x"18",x"1F",x"C1",x"91",x"0B",x"4C",x"24",x"05",x"56",x"41",x"18",x"1F",x"CC",x"81",x"17",
    x"4C",x"18",x"1F",x"56",x"41",x"24",x"02",x"C6",x"91",x"36",x"41",x"24",x"02",x"18",x"1F",x"56",
    x"4C",x"24",x"05",x"C6",x"91",x"2A",x"4D",x"4C",x"18",x"1F",x"56",x"42",x"C6",x"91",x"0B",x"42",
    x"18",x"1F",x"56",x"4C",x"24",x"05",x"C6",x"81",x"1D",x"4C",x"18",x"1F",x"56",x"42",x"24",x"02",
    x"C6",x"91",x"0D",x"42",x"24",x"02",x"18",x"1F",x"56",x"4C",x"24",x"05",x"C6",x"81",x"07",x"70",
    x"50",x"28",x"01",x"1E",x"0C",x"71",x"90",x"F9",x"2A",x"06",x"74",x"64",x"6D",x"4C",x"21",x"20",
    x"84",x"12",x"66",x"6F",x"3C",x"94",x"0D",x"63",x"6C",x"4C",x"12",x"8E",x"16",x"66",x"6F",x"5D",
    x"67",x"71",x"5C",x"1C",x"09",x"0D",x"15",x"1C",x"1C",x"2A",x"07",x"67",x"08",x"28",x"01",x"07",
    x"0A",x"66",x"6C",x"5D",x"43",x"5D",x"44",x"5C",x"75",x"54",x"20",x"C0",x"F0",x"53",x"20",x"3F",
    x"F0",x"50",x"25",x"15",x"94",x"1F",x"64",x"68",x"72",x"54",x"28",x"06",x"EC",x"20",x"15",x"50",
    x"28",x"07",x"18",x"41",x"24",x"06",x"51",x"66",x"6D",x"4D",x"53",x"4C",x"54",x"6C",x"4C",x"0B",
    x"28",x"01",x"1E",x"0C",x"25",x"30",x"94",x"0B",x"62",x"69",x"28",x"06",x"EC",x"68",x"4D",x"50",
    x"90",x"DF",x"25",x"31",x"94",x"0B",x"62",x"6C",x"28",x"06",x"EC",x"6B",x"4D",x"50",x"90",x"D1",
    x"25",x"32",x"94",x"0B",x"63",x"68",x"28",x"06",x"EC",x"20",x"14",x"50",x"90",x"C3",x"25",x"33",
    x"94",x"BF",x"63",x"6A",x"28",x"06",x"EC",x"20",x"14",x"50",x"90",x"B5",x"08",x"28",x"01",x"07",
    x"4C",x"E1",x"94",x"06",x"4D",x"4E",x"E2",x"84",x"1C",x"41",x"55",x"42",x"56",x"4C",x"51",x"45",
    x"5D",x"4C",x"52",x"46",x"5E",x"7D",x"50",x"2A",x"07",x"67",x"28",x"07",x"18",x"2A",x"07",x"67",
    x"4D",x"51",x"4E",x"52",x"28",x"01",x"1E",x"0C",x"40",x"13",x"8E",x"C0",x"8E",x"20",x"40",x"B0",
    x"44",x"56",x"55",x"16",x"57",x"42",x"24",x"00",x"18",x"21",x"3F",x"58",x"A5",x"21",x"C0",x"C8",
    x"B5",x"41",x"24",x"FC",x"18",x"B4",x"47",x"22",x"00",x"43",x"91",x"02",x"70",x"18",x"B1",x"47",
    x"13",x"57",x"20",x"60",x"B0",x"20",x"50",x"B0",x"41",x"1F",x"51",x"74",x"58",x"38",x"94",x"FE",
    x"35",x"94",x"DF",x"42",x"1F",x"52",x"44",x"18",x"1F",x"C1",x"51",x"44",x"36",x"94",x"C4",x"44",
    x"18",x"1F",x"C2",x"52",x"70",x"B0",x"1C",x"F8",x"88",x"88",x"88",x"F8",x"20",x"20",x"20",x"20",
    x"20",x"F8",x"08",x"F8",x"80",x"F8",x"F8",x"08",x"F8",x"08",x"F8",x"88",x"88",x"F8",x"08",x"08",
    x"F8",x"80",x"F8",x"08",x"F8",x"F8",x"80",x"F8",x"88",x"F8",x"F8",x"08",x"10",x"10",x"10",x"F8",
    x"88",x"F8",x"88",x"F8",x"F8",x"88",x"F8",x"08",x"F8",x"F8",x"80",x"98",x"88",x"F8",x"F8",x"08",
    x"38",x"00",x"20",x"F8",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"F8",x"A8",x"A8",
    x"A8",x"A8",x"88",x"50",x"20",x"50",x"88",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"20",x"00",x"20",
    x"00",x"00",x"00",x"F8",x"00",x"00",x"50",x"50",x"50",x"50",x"50",x"A0",x"A0",x"A0",x"A0",x"A0",
    x"C0",x"C0",x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"20",x"20",x"20",x"20",x"20",x"10",
    x"10",x"20",x"40",x"40",x"08",x"10",x"20",x"40",x"80",x"00",x"18",x"20",x"C0",x"00",x"00",x"C0",
    x"20",x"18",x"00",x"80",x"40",x"20",x"10",x"08",x"40",x"40",x"20",x"10",x"10",x"00",x"00",x"00");

END PACKAGE; 