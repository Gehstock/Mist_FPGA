library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity monitor is
    generic(
        AddrWidth   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end monitor;

architecture rtl of monitor is
    type rom8192x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"31",  x"c0",  x"eb",  x"21",  x"54",  x"00",  x"11",  x"00", -- 0000
         x"80",  x"cd",  x"0f",  x"00",  x"c3",  x"10",  x"80",  x"3e", -- 0008
         x"80",  x"ed",  x"a0",  x"cd",  x"4e",  x"00",  x"30",  x"f9", -- 0010
         x"d5",  x"01",  x"00",  x"00",  x"50",  x"14",  x"cd",  x"4e", -- 0018
         x"00",  x"30",  x"fa",  x"d4",  x"4e",  x"00",  x"cb",  x"11", -- 0020
         x"cb",  x"10",  x"38",  x"1f",  x"15",  x"20",  x"f4",  x"03", -- 0028
         x"5e",  x"23",  x"cb",  x"33",  x"30",  x"0c",  x"16",  x"10", -- 0030
         x"cd",  x"4e",  x"00",  x"cb",  x"12",  x"30",  x"f9",  x"14", -- 0038
         x"cb",  x"3a",  x"cb",  x"1b",  x"e3",  x"e5",  x"ed",  x"52", -- 0040
         x"d1",  x"ed",  x"b0",  x"e1",  x"30",  x"c5",  x"87",  x"c0", -- 0048
         x"7e",  x"23",  x"17",  x"c9",  x"c3",  x"04",  x"0c",  x"80", -- 0050
         x"53",  x"44",  x"20",  x"80",  x"00",  x"00",  x"3e",  x"01", -- 0058
         x"d3",  x"02",  x"00",  x"31",  x"00",  x"c0",  x"cd",  x"0d", -- 0060
         x"af",  x"cd",  x"2a",  x"07",  x"87",  x"c3",  x"03",  x"f0", -- 0068
         x"00",  x"00",  x"80",  x"13",  x"02",  x"cf",  x"c9",  x"3e", -- 0070
         x"00",  x"cf",  x"76",  x"03",  x"18",  x"fd",  x"dd",  x"e5", -- 0078
         x"dd",  x"21",  x"0f",  x"00",  x"dd",  x"39",  x"f5",  x"dd", -- 0080
         x"7e",  x"04",  x"dd",  x"77",  x"6c",  x"fe",  x"05",  x"05", -- 0088
         x"05",  x"ff",  x"e1",  x"00",  x"e5",  x"56",  x"23",  x"66", -- 0090
         x"dd",  x"4e",  x"06",  x"06",  x"00",  x"00",  x"7a",  x"a9", -- 0098
         x"5f",  x"7c",  x"a8",  x"57",  x"26",  x"00",  x"00",  x"cb", -- 00A0
         x"7c",  x"28",  x"19",  x"6b",  x"42",  x"cb",  x"00",  x"28", -- 00A8
         x"cb",  x"1d",  x"cb",  x"43",  x"28",  x"0a",  x"7d",  x"00", -- 00B0
         x"ee",  x"01",  x"5f",  x"78",  x"ee",  x"a0",  x"57",  x"18", -- 00B8
         x"03",  x"02",  x"5d",  x"50",  x"24",  x"18",  x"e3",  x"2e", -- 00C0
         x"00",  x"73",  x"23",  x"72",  x"f1",  x"dd",  x"e1",  x"c9", -- 00C8
         x"f5",  x"00",  x"21",  x"04",  x"00",  x"39",  x"4e",  x"23", -- 00D0
         x"46",  x"c5",  x"00",  x"cd",  x"82",  x"a2",  x"f1",  x"55", -- 00D8
         x"7a",  x"b7",  x"20",  x"78",  x"3e",  x"5b",  x"10",  x"e5", -- 00E0
         x"21",  x"0a",  x"96",  x"15",  x"70",  x"07",  x"cd",  x"79", -- 00E8
         x"a3",  x"f1",  x"d6",  x"00",  x"55",  x"1b",  x"7e",  x"00", -- 00F0
         x"fd",  x"21",  x"08",  x"00",  x"fd",  x"39",  x"fd",  x"96", -- 00F8
         x"04",  x"00",  x"20",  x"10",  x"21",  x"01",  x"50",  x"0f", -- 0100
         x"01",  x"28",  x"02",  x"04",  x"16",  x"01",  x"6a",  x"f1", -- 0108
         x"c9",  x"40",  x"9f",  x"60",  x"00",  x"21",  x"26",  x"b2", -- 0110
         x"36",  x"00",  x"2d",  x"21",  x"27",  x"04",  x"2a",  x"6b", -- 0118
         x"04",  x"2b",  x"04",  x"5a",  x"28",  x"04",  x"29",  x"d6", -- 0120
         x"04",  x"15",  x"04",  x"1e",  x"f6",  x"04",  x"2c",  x"6e", -- 0128
         x"c9",  x"02",  x"66",  x"05",  x"e5",  x"c0",  x"83",  x"dd", -- 0130
         x"75",  x"02",  x"fc",  x"7d",  x"b7",  x"c2",  x"64",  x"84", -- 0138
         x"fc",  x"6a",  x"0b",  x"dd",  x"00",  x"74",  x"ff",  x"eb", -- 0140
         x"21",  x"1a",  x"b1",  x"07",  x"d5",  x"01",  x"10",  x"00", -- 0148
         x"c5",  x"1f",  x"61",  x"85",  x"13",  x"21",  x"d8",  x"16", -- 0150
         x"15",  x"01",  x"85",  x"84",  x"a2",  x"19",  x"a7",  x"ac", -- 0158
         x"20",  x"19",  x"46",  x"83",  x"32",  x"dd",  x"5e",  x"37", -- 0160
         x"56",  x"ff",  x"44",  x"36",  x"81",  x"69",  x"36",  x"28", -- 0168
         x"0e",  x"88",  x"ae",  x"fa",  x"d6",  x"81",  x"31",  x"20", -- 0170
         x"07",  x"06",  x"fb",  x"b7",  x"ca",  x"bc",  x"29",  x"3a", -- 0178
         x"23",  x"bc",  x"40",  x"fd",  x"3d",  x"c2",  x"69",  x"82", -- 0180
         x"3a",  x"0b",  x"1b",  x"b1",  x"d6",  x"d3",  x"07",  x"4c", -- 0188
         x"1c",  x"07",  x"1d",  x"94",  x"07",  x"21",  x"96",  x"62", -- 0190
         x"84",  x"40",  x"c1",  x"8b",  x"f1",  x"c0",  x"a7",  x"01", -- 0198
         x"1e",  x"c2",  x"e8",  x"80",  x"b4",  x"d5",  x"16",  x"c2", -- 01A0
         x"06",  x"19",  x"d1",  x"4b",  x"0c",  x"ab",  x"00",  x"63", -- 01A8
         x"f1",  x"16",  x"09",  x"82",  x"20",  x"77",  x"00",  x"1c", -- 01B0
         x"7b",  x"d6",  x"15",  x"08",  x"38",  x"e1",  x"1d",  x"a4", -- 01B8
         x"1c",  x"19",  x"da",  x"0b",  x"35",  x"00",  x"26",  x"0a", -- 01C0
         x"e3",  x"33",  x"cd",  x"ab",  x"8b",  x"33",  x"b1",  x"87", -- 01C8
         x"58",  x"01",  x"87",  x"8b",  x"04",  x"21",  x"13",  x"09", -- 01D0
         x"50",  x"14",  x"09",  x"3a",  x"27",  x"b1",  x"60",  x"47", -- 01D8
         x"2b",  x"3a",  x"26",  x"b1",  x"67",  x"2e",  x"c9",  x"b3", -- 01E0
         x"b4",  x"91",  x"9c",  x"b5",  x"57",  x"88",  x"cd",  x"04", -- 01E8
         x"19",  x"22",  x"c4",  x"9d",  x"21",  x"9d",  x"95",  x"71", -- 01F0
         x"2a",  x"e0",  x"34",  x"07",  x"17",  x"8c",  x"21",  x"ac", -- 01F8
         x"84",  x"49",  x"e3",  x"0e",  x"dc",  x"19",  x"0e",  x"f8", -- 0200
         x"52",  x"c0",  x"32",  x"06",  x"ac",  x"13",  x"1c",  x"21", -- 0208
         x"ba",  x"77",  x"2b",  x"56",  x"1c",  x"60",  x"07",  x"11", -- 0210
         x"28",  x"b1",  x"eb",  x"01",  x"01",  x"73",  x"00",  x"ed", -- 0218
         x"b0",  x"3e",  x"0a",  x"f5",  x"2e",  x"7c",  x"13",  x"7e", -- 0220
         x"00",  x"c6",  x"73",  x"77",  x"23",  x"7e",  x"ce",  x"00", -- 0228
         x"77",  x"50",  x"c3",  x"9c",  x"e1",  x"ad",  x"62",  x"a3", -- 0230
         x"21",  x"44",  x"c8",  x"83",  x"d7",  x"02",  x"d7",  x"00", -- 0238
         x"3e",  x"15",  x"83",  x"4f",  x"37",  x"3e",  x"b2",  x"21", -- 0240
         x"47",  x"52",  x"85",  x"d2",  x"01",  x"c2",  x"7e",  x"02", -- 0248
         x"60",  x"cf",  x"e9",  x"85",  x"83",  x"cf",  x"13",  x"09", -- 0250
         x"7a",  x"c6",  x"09",  x"4f",  x"40",  x"fc",  x"66",  x"d5", -- 0258
         x"48",  x"e5",  x"13",  x"d1",  x"02",  x"14",  x"7a",  x"d6", -- 0260
         x"03",  x"38",  x"e7",  x"70",  x"75",  x"3a",  x"2d",  x"b1", -- 0268
         x"57",  x"cc",  x"56",  x"3a",  x"2c",  x"e4",  x"01",  x"0e", -- 0270
         x"00",  x"7b",  x"b0",  x"32",  x"80",  x"cb",  x"7a",  x"b1", -- 0278
         x"32",  x"c6",  x"80",  x"81",  x"d3",  x"22",  x"81",  x"8e", -- 0280
         x"3a",  x"2f",  x"22",  x"1b",  x"2e",  x"65",  x"1b",  x"28", -- 0288
         x"b4",  x"1b",  x"29",  x"15",  x"31",  x"89",  x"15",  x"30", -- 0290
         x"96",  x"15",  x"2a",  x"15",  x"2b",  x"87",  x"84",  x"8d", -- 0298
         x"21",  x"d0",  x"99",  x"0e",  x"2a",  x"28",  x"ff",  x"4e", -- 02A0
         x"7d",  x"26",  x"28",  x"10",  x"e5",  x"95",  x"0c",  x"67", -- 02A8
         x"8c",  x"03",  x"a9",  x"8d",  x"00",  x"e1",  x"24",  x"7c", -- 02B0
         x"d6",  x"17",  x"38",  x"ef",  x"3e",  x"76",  x"10",  x"1a", -- 02B8
         x"11",  x"3a",  x"e9",  x"69",  x"82",  x"01",  x"b6",  x"20", -- 02C0
         x"12",  x"21",  x"e0",  x"25",  x"59",  x"6d",  x"06",  x"42", -- 02C8
         x"cc",  x"3a",  x"c3",  x"9d",  x"d1",  x"85",  x"e5",  x"b1", -- 02D0
         x"0a",  x"3a",  x"93",  x"02",  x"3d",  x"20",  x"08",  x"21", -- 02D8
         x"f9",  x"84",  x"72",  x"0d",  x"d6",  x"02",  x"89",  x"0e", -- 02E0
         x"00",  x"85",  x"34",  x"0e",  x"ed",  x"93",  x"07",  x"97", -- 02E8
         x"09",  x"64",  x"36",  x"97",  x"03",  x"51",  x"8d",  x"97", -- 02F0
         x"09",  x"92",  x"0e",  x"28",  x"a6",  x"0e",  x"d0",  x"0e", -- 02F8
         x"48",  x"2a",  x"0e",  x"f1",  x"b2",  x"ad",  x"b4",  x"b2", -- 0300
         x"4a",  x"0a",  x"43",  x"dd",  x"68",  x"46",  x"a0",  x"4e", -- 0308
         x"51",  x"ff",  x"fc",  x"81",  x"3c",  x"28",  x"6b",  x"68", -- 0310
         x"61",  x"11",  x"e8",  x"07",  x"a4",  x"21",  x"d0",  x"a9", -- 0318
         x"e5",  x"d5",  x"95",  x"a9",  x"14",  x"c1",  x"aa",  x"92", -- 0320
         x"a2",  x"a6",  x"4e",  x"d0",  x"a6",  x"20",  x"48",  x"db", -- 0328
         x"05",  x"fc",  x"05",  x"42",  x"c7",  x"27",  x"85",  x"26", -- 0330
         x"60",  x"ec",  x"c1",  x"a2",  x"e5",  x"58",  x"c5",  x"ee", -- 0338
         x"4f",  x"09",  x"56",  x"60",  x"09",  x"11",  x"79",  x"1b", -- 0340
         x"47",  x"fa",  x"22",  x"80",  x"89",  x"fa",  x"c1",  x"21", -- 0348
         x"fb",  x"25",  x"80",  x"fb",  x"22",  x"18",  x"8f",  x"7a", -- 0350
         x"16",  x"4f",  x"a7",  x"08",  x"f8",  x"08",  x"10",  x"10", -- 0358
         x"6e",  x"d4",  x"70",  x"f9",  x"8d",  x"e0",  x"c3",  x"4b", -- 0360
         x"43",  x"2d",  x"54",  x"00",  x"41",  x"50",  x"45",  x"20", -- 0368
         x"62",  x"79",  x"20",  x"41",  x"38",  x"46",  x"2e",  x"89", -- 0370
         x"06",  x"42",  x"61",  x"73",  x"69",  x"63",  x"83",  x"e0", -- 0378
         x"0a",  x"4c",  x"61",  x"64",  x"65",  x"c0",  x"02",  x"72", -- 0380
         x"65",  x"73",  x"73",  x"65",  x"3a",  x"c2",  x"15",  x"0a", -- 0388
         x"45",  x"6e",  x"64",  x"24",  x"0d",  x"63",  x"6f",  x"60", -- 0390
         x"70",  x"2d",  x"31",  x"34",  x"2d",  x"31",  x"32",  x"50", -- 0398
         x"38",  x"0d",  x"53",  x"79",  x"73",  x"14",  x"74",  x"65", -- 03A0
         x"6d",  x"32",  x"53",  x"08",  x"74",  x"61",  x"72",  x"74", -- 03A8
         x"a0",  x"33",  x"46",  x"65",  x"68",  x"6c",  x"00",  x"65", -- 03B0
         x"72",  x"21",  x"20",  x"4b",  x"65",  x"69",  x"6e",  x"01", -- 03B8
         x"20",  x"54",  x"61",  x"70",  x"2d",  x"46",  x"69",  x"d3", -- 03C0
         x"0f",  x"df",  x"a4",  x"09",  x"63",  x"e5",  x"06",  x"38", -- 03C8
         x"fb",  x"27",  x"01",  x"6d",  x"89",  x"58",  x"a5",  x"57", -- 03D0
         x"39",  x"4e",  x"0c",  x"d5",  x"e1",  x"21",  x"e4",  x"ff", -- 03D8
         x"39",  x"81",  x"aa",  x"36",  x"ff",  x"53",  x"a4",  x"29", -- 03E0
         x"cf",  x"4a",  x"a8",  x"fc",  x"95",  x"9a",  x"74",  x"fe", -- 03E8
         x"15",  x"fa",  x"9d",  x"c9",  x"fa",  x"c2",  x"fa",  x"29", -- 03F0
         x"80",  x"00",  x"3e",  x"3a",  x"85",  x"5f",  x"3e",  x"b0", -- 03F8
         x"19",  x"8c",  x"57",  x"af",  x"e7",  x"34",  x"0f",  x"c1", -- 0400
         x"db",  x"20",  x"fb",  x"20",  x"fc",  x"1c",  x"cd",  x"05", -- 0408
         x"66",  x"fc",  x"cd",  x"14",  x"d5",  x"95",  x"6c",  x"d1", -- 0410
         x"80",  x"bc",  x"33",  x"86",  x"b8",  x"97",  x"28",  x"b0", -- 0418
         x"d5",  x"c1",  x"4c",  x"d0",  x"a7",  x"f6",  x"4c",  x"7d", -- 0420
         x"d1",  x"e4",  x"54",  x"51",  x"9d",  x"b4",  x"d9",  x"9a", -- 0428
         x"05",  x"fe",  x"95",  x"8a",  x"0a",  x"ba",  x"ae",  x"41", -- 0430
         x"8a",  x"87",  x"a4",  x"dd",  x"69",  x"60",  x"00",  x"c5", -- 0438
         x"af",  x"be",  x"ed",  x"a0",  x"20",  x"fb",  x"c1",  x"a9", -- 0440
         x"09",  x"0a",  x"c1",  x"cc",  x"b8",  x"f3",  x"85",  x"90", -- 0448
         x"fb",  x"fc",  x"55",  x"48",  x"66",  x"fe",  x"30",  x"11", -- 0450
         x"08",  x"65",  x"cb",  x"66",  x"28",  x"10",  x"9b",  x"63", -- 0458
         x"e3",  x"64",  x"f5",  x"c6",  x"ae",  x"f3",  x"98",  x"f2", -- 0460
         x"8b",  x"34",  x"fa",  x"d3",  x"20",  x"0e",  x"da",  x"47", -- 0468
         x"85",  x"d2",  x"22",  x"ff",  x"0d",  x"ed",  x"00",  x"fb", -- 0470
         x"3c",  x"44",  x"49",  x"22",  x"52",  x"3e",  x"41",  x"db", -- 0478
         x"ea",  x"41",  x"db",  x"40",  x"91",  x"01",  x"29",  x"9b", -- 0480
         x"b1",  x"65",  x"27",  x"41",  x"93",  x"61",  x"dc",  x"a8", -- 0488
         x"ec",  x"5a",  x"14",  x"7b",  x"06",  x"dd",  x"96",  x"04", -- 0490
         x"30",  x"1a",  x"9d",  x"a6",  x"4d",  x"44",  x"a4",  x"7c", -- 0498
         x"f1",  x"69",  x"21",  x"c5",  x"00",  x"b1",  x"d1",  x"e1", -- 04A0
         x"df",  x"f5",  x"51",  x"09",  x"38",  x"ea",  x"18",  x"de", -- 04A8
         x"04",  x"4f",  x"21",  x"dd",  x"86",  x"89",  x"d0",  x"d9", -- 04B0
         x"06",  x"fb",  x"f2",  x"4c",  x"7f",  x"06",  x"42",  x"07", -- 04B8
         x"a5",  x"4f",  x"28",  x"34",  x"cf",  x"ba",  x"53",  x"28", -- 04C0
         x"77",  x"80",  x"df",  x"ea",  x"86",  x"44",  x"11",  x"21", -- 04C8
         x"fd",  x"a9",  x"2b",  x"fd",  x"41",  x"24",  x"18",  x"0f", -- 04D0
         x"21",  x"07",  x"87",  x"27",  x"10",  x"06",  x"2a",  x"35", -- 04D8
         x"0d",  x"5e",  x"0e",  x"06",  x"44",  x"4b",  x"17",  x"de", -- 04E0
         x"15",  x"07",  x"47",  x"10",  x"a4",  x"4b",  x"f0",  x"52", -- 04E8
         x"4b",  x"10",  x"39",  x"4b",  x"c9",  x"1c",  x"4a",  x"c3", -- 04F0
         x"2c",  x"c3",  x"8d",  x"d0",  x"92",  x"20",  x"13",  x"e7", -- 04F8
         x"3a",  x"f4",  x"00",  x"2f",  x"52",  x"4f",  x"4d",  x"00", -- 0500
         x"53",  x"2f",  x"42",  x"41",  x"53",  x"49",  x"43",  x"5f", -- 0508
         x"02",  x"43",  x"30",  x"2e",  x"38",  x"37",  x"42",  x"20", -- 0510
         x"9c",  x"e8",  x"fc",  x"8a",  x"4f",  x"6b",  x"05",  x"90", -- 0518
         x"2f",  x"4f",  x"53",  x"88",  x"2c",  x"d4",  x"0a",  x"5f", -- 0520
         x"00",  x"46",  x"96",  x"2c",  x"20",  x"ad",  x"52",  x"f6", -- 0528
         x"1b",  x"89",  x"f7",  x"0a",  x"03",  x"36",  x"f6",  x"01", -- 0530
         x"cd",  x"47",  x"8c",  x"c2",  x"8a",  x"90",  x"36",  x"70", -- 0538
         x"90",  x"64",  x"2a",  x"22",  x"ad",  x"c5",  x"76",  x"07", -- 0540
         x"86",  x"06",  x"00",  x"b0",  x"86",  x"00",  x"3e",  x"9e", -- 0548
         x"f1",  x"65",  x"7c",  x"cb",  x"de",  x"f6",  x"02",  x"98", -- 0550
         x"8a",  x"4e",  x"13",  x"06",  x"50",  x"f6",  x"1a",  x"16", -- 0558
         x"11",  x"a6",  x"10",  x"d5",  x"ca",  x"c5",  x"31",  x"8f", -- 0560
         x"4b",  x"21",  x"b2",  x"26",  x"ce",  x"14",  x"db",  x"02", -- 0568
         x"01",  x"35",  x"a9",  x"7c",  x"0f",  x"45",  x"07",  x"3e", -- 0570
         x"7c",  x"03",  x"9f",  x"cd",  x"2d",  x"43",  x"86",  x"06", -- 0578
         x"21",  x"96",  x"aa",  x"cf",  x"73",  x"bc",  x"da",  x"61", -- 0580
         x"ba",  x"5a",  x"6f",  x"18",  x"74",  x"a4",  x"25",  x"3e", -- 0588
         x"0c",  x"9b",  x"03",  x"cd",  x"20",  x"fd",  x"20",  x"75", -- 0590
         x"ff",  x"18",  x"10",  x"2f",  x"11",  x"bf",  x"76",  x"81", -- 0598
         x"09",  x"5a",  x"76",  x"18",  x"86",  x"3b",  x"e7",  x"0f", -- 05A0
         x"e7",  x"12",  x"29",  x"8b",  x"40",  x"97",  x"1a",  x"cd", -- 05A8
         x"38",  x"8c",  x"26",  x"f8",  x"85",  x"db",  x"f6",  x"83", -- 05B0
         x"db",  x"fe",  x"df",  x"02",  x"7e",  x"f6",  x"29",  x"45", -- 05B8
         x"9e",  x"e0",  x"07",  x"10",  x"f8",  x"d6",  x"0a",  x"28", -- 05C0
         x"6a",  x"a2",  x"17",  x"c6",  x"ff",  x"b2",  x"be",  x"c2", -- 05C8
         x"0e",  x"0b",  x"ca",  x"c3",  x"88",  x"c2",  x"07",  x"0d", -- 05D0
         x"ca",  x"19",  x"89",  x"c5",  x"07",  x"1b",  x"28",  x"42", -- 05D8
         x"89",  x"06",  x"1f",  x"ca",  x"d1",  x"04",  x"0e",  x"20", -- 05E0
         x"ca",  x"15",  x"82",  x"07",  x"42",  x"ca",  x"f3",  x"40", -- 05E8
         x"26",  x"44",  x"ca",  x"1e",  x"8a",  x"b1",  x"07",  x"52", -- 05F0
         x"ca",  x"6b",  x"20",  x"07",  x"62",  x"28",  x"72",  x"b4", -- 05F8
         x"06",  x"64",  x"ca",  x"16",  x"72",  x"16",  x"14",  x"c3", -- 0600
         x"73",  x"8a",  x"d4",  x"20",  x"cd",  x"d9",  x"8d",  x"c3", -- 0608
         x"84",  x"fc",  x"13",  x"69",  x"e7",  x"cf",  x"30",  x"0f", -- 0610
         x"06",  x"6e",  x"14",  x"96",  x"f6",  x"da",  x"0f",  x"34", -- 0618
         x"54",  x"f6",  x"15",  x"a1",  x"cc",  x"63",  x"fd",  x"ab", -- 0620
         x"0f",  x"f7",  x"0f",  x"ec",  x"0a",  x"1d",  x"29",  x"30", -- 0628
         x"09",  x"c2",  x"70",  x"94",  x"bd",  x"1f",  x"08",  x"f7", -- 0630
         x"ed",  x"e3",  x"7e",  x"06",  x"20",  x"f5",  x"95",  x"35", -- 0638
         x"f7",  x"0d",  x"40",  x"bd",  x"fc",  x"4c",  x"85",  x"83", -- 0640
         x"34",  x"1f",  x"21",  x"10",  x"76",  x"8b",  x"e5",  x"96", -- 0648
         x"d9",  x"48",  x"0e",  x"e7",  x"e2",  x"d2",  x"f0",  x"41", -- 0650
         x"fd",  x"55",  x"01",  x"e5",  x"e3",  x"e1",  x"28",  x"d6", -- 0658
         x"98",  x"4a",  x"ad",  x"d6",  x"df",  x"f5",  x"13",  x"86", -- 0660
         x"8b",  x"52",  x"0c",  x"fa",  x"ca",  x"ed",  x"d2",  x"b6", -- 0668
         x"df",  x"f3",  x"da",  x"fa",  x"66",  x"07",  x"77",  x"fb", -- 0670
         x"f7",  x"c3",  x"dd",  x"8e",  x"fc",  x"07",  x"a9",  x"c4", -- 0678
         x"a7",  x"0d",  x"f9",  x"05",  x"4a",  x"0b",  x"fa",  x"37", -- 0680
         x"db",  x"f1",  x"0b",  x"25",  x"46",  x"fa",  x"3a",  x"a4", -- 0688
         x"0e",  x"e3",  x"56",  x"d0",  x"4a",  x"b5",  x"ca",  x"11", -- 0690
         x"a9",  x"76",  x"7e",  x"f4",  x"22",  x"34",  x"21",  x"88", -- 0698
         x"50",  x"98",  x"a7",  x"24",  x"11",  x"78",  x"2b",  x"f9", -- 06A0
         x"51",  x"e8",  x"49",  x"13",  x"39",  x"f0",  x"a3",  x"af", -- 06A8
         x"82",  x"cc",  x"aa",  x"c4",  x"9f",  x"b5",  x"14",  x"c9", -- 06B0
         x"d5",  x"ca",  x"aa",  x"97",  x"33",  x"a4",  x"10",  x"30", -- 06B8
         x"60",  x"75",  x"69",  x"5d",  x"cb",  x"7b",  x"20",  x"13", -- 06C0
         x"ab",  x"0c",  x"d4",  x"d0",  x"d6",  x"2f",  x"20",  x"03", -- 06C8
         x"e9",  x"87",  x"05",  x"81",  x"cf",  x"1d",  x"18",  x"ea", -- 06D0
         x"da",  x"8c",  x"4e",  x"64",  x"19",  x"34",  x"88",  x"21", -- 06D8
         x"32",  x"5e",  x"18",  x"66",  x"5d",  x"b7",  x"31",  x"ed", -- 06E0
         x"5b",  x"9a",  x"67",  x"3a",  x"06",  x"93",  x"3a",  x"bf", -- 06E8
         x"e2",  x"9a",  x"30",  x"52",  x"6e",  x"f3",  x"27",  x"26", -- 06F0
         x"20",  x"93",  x"ea",  x"10",  x"55",  x"46",  x"f0",  x"1f", -- 06F8
         x"34",  x"20",  x"e5",  x"ed",  x"20",  x"34",  x"a7",  x"ec", -- 0700
         x"db",  x"ef",  x"96",  x"80",  x"ee",  x"80",  x"d6",  x"90", -- 0708
         x"38",  x"e2",  x"9d",  x"c1",  x"0b",  x"18",  x"b9",  x"d6", -- 0710
         x"2d",  x"bd",  x"0a",  x"18",  x"11",  x"e9",  x"28",  x"eb", -- 0718
         x"86",  x"ca",  x"e6",  x"35",  x"ae",  x"00",  x"c3",  x"0d", -- 0720
         x"88",  x"46",  x"53",  x"20",  x"74",  x"67",  x"96",  x"6f", -- 0728
         x"3a",  x"75",  x"6e",  x"9c",  x"6d",  x"74",  x"8e",  x"52", -- 0730
         x"0d",  x"b4",  x"aa",  x"b5",  x"e9",  x"d6",  x"a1",  x"16", -- 0738
         x"72",  x"2e",  x"6f",  x"6c",  x"de",  x"87",  x"53",  x"44", -- 0740
         x"43",  x"ef",  x"43",  x"64",  x"20",  x"6b",  x"11",  x"a3", -- 0748
         x"29",  x"20",  x"6e",  x"e9",  x"62",  x"68",  x"74",  x"81", -- 0750
         x"38",  x"6f",  x"65",  x"66",  x"66",  x"6e",  x"9e",  x"38", -- 0758
         x"20",  x"77",  x"31",  x"d1",  x"cb",  x"6e",  x"df",  x"60", -- 0760
         x"2a",  x"20",  x"43",  x"75",  x"15",  x"72",  x"73",  x"6f", -- 0768
         x"9a",  x"7d",  x"ee",  x"78",  x"11",  x"39",  x"4e",  x"61", -- 0770
         x"76",  x"07",  x"69",  x"67",  x"61",  x"74",  x"69",  x"37", -- 0778
         x"4e",  x"1a",  x"45",  x"3b",  x"c1",  x"5a",  x"41",  x"75", -- 0780
         x"73",  x"77",  x"61",  x"d0",  x"65",  x"10",  x"53",  x"70", -- 0788
         x"61",  x"55",  x"63",  x"8a",  x"8d",  x"49",  x"6e",  x"66", -- 0790
         x"31",  x"6d",  x"25",  x"25",  x"b2",  x"41",  x"42",  x"14", -- 0798
         x"6b",  x"73",  x"56",  x"19",  x"56",  x"2f",  x"7a",  x"56", -- 07A0
         x"65",  x"6c",  x"70",  x"73",  x"1d",  x"20",  x"68",  x"6f", -- 07A8
         x"07",  x"e1",  x"44",  x"96",  x"b6",  x"17",  x"76",  x"17", -- 07B0
         x"6c",  x"61",  x"73",  x"ed",  x"61",  x"2e",  x"3a",  x"2b", -- 07B8
         x"fb",  x"98",  x"2d",  x"50",  x"ab",  x"00",  x"67",  x"72", -- 07C0
         x"61",  x"6d",  x"6d",  x"20",  x"73",  x"bc",  x"9b",  x"ae", -- 07C8
         x"1b",  x"4c",  x"59",  x"09",  x"7d",  x"1f",  x"26",  x"ee", -- 07D0
         x"c7",  x"00",  x"43",  x"44",  x"15",  x"8a",  x"03",  x"20", -- 07D8
         x"55",  x"70",  x"0d",  x"fb",  x"bd",  x"3c",  x"98",  x"d7", -- 07E0
         x"1b",  x"56",  x"fb",  x"85",  x"30",  x"30",  x"31",  x"20", -- 07E8
         x"62",  x"11",  x"1e",  x"db",  x"00",  x"b7",  x"8d",  x"8f", -- 07F0
         x"02",  x"d0",  x"99",  x"7e",  x"d3",  x"00",  x"19",  x"c9", -- 07F8
         x"db",  x"01",  x"b0",  x"80",  x"02",  x"d3",  x"01",  x"6f", -- 0800
         x"c9",  x"c1",  x"e1",  x"33",  x"e5",  x"c5",  x"bc",  x"12", -- 0808
         x"c8",  x"23",  x"e5",  x"88",  x"cb",  x"e1",  x"18",  x"f2", -- 0810
         x"28",  x"c9",  x"fd",  x"24",  x"fd",  x"39",  x"33",  x"fd", -- 0818
         x"56",  x"04",  x"7e",  x"00",  x"b0",  x"60",  x"30",  x"0a", -- 0820
         x"7a",  x"c6",  x"4a",  x"30",  x"1c",  x"c9",  x"d3",  x"09", -- 0828
         x"37",  x"48",  x"09",  x"47",  x"07",  x"a2",  x"00",  x"e6", -- 0830
         x"0f",  x"9c",  x"11",  x"d4",  x"11",  x"93",  x"10",  x"ce", -- 0838
         x"0c",  x"42",  x"66",  x"3f",  x"01",  x"2e",  x"9e",  x"90", -- 0840
         x"ab",  x"a7",  x"10",  x"9b",  x"0e",  x"3f",  x"0c",  x"25", -- 0848
         x"00",  x"56",  x"7a",  x"82",  x"15",  x"05",  x"07",  x"9b", -- 0850
         x"d6",  x"6a",  x"0e",  x"3e",  x"2c",  x"b2",  x"06",  x"f2", -- 0858
         x"00",  x"ec",  x"36",  x"20",  x"5d",  x"54",  x"13",  x"1f", -- 0860
         x"01",  x"bf",  x"03",  x"8b",  x"e8",  x"0c",  x"e8",  x"99", -- 0868
         x"0c",  x"5a",  x"6e",  x"32",  x"24",  x"c9",  x"79",  x"c5", -- 0870
         x"33",  x"ed",  x"4b",  x"0c",  x"06",  x"00",  x"d6",  x"cd", -- 0878
         x"c3",  x"54",  x"09",  x"c7",  x"af",  x"11",  x"2c",  x"ab", -- 0880
         x"d3",  x"5e",  x"04",  x"cb",  x"33",  x"d5",  x"01",  x"28", -- 0888
         x"a5",  x"a9",  x"69",  x"1f",  x"bf",  x"f7",  x"00",  x"da", -- 0890
         x"04",  x"28",  x"2d",  x"20",  x"4d",  x"2d",  x"3b",  x"1e", -- 0898
         x"2e",  x"ec",  x"61",  x"19",  x"88",  x"b3",  x"85",  x"04", -- 08A0
         x"85",  x"65",  x"05",  x"69",  x"db",  x"4a",  x"03",  x"5a", -- 08A8
         x"d9",  x"d6",  x"14",  x"09",  x"28",  x"21",  x"d6",  x"f8", -- 08B0
         x"9d",  x"b5",  x"20",  x"f5",  x"da",  x"2b",  x"34",  x"e1", -- 08B8
         x"79",  x"04",  x"4e",  x"6b",  x"62",  x"a2",  x"2c",  x"19", -- 08C0
         x"08",  x"30",  x"18",  x"d3",  x"46",  x"15",  x"da",  x"a9", -- 08C8
         x"94",  x"19",  x"b9",  x"3a",  x"12",  x"02",  x"13",  x"18", -- 08D0
         x"b2",  x"3e",  x"17",  x"fd",  x"81",  x"3d",  x"fd",  x"96", -- 08D8
         x"00",  x"30",  x"05",  x"20",  x"80",  x"a1",  x"33",  x"d0", -- 08E0
         x"84",  x"3d",  x"01",  x"12",  x"f9",  x"bf",  x"c2",  x"d8", -- 08E8
         x"3d",  x"04",  x"e8",  x"b1",  x"4f",  x"47",  x"1b",  x"79", -- 08F0
         x"47",  x"44",  x"9e",  x"07",  x"64",  x"78",  x"9e",  x"77", -- 08F8
         x"6d",  x"eb",  x"9d",  x"b6",  x"06",  x"37",  x"06",  x"06", -- 0900
         x"a4",  x"03",  x"cb",  x"05",  x"3e",  x"03",  x"1d",  x"04", -- 0908
         x"1e",  x"10",  x"83",  x"16",  x"34",  x"ff",  x"a2",  x"02", -- 0910
         x"04",  x"38",  x"cf",  x"e1",  x"57",  x"13",  x"4e",  x"06", -- 0918
         x"28",  x"e0",  x"10",  x"23",  x"10",  x"fb",  x"c9",  x"14", -- 0920
         x"01",  x"07",  x"00",  x"0e",  x"21",  x"31",  x"d1",  x"8d", -- 0928
         x"e7",  x"67",  x"c3",  x"07",  x"3e",  x"05",  x"9d",  x"79", -- 0930
         x"06",  x"f0",  x"c9",  x"55",  x"cb",  x"66",  x"0a",  x"31", -- 0938
         x"00",  x"0d",  x"89",  x"ec",  x"0d",  x"0a",  x"c1",  x"d1", -- 0940
         x"01",  x"ed",  x"53",  x"d7",  x"03",  x"21",  x"bd",  x"c0", -- 0948
         x"86",  x"2d",  x"03",  x"01",  x"67",  x"00",  x"2d",  x"eb", -- 0950
         x"00",  x"f9",  x"af",  x"32",  x"ab",  x"03",  x"32",  x"00", -- 0958
         x"04",  x"28",  x"2a",  x"36",  x"41",  x"ff",  x"22",  x"01", -- 0960
         x"b0",  x"03",  x"19",  x"22",  x"56",  x"03",  x"3e",  x"80", -- 0968
         x"14",  x"fc",  x"03",  x"cd",  x"4f",  x"c6",  x"23",  x"eb", -- 0970
         x"00",  x"cd",  x"93",  x"c4",  x"cd",  x"69",  x"c6",  x"c3", -- 0978
         x"54",  x"21",  x"c8",  x"c9",  x"21",  x"3a",  x"21",  x"c0", -- 0980
         x"01",  x"55",  x"2c",  x"1f",  x"09",  x"6b",  x"42",  x"41", -- 0988
         x"5e",  x"41",  x"90",  x"49",  x"31",  x"67",  x"ba",  x"24", -- 0990
         x"0d",  x"b0",  x"47",  x"3e",  x"ff",  x"d3",  x"04",  x"29", -- 0998
         x"db",  x"05",  x"c6",  x"06",  x"db",  x"04",  x"6f",  x"0c", -- 09A0
         x"3c",  x"25",  x"d3",  x"07",  x"98",  x"3a",  x"07",  x"93", -- 09A8
         x"15",  x"c9",  x"a0",  x"d3",  x"06",  x"c3",  x"6e",  x"49", -- 09B0
         x"8e",  x"0b",  x"cb",  x"09",  x"13",  x"28",  x"20",  x"04", -- 09B8
         x"c9",  x"16",  x"22",  x"5a",  x"00",  x"4d",  x"00",  x"15", -- 09C0
         x"7a",  x"19",  x"f0",  x"10",  x"ea",  x"34",  x"ae",  x"2a", -- 09C8
         x"7e",  x"ce",  x"2d",  x"05",  x"be",  x"8b",  x"af",  x"09", -- 09D0
         x"c0",  x"4a",  x"13",  x"59",  x"e5",  x"03",  x"3e",  x"77", -- 09D8
         x"48",  x"cc",  x"bc",  x"51",  x"8e",  x"9b",  x"e0",  x"57", -- 09E0
         x"95",  x"da",  x"98",  x"8f",  x"cd",  x"28",  x"94",  x"8e", -- 09E8
         x"f9",  x"68",  x"13",  x"9c",  x"8e",  x"39",  x"33",  x"f5", -- 09F0
         x"f6",  x"72",  x"05",  x"fc",  x"06",  x"19",  x"dd",  x"56", -- 09F8
         x"07",  x"c8",  x"80",  x"08",  x"f1",  x"06",  x"18",  x"cb", -- 0A00
         x"3b",  x"cb",  x"06",  x"1a",  x"cb",  x"1d",  x"cb",  x"1c", -- 0A08
         x"f5",  x"28",  x"e5",  x"4d",  x"1f",  x"10",  x"0f",  x"23", -- 0A10
         x"1f",  x"08",  x"ea",  x"1f",  x"1e",  x"52",  x"08",  x"26", -- 0A18
         x"01",  x"80",  x"73",  x"d6",  x"40",  x"20",  x"02",  x"26", -- 0A20
         x"95",  x"b5",  x"08",  x"48",  x"25",  x"08",  x"87",  x"19", -- 0A28
         x"3a",  x"16",  x"0a",  x"b3",  x"c0",  x"eb",  x"d1",  x"cb", -- 0A30
         x"6b",  x"7d",  x"c4",  x"60",  x"ce",  x"f2",  x"a0",  x"bb", -- 0A38
         x"d1",  x"9c",  x"08",  x"a1",  x"cd",  x"88",  x"8e",  x"40", -- 0A40
         x"a8",  x"e1",  x"8a",  x"c9",  x"30",  x"f5",  x"f5",  x"3b", -- 0A48
         x"cd",  x"0d",  x"7b",  x"8e",  x"26",  x"64",  x"1a",  x"a9", -- 0A50
         x"ab",  x"17",  x"25",  x"de",  x"9d",  x"f6",  x"b5",  x"5c", -- 0A58
         x"26",  x"b6",  x"0b",  x"d0",  x"78",  x"df",  x"45",  x"02", -- 0A60
         x"f5",  x"40",  x"70",  x"f5",  x"09",  x"2d",  x"c2",  x"25", -- 0A68
         x"91",  x"53",  x"4d",  x"af",  x"1a",  x"1e",  x"aa",  x"01", -- 0A70
         x"1e",  x"48",  x"24",  x"1e",  x"ad",  x"90",  x"a6",  x"15", -- 0A78
         x"39",  x"f3",  x"67",  x"00",  x"68",  x"cd",  x"8d",  x"19", -- 0A80
         x"c5",  x"ec",  x"8e",  x"0d",  x"7d",  x"d1",  x"cf",  x"c5", -- 0A88
         x"77",  x"04",  x"78",  x"19",  x"f4",  x"eb",  x"d5",  x"2b", -- 0A90
         x"3b",  x"d1",  x"ff",  x"40",  x"23",  x"23",  x"7e",  x"3d", -- 0A98
         x"a1",  x"4b",  x"d5",  x"fd",  x"e1",  x"b8",  x"d0",  x"03", -- 0AA0
         x"d6",  x"aa",  x"a0",  x"0a",  x"01",  x"10",  x"27",  x"78", -- 0AA8
         x"1c",  x"b1",  x"28",  x"28",  x"32",  x"a9",  x"79",  x"40", -- 0AB0
         x"53",  x"79",  x"e9",  x"d6",  x"5a",  x"45",  x"ca",  x"0a", -- 0AB8
         x"0a",  x"50",  x"c3",  x"b0",  x"09",  x"1a",  x"0b",  x"18", -- 0AC0
         x"d4",  x"2b",  x"ca",  x"91",  x"3e",  x"af",  x"40",  x"a4", -- 0AC8
         x"7a",  x"89",  x"2a",  x"52",  x"b7",  x"4f",  x"47",  x"14", -- 0AD0
         x"81",  x"0c",  x"d1",  x"47",  x"77",  x"28",  x"04",  x"93", -- 0AD8
         x"61",  x"18",  x"02",  x"3e",  x"04",  x"4c",  x"b2",  x"c3", -- 0AE0
         x"e3",  x"26",  x"01",  x"e7",  x"e9",  x"14",  x"dd",  x"45", -- 0AE8
         x"38",  x"08",  x"08",  x"86",  x"02",  x"16",  x"e9",  x"28", -- 0AF0
         x"18",  x"06",  x"07",  x"01",  x"16",  x"4a",  x"41",  x"9f", -- 0AF8
         x"0e",  x"26",  x"50",  x"2d",  x"31",  x"d5",  x"0a",  x"82", -- 0B00
         x"9d",  x"d6",  x"91",  x"29",  x"1a",  x"2d",  x"27",  x"02", -- 0B08
         x"59",  x"50",  x"10",  x"9c",  x"1a",  x"27",  x"04",  x"56", -- 0B10
         x"b0",  x"0a",  x"ff",  x"32",  x"1f",  x"b2",  x"8f",  x"12", -- 0B18
         x"3e",  x"02",  x"94",  x"1a",  x"80",  x"de",  x"5d",  x"10", -- 0B20
         x"73",  x"1a",  x"9b",  x"83",  x"9a",  x"2e",  x"df",  x"24", -- 0B28
         x"f9",  x"59",  x"ab",  x"18",  x"3b",  x"21",  x"28",  x"cb", -- 0B30
         x"5e",  x"20",  x"33",  x"16",  x"f5",  x"94",  x"d8",  x"eb", -- 0B38
         x"cb",  x"06",  x"66",  x"26",  x"03",  x"07",  x"16",  x"03", -- 0B40
         x"08",  x"a0",  x"03",  x"09",  x"16",  x"10",  x"ee",  x"ab", -- 0B48
         x"4c",  x"e2",  x"dc",  x"b9",  x"f0",  x"af",  x"16",  x"66", -- 0B50
         x"09",  x"e5",  x"c0",  x"66",  x"66",  x"07",  x"6f",  x"51", -- 0B58
         x"89",  x"6f",  x"04",  x"20",  x"74",  x"11",  x"40",  x"9c", -- 0B60
         x"86",  x"97",  x"7d",  x"03",  x"3c",  x"20",  x"05",  x"1b", -- 0B68
         x"7a",  x"b3",  x"97",  x"30",  x"7d",  x"d6",  x"fe",  x"20", -- 0B70
         x"61",  x"5e",  x"78",  x"dd",  x"96",  x"0a",  x"67",  x"41", -- 0B78
         x"05",  x"9e",  x"0b",  x"6f",  x"7c",  x"8d",  x"0a",  x"0c", -- 0B80
         x"67",  x"7d",  x"09",  x"0d",  x"fb",  x"fa",  x"fd",  x"97", -- 0B88
         x"16",  x"fe",  x"8b",  x"00",  x"0b",  x"dd",  x"b6",  x"0a", -- 0B90
         x"28",  x"6c",  x"10",  x"4d",  x"0a",  x"4d",  x"0b",  x"e5", -- 0B98
         x"a0",  x"3b",  x"e1",  x"2b",  x"7c",  x"b5",  x"cf",  x"98", -- 0BA0
         x"0f",  x"5a",  x"04",  x"a4",  x"1a",  x"5e",  x"0c",  x"a4", -- 0BA8
         x"12",  x"0d",  x"e5",  x"8e",  x"d9",  x"d8",  x"2b",  x"23", -- 0BB0
         x"52",  x"77",  x"f1",  x"b2",  x"15",  x"26",  x"41",  x"df", -- 0BB8
         x"41",  x"d9",  x"a3",  x"2d",  x"ff",  x"02",  x"c8",  x"76", -- 0BC0
         x"3d",  x"08",  x"3d",  x"09",  x"38",  x"43",  x"4a",  x"a9", -- 0BC8
         x"1b",  x"b0",  x"28",  x"07",  x"68",  x"06",  x"3f",  x"ee", -- 0BD0
         x"de",  x"31",  x"99",  x"29",  x"d3",  x"24",  x"82",  x"0f", -- 0BD8
         x"29",  x"a0",  x"2a",  x"1f",  x"de",  x"05",  x"fc",  x"05", -- 0BE0
         x"28",  x"77",  x"5b",  x"fd",  x"1e",  x"4e",  x"3b",  x"00", -- 0BE8
         x"46",  x"09",  x"51",  x"58",  x"0b",  x"7b",  x"b2",  x"28", -- 0BF0
         x"78",  x"2e",  x"4e",  x"24",  x"66",  x"ff",  x"7e",  x"e3", -- 0BF8
         x"d2",  x"cb",  x"05",  x"03",  x"40",  x"d7",  x"5f",  x"17", -- 0C00
         x"9f",  x"61",  x"57",  x"84",  x"4b",  x"0e",  x"fc",  x"0e", -- 0C08
         x"30",  x"fd",  x"67",  x"0e",  x"6f",  x"7b",  x"94",  x"5f", -- 0C10
         x"00",  x"7a",  x"9d",  x"57",  x"6b",  x"7a",  x"67",  x"b3", -- 0C18
         x"28",  x"46",  x"cb",  x"00",  x"89",  x"21",  x"ef",  x"ff", -- 0C20
         x"3a",  x"39",  x"f9",  x"8a",  x"2d",  x"20",  x"b2",  x"bf", -- 0C28
         x"54",  x"02",  x"6a",  x"de",  x"fb",  x"14",  x"69",  x"04", -- 0C30
         x"65",  x"07",  x"04",  x"38",  x"21",  x"a0",  x"95",  x"66", -- 0C38
         x"06",  x"fd",  x"00",  x"6e",  x"07",  x"fd",  x"46",  x"08", -- 0C40
         x"fd",  x"4e",  x"09",  x"a5",  x"24",  x"94",  x"29",  x"23", -- 0C48
         x"9d",  x"22",  x"98",  x"40",  x"21",  x"99",  x"38",  x"09", -- 0C50
         x"21",  x"01",  x"e3",  x"99",  x"47",  x"00",  x"c3",  x"3e", -- 0C58
         x"95",  x"1a",  x"67",  x"d6",  x"01",  x"da",  x"05",  x"38", -- 0C60
         x"95",  x"3e",  x"03",  x"94",  x"0b",  x"05",  x"7c",  x"c6", -- 0C68
         x"ff",  x"b2",  x"09",  x"2e",  x"94",  x"bd",  x"9f",  x"19", -- 0C70
         x"a0",  x"ee",  x"c5",  x"21",  x"10",  x"a5",  x"8c",  x"2a", -- 0C78
         x"01",  x"04",  x"dd",  x"18",  x"c1",  x"f7",  x"3a",  x"ff", -- 0C80
         x"f8",  x"0c",  x"21",  x"23",  x"93",  x"19",  x"00",  x"d1", -- 0C88
         x"e9",  x"00",  x"c3",  x"2c",  x"93",  x"c3",  x"41",  x"94", -- 0C90
         x"c3",  x"b9",  x"72",  x"94",  x"fc",  x"cb",  x"6c",  x"3c", -- 0C98
         x"e4",  x"09",  x"00",  x"4d",  x"7c",  x"e6",  x"01",  x"47", -- 0CA0
         x"7c",  x"cb",  x"3f",  x"d8",  x"3f",  x"f7",  x"bc",  x"9a", -- 0CA8
         x"f8",  x"00",  x"03",  x"f9",  x"94",  x"03",  x"fa",  x"8f", -- 0CB0
         x"03",  x"fb",  x"dd",  x"86",  x"11",  x"3c",  x"77",  x"f3", -- 0CB8
         x"08",  x"84",  x"4d",  x"8e",  x"f8",  x"08",  x"f4",  x"b7", -- 0CC0
         x"08",  x"fd",  x"08",  x"f9",  x"08",  x"42",  x"a5",  x"fe", -- 0CC8
         x"d9",  x"08",  x"fa",  x"08",  x"f6",  x"79",  x"96",  x"d4", -- 0CD0
         x"da",  x"82",  x"3d",  x"28",  x"2c",  x"45",  x"f7",  x"a8", -- 0CD8
         x"d9",  x"d3",  x"f2",  x"98",  x"1a",  x"ca",  x"7d",  x"b4", -- 0CE0
         x"fc",  x"06",  x"36",  x"66",  x"f4",  x"a2",  x"a6",  x"31", -- 0CE8
         x"47",  x"91",  x"bb",  x"5e",  x"0a",  x"e9",  x"b3",  x"f9", -- 0CF0
         x"8c",  x"3c",  x"ca",  x"1f",  x"75",  x"a9",  x"2c",  x"2b", -- 0CF8
         x"4d",  x"44",  x"61",  x"c5",  x"e6",  x"a5",  x"b1",  x"06", -- 0D00
         x"ca",  x"a1",  x"99",  x"c1",  x"a3",  x"e5",  x"48",  x"34", -- 0D08
         x"fd",  x"e5",  x"ba",  x"35",  x"dc",  x"46",  x"c2",  x"34", -- 0D10
         x"eb",  x"14",  x"5e",  x"23",  x"56",  x"b6",  x"c1",  x"2b", -- 0D18
         x"6e",  x"67",  x"7b",  x"41",  x"94",  x"8d",  x"d9",  x"01", -- 0D20
         x"90",  x"57",  x"7d",  x"41",  x"8c",  x"47",  x"bc",  x"80", -- 0D28
         x"88",  x"67",  x"1c",  x"20",  x"30",  x"07",  x"14",  x"88", -- 0D30
         x"05",  x"2c",  x"20",  x"01",  x"24",  x"03",  x"37",  x"57", -- 0D38
         x"01",  x"55",  x"c5",  x"02",  x"f1",  x"03",  x"7d",  x"b7", -- 0D40
         x"49",  x"47",  x"61",  x"7c",  x"7e",  x"23",  x"66",  x"6f", -- 0D48
         x"52",  x"dc",  x"46",  x"d7",  x"b3",  x"9d",  x"cb",  x"80", -- 0D50
         x"10",  x"10",  x"fa",  x"18",  x"04",  x"c4",  x"82",  x"0f", -- 0D58
         x"67",  x"94",  x"d5",  x"5b",  x"69",  x"b9",  x"14",  x"29", -- 0D60
         x"eb",  x"8e",  x"18",  x"c8",  x"b3",  x"6e",  x"84",  x"66", -- 0D68
         x"46",  x"81",  x"4e",  x"6d",  x"07",  x"90",  x"c8",  x"8e", -- 0D70
         x"39",  x"cb",  x"18",  x"b9",  x"8e",  x"3c",  x"3d",  x"20", -- 0D78
         x"19",  x"96",  x"52",  x"84",  x"8a",  x"94",  x"8d",  x"51", -- 0D80
         x"92",  x"4a",  x"88",  x"90",  x"2a",  x"89",  x"8e",  x"18", -- 0D88
         x"90",  x"da",  x"b1",  x"8b",  x"43",  x"d5",  x"61",  x"d6", -- 0D90
         x"20",  x"d5",  x"65",  x"80",  x"61",  x"8b",  x"31",  x"77", -- 0D98
         x"cb",  x"bd",  x"50",  x"79",  x"82",  x"7a",  x"07",  x"0c", -- 0DA0
         x"50",  x"7a",  x"04",  x"40",  x"7a",  x"20",  x"78",  x"11", -- 0DA8
         x"79",  x"ce",  x"98",  x"46",  x"23",  x"d4",  x"86",  x"4e", -- 0DB0
         x"6a",  x"60",  x"79",  x"fa",  x"0d",  x"57",  x"e7",  x"e5", -- 0DB8
         x"d5",  x"38",  x"d6",  x"fb",  x"4c",  x"f5",  x"a5",  x"86", -- 0DC0
         x"c6",  x"fe",  x"60",  x"04",  x"a4",  x"84",  x"51",  x"ce", -- 0DC8
         x"e2",  x"a9",  x"05",  x"88",  x"2d",  x"07",  x"06",  x"49", -- 0DD0
         x"8c",  x"6b",  x"07",  x"07",  x"af",  x"4d",  x"f7",  x"b4", -- 0DD8
         x"b2",  x"99",  x"af",  x"1e",  x"7d",  x"2c",  x"93",  x"59", -- 0DE0
         x"18",  x"67",  x"78",  x"9a",  x"03",  x"47",  x"79",  x"03", -- 0DE8
         x"4f",  x"94",  x"3e",  x"95",  x"3a",  x"9c",  x"88",  x"bf", -- 0DF0
         x"45",  x"07",  x"57",  x"5b",  x"f2",  x"ae",  x"4e",  x"86", -- 0DF8
         x"9d",  x"4e",  x"aa",  x"53",  x"0d",  x"d5",  x"b5",  x"39", -- 0E00
         x"9e",  x"b9",  x"56",  x"a4",  x"c0",  x"ac",  x"53",  x"a8", -- 0E08
         x"51",  x"f1",  x"00",  x"dd",  x"72",  x"96",  x"5f",  x"73", -- 0E10
         x"fe",  x"94",  x"e1",  x"75",  x"fc",  x"e1",  x"11",  x"f9", -- 0E18
         x"eb",  x"19",  x"56",  x"61",  x"b0",  x"85",  x"b6",  x"01", -- 0E20
         x"ff",  x"82",  x"6f",  x"40",  x"fd",  x"8b",  x"58",  x"67", -- 0E28
         x"fb",  x"2a",  x"5f",  x"bb",  x"08",  x"88",  x"57",  x"e0", -- 0E30
         x"b8",  x"61",  x"2a",  x"b7",  x"41",  x"cd",  x"46",  x"84", -- 0E38
         x"7e",  x"0b",  x"d6",  x"03",  x"20",  x"1f",  x"c2",  x"02", -- 0E40
         x"14",  x"6f",  x"c0",  x"c0",  x"00",  x"67",  x"a3",  x"c7", -- 0E48
         x"a7",  x"16",  x"3e",  x"80",  x"a0",  x"23",  x"cb",  x"12", -- 0E50
         x"cb",  x"11",  x"24",  x"cb",  x"10",  x"d6",  x"1d",  x"1e", -- 0E58
         x"1a",  x"36",  x"1e",  x"8f",  x"4b",  x"6e",  x"f3",  x"66", -- 0E60
         x"75",  x"73",  x"36",  x"2d",  x"fe",  x"00",  x"ca",  x"f3", -- 0E68
         x"ee",  x"0f",  x"b6",  x"fc",  x"6f",  x"7a",  x"04",  x"d3", -- 0E70
         x"66",  x"79",  x"04",  x"fe",  x"34",  x"5f",  x"78",  x"04", -- 0E78
         x"ff",  x"7c",  x"6c",  x"89",  x"6e",  x"e3",  x"57",  x"fa", -- 0E80
         x"d7",  x"16",  x"af",  x"d3",  x"e5",  x"77",  x"c5",  x"dd", -- 0E88
         x"d9",  x"39",  x"c8",  x"fa",  x"fd",  x"6e",  x"c8",  x"fb", -- 0E90
         x"ed",  x"05",  x"c8",  x"fb",  x"05",  x"c8",  x"7d",  x"66", -- 0E98
         x"fa",  x"a8",  x"72",  x"12",  x"c9",  x"b2",  x"84",  x"50", -- 0EA0
         x"0c",  x"c8",  x"7e",  x"05",  x"1a",  x"c9",  x"1c",  x"fb", -- 0EA8
         x"b7",  x"21",  x"bd",  x"25",  x"11",  x"06",  x"e1",  x"0a", -- 0EB0
         x"e5",  x"4a",  x"9f",  x"4d",  x"26",  x"92",  x"4a",  x"24", -- 0EB8
         x"9b",  x"22",  x"50",  x"9c",  x"20",  x"9d",  x"38",  x"05", -- 0EC0
         x"e8",  x"98",  x"c3",  x"65",  x"62",  x"97",  x"0a",  x"f8", -- 0EC8
         x"c6",  x"0e",  x"81",  x"f1",  x"f9",  x"82",  x"aa",  x"57", -- 0ED0
         x"a8",  x"16",  x"9b",  x"36",  x"02",  x"fb",  x"02",  x"fa", -- 0ED8
         x"3b",  x"20",  x"15",  x"3f",  x"ea",  x"05",  x"0e",  x"37", -- 0EE0
         x"f5",  x"46",  x"3b",  x"f5",  x"03",  x"d1",  x"21",  x"08", -- 0EE8
         x"00",  x"09",  x"11",  x"5c",  x"eb",  x"12",  x"ef",  x"11", -- 0EF0
         x"0c",  x"11",  x"dd",  x"0a",  x"d4",  x"14",  x"ff",  x"59", -- 0EF8
         x"3e",  x"28",  x"17",  x"8e",  x"f9",  x"0a",  x"66",  x"cf", -- 0F00
         x"a6",  x"06",  x"6c",  x"fa",  x"06",  x"fb",  x"80",  x"8c", -- 0F08
         x"43",  x"95",  x"fe",  x"73",  x"cd",  x"09",  x"18",  x"08", -- 0F10
         x"eb",  x"4e",  x"0d",  x"a5",  x"56",  x"2c",  x"ee",  x"00", -- 0F18
         x"71",  x"23",  x"70",  x"23",  x"73",  x"23",  x"72",  x"ee", -- 0F20
         x"a6",  x"36",  x"cf",  x"15",  x"f0",  x"cf",  x"16",  x"81", -- 0F28
         x"31",  x"93",  x"bb",  x"25",  x"30",  x"32",  x"39",  x"13", -- 0F30
         x"c2",  x"e4",  x"e1",  x"72",  x"f3",  x"a1",  x"c1",  x"14", -- 0F38
         x"f2",  x"28",  x"23",  x"af",  x"44",  x"c6",  x"0c",  x"92", -- 0F40
         x"d3",  x"ff",  x"c2",  x"c0",  x"c6",  x"8c",  x"49",  x"75", -- 0F48
         x"8b",  x"d6",  x"b6",  x"c3",  x"b3",  x"b2",  x"a2",  x"b0", -- 0F50
         x"2e",  x"03",  x"c3",  x"ce",  x"a3",  x"a8",  x"68",  x"f2", -- 0F58
         x"94",  x"c2",  x"36",  x"bd",  x"98",  x"d4",  x"6c",  x"07", -- 0F60
         x"da",  x"04",  x"6c",  x"0c",  x"d7",  x"04",  x"95",  x"29", -- 0F68
         x"72",  x"54",  x"7e",  x"84",  x"16",  x"46",  x"08",  x"a1", -- 0F70
         x"dd",  x"99",  x"46",  x"fb",  x"28",  x"b5",  x"54",  x"6c", -- 0F78
         x"ae",  x"46",  x"b2",  x"91",  x"d4",  x"19",  x"ce",  x"2b", -- 0F80
         x"04",  x"ce",  x"15",  x"66",  x"50",  x"4a",  x"c8",  x"8e", -- 0F88
         x"f3",  x"9c",  x"da",  x"4d",  x"7d",  x"5a",  x"31",  x"f8", -- 0F90
         x"5a",  x"11",  x"05",  x"f9",  x"b9",  x"86",  x"cb",  x"e5", -- 0F98
         x"04",  x"03",  x"f8",  x"1e",  x"1f",  x"85",  x"31",  x"8b", -- 0FA0
         x"f9",  x"6e",  x"81",  x"66",  x"2b",  x"d5",  x"e6",  x"a6", -- 0FA8
         x"f8",  x"c1",  x"9b",  x"04",  x"f9",  x"cb",  x"b5",  x"70", -- 0FB0
         x"69",  x"d3",  x"9a",  x"92",  x"63",  x"89",  x"e8",  x"ce", -- 0FB8
         x"b9",  x"3e",  x"00",  x"6c",  x"98",  x"02",  x"9b",  x"02", -- 0FC0
         x"9a",  x"38",  x"f4",  x"a7",  x"01",  x"18",  x"51",  x"66", -- 0FC8
         x"e1",  x"24",  x"e5",  x"d7",  x"24",  x"f4",  x"84",  x"d7", -- 0FD0
         x"f5",  x"e8",  x"05",  x"91",  x"1a",  x"f6",  x"05",  x"09", -- 0FD8
         x"a7",  x"c5",  x"a9",  x"33",  x"96",  x"f4",  x"a8",  x"31", -- 0FE0
         x"9e",  x"f5",  x"7b",  x"9b",  x"03",  x"f6",  x"7a",  x"03", -- 0FE8
         x"f7",  x"31",  x"c9",  x"7a",  x"18",  x"34",  x"42",  x"a5", -- 0FF0
         x"61",  x"c3",  x"ca",  x"95",  x"41",  x"e3",  x"25",  x"45", -- 0FF8
         x"4c",  x"d8",  x"0d",  x"13",  x"71",  x"72",  x"15",  x"8d", -- 1000
         x"b5",  x"06",  x"a2",  x"c3",  x"74",  x"a1",  x"0c",  x"77", -- 1008
         x"e8",  x"63",  x"ce",  x"e9",  x"75",  x"a0",  x"2b",  x"69", -- 1010
         x"96",  x"db",  x"44",  x"c2",  x"a8",  x"99",  x"6e",  x"ae", -- 1018
         x"25",  x"fe",  x"da",  x"19",  x"06",  x"d8",  x"e8",  x"48", -- 1020
         x"fe",  x"18",  x"7a",  x"c7",  x"ad",  x"6f",  x"d6",  x"e9", -- 1028
         x"00",  x"e3",  x"2b",  x"6a",  x"11",  x"81",  x"34",  x"19", -- 1030
         x"c2",  x"aa",  x"21",  x"27",  x"20",  x"00",  x"f1",  x"2c", -- 1038
         x"e9",  x"26",  x"82",  x"68",  x"c9",  x"b0",  x"fd",  x"92", -- 1040
         x"16",  x"83",  x"ea",  x"02",  x"b9",  x"b6",  x"7a",  x"a6", -- 1048
         x"89",  x"4e",  x"5f",  x"1f",  x"7e",  x"09",  x"13",  x"80", -- 1050
         x"cc",  x"40",  x"01",  x"0b",  x"ce",  x"c7",  x"bd",  x"96", -- 1058
         x"27",  x"2a",  x"68",  x"23",  x"e9",  x"4d",  x"f4",  x"25", -- 1060
         x"23",  x"57",  x"d5",  x"1c",  x"0c",  x"5c",  x"92",  x"35", -- 1068
         x"c7",  x"bb",  x"00",  x"7c",  x"d1",  x"94",  x"28",  x"4b", -- 1070
         x"11",  x"26",  x"86",  x"11",  x"6a",  x"97",  x"f1",  x"55", -- 1078
         x"4c",  x"ca",  x"11",  x"06",  x"99",  x"6a",  x"e0",  x"d9", -- 1080
         x"3b",  x"ab",  x"f6",  x"47",  x"03",  x"04",  x"ce",  x"24", -- 1088
         x"ab",  x"73",  x"27",  x"8f",  x"f4",  x"c0",  x"b0",  x"b1", -- 1090
         x"ca",  x"6e",  x"9a",  x"96",  x"56",  x"a6",  x"c3",  x"24", -- 1098
         x"e5",  x"34",  x"dc",  x"c0",  x"cf",  x"74",  x"fb",  x"8a", -- 10A0
         x"d9",  x"0c",  x"e9",  x"61",  x"50",  x"d9",  x"50",  x"3e", -- 10A8
         x"d9",  x"29",  x"3e",  x"58",  x"f9",  x"82",  x"d1",  x"39", -- 10B0
         x"5e",  x"21",  x"55",  x"da",  x"8d",  x"80",  x"86",  x"18", -- 10B8
         x"28",  x"b0",  x"de",  x"00",  x"7e",  x"e6",  x"3f",  x"67", -- 10C0
         x"7a",  x"fe",  x"e5",  x"28",  x"18",  x"08",  x"d6",  x"2e", -- 10C8
         x"2d",  x"cb",  x"5c",  x"28",  x"45",  x"13",  x"07",  x"c4", -- 10D0
         x"65",  x"78",  x"ce",  x"d9",  x"a1",  x"ff",  x"c9",  x"3e", -- 10D8
         x"28",  x"0f",  x"42",  x"9a",  x"d9",  x"f8",  x"23",  x"7a", -- 10E0
         x"04",  x"0e",  x"f9",  x"38",  x"dd",  x"12",  x"3b",  x"95", -- 10E8
         x"b7",  x"35",  x"da",  x"25",  x"ad",  x"f0",  x"04",  x"cf", -- 10F0
         x"e5",  x"b1",  x"a4",  x"3d",  x"01",  x"20",  x"03",  x"4f", -- 10F8
         x"10",  x"63",  x"a6",  x"bd",  x"77",  x"fd",  x"2a",  x"f3", -- 1100
         x"f3",  x"c4",  x"e7",  x"93",  x"c6",  x"75",  x"07",  x"bb", -- 1108
         x"c0",  x"5e",  x"aa",  x"0e",  x"aa",  x"36",  x"b9",  x"18", -- 1110
         x"60",  x"04",  x"6c",  x"da",  x"03",  x"19",  x"4e",  x"3e", -- 1118
         x"20",  x"91",  x"ad",  x"05",  x"17",  x"0e",  x"97",  x"6f", -- 1120
         x"42",  x"06",  x"79",  x"fe",  x"2f",  x"28",  x"3d",  x"95", -- 1128
         x"0b",  x"20",  x"c3",  x"01",  x"01",  x"af",  x"67",  x"82", -- 1130
         x"b5",  x"08",  x"d8",  x"cc",  x"96",  x"fe",  x"28",  x"38", -- 1138
         x"14",  x"b4",  x"40",  x"d6",  x"08",  x"20",  x"21",  x"b4", -- 1140
         x"28",  x"57",  x"1e",  x"4f",  x"15",  x"8f",  x"4f",  x"0b", -- 1148
         x"18",  x"bf",  x"78",  x"1b",  x"34",  x"34",  x"fd",  x"d1", -- 1150
         x"1f",  x"86",  x"fb",  x"6f",  x"41",  x"ad",  x"a0",  x"fc", -- 1158
         x"67",  x"71",  x"18",  x"ab",  x"51",  x"68",  x"52",  x"fd", -- 1160
         x"75",  x"94",  x"60",  x"74",  x"01",  x"e4",  x"e5",  x"c6", -- 1168
         x"0b",  x"3a",  x"d1",  x"fc",  x"47",  x"d1",  x"7f",  x"ff", -- 1170
         x"d1",  x"51",  x"65",  x"02",  x"9d",  x"12",  x"84",  x"13", -- 1178
         x"81",  x"22",  x"ec",  x"55",  x"a1",  x"93",  x"09",  x"12", -- 1180
         x"a1",  x"09",  x"30",  x"a1",  x"ac",  x"e4",  x"2c",  x"df", -- 1188
         x"e5",  x"a5",  x"25",  x"7e",  x"90",  x"a4",  x"5d",  x"9c", -- 1190
         x"c1",  x"12",  x"c5",  x"1e",  x"00",  x"8a",  x"e0",  x"16", -- 1198
         x"9b",  x"91",  x"d1",  x"16",  x"20",  x"b0",  x"23",  x"d6", -- 11A0
         x"05",  x"20",  x"d5",  x"30",  x"e5",  x"7a",  x"02",  x"03", -- 11A8
         x"30",  x"1c",  x"7b",  x"ae",  x"09",  x"38",  x"e2",  x"33", -- 11B0
         x"33",  x"88",  x"a3",  x"11",  x"08",  x"f8",  x"21",  x"c6", -- 11B8
         x"c6",  x"20",  x"1f",  x"3e",  x"2e",  x"1b",  x"1e",  x"e7", -- 11C0
         x"69",  x"35",  x"f4",  x"68",  x"13",  x"08",  x"82",  x"2d", -- 11C8
         x"0b",  x"38",  x"ea",  x"ed",  x"2d",  x"80",  x"ee",  x"f8", -- 11D0
         x"ac",  x"b4",  x"24",  x"24",  x"90",  x"b0",  x"aa",  x"d6", -- 11D8
         x"42",  x"06",  x"c6",  x"1c",  x"6f",  x"f3",  x"99",  x"c9", -- 11E0
         x"ab",  x"d5",  x"7c",  x"85",  x"12",  x"4e",  x"95",  x"b4", -- 11E8
         x"bd",  x"b8",  x"2d",  x"e3",  x"bb",  x"37",  x"04",  x"31", -- 11F0
         x"37",  x"5a",  x"5f",  x"2b",  x"18",  x"6a",  x"2b",  x"27", -- 11F8
         x"26",  x"6a",  x"63",  x"1f",  x"45",  x"06",  x"23",  x"1f", -- 1200
         x"16",  x"b2",  x"1f",  x"b5",  x"47",  x"36",  x"42",  x"fb", -- 1208
         x"f6",  x"a3",  x"fb",  x"62",  x"67",  x"08",  x"62",  x"09", -- 1210
         x"46",  x"d4",  x"86",  x"13",  x"78",  x"bb",  x"07",  x"20", -- 1218
         x"0a",  x"d8",  x"9c",  x"f2",  x"61",  x"10",  x"72",  x"09", -- 1220
         x"18",  x"ed",  x"9e",  x"a5",  x"07",  x"74",  x"6c",  x"09", -- 1228
         x"14",  x"2f",  x"d6",  x"e5",  x"12",  x"96",  x"a3",  x"fe", -- 1230
         x"a0",  x"9e",  x"83",  x"a5",  x"9c",  x"08",  x"a3",  x"b8", -- 1238
         x"ba",  x"48",  x"80",  x"11",  x"30",  x"11",  x"c5",  x"6c", -- 1240
         x"e2",  x"55",  x"94",  x"db",  x"30",  x"73",  x"c3",  x"62", -- 1248
         x"9d",  x"dd",  x"62",  x"71",  x"e7",  x"70",  x"ab",  x"bd", -- 1250
         x"5c",  x"06",  x"f7",  x"5b",  x"f1",  x"e9",  x"e3",  x"eb", -- 1258
         x"91",  x"39",  x"bd",  x"3c",  x"28",  x"8b",  x"9a",  x"cd", -- 1260
         x"bd",  x"c1",  x"4a",  x"d5",  x"20",  x"4e",  x"66",  x"e9", -- 1268
         x"99",  x"13",  x"d3",  x"98",  x"32",  x"13",  x"52",  x"54", -- 1270
         x"9b",  x"ce",  x"f9",  x"fd",  x"e8",  x"c5",  x"62",  x"a5", -- 1278
         x"c1",  x"a6",  x"c2",  x"4a",  x"3c",  x"9b",  x"ac",  x"11", -- 1280
         x"0e",  x"19",  x"cb",  x"48",  x"66",  x"d0",  x"c8",  x"2a", -- 1288
         x"85",  x"a5",  x"2b",  x"fc",  x"95",  x"f8",  x"70",  x"d3", -- 1290
         x"72",  x"73",  x"a3",  x"74",  x"60",  x"f7",  x"a5",  x"f6", -- 1298
         x"30",  x"dd",  x"5e",  x"a2",  x"09",  x"56",  x"ff",  x"21", -- 12A0
         x"02",  x"ec",  x"c1",  x"18",  x"88",  x"8d",  x"ba",  x"6a", -- 12A8
         x"19",  x"04",  x"e5",  x"21",  x"fe",  x"01",  x"e5",  x"a0", -- 12B0
         x"bb",  x"e5",  x"8e",  x"c8",  x"e8",  x"c5",  x"f2",  x"ba", -- 12B8
         x"db",  x"3c",  x"3b",  x"9e",  x"4d",  x"1a",  x"5e",  x"05", -- 12C0
         x"c7",  x"ce",  x"d3",  x"16",  x"66",  x"99",  x"2e",  x"55", -- 12C8
         x"f0",  x"85",  x"7c",  x"d6",  x"aa",  x"29",  x"19",  x"02", -- 12D0
         x"19",  x"d5",  x"64",  x"4b",  x"2e",  x"36",  x"10",  x"b0", -- 12D8
         x"4a",  x"d1",  x"c1",  x"4c",  x"12",  x"40",  x"46",  x"d3", -- 12E0
         x"fb",  x"40",  x"02",  x"41",  x"20",  x"03",  x"6f",  x"18", -- 12E8
         x"41",  x"54",  x"3e",  x"52",  x"13",  x"dc",  x"3e",  x"9c", -- 12F0
         x"c5",  x"3a",  x"3e",  x"02",  x"d4",  x"8b",  x"d5",  x"05", -- 12F8
         x"be",  x"16",  x"d7",  x"c4",  x"ec",  x"b2",  x"fa",  x"4a", -- 1300
         x"21",  x"21",  x"04",  x"02",  x"cd",  x"9b",  x"8f",  x"7d", -- 1308
         x"0f",  x"30",  x"c0",  x"a5",  x"7d",  x"a2",  x"62",  x"af", -- 1310
         x"fa",  x"c2",  x"db",  x"02",  x"c3",  x"02",  x"c4",  x"02", -- 1318
         x"56",  x"c5",  x"e0",  x"a5",  x"39",  x"ca",  x"27",  x"eb", -- 1320
         x"37",  x"df",  x"7d",  x"03",  x"b2",  x"65",  x"68",  x"9d", -- 1328
         x"32",  x"cf",  x"55",  x"43",  x"eb",  x"8a",  x"9d",  x"57", -- 1330
         x"7a",  x"e3",  x"6c",  x"68",  x"ff",  x"b3",  x"2a",  x"46", -- 1338
         x"ff",  x"a8",  x"07",  x"10",  x"26",  x"e3",  x"61",  x"b3", -- 1340
         x"3a",  x"32",  x"c5",  x"34",  x"9d",  x"16",  x"28",  x"90", -- 1348
         x"49",  x"3c",  x"49",  x"b8",  x"7e",  x"a2",  x"0d",  x"32", -- 1350
         x"d3",  x"ed",  x"bb",  x"39",  x"fa",  x"dd",  x"52",  x"98", -- 1358
         x"de",  x"25",  x"c4",  x"25",  x"85",  x"7b",  x"06",  x"c2", -- 1360
         x"06",  x"44",  x"c3",  x"2b",  x"7b",  x"7a",  x"8a",  x"ef", -- 1368
         x"b0",  x"f0",  x"ad",  x"58",  x"7a",  x"f6",  x"aa",  x"06", -- 1370
         x"08",  x"62",  x"c7",  x"50",  x"24",  x"a2",  x"91",  x"0d", -- 1378
         x"e5",  x"f1",  x"35",  x"c5",  x"a6",  x"72",  x"38",  x"32", -- 1380
         x"dc",  x"6f",  x"45",  x"74",  x"67",  x"33",  x"ce",  x"11", -- 1388
         x"a6",  x"0b",  x"f3",  x"92",  x"20",  x"13",  x"d3",  x"17", -- 1390
         x"17",  x"c5",  x"17",  x"fa",  x"9c",  x"23",  x"48",  x"dd", -- 1398
         x"54",  x"f8",  x"bf",  x"d4",  x"c7",  x"28",  x"fa",  x"03", -- 13A0
         x"fb",  x"00",  x"9a",  x"81",  x"bc",  x"06",  x"15",  x"66", -- 13A8
         x"f9",  x"f0",  x"66",  x"e6",  x"28",  x"53",  x"a8",  x"9d", -- 13B0
         x"2a",  x"bc",  x"58",  x"be",  x"b0",  x"f0",  x"96",  x"73", -- 13B8
         x"66",  x"c0",  x"e7",  x"c1",  x"92",  x"f1",  x"bb",  x"1e", -- 13C0
         x"f1",  x"a6",  x"f9",  x"05",  x"f8",  x"2b",  x"c6",  x"0a", -- 13C8
         x"c4",  x"6a",  x"d4",  x"6c",  x"b1",  x"49",  x"f7",  x"e5", -- 13D0
         x"bd",  x"58",  x"e7",  x"56",  x"e1",  x"ec",  x"aa",  x"e1", -- 13D8
         x"6d",  x"c8",  x"9b",  x"7e",  x"c2",  x"53",  x"81",  x"a1", -- 13E0
         x"14",  x"c3",  x"88",  x"90",  x"23",  x"c4",  x"8d",  x"4f", -- 13E8
         x"04",  x"1e",  x"c5",  x"8c",  x"47",  x"27",  x"33",  x"66", -- 13F0
         x"44",  x"f7",  x"7e",  x"9c",  x"45",  x"02",  x"ae",  x"96", -- 13F8
         x"99",  x"45",  x"f5",  x"35",  x"a3",  x"f8",  x"06",  x"11", -- 1400
         x"66",  x"f5",  x"77",  x"ba",  x"1d",  x"71",  x"4c",  x"f2", -- 1408
         x"1d",  x"f3",  x"94",  x"e5",  x"69",  x"ab",  x"fc",  x"08", -- 1410
         x"13",  x"66",  x"f3",  x"a9",  x"43",  x"1e",  x"83",  x"30", -- 1418
         x"f8",  x"09",  x"7b",  x"b2",  x"c1",  x"f8",  x"13",  x"14", -- 1420
         x"f8",  x"14",  x"33",  x"fd",  x"62",  x"66",  x"b3",  x"6e", -- 1428
         x"cc",  x"b6",  x"74",  x"ee",  x"c1",  x"d1",  x"ef",  x"82", -- 1430
         x"ef",  x"f0",  x"80",  x"f3",  x"f1",  x"00",  x"ae",  x"fb", -- 1438
         x"2b",  x"ee",  x"6f",  x"fc",  x"9d",  x"ef",  x"bb",  x"e5", -- 1440
         x"04",  x"f0",  x"4f",  x"78",  x"82",  x"f1",  x"47",  x"7d", -- 1448
         x"d9",  x"13",  x"be",  x"6b",  x"ee",  x"7c",  x"b6",  x"0b", -- 1450
         x"bf",  x"06",  x"ef",  x"21",  x"9e",  x"6a",  x"c0",  x"06", -- 1458
         x"f0",  x"23",  x"69",  x"c1",  x"06",  x"f1",  x"71",  x"77", -- 1460
         x"c5",  x"3b",  x"66",  x"06",  x"e3",  x"02",  x"3c",  x"cb", -- 1468
         x"1b",  x"10",  x"fa",  x"01",  x"c0",  x"e3",  x"ee",  x"93", -- 1470
         x"ac",  x"2f",  x"06",  x"ef",  x"9c",  x"ac",  x"2f",  x"06", -- 1478
         x"f0",  x"99",  x"ac",  x"2f",  x"06",  x"f1",  x"98",  x"92", -- 1480
         x"2f",  x"c1",  x"c7",  x"5e",  x"cc",  x"94",  x"87",  x"eb", -- 1488
         x"e5",  x"0d",  x"17",  x"66",  x"f1",  x"0e",  x"a8",  x"2c", -- 1490
         x"66",  x"68",  x"ef",  x"e4",  x"5f",  x"90",  x"df",  x"58", -- 1498
         x"7d",  x"ff",  x"14",  x"6f",  x"7c",  x"a5",  x"0a",  x"7b", -- 14A0
         x"c5",  x"85",  x"7a",  x"1e",  x"b3",  x"db",  x"4d",  x"06", -- 14A8
         x"52",  x"4e",  x"88",  x"e4",  x"46",  x"f9",  x"fd",  x"4b", -- 14B0
         x"09",  x"f4",  x"40",  x"fd",  x"73",  x"02",  x"fd",  x"72", -- 14B8
         x"60",  x"03",  x"15",  x"7d",  x"d6",  x"f7",  x"7c",  x"de", -- 14C0
         x"19",  x"0f",  x"7b",  x"de",  x"db",  x"61",  x"02",  x"30", -- 14C8
         x"02",  x"06",  x"01",  x"22",  x"0f",  x"ff",  x"5a",  x"0f", -- 14D0
         x"87",  x"b6",  x"4f",  x"0f",  x"f8",  x"88",  x"1f",  x"19", -- 14D8
         x"38",  x"06",  x"79",  x"9b",  x"ed",  x"23",  x"02",  x"05", -- 14E0
         x"20",  x"9c",  x"05",  x"03",  x"78",  x"05",  x"c7",  x"d7", -- 14E8
         x"21",  x"dc",  x"48",  x"f5",  x"2b",  x"0e",  x"b3",  x"09", -- 14F0
         x"44",  x"d7",  x"ef",  x"78",  x"a4",  x"81",  x"58",  x"31", -- 14F8
         x"b2",  x"a4",  x"1f",  x"8a",  x"24",  x"ff",  x"a4",  x"8a", -- 1500
         x"5e",  x"c2",  x"0a",  x"56",  x"f5",  x"21",  x"2c",  x"25", -- 1508
         x"c2",  x"32",  x"2f",  x"56",  x"ef",  x"e4",  x"0f",  x"0e", -- 1510
         x"36",  x"18",  x"43",  x"10",  x"f6",  x"10",  x"f7",  x"8a", -- 1518
         x"20",  x"3c",  x"7e",  x"ea",  x"b6",  x"a1",  x"ba",  x"cf", -- 1520
         x"05",  x"7e",  x"eb",  x"b9",  x"28",  x"bc",  x"73",  x"05", -- 1528
         x"7e",  x"ec",  x"08",  x"a1",  x"be",  x"ce",  x"05",  x"7e", -- 1530
         x"ed",  x"08",  x"85",  x"c0",  x"ed",  x"1c",  x"44",  x"fd", -- 1538
         x"a9",  x"96",  x"de",  x"12",  x"f8",  x"12",  x"ec",  x"09", -- 1540
         x"19",  x"4e",  x"97",  x"5b",  x"88",  x"da",  x"ec",  x"54", -- 1548
         x"49",  x"7b",  x"a9",  x"47",  x"78",  x"53",  x"45",  x"7c", -- 1550
         x"4c",  x"43",  x"84",  x"4a",  x"56",  x"84",  x"25",  x"3a", -- 1558
         x"95",  x"84",  x"9e",  x"e8",  x"7b",  x"83",  x"51",  x"5f", -- 1560
         x"77",  x"8a",  x"57",  x"45",  x"73",  x"8c",  x"67",  x"18", -- 1568
         x"6f",  x"8d",  x"6f",  x"b7",  x"e2",  x"bd",  x"72",  x"c5", -- 1570
         x"bd",  x"74",  x"89",  x"bd",  x"75",  x"03",  x"28",  x"f8", -- 1578
         x"37",  x"23",  x"9c",  x"95",  x"08",  x"22",  x"bc",  x"ac", -- 1580
         x"76",  x"ac",  x"94",  x"21",  x"ba",  x"c3",  x"e6",  x"ed", -- 1588
         x"4b",  x"17",  x"78",  x"50",  x"b1",  x"ab",  x"81",  x"05", -- 1590
         x"c3",  x"74",  x"a3",  x"21",  x"01",  x"1b",  x"f8",  x"5d", -- 1598
         x"3b",  x"86",  x"b6",  x"11",  x"fc",  x"c3",  x"11",  x"fd", -- 15A0
         x"eb",  x"13",  x"13",  x"ef",  x"7b",  x"0c",  x"6c",  x"fa", -- 15A8
         x"0c",  x"fb",  x"6c",  x"fa",  x"12",  x"a3",  x"f0",  x"2b", -- 15B0
         x"fb",  x"12",  x"48",  x"8a",  x"16",  x"d5",  x"ff",  x"9e", -- 15B8
         x"2c",  x"23",  x"6e",  x"78",  x"fd",  x"19",  x"1c",  x"75", -- 15C0
         x"fb",  x"c5",  x"4d",  x"d5",  x"d3",  x"1a",  x"93",  x"cc", -- 15C8
         x"e0",  x"a2",  x"cd",  x"66",  x"9c",  x"88",  x"f6",  x"d1", -- 15D0
         x"c1",  x"d8",  x"bc",  x"20",  x"74",  x"64",  x"1a",  x"a4", -- 15D8
         x"09",  x"a0",  x"30",  x"fd",  x"cb",  x"0b",  x"66",  x"df", -- 15E0
         x"c7",  x"f0",  x"91",  x"18",  x"63",  x"21",  x"ed",  x"fd", -- 15E8
         x"ef",  x"10",  x"e4",  x"c2",  x"04",  x"15",  x"dc",  x"b6", -- 15F0
         x"32",  x"e1",  x"95",  x"e1",  x"b9",  x"40",  x"3d",  x"dc", -- 15F8
         x"31",  x"d1",  x"bd",  x"60",  x"1a",  x"e1",  x"09",  x"3b", -- 1600
         x"21",  x"1c",  x"97",  x"b1",  x"b5",  x"d9",  x"d0",  x"2b", -- 1608
         x"de",  x"b4",  x"f0",  x"1a",  x"11",  x"73",  x"60",  x"f3", -- 1610
         x"38",  x"21",  x"16",  x"4b",  x"ac",  x"ad",  x"90",  x"c3", -- 1618
         x"11",  x"01",  x"e0",  x"f6",  x"da",  x"bd",  x"92",  x"b6", -- 1620
         x"d6",  x"5b",  x"dc",  x"d6",  x"6c",  x"26",  x"2a",  x"81", -- 1628
         x"51",  x"e3",  x"9f",  x"b6",  x"11",  x"f4",  x"98",  x"0f", -- 1630
         x"db",  x"dd",  x"b6",  x"48",  x"da",  x"9c",  x"26",  x"22", -- 1638
         x"a7",  x"0c",  x"da",  x"2e",  x"c6",  x"01",  x"af",  x"79", -- 1640
         x"14",  x"be",  x"cd",  x"48",  x"ff",  x"35",  x"0f",  x"38", -- 1648
         x"1e",  x"04",  x"60",  x"1e",  x"c0",  x"11",  x"4f",  x"1a", -- 1650
         x"d8",  x"eb",  x"56",  x"2b",  x"5e",  x"16",  x"88",  x"ca", -- 1658
         x"2b",  x"fb",  x"c3",  x"c4",  x"f2",  x"2c",  x"0c",  x"56", -- 1660
         x"fb",  x"b1",  x"c1",  x"4c",  x"eb",  x"ca",  x"14",  x"88", -- 1668
         x"c5",  x"f6",  x"4f",  x"29",  x"e4",  x"f7",  x"47",  x"4c", -- 1670
         x"83",  x"f8",  x"d7",  x"88",  x"04",  x"24",  x"f9",  x"67", -- 1678
         x"be",  x"d4",  x"f6",  x"9b",  x"be",  x"80",  x"fe",  x"36", -- 1680
         x"f8",  x"00",  x"b8",  x"ac",  x"bb",  x"27",  x"26",  x"b5", -- 1688
         x"25",  x"7c",  x"36",  x"24",  x"30",  x"22",  x"71",  x"02", -- 1690
         x"70",  x"5a",  x"07",  x"63",  x"22",  x"e5",  x"2d",  x"63", -- 1698
         x"fb",  x"2f",  x"0f",  x"ca",  x"4e",  x"0d",  x"d2",  x"c8", -- 16A0
         x"d2",  x"0b",  x"f2",  x"2d",  x"0b",  x"f3",  x"27",  x"26", -- 16A8
         x"6d",  x"9f",  x"2a",  x"27",  x"f1",  x"c0",  x"f4",  x"b6", -- 16B0
         x"04",  x"29",  x"d6",  x"01",  x"bf",  x"6d",  x"bc",  x"bc", -- 16B8
         x"6b",  x"0d",  x"06",  x"ca",  x"26",  x"20",  x"a7",  x"a0", -- 16C0
         x"04",  x"11",  x"4a",  x"da",  x"00",  x"eb",  x"b7",  x"c2", -- 16C8
         x"f9",  x"a5",  x"dd",  x"cb",  x"2a",  x"ec",  x"46",  x"06", -- 16D0
         x"95",  x"9a",  x"eb",  x"e8",  x"1e",  x"d4",  x"4e",  x"d0", -- 16D8
         x"8a",  x"46",  x"ee",  x"03",  x"f1",  x"3e",  x"09",  x"cb", -- 16E0
         x"38",  x"cb",  x"99",  x"e6",  x"1a",  x"89",  x"9d",  x"b3", -- 16E8
         x"a5",  x"f5",  x"9b",  x"4c",  x"8b",  x"8c",  x"66",  x"25", -- 16F0
         x"b3",  x"98",  x"e7",  x"b0",  x"28",  x"e8",  x"b4",  x"14", -- 16F8
         x"e9",  x"03",  x"ea",  x"e0",  x"96",  x"dd",  x"a6",  x"6f", -- 1700
         x"e7",  x"e4",  x"99",  x"04",  x"e8",  x"79",  x"03",  x"e9", -- 1708
         x"78",  x"b3",  x"03",  x"ea",  x"1f",  x"de",  x"7c",  x"53", -- 1710
         x"7b",  x"9f",  x"53",  x"be",  x"fb",  x"73",  x"48",  x"b6", -- 1718
         x"4e",  x"09",  x"b6",  x"eb",  x"20",  x"1f",  x"5d",  x"b0", -- 1720
         x"11",  x"9a",  x"85",  x"19",  x"a9",  x"9e",  x"e1",  x"74", -- 1728
         x"a3",  x"e2",  x"b5",  x"04",  x"e3",  x"89",  x"04",  x"e4", -- 1730
         x"18",  x"3d",  x"95",  x"f2",  x"0d",  x"38",  x"97",  x"6d", -- 1738
         x"2e",  x"e9",  x"2e",  x"ea",  x"47",  x"d9",  x"99",  x"6b", -- 1740
         x"66",  x"e8",  x"b0",  x"95",  x"9a",  x"92",  x"af",  x"4d", -- 1748
         x"72",  x"5a",  x"73",  x"99",  x"15",  x"74",  x"e8",  x"b1", -- 1750
         x"8a",  x"e7",  x"21",  x"07",  x"28",  x"b9",  x"2d",  x"19", -- 1758
         x"2c",  x"3e",  x"b0",  x"18",  x"be",  x"e1",  x"e8",  x"62", -- 1760
         x"b5",  x"e2",  x"b5",  x"04",  x"e3",  x"89",  x"04",  x"e4", -- 1768
         x"38",  x"0d",  x"4b",  x"b9",  x"dc",  x"4e",  x"c7",  x"ec", -- 1770
         x"d6",  x"a5",  x"5f",  x"4d",  x"07",  x"31",  x"2b",  x"92", -- 1778
         x"51",  x"c2",  x"28",  x"23",  x"ca",  x"b4",  x"92",  x"1f", -- 1780
         x"cd",  x"43",  x"95",  x"5f",  x"d8",  x"62",  x"b4",  x"b5", -- 1788
         x"20",  x"38",  x"35",  x"7e",  x"de",  x"c2",  x"9d",  x"30", -- 1790
         x"ed",  x"39",  x"c3",  x"14",  x"86",  x"e7",  x"47",  x"ae", -- 1798
         x"ce",  x"e8",  x"d2",  x"76",  x"04",  x"e9",  x"ce",  x"59", -- 17A0
         x"04",  x"ea",  x"57",  x"2c",  x"fd",  x"2a",  x"70",  x"f5", -- 17A8
         x"ba",  x"f9",  x"4a",  x"72",  x"8b",  x"b3",  x"36",  x"ec", -- 17B0
         x"b2",  x"02",  x"e7",  x"7b",  x"e6",  x"8d",  x"cd",  x"e8", -- 17B8
         x"f3",  x"ad",  x"96",  x"46",  x"1d",  x"77",  x"df",  x"3e", -- 17C0
         x"91",  x"9a",  x"9e",  x"e8",  x"07",  x"e0",  x"cc",  x"80", -- 17C8
         x"96",  x"df",  x"b2",  x"94",  x"09",  x"9e",  x"e0",  x"30", -- 17D0
         x"0c",  x"0e",  x"8e",  x"ed",  x"0d",  x"19",  x"5e",  x"91", -- 17D8
         x"4b",  x"56",  x"f1",  x"64",  x"9f",  x"ef",  x"d5",  x"c9", -- 17E0
         x"0a",  x"a8",  x"79",  x"e5",  x"7d",  x"e6",  x"00",  x"53", -- 17E8
         x"18",  x"2b",  x"dc",  x"25",  x"6d",  x"e5",  x"05",  x"dd", -- 17F0
         x"05",  x"e6",  x"e4",  x"6a",  x"34",  x"66",  x"e0",  x"e3", -- 17F8
         x"a3",  x"b5",  x"06",  x"ed",  x"06",  x"ee",  x"35",  x"06", -- 1800
         x"eb",  x"06",  x"ec",  x"62",  x"06",  x"02",  x"66",  x"e6", -- 1808
         x"e5",  x"37",  x"d2",  x"63",  x"c6",  x"92",  x"ce",  x"8a", -- 1810
         x"28",  x"f2",  x"58",  x"66",  x"4e",  x"6e",  x"e0",  x"11", -- 1818
         x"b7",  x"f2",  x"2b",  x"e7",  x"84",  x"d1",  x"06",  x"e8", -- 1820
         x"8d",  x"47",  x"04",  x"e9",  x"53",  x"8b",  x"fc",  x"b7", -- 1828
         x"ea",  x"fc",  x"94",  x"d6",  x"2b",  x"d7",  x"2c",  x"e3", -- 1830
         x"2c",  x"84",  x"1d",  x"86",  x"2c",  x"ae",  x"d9",  x"87", -- 1838
         x"05",  x"8e",  x"e0",  x"2c",  x"dc",  x"c0",  x"d0",  x"77", -- 1840
         x"4a",  x"06",  x"d3",  x"1a",  x"08",  x"07",  x"55",  x"de", -- 1848
         x"5c",  x"56",  x"f0",  x"65",  x"2a",  x"57",  x"7c",  x"25", -- 1850
         x"26",  x"5f",  x"12",  x"ac",  x"db",  x"11",  x"c3",  x"8f", -- 1858
         x"a4",  x"ec",  x"ad",  x"d1",  x"a6",  x"ad",  x"a6",  x"a1", -- 1860
         x"65",  x"7c",  x"81",  x"9b",  x"39",  x"36",  x"fd",  x"88", -- 1868
         x"12",  x"c8",  x"a7",  x"37",  x"bb",  x"30",  x"6c",  x"bb", -- 1870
         x"ff",  x"97",  x"b5",  x"e5",  x"9a",  x"81",  x"45",  x"4c", -- 1878
         x"78",  x"c2",  x"94",  x"79",  x"48",  x"92",  x"38",  x"5d", -- 1880
         x"54",  x"83",  x"62",  x"4e",  x"72",  x"46",  x"07",  x"c5", -- 1888
         x"6e",  x"a3",  x"9e",  x"82",  x"33",  x"a1",  x"54",  x"fd", -- 1890
         x"84",  x"2a",  x"43",  x"84",  x"13",  x"2b",  x"c2",  x"84", -- 1898
         x"1e",  x"ed",  x"85",  x"04",  x"36",  x"b8",  x"f9",  x"b1", -- 18A0
         x"70",  x"82",  x"4d",  x"26",  x"44",  x"e1",  x"d0",  x"07", -- 18A8
         x"18",  x"6a",  x"b6",  x"74",  x"03",  x"1b",  x"fd",  x"34", -- 18B0
         x"0e",  x"9c",  x"49",  x"69",  x"96",  x"55",  x"f1",  x"46", -- 18B8
         x"c4",  x"ee",  x"60",  x"a8",  x"22",  x"d2",  x"67",  x"cd", -- 18C0
         x"d7",  x"81",  x"05",  x"18",  x"65",  x"86",  x"9a",  x"3b", -- 18C8
         x"56",  x"05",  x"05",  x"4b",  x"42",  x"03",  x"03",  x"84", -- 18D0
         x"9c",  x"d3",  x"d6",  x"bd",  x"6a",  x"02",  x"4d",  x"69", -- 18D8
         x"02",  x"2a",  x"f6",  x"e0",  x"d2",  x"d5",  x"b2",  x"4d", -- 18E0
         x"18",  x"39",  x"c3",  x"b3",  x"7a",  x"a2",  x"7c",  x"ad", -- 18E8
         x"99",  x"49",  x"a7",  x"ac",  x"9c",  x"28",  x"01",  x"6f", -- 18F0
         x"a8",  x"1b",  x"20",  x"65",  x"06",  x"73",  x"73",  x"07", -- 18F8
         x"9b",  x"94",  x"19",  x"55",  x"9b",  x"bf",  x"13",  x"48", -- 1900
         x"d8",  x"cd",  x"6a",  x"97",  x"4b",  x"f1",  x"23",  x"20", -- 1908
         x"82",  x"00",  x"c3",  x"84",  x"ad",  x"c3",  x"f6",  x"a9", -- 1910
         x"c3",  x"00",  x"9a",  x"aa",  x"c3",  x"57",  x"ab",  x"c3", -- 1918
         x"29",  x"ac",  x"04",  x"3e",  x"05",  x"cf",  x"c3",  x"0d", -- 1920
         x"85",  x"05",  x"df",  x"a8",  x"96",  x"05",  x"27",  x"a9", -- 1928
         x"05",  x"e3",  x"91",  x"05",  x"e8",  x"22",  x"11",  x"a4", -- 1930
         x"44",  x"0b",  x"bd",  x"89",  x"05",  x"2f",  x"12",  x"05", -- 1938
         x"c8",  x"24",  x"17",  x"cf",  x"0b",  x"48",  x"89",  x"05", -- 1940
         x"68",  x"91",  x"05",  x"d9",  x"22",  x"05",  x"95",  x"44", -- 1948
         x"05",  x"77",  x"89",  x"05",  x"b1",  x"03",  x"05",  x"d4", -- 1950
         x"a8",  x"21",  x"03",  x"b2",  x"00",  x"5e",  x"2b",  x"6e", -- 1958
         x"cd",  x"01",  x"36",  x"a9",  x"eb",  x"c9",  x"f1",  x"e1", -- 1960
         x"d1",  x"80",  x"bc",  x"f5",  x"cd",  x"39",  x"88",  x"0a", -- 1968
         x"27",  x"c3",  x"f7",  x"1f",  x"1f",  x"7d",  x"07",  x"9f", -- 1970
         x"e7",  x"79",  x"03",  x"e7",  x"03",  x"aa",  x"17",  x"7c", -- 1978
         x"f5",  x"17",  x"bb",  x"80",  x"97",  x"95",  x"6f",  x"9f", -- 1980
         x"06",  x"94",  x"67",  x"cb",  x"7a",  x"28",  x"09",  x"93", -- 1988
         x"0a",  x"5f",  x"9f",  x"92",  x"57",  x"34",  x"12",  x"f1", -- 1990
         x"d0",  x"47",  x"82",  x"15",  x"78",  x"c9",  x"17",  x"eb", -- 1998
         x"d0",  x"59",  x"0a",  x"89",  x"47",  x"18",  x"0a",  x"86", -- 19A0
         x"46",  x"26",  x"00",  x"54",  x"af",  x"a0",  x"80",  x"b2", -- 19A8
         x"20",  x"10",  x"06",  x"00",  x"10",  x"ed",  x"6a",  x"17", -- 19B0
         x"93",  x"30",  x"01",  x"83",  x"60",  x"3f",  x"07",  x"10", -- 19B8
         x"f6",  x"5f",  x"c9",  x"06",  x"19",  x"09",  x"7d",  x"6c", -- 19C0
         x"1c",  x"cb",  x"1d",  x"98",  x"0d",  x"ed",  x"52",  x"15", -- 19C8
         x"19",  x"3f",  x"17",  x"03",  x"10",  x"f5",  x"cb",  x"10", -- 19D0
         x"50",  x"5f",  x"88",  x"08",  x"80",  x"38",  x"cd",  x"f3", -- 19D8
         x"a8",  x"c3",  x"3e",  x"1d",  x"a9",  x"0e",  x"41",  x"70", -- 19E0
         x"8f",  x"26",  x"cd",  x"f7",  x"11",  x"95",  x"20",  x"c3", -- 19E8
         x"c5",  x"20",  x"c4",  x"1d",  x"81",  x"bb",  x"cd",  x"ef", -- 19F0
         x"73",  x"27",  x"02",  x"dc",  x"f7",  x"28",  x"45",  x"66", -- 19F8
         x"6a",  x"15",  x"06",  x"08",  x"29",  x"6d",  x"f5",  x"87", -- 1A00
         x"a8",  x"66",  x"44",  x"11",  x"4e",  x"18",  x"16",  x"16", -- 1A08
         x"21",  x"02",  x"09",  x"23",  x"d3",  x"09",  x"0c",  x"07", -- 1A10
         x"3e",  x"4d",  x"7d",  x"17",  x"9f",  x"db",  x"58",  x"03", -- 1A18
         x"57",  x"c3",  x"15",  x"4e",  x"ac",  x"a5",  x"62",  x"f5", -- 1A20
         x"f5",  x"3b",  x"89",  x"fa",  x"07",  x"6c",  x"fa",  x"fb", -- 1A28
         x"d1",  x"83",  x"19",  x"4d",  x"fd",  x"9d",  x"f9",  x"c1", -- 1A30
         x"95",  x"05",  x"67",  x"65",  x"05",  x"06",  x"5f",  x"9c", -- 1A38
         x"05",  x"07",  x"57",  x"42",  x"a5",  x"e8",  x"9e",  x"c2", -- 1A40
         x"fd",  x"44",  x"56",  x"07",  x"bb",  x"ff",  x"c6",  x"e1", -- 1A48
         x"c0",  x"6c",  x"72",  x"c0",  x"f4",  x"b1",  x"48",  x"7e", -- 1A50
         x"36",  x"08",  x"59",  x"4f",  x"2a",  x"09",  x"47",  x"69", -- 1A58
         x"05",  x"0a",  x"0a",  x"42",  x"0b",  x"67",  x"36",  x"78", -- 1A60
         x"4e",  x"c6",  x"46",  x"6d",  x"09",  x"3c",  x"0a",  x"3c", -- 1A68
         x"0b",  x"9c",  x"b4",  x"c9",  x"b0",  x"2b",  x"db",  x"66", -- 1A70
         x"b4",  x"59",  x"2b",  x"a8",  x"f1",  x"00",  x"7e",  x"a1", -- 1A78
         x"78",  x"0f",  x"af",  x"95",  x"4a",  x"33",  x"9c",  x"74", -- 1A80
         x"51",  x"9b",  x"72",  x"9a",  x"57",  x"18",  x"c9",  x"92", -- 1A88
         x"31",  x"e8",  x"0b",  x"cb",  x"40",  x"a4",  x"20",  x"31", -- 1A90
         x"44",  x"f5",  x"2f",  x"cb",  x"08",  x"26",  x"9b",  x"03", -- 1A98
         x"09",  x"16",  x"03",  x"0a",  x"03",  x"d6",  x"7d",  x"16", -- 1AA0
         x"fd",  x"bd",  x"7d",  x"af",  x"fd",  x"7d",  x"6d",  x"dc", -- 1AA8
         x"da",  x"7d",  x"cb",  x"65",  x"7d",  x"30",  x"14",  x"94", -- 1AB0
         x"2b",  x"0b",  x"3e",  x"27",  x"1e",  x"af",  x"2f",  x"03", -- 1AB8
         x"37",  x"6a",  x"1e",  x"bd",  x"1c",  x"10",  x"53",  x"18", -- 1AC0
         x"b3",  x"b9",  x"31",  x"38",  x"24",  x"31",  x"19",  x"77", -- 1AC8
         x"04",  x"31",  x"1c",  x"77",  x"05",  x"34",  x"1f",  x"ce", -- 1AD0
         x"ae",  x"0b",  x"a7",  x"ae",  x"84",  x"4e",  x"55",  x"62", -- 1AD8
         x"15",  x"c5",  x"c8",  x"20",  x"aa",  x"c1",  x"a1",  x"8a", -- 1AE0
         x"86",  x"65",  x"fa",  x"f4",  x"dd",  x"c2",  x"e2",  x"ff", -- 1AE8
         x"98",  x"e2",  x"64",  x"ab",  x"12",  x"05",  x"47",  x"38", -- 1AF0
         x"e2",  x"5a",  x"4e",  x"40",  x"46",  x"7c",  x"40",  x"ef", -- 1AF8
         x"24",  x"30",  x"6b",  x"fe",  x"30",  x"21",  x"dc",  x"1a", -- 1B00
         x"ba",  x"e9",  x"06",  x"de",  x"8a",  x"a5",  x"41",  x"e0", -- 1B08
         x"ae",  x"f6",  x"90",  x"e2",  x"6b",  x"f6",  x"8e",  x"18", -- 1B10
         x"18",  x"2c",  x"fb",  x"1f",  x"05",  x"1d",  x"ef",  x"05", -- 1B18
         x"1b",  x"05",  x"b9",  x"19",  x"86",  x"e7",  x"59",  x"90", -- 1B20
         x"d8",  x"cb",  x"c5",  x"cd",  x"4c",  x"5f",  x"f0",  x"39", -- 1B28
         x"b5",  x"10",  x"ae",  x"fe",  x"a8",  x"f2",  x"ca",  x"db", -- 1B30
         x"60",  x"44",  x"4d",  x"af",  x"6f",  x"b0",  x"d3",  x"d8", -- 1B38
         x"b6",  x"7c",  x"d5",  x"c1",  x"79",  x"29",  x"cb",  x"11", -- 1B40
         x"17",  x"66",  x"d9",  x"f7",  x"88",  x"d1",  x"03",  x"3b", -- 1B48
         x"01",  x"05",  x"b2",  x"92",  x"14",  x"36",  x"ff",  x"20", -- 1B50
         x"d7",  x"16",  x"96",  x"4b",  x"67",  x"93",  x"15",  x"04", -- 1B58
         x"12",  x"95",  x"05",  x"89",  x"91",  x"06",  x"e3",  x"03", -- 1B60
         x"13",  x"16",  x"cb",  x"20",  x"37",  x"00",  x"cb",  x"13", -- 1B68
         x"cb",  x"12",  x"cb",  x"44",  x"28",  x"02",  x"3d",  x"cb", -- 1B70
         x"c0",  x"ec",  x"74",  x"96",  x"49",  x"be",  x"15",  x"b2", -- 1B78
         x"e5",  x"0a",  x"7a",  x"8a",  x"e9",  x"18",  x"d6",  x"11", -- 1B80
         x"47",  x"12",  x"4f",  x"b5",  x"13",  x"5f",  x"a8",  x"14", -- 1B88
         x"57",  x"43",  x"c6",  x"dd",  x"54",  x"35",  x"93",  x"62", -- 1B90
         x"a6",  x"20",  x"45",  x"a5",  x"8a",  x"ce",  x"33",  x"28", -- 1B98
         x"cf",  x"74",  x"b0",  x"b0",  x"e8",  x"0a",  x"b6",  x"08", -- 1BA0
         x"20",  x"05",  x"0e",  x"23",  x"18",  x"5c",  x"45",  x"b4", -- 1BA8
         x"08",  x"75",  x"87",  x"62",  x"87",  x"ff",  x"94",  x"ea", -- 1BB0
         x"d2",  x"2b",  x"c5",  x"e5",  x"09",  x"92",  x"fd",  x"1a", -- 1BB8
         x"63",  x"96",  x"f8",  x"59",  x"39",  x"f9",  x"2e",  x"12", -- 1BC0
         x"be",  x"4a",  x"28",  x"0c",  x"05",  x"c1",  x"84",  x"fc", -- 1BC8
         x"80",  x"e4",  x"03",  x"13",  x"18",  x"5c",  x"d1",  x"bc", -- 1BD0
         x"fa",  x"0e",  x"9a",  x"ba",  x"67",  x"49",  x"25",  x"52", -- 1BD8
         x"fc",  x"a3",  x"b6",  x"bf",  x"be",  x"8c",  x"84",  x"49", -- 1BE0
         x"82",  x"8f",  x"44",  x"cf",  x"02",  x"51",  x"58",  x"0b", -- 1BE8
         x"7b",  x"b2",  x"28",  x"81",  x"6f",  x"06",  x"77",  x"23", -- 1BF0
         x"18",  x"f2",  x"34",  x"19",  x"54",  x"2a",  x"80",  x"93", -- 1BF8
         x"0a",  x"f9",  x"62",  x"e9",  x"25",  x"18",  x"f9",  x"9a", -- 1C00
         x"03",  x"1a",  x"13",  x"e6",  x"9c",  x"d4",  x"39",  x"0c", -- 1C08
         x"cd",  x"2a",  x"c1",  x"e1",  x"8d",  x"40",  x"af",  x"47", -- 1C10
         x"4f",  x"ed",  x"b1",  x"21",  x"08",  x"ff",  x"ff",  x"ed", -- 1C18
         x"42",  x"d3",  x"ac",  x"ad",  x"85",  x"74",  x"39",  x"f0", -- 1C20
         x"23",  x"4a",  x"23",  x"bb",  x"07",  x"69",  x"60",  x"09", -- 1C28
         x"5c",  x"fd",  x"21",  x"73",  x"0e",  x"14",  x"2c",  x"f7", -- 1C30
         x"84",  x"d5",  x"7e",  x"f0",  x"ae",  x"6f",  x"c5",  x"aa", -- 1C38
         x"9f",  x"e7",  x"d7",  x"d0",  x"21",  x"55",  x"5c",  x"c1", -- 1C40
         x"11",  x"b0",  x"9c",  x"2e",  x"5a",  x"38",  x"7e",  x"8e", -- 1C48
         x"97",  x"cd",  x"04",  x"fb",  x"d1",  x"6f",  x"d5",  x"27", -- 1C50
         x"47",  x"15",  x"17",  x"39",  x"85",  x"37",  x"7e",  x"fa", -- 1C58
         x"85",  x"57",  x"31",  x"81",  x"8c",  x"5f",  x"18",  x"41", -- 1C60
         x"e3",  x"9b",  x"75",  x"06",  x"b4",  x"3d",  x"fe",  x"be", -- 1C68
         x"72",  x"37",  x"c2",  x"75",  x"de",  x"9e",  x"8f",  x"a7", -- 1C70
         x"55",  x"ec",  x"70",  x"c1",  x"d1",  x"19",  x"eb",  x"eb", -- 1C78
         x"58",  x"95",  x"2d",  x"5e",  x"5e",  x"e8",  x"2c",  x"21", -- 1C80
         x"c5",  x"b4",  x"1d",  x"eb",  x"cf",  x"37",  x"e5",  x"d8", -- 1C88
         x"3b",  x"1b",  x"8a",  x"09",  x"9e",  x"0f",  x"7e",  x"47", -- 1C90
         x"6e",  x"66",  x"46",  x"fa",  x"1f",  x"48",  x"fd",  x"75", -- 1C98
         x"fa",  x"13",  x"74",  x"01",  x"50",  x"20",  x"80",  x"44", -- 1CA0
         x"cf",  x"3a",  x"34",  x"40",  x"b6",  x"19",  x"96",  x"25", -- 1CA8
         x"8b",  x"9a",  x"b0",  x"46",  x"17",  x"72",  x"77",  x"09", -- 1CB0
         x"59",  x"50",  x"0a",  x"4f",  x"70",  x"1e",  x"9a",  x"45", -- 1CB8
         x"59",  x"31",  x"4e",  x"d1",  x"be",  x"f5",  x"f6",  x"13", -- 1CC0
         x"ed",  x"fc",  x"8f",  x"e5",  x"c2",  x"f6",  x"d4",  x"c2", -- 1CC8
         x"86",  x"08",  x"6f",  x"d8",  x"d2",  x"8e",  x"09",  x"5b", -- 1CD0
         x"67",  x"d0",  x"33",  x"8e",  x"f0",  x"b6",  x"ce",  x"25", -- 1CD8
         x"8e",  x"0b",  x"f4",  x"41",  x"94",  x"8b",  x"00",  x"38", -- 1CE0
         x"00",  x"01",  x"0b",  x"00",  x"f4",  x"ae",  x"28",  x"08", -- 1CE8
         x"1c",  x"11",  x"22",  x"b2",  x"bd",  x"bf",  x"af",  x"e8", -- 1CF0
         x"40",  x"c9",  x"00",  x"20",  x"00",  x"00",  x"00",  x"00", -- 1CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
