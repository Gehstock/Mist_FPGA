library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity exerion_03 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of exerion_03 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"C0",X"F0",X"10",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"CC",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"68",X"87",X"30",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"73",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"3E",X"0F",X"3D",X"F0",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"73",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",
		X"00",X"00",X"FF",X"FF",X"3F",X"F0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"CE",X"73",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",
		X"00",X"00",X"7F",X"8F",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"AE",X"73",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",
		X"00",X"00",X"3F",X"0F",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"73",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"3C",
		X"00",X"00",X"7F",X"8F",X"3F",X"FF",X"F0",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"1E",
		X"00",X"00",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"13",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"87",
		X"00",X"00",X"3F",X"0F",X"33",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"13",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"78",X"E1",
		X"00",X"00",X"6E",X"8F",X"11",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"EF",X"13",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"F0",X"96",X"F0",
		X"00",X"00",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"01",X"00",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"88",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"01",X"00",
		X"00",X"08",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"00",X"3C",X"C3",X"F0",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F1",X"F4",X"F0",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F5",X"F6",X"F8",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FD",X"FE",X"F8",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F3",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"77",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"3B",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"1D",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"0E",X"F0",X"F0",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"10",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"77",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0F",X"F0",X"F0",X"00",X"00",X"1F",X"0F",X"0F",X"87",X"0F",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"F0",X"F0",X"00",X"00",X"2F",X"0F",X"0F",X"87",X"0F",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"3D",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"F0",X"F0",X"00",X"08",X"2F",X"0F",X"1E",X"A5",X"4B",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3D",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"F0",X"F0",X"00",X"08",X"2F",X"1E",X"3C",X"E1",X"E1",X"61",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"00",X"FF",X"FB",X"17",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"0F",X"F0",X"F0",X"00",X"08",X"6B",X"96",X"3C",X"F0",X"F4",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F0",X"00",X"00",X"00",X"FF",X"FB",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"3F",X"F0",X"F0",X"00",X"08",X"E3",X"D2",X"78",X"F0",X"F4",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"88",X"FF",X"FB",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"F0",X"F0",X"00",X"08",X"E3",X"F8",X"78",X"F4",X"F4",X"F6",
		X"00",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"00",X"00",X"88",X"FF",X"FB",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"F0",X"F0",X"00",X"08",X"E3",X"FC",X"F4",X"FD",X"FF",X"F7",
		X"00",X"00",X"00",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FB",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"00",X"08",X"E3",X"FF",X"FE",X"FD",X"F9",X"F7",
		X"00",X"00",X"00",X"E0",X"10",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FD",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"F0",X"F0",X"00",X"08",X"EB",X"FF",X"FF",X"FD",X"FD",X"FE",
		X"00",X"00",X"80",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"F0",X"F0",X"00",X"00",X"E3",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"00",X"00",X"C0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"F0",X"F0",X"00",X"00",X"F1",X"FA",X"FF",X"FE",X"FF",X"F3",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"FA",X"FA",X"FF",X"F3",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"17",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"E0",X"F8",X"F0",X"FC",X"FB",
		X"00",X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"25",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F8",X"F0",X"FC",X"F3",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"71",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F7",
		X"00",X"C0",X"00",X"80",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"73",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"FF",
		X"00",X"60",X"00",X"84",X"F0",X"34",X"00",X"0C",X"00",X"00",X"00",X"CC",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FE",
		X"00",X"60",X"00",X"A4",X"F0",X"B4",X"00",X"0E",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",
		X"00",X"30",X"00",X"A5",X"F0",X"B4",X"01",X"0F",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"30",X"80",X"A5",X"F0",X"B4",X"21",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"F1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"30",X"84",X"A5",X"F0",X"B4",X"29",X"01",X"00",X"00",X"00",X"FF",X"FF",X"43",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"80",X"10",X"A4",X"A5",X"F0",X"B4",X"2D",X"00",X"00",X"00",X"00",X"FF",X"CF",X"37",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",
		X"80",X"10",X"B4",X"A5",X"F0",X"B4",X"2D",X"00",X"00",X"00",X"00",X"FF",X"8C",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",
		X"80",X"10",X"AE",X"A5",X"F0",X"B4",X"2F",X"00",X"00",X"00",X"00",X"FF",X"3B",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",
		X"C0",X"00",X"8C",X"A7",X"F0",X"BC",X"2B",X"01",X"00",X"00",X"00",X"FF",X"7F",X"7F",X"01",X"00",
		X"00",X"00",X"00",X"00",X"2E",X"0F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"C0",X"00",X"88",X"AF",X"FF",X"BF",X"23",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"01",X"00",
		X"00",X"00",X"00",X"00",X"6E",X"0F",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"C0",X"00",X"00",X"AF",X"FF",X"BF",X"01",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"C0",X"00",X"00",X"AE",X"FF",X"BF",X"00",X"0E",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"C0",X"00",X"00",X"8C",X"FF",X"37",X"00",X"0C",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"60",X"00",X"00",X"88",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"CC",X"F7",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",
		X"60",X"00",X"00",X"00",X"00",X"F0",X"10",X"0E",X"00",X"00",X"00",X"CC",X"F7",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"60",X"00",X"00",X"00",X"08",X"F0",X"12",X"07",X"00",X"00",X"00",X"C8",X"FB",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",
		X"60",X"00",X"00",X"00",X"48",X"F0",X"5A",X"00",X"00",X"00",X"00",X"80",X"39",X"7F",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"60",X"00",X"00",X"00",X"4A",X"F0",X"D2",X"00",X"00",X"00",X"00",X"80",X"18",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",
		X"30",X"00",X"00",X"00",X"5A",X"F0",X"D2",X"0C",X"00",X"00",X"00",X"00",X"00",X"AF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",
		X"30",X"00",X"00",X"80",X"5B",X"F0",X"DA",X"0F",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",
		X"30",X"00",X"00",X"00",X"5F",X"F0",X"DE",X"0C",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",
		X"30",X"00",X"00",X"E0",X"4E",X"FF",X"DF",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"30",X"00",X"00",X"E1",X"5C",X"FF",X"5F",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"30",X"00",X"80",X"E1",X"38",X"FF",X"13",X"07",X"00",X"00",X"B3",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",
		X"30",X"00",X"C0",X"E1",X"70",X"FF",X"51",X"0E",X"00",X"88",X"F7",X"31",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FD",
		X"30",X"00",X"C2",X"E1",X"F0",X"00",X"42",X"08",X"00",X"88",X"FF",X"31",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"F0",X"00",X"FF",X"FF",X"FF",X"FD",X"FF",X"FB",X"FD",
		X"30",X"00",X"D2",X"E1",X"F0",X"B4",X"52",X"00",X"00",X"88",X"FF",X"31",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F0",X"08",X"FF",X"FF",X"FF",X"FD",X"FF",X"F3",X"FD",
		X"30",X"80",X"D2",X"E1",X"F0",X"B4",X"52",X"00",X"00",X"88",X"FF",X"31",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"F3",X"F0",X"08",X"FF",X"FF",X"FF",X"FD",X"FF",X"F1",X"FD",
		X"30",X"84",X"D2",X"E1",X"F0",X"B4",X"52",X"0C",X"00",X"CC",X"FF",X"31",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"F3",X"F0",X"08",X"FF",X"FF",X"F5",X"F9",X"FF",X"F1",X"FD",
		X"30",X"A4",X"D2",X"E1",X"F0",X"B4",X"1E",X"0F",X"00",X"CC",X"FF",X"73",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",X"F0",X"08",X"FF",X"FF",X"F5",X"F9",X"FE",X"F1",X"FD",
		X"30",X"B4",X"D2",X"E1",X"F0",X"B4",X"1E",X"0F",X"00",X"EE",X"FF",X"73",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F3",X"F0",X"08",X"FF",X"FE",X"F1",X"F8",X"FE",X"F0",X"F8",
		X"30",X"A6",X"D2",X"E1",X"F0",X"B4",X"52",X"0C",X"00",X"EE",X"FF",X"71",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"F7",X"F0",X"08",X"F6",X"FC",X"F0",X"F0",X"FC",X"F0",X"F8",
		X"30",X"8C",X"D3",X"E1",X"F0",X"B4",X"56",X"00",X"00",X"FF",X"FF",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"F7",X"F0",X"08",X"F6",X"FC",X"F0",X"F0",X"FC",X"F0",X"F8",
		X"30",X"88",X"DF",X"E1",X"F0",X"BC",X"57",X"00",X"00",X"FF",X"F7",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"F0",X"08",X"E3",X"F8",X"96",X"F0",X"F8",X"C3",X"F0",
		X"60",X"00",X"DF",X"EF",X"FF",X"BF",X"57",X"00",X"00",X"FF",X"F3",X"17",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"F7",X"F0",X"08",X"E1",X"5A",X"4B",X"B4",X"F8",X"C3",X"D2",
		X"60",X"00",X"CE",X"EF",X"FF",X"BF",X"17",X"00",X"00",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"F7",X"F0",X"08",X"69",X"5A",X"4B",X"B4",X"F0",X"E1",X"D2",
		X"60",X"00",X"CC",X"EF",X"FF",X"BF",X"1F",X"00",X"00",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"F7",X"F0",X"08",X"69",X"0F",X"0F",X"0F",X"F0",X"B4",X"D2",
		X"60",X"00",X"88",X"EF",X"FF",X"BF",X"0C",X"03",X"00",X"FE",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"FF",X"FF",X"F7",X"F0",X"08",X"3D",X"87",X"3C",X"0F",X"87",X"B4",X"C3",
		X"60",X"00",X"00",X"EF",X"FF",X"37",X"08",X"0F",X"00",X"EC",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"08",X"1F",X"0F",X"3C",X"0F",X"0F",X"A5",X"C3",
		X"60",X"00",X"00",X"EE",X"FF",X"33",X"00",X"0F",X"00",X"EC",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"F0",X"08",X"1F",X"0F",X"96",X"4B",X"0F",X"C3",X"96",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"C8",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"78",X"1E",X"87",X"4B",X"0F",X"B4",X"96",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"E8",X"FD",X"17",X"00",X"00",X"08",X"00",
		X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"F0",X"F0",X"0F",X"4B",X"0F",X"78",X"96",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"FE",X"17",X"00",X"00",X"08",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"F0",X"A5",X"F0",X"0F",X"78",X"96",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"FF",X"12",X"00",X"00",X"4C",X"00",
		X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"A5",X"F0",X"0F",X"78",X"3C",
		X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"FF",X"10",X"00",X"00",X"CC",X"01",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"80",X"F0",X"5A",X"69",X"78",
		X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"FF",X"10",X"00",X"00",X"CC",X"01",
		X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"00",X"C0",X"F0",X"1E",X"69",
		X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"F7",X"00",X"00",X"00",X"EE",X"13",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"00",X"00",X"E0",X"1E",X"69",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F3",X"00",X"00",X"00",X"EE",X"13",
		X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"00",X"00",X"80",X"1E",X"4B",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"00",X"00",X"00",X"FF",X"13",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"87",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"37",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"1E",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",
		X"0E",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"3C",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"F0",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",
		X"0C",X"0F",X"8F",X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"78",
		X"00",X"C0",X"00",X"00",X"00",X"78",X"F0",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",
		X"08",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",
		X"00",X"80",X"10",X"00",X"78",X"78",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",
		X"00",X"0F",X"0F",X"0F",X"0F",X"EF",X"FF",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",
		X"00",X"80",X"10",X"00",X"7F",X"7F",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",
		X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"CF",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"30",X"00",X"00",X"7F",X"FF",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",
		X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"60",X"00",X"00",X"00",X"FF",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",
		X"00",X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"17",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"21",
		X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"71",
		X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"E0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"71",
		X"00",X"00",X"08",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",
		X"00",X"00",X"00",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"88",X"FF",X"73",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"00",X"00",X"13",X"00",X"00",X"88",X"FF",X"F3",
		X"00",X"00",X"00",X"0E",X"0F",X"0F",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"E1",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"37",X"00",X"00",X"88",X"FF",X"F7",
		X"00",X"00",X"00",X"0C",X"0F",X"0F",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"E9",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F0",X"00",X"00",X"37",X"00",X"00",X"88",X"FF",X"F7",
		X"00",X"00",X"00",X"08",X"0F",X"0F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"E9",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"88",X"37",X"00",X"00",X"00",X"FD",X"F7",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"ED",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"37",X"00",X"00",X"00",X"EC",X"F7",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"EF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"3F",X"00",X"00",X"00",X"E8",X"73",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",X"00",X"00",X"00",X"C0",X"70",
		X"00",X"00",X"00",X"00",X"08",X"0F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F3",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",
		X"00",X"00",X"E0",X"30",X"F0",X"90",X"F0",X"70",X"00",X"88",X"F5",X"12",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"3C",
		X"00",X"00",X"E0",X"B4",X"F0",X"96",X"F0",X"78",X"00",X"88",X"FF",X"12",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"1E",
		X"00",X"30",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"00",X"88",X"FF",X"71",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"87",
		X"80",X"3C",X"E1",X"B4",X"F0",X"F0",X"F0",X"78",X"00",X"CC",X"FF",X"71",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"78",X"E1",
		X"C0",X"3C",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"00",X"CC",X"FF",X"73",X"00",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"F0",X"96",X"F0",
		X"C0",X"3C",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"00",X"CE",X"FF",X"73",X"00",X"00",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"3C",X"E1",X"B4",X"F0",X"F0",X"F0",X"78",X"00",X"CE",X"FF",X"73",X"00",X"88",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"3C",X"C3",X"F0",X"F9",
		X"C0",X"3C",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"00",X"CE",X"FF",X"73",X"00",X"88",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F1",X"F4",X"F0",X"F9",
		X"C4",X"3C",X"E1",X"BC",X"FF",X"97",X"F0",X"78",X"00",X"8E",X"FF",X"73",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F5",X"F6",X"F8",X"FF",
		X"CC",X"3C",X"E1",X"BC",X"FF",X"F9",X"FF",X"7F",X"00",X"8E",X"FF",X"43",X"00",X"88",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FD",X"FE",X"F8",X"7F",
		X"CC",X"3F",X"EF",X"BF",X"FF",X"9F",X"FF",X"7F",X"00",X"0C",X"FF",X"37",X"00",X"88",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F3",X"7F",
		X"88",X"3F",X"EF",X"BF",X"FF",X"9F",X"FF",X"7F",X"00",X"0C",X"FF",X"7F",X"00",X"CC",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",
		X"00",X"33",X"EF",X"BF",X"FF",X"F9",X"FF",X"7F",X"00",X"08",X"6F",X"7F",X"00",X"CC",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"08",X"E1",X"F0",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"1F",
		X"00",X"00",X"EE",X"BF",X"FF",X"9F",X"FF",X"7F",X"00",X"00",X"8F",X"7F",X"00",X"CC",X"5F",X"10",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"0F",
		X"00",X"00",X"EE",X"33",X"FF",X"99",X"FF",X"77",X"00",X"00",X"CC",X"7F",X"00",X"CC",X"BF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"0F",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"88",X"CC",X"3F",X"00",X"88",X"EF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"88",X"88",X"37",X"00",X"88",X"C7",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0F",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"CC",X"98",X"17",X"00",X"00",X"C1",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"CC",X"10",X"07",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"CC",X"31",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"87",
		X"00",X"00",X"C0",X"F0",X"AE",X"C0",X"10",X"F0",X"00",X"EE",X"31",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0F",X"0F",X"0F",X"C3",X"00",X"00",X"1F",X"0F",X"0F",X"87",X"0F",X"87",
		X"00",X"00",X"E0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"EE",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"87",X"00",X"00",X"2F",X"0F",X"0F",X"87",X"0F",X"C3",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"E6",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"0F",X"0F",X"FF",X"F7",X"00",X"08",X"2F",X"0F",X"1E",X"A5",X"4B",X"C3",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"1E",X"F0",X"00",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"FF",X"FF",X"F7",X"00",X"08",X"2F",X"1E",X"3C",X"E1",X"E1",X"E1",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"8F",X"FF",X"FF",X"FF",X"F7",X"00",X"08",X"6B",X"96",X"3C",X"F0",X"F0",X"E1",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"08",X"E3",X"D2",X"78",X"F0",X"F0",X"E1",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"1E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"08",X"E3",X"F0",X"78",X"F0",X"F0",X"F0",
		X"00",X"00",X"F3",X"F0",X"EF",X"D3",X"5A",X"FF",X"00",X"00",X"00",X"00",X"22",X"01",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"F1",X"00",X"08",X"E3",X"FF",X"F7",X"F0",X"FF",X"F1",
		X"00",X"00",X"EE",X"FF",X"EF",X"DF",X"5B",X"FF",X"00",X"00",X"00",X"00",X"3B",X"03",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"E3",X"F8",X"FF",X"F1",X"F8",X"F7",
		X"00",X"00",X"CC",X"FF",X"AE",X"CC",X"11",X"FF",X"00",X"00",X"00",X"88",X"3F",X"13",X"00",X"00",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"F1",X"F0",X"F8",X"F7",X"F0",X"FE",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"BF",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"F0",
		X"00",X"00",X"00",X"E0",X"F0",X"30",X"F0",X"0C",X"00",X"00",X"00",X"CC",X"FF",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F3",
		X"00",X"00",X"80",X"E1",X"F0",X"3C",X"F0",X"2E",X"00",X"00",X"00",X"CC",X"FF",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F6",
		X"00",X"00",X"E0",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"CC",X"FF",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FC",
		X"00",X"C0",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"CC",X"FF",X"37",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"80",X"D2",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"CC",X"FF",X"37",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"A4",X"D2",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"CE",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"B4",X"D2",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"CE",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"B4",X"D2",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"CE",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"B7",X"D2",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"8C",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"AE",X"D3",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"6E",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"88",X"DF",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"EE",X"CF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"CC",X"EF",X"EF",X"FF",X"3F",X"FF",X"2F",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"EE",X"EF",X"FF",X"3F",X"FF",X"2F",X"00",X"00",X"00",X"FF",X"FF",X"37",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"E0",X"98",X"EF",X"FF",X"3F",X"FF",X"2E",X"00",X"00",X"00",X"FF",X"FF",X"37",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"00",X"F0",X"70",X"EE",X"FF",X"33",X"FF",X"0C",X"00",X"00",X"00",X"FF",X"FF",X"03",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"AE",X"FF",X"FF",
		X"00",X"F0",X"F0",X"10",X"00",X"C0",X"00",X"30",X"00",X"00",X"00",X"FF",X"FF",X"73",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"6E",X"FF",X"FF",
		X"00",X"F0",X"F0",X"B4",X"F0",X"D2",X"F0",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FD",
		X"00",X"F0",X"F0",X"B4",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FD",
		X"00",X"F0",X"F0",X"B4",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"FD",X"F8",
		X"00",X"F0",X"F0",X"B4",X"F0",X"D2",X"F0",X"F0",X"00",X"00",X"00",X"EE",X"77",X"E7",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"FC",X"F8",
		X"00",X"F0",X"F0",X"B4",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"EE",X"77",X"E7",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"F4",X"F8",
		X"00",X"F1",X"F0",X"B4",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"CC",X"3B",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"F0",X"F8",
		X"00",X"F3",X"F0",X"BC",X"FF",X"D3",X"F8",X"FF",X"00",X"00",X"00",X"CC",X"BF",X"71",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"F0",X"F8",
		X"00",X"EE",X"FF",X"BF",X"FF",X"DF",X"8F",X"FF",X"00",X"00",X"00",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"F0",X"F0",
		X"00",X"CC",X"FF",X"BF",X"FF",X"DF",X"8F",X"FF",X"00",X"00",X"00",X"CC",X"FE",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"F0",X"F0",
		X"00",X"88",X"FF",X"33",X"00",X"CC",X"88",X"FF",X"00",X"00",X"00",X"88",X"F0",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"7F",X"F0",X"F0",
		X"00",X"00",X"00",X"E0",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"88",X"D0",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"6E",X"F0",X"F0",
		X"00",X"00",X"00",X"E1",X"F0",X"3C",X"00",X"0E",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"A6",X"F0",X"F0",
		X"00",X"00",X"80",X"E1",X"F0",X"3C",X"10",X"0F",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",
		X"00",X"00",X"C0",X"E1",X"F0",X"3C",X"38",X"01",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"C2",X"E1",X"F0",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",
		X"00",X"00",X"D2",X"E1",X"F0",X"3C",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"80",X"D2",X"E1",X"F0",X"3C",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"84",X"D2",X"E1",X"F0",X"3C",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"A4",X"D2",X"E1",X"F0",X"00",X"24",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"B4",X"D2",X"E1",X"70",X"F0",X"14",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"A6",X"D2",X"E1",X"38",X"F0",X"12",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",
		X"00",X"8C",X"D3",X"E1",X"58",X"F0",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F7",X"10",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",
		X"00",X"88",X"DF",X"E1",X"4A",X"F0",X"D2",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"FB",X"31",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",
		X"00",X"00",X"DF",X"67",X"5A",X"F0",X"D2",X"0C",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",X"31",
		X"00",X"00",X"00",X"88",X"FF",X"1F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"CE",X"A3",X"5B",X"F0",X"DA",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",X"31",
		X"00",X"00",X"00",X"CC",X"1F",X"0F",X"C3",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"CC",X"67",X"5F",X"F0",X"DE",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"31",
		X"00",X"00",X"00",X"08",X"0F",X"0F",X"C3",X"F0",X"00",X"00",X"CE",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"00",X"00",X"88",X"EF",X"4E",X"FF",X"DF",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"DF",X"31",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"AE",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"00",X"00",X"00",X"EF",X"5D",X"FF",X"5F",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"FF",X"30",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"E1",X"F0",X"00",X"00",X"BF",X"FB",X"F7",X"FB",X"FF",X"FB",
		X"00",X"00",X"00",X"EE",X"3B",X"FF",X"13",X"07",X"00",X"00",X"3B",X"01",X"00",X"00",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"E1",X"F0",X"00",X"00",X"B7",X"F3",X"F7",X"F1",X"FF",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"0E",X"00",X"88",X"7F",X"13",X"00",X"00",X"EE",X"01",
		X"00",X"00",X"00",X"00",X"08",X"0F",X"E1",X"F0",X"00",X"00",X"B7",X"F2",X"F5",X"F0",X"F7",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"88",X"FF",X"13",X"00",X"00",X"EE",X"01",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"00",X"00",X"B7",X"F2",X"F4",X"F0",X"F6",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"13",X"00",X"00",X"CC",X"01",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"00",X"00",X"B7",X"F0",X"F0",X"F0",X"F6",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"13",X"00",X"00",X"8C",X"01",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"F0",X"F0",X"00",X"00",X"B7",X"3C",X"E1",X"F0",X"F2",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"13",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"F0",X"00",X"00",X"A6",X"F0",X"1E",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",X"CC",X"FF",X"37",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"C2",X"F0",X"F0",X"F0",X"C3",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"02",X"E0",X"E0",X"00",X"EE",X"FF",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"3C",X"F0",
		X"00",X"00",X"00",X"00",X"80",X"30",X"E1",X"E1",X"00",X"EE",X"FF",X"17",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E1",
		X"00",X"00",X"00",X"70",X"B0",X"78",X"E1",X"E1",X"00",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"D2",
		X"00",X"08",X"80",X"78",X"B4",X"78",X"E1",X"E1",X"00",X"FF",X"7F",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"F1",X"B4",
		X"00",X"48",X"C1",X"78",X"B4",X"78",X"E1",X"E1",X"00",X"FF",X"3F",X"71",X"00",X"00",X"13",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"F7",X"F0",
		X"00",X"68",X"C3",X"7F",X"BC",X"7F",X"E1",X"EF",X"00",X"FF",X"FF",X"F3",X"00",X"88",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"F0",
		X"00",X"6E",X"CF",X"7F",X"BF",X"7F",X"EF",X"EF",X"00",X"FF",X"FF",X"F3",X"00",X"88",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"F1",
		X"00",X"4C",X"CD",X"7F",X"BF",X"7F",X"EF",X"EF",X"00",X"FF",X"FF",X"F3",X"00",X"CC",X"3F",X"00",
		X"00",X"2F",X"0F",X"0F",X"0F",X"0F",X"E1",X"F0",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"F1",
		X"00",X"08",X"88",X"7F",X"BF",X"7F",X"EF",X"EF",X"00",X"EE",X"FF",X"F3",X"00",X"CC",X"3F",X"00",
		X"00",X"4F",X"0F",X"0F",X"0F",X"0F",X"C3",X"F0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",
		X"00",X"00",X"00",X"77",X"BB",X"7F",X"EF",X"EF",X"00",X"EE",X"FF",X"F3",X"00",X"88",X"3F",X"00",
		X"00",X"8F",X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"33",X"EF",X"EF",X"00",X"8C",X"FF",X"F3",X"00",X"88",X"3F",X"00",
		X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"F7",X"F0",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"02",X"EE",X"EE",X"00",X"8E",X"DF",X"71",X"00",X"88",X"7F",X"01",
		X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"F7",X"F0",X"88",X"EF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F7",
		X"00",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",X"4E",X"EF",X"71",X"00",X"88",X"7F",X"01",
		X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"F7",X"F0",X"CC",X"EF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"FF",X"21",X"00",X"CC",X"7F",X"01",
		X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F0",X"CC",X"EF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"FF",X"01",X"00",X"CC",X"7F",X"01",
		X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F0",X"CC",X"EF",X"FF",X"F5",X"FF",X"FF",X"F9",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"FF",X"01",X"00",X"CC",X"3F",X"00",
		X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F0",X"CC",X"EF",X"FF",X"F5",X"FE",X"FF",X"F8",X"FF",
		X"00",X"00",X"00",X"80",X"F0",X"30",X"00",X"00",X"00",X"8C",X"7F",X"00",X"00",X"EE",X"3F",X"00",
		X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F0",X"CC",X"EF",X"FE",X"F1",X"FE",X"FE",X"F0",X"FF",
		X"00",X"00",X"00",X"84",X"F0",X"34",X"00",X"0C",X"00",X"08",X"3F",X"00",X"00",X"EE",X"17",X"00",
		X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F0",X"CC",X"E7",X"FC",X"F0",X"FE",X"FE",X"F0",X"FF",
		X"00",X"00",X"00",X"A4",X"F0",X"B4",X"00",X"0E",X"00",X"08",X"07",X"00",X"00",X"EE",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"CC",X"E7",X"FC",X"F0",X"FC",X"FC",X"F0",X"FF",
		X"00",X"00",X"00",X"A5",X"F0",X"B4",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"EE",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"CC",X"E3",X"F8",X"F0",X"F4",X"FC",X"F0",X"F7",
		X"00",X"00",X"80",X"A5",X"F0",X"B4",X"21",X"0F",X"00",X"00",X"00",X"00",X"00",X"EE",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"CC",X"E1",X"F0",X"F0",X"F0",X"F4",X"F0",X"F6",
		X"00",X"00",X"84",X"A5",X"F0",X"B4",X"29",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"23",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"F0",X"CC",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F6",
		X"00",X"00",X"A4",X"A5",X"F0",X"B4",X"2D",X"08",X"00",X"00",X"00",X"00",X"00",X"FF",X"63",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"CC",X"E1",X"78",X"0F",X"0F",X"F0",X"F0",X"F6",
		X"00",X"00",X"B4",X"A5",X"F0",X"B4",X"2D",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"73",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"C3",X"F0",X"CC",X"E1",X"F0",X"78",X"0F",X"87",X"F0",X"F4",
		X"00",X"00",X"AE",X"A5",X"F0",X"B4",X"2F",X"08",X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"C3",X"F0",X"CC",X"87",X"F0",X"F0",X"F0",X"0F",X"E1",X"F0",
		X"00",X"00",X"8C",X"A7",X"F0",X"BC",X"2B",X"01",X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0F",X"87",X"F0",X"CC",X"0F",X"E1",X"F0",X"F0",X"F0",X"C3",X"F0",
		X"00",X"00",X"88",X"AF",X"FF",X"BF",X"23",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"F3",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"87",X"F0",X"08",X"F0",X"1E",X"E1",X"F0",X"F0",X"B4",X"F0",
		X"00",X"00",X"00",X"AF",X"FF",X"BF",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"F3",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"F0",X"80",X"F0",X"F0",X"1E",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"AE",X"FF",X"BF",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"8C",X"FF",X"37",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"00",X"00",X"08",X"0F",X"0F",X"0F",X"C3",X"00",X"00",X"00",X"F0",X"F0",X"96",X"F0",X"F0",
		X"00",X"00",X"00",X"88",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F5",X"10",
		X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"E7",X"00",X"00",X"00",X"80",X"F0",X"78",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"CE",X"F7",X"10",
		X"00",X"00",X"00",X"0E",X"0F",X"0F",X"EF",X"F3",X"00",X"00",X"00",X"00",X"C0",X"F0",X"96",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"0E",X"00",X"00",X"00",X"00",X"00",X"8E",X"F7",X"10",
		X"00",X"00",X"00",X"0F",X"0F",X"EF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"00",X"E0",X"3C",X"E1",
		X"00",X"00",X"00",X"00",X"08",X"F0",X"12",X"07",X"00",X"00",X"00",X"00",X"00",X"8E",X"FF",X"10",
		X"00",X"00",X"08",X"0F",X"EF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"00",X"00",X"80",X"78",X"C3",
		X"00",X"00",X"00",X"00",X"48",X"F0",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"F7",X"30",
		X"00",X"00",X"0C",X"CF",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"87",
		X"00",X"00",X"00",X"00",X"4A",X"F0",X"D2",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"FB",X"31",
		X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"5A",X"F0",X"D2",X"0C",X"00",X"00",X"00",X"00",X"00",X"4C",X"FF",X"31",
		X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",
		X"00",X"00",X"00",X"00",X"5B",X"F0",X"DA",X"0F",X"00",X"00",X"00",X"00",X"00",X"4C",X"FF",X"31",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",
		X"00",X"00",X"00",X"00",X"5F",X"F0",X"DE",X"0C",X"00",X"00",X"00",X"00",X"00",X"88",X"EF",X"31",
		X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",
		X"00",X"00",X"00",X"00",X"4E",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"DF",X"31",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"4C",X"FF",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"30",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"08",X"FF",X"13",X"07",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"01",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"01",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
