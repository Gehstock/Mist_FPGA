library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_2 is
	type rom is array(0 to  6655) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"20",X"38",X"F4",X"FF",X"F8",X"FC",X"F8",X"F0",X"7E",X"30",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"18",X"60",X"01",X"03",X"03",X"03",X"03",X"01",X"60",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"C8",X"C0",X"E2",X"C0",X"C8",X"C0",X"E0",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",
		X"00",X"80",X"B0",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"B0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"31",X"31",X"61",X"61",X"61",X"31",X"31",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"6C",X"EE",X"EE",X"EE",X"EE",X"EE",X"6C",X"00",X"64",X"F6",X"A2",X"A2",X"82",X"F6",X"64",
		X"00",X"54",X"82",X"F6",X"82",X"B2",X"82",X"54",X"00",X"00",X"0C",X"0E",X"0E",X"4E",X"6C",X"00",
		X"00",X"00",X"60",X"E0",X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"00",X"44",X"60",X"61",X"20",X"20",X"20",X"60",X"64",X"E8",X"C0",X"48",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"60",X"60",X"66",X"78",X"18",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"4C",X"68",X"69",X"28",X"24",X"20",X"20",X"60",X"60",X"60",X"08",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0C",X"00",X"61",X"61",X"01",X"01",X"11",X"11",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"11",X"11",X"01",X"01",X"61",X"61",X"00",X"0C",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"61",X"61",X"01",X"01",X"61",X"61",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"10",X"10",
		X"00",X"C0",X"00",X"00",X"E0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"01",X"60",X"60",X"66",X"78",X"78",X"68",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"61",X"61",X"01",X"01",X"21",X"61",X"60",X"00",X"00",X"10",X"10",
		X"00",X"70",X"30",X"40",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"60",X"E0",X"C0",X"00",X"00",X"10",X"10",
		X"20",X"20",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"20",X"20",
		X"00",X"00",X"00",X"00",X"10",X"70",X"70",X"10",X"10",X"70",X"70",X"10",X"00",X"00",X"00",X"00",
		X"20",X"20",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"20",X"20",
		X"00",X"00",X"00",X"00",X"10",X"70",X"70",X"10",X"10",X"70",X"70",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"08",X"F1",X"FA",X"F8",X"FB",X"F8",X"F8",X"FA",X"F1",X"08",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"70",X"70",X"10",X"10",X"70",X"70",X"10",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"78",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"78",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"06",X"0F",X"01",X"01",X"07",X"07",X"01",X"01",X"0F",X"06",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"F0",X"F0",X"00",X"00",X"00",
		X"03",X"03",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"03",X"03",X"00",X"7F",X"FF",X"FD",X"FC",X"F8",X"F8",X"FC",X"FD",X"FF",X"7F",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"0F",X"7F",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"7F",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"4C",X"40",X"40",X"4C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"4C",X"40",X"40",X"4C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"50",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"90",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"24",X"00",X"00",X"10",X"20",X"00",X"10",X"00",X"00",X"08",X"20",X"10",X"40",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F8",X"D4",X"FC",X"E8",X"B8",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"3D",X"7F",X"FE",X"FF",X"FF",X"7F",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"DE",X"F4",X"EF",X"B6",X"FC",X"E8",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"1F",X"3C",X"3F",X"37",X"1A",X"0E",X"03",X"00",X"00",X"00",X"00",
		X"E0",X"10",X"04",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"04",X"18",X"E0",
		X"01",X"06",X"08",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"10",X"10",X"08",X"06",X"01",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"E0",X"18",X"04",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"04",X"18",X"E0",
		X"01",X"06",X"08",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"10",X"10",X"08",X"06",X"01",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"E0",X"18",X"04",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"04",X"18",X"E0",
		X"01",X"06",X"08",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"10",X"10",X"08",X"06",X"01",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"C0",X"20",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"08",X"10",X"10",X"20",X"C0",X"00",
		X"07",X"18",X"20",X"40",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"40",X"40",X"20",X"18",X"07",
		X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"80",X"00",X"00",X"00",
		X"18",X"26",X"41",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"40",X"41",X"26",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"10",X"10",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"F0",X"F0",X"68",X"F8",X"78",X"F8",X"D8",X"78",X"E0",X"F0",X"E0",X"80",X"00",
		X"00",X"07",X"1F",X"3F",X"3A",X"7F",X"7F",X"7F",X"7F",X"7B",X"7F",X"3E",X"3F",X"1E",X"07",X"00",
		X"00",X"E0",X"B8",X"F4",X"A8",X"1E",X"B4",X"FE",X"DA",X"BC",X"1E",X"AC",X"DC",X"F0",X"A0",X"00",
		X"00",X"00",X"07",X"0F",X"0E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0E",X"0E",X"07",X"01",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"00",X"04",X"18",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"04",X"18",X"20",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C4",X"C0",X"98",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E2",X"E4",X"E8",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"07",X"07",X"07",X"07",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"09",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"08",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"30",X"78",X"78",X"78",X"78",X"30",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"50",X"F8",X"D8",X"FC",X"F4",X"FC",X"D8",X"F8",X"F0",X"C0",X"80",X"00",X"00",
		X"8E",X"9F",X"7F",X"7F",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7F",X"BF",X"9C",
		X"80",X"40",X"C0",X"F8",X"FC",X"FC",X"FA",X"FE",X"FF",X"F7",X"FE",X"FE",X"EC",X"78",X"E0",X"C0",
		X"01",X"03",X"07",X"97",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"9F",X"0B",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"00",
		X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",
		X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"1C",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",X"00",
		X"38",X"3C",X"3E",X"3E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3E",X"3E",X"3C",X"00",
		X"70",X"78",X"7C",X"7C",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7C",X"7C",X"78",X"00",
		X"1E",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"00",
		X"3C",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",
		X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",
		X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",
		X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",
		X"03",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",
		X"07",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"00",
		X"0F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"00",
		X"00",X"00",X"78",X"FC",X"CC",X"84",X"84",X"B4",X"B4",X"B4",X"F4",X"B4",X"F4",X"F4",X"F4",X"F4",
		X"FC",X"FC",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"B4",X"BC",X"CC",X"FC",X"FC",X"78",X"00",X"00",
		X"00",X"00",X"F0",X"F8",X"98",X"08",X"08",X"68",X"68",X"68",X"E8",X"68",X"E8",X"E8",X"E8",X"E8",
		X"F8",X"F8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"68",X"78",X"98",X"F8",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"30",X"10",X"10",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"F0",X"F0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"F0",X"30",X"F0",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"60",X"20",X"20",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"E0",X"E0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"E0",X"60",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"C0",X"C0",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"02",X"02",X"02",X"02",X"02",X"03",X"02",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"02",X"02",X"03",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"03",X"07",X"06",X"04",X"04",X"05",X"05",X"05",X"07",X"05",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"05",X"05",X"06",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"0C",X"08",X"08",X"0B",X"0B",X"0B",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"0B",X"0C",X"0F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"0F",X"1F",X"19",X"10",X"10",X"16",X"16",X"16",X"1E",X"16",X"1E",X"1E",X"1E",X"1E",
		X"1F",X"1F",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"16",X"17",X"19",X"1F",X"1F",X"0F",X"00",X"00",
		X"00",X"00",X"1E",X"3F",X"33",X"21",X"21",X"2D",X"2D",X"2D",X"3D",X"2D",X"3D",X"3D",X"3D",X"3D",
		X"3F",X"3F",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"2D",X"2F",X"33",X"3F",X"3F",X"1E",X"00",X"00",
		X"00",X"00",X"3C",X"7E",X"66",X"42",X"42",X"5A",X"5A",X"5A",X"7A",X"5A",X"7A",X"7A",X"7A",X"7A",
		X"7E",X"7E",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"5A",X"5E",X"66",X"7E",X"7E",X"3C",X"00",X"00",
		X"00",X"00",X"38",X"7C",X"54",X"FE",X"EA",X"FE",X"B6",X"FE",X"EE",X"FE",X"BA",X"EE",X"FE",X"B6",
		X"B6",X"FE",X"EE",X"BA",X"FE",X"EE",X"FE",X"B6",X"FE",X"EA",X"FE",X"54",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"70",X"F8",X"A8",X"FC",X"D4",X"FC",X"6C",X"FC",X"DC",X"FC",X"74",X"DC",X"FC",X"6C",
		X"6C",X"FC",X"DC",X"74",X"FC",X"DC",X"FC",X"6C",X"FC",X"D4",X"FC",X"A8",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"50",X"F8",X"A8",X"F8",X"D8",X"F8",X"B8",X"F8",X"E8",X"B8",X"F8",X"D8",
		X"D8",X"F8",X"B8",X"E8",X"F8",X"B8",X"F8",X"D8",X"F8",X"A8",X"F8",X"50",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"A0",X"F0",X"50",X"F0",X"B0",X"F0",X"70",X"F0",X"D0",X"70",X"F0",X"B0",
		X"B0",X"F0",X"70",X"D0",X"F0",X"70",X"F0",X"B0",X"F0",X"50",X"F0",X"A0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"40",X"E0",X"A0",X"E0",X"60",X"E0",X"E0",X"E0",X"A0",X"E0",X"E0",X"60",
		X"60",X"E0",X"E0",X"A0",X"E0",X"E0",X"E0",X"60",X"E0",X"A0",X"E0",X"40",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"02",
		X"02",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"02",X"07",X"07",X"07",X"05",X"07",X"07",X"07",X"05",X"07",X"07",X"05",
		X"05",X"07",X"07",X"05",X"07",X"07",X"07",X"05",X"07",X"07",X"07",X"02",X"03",X"01",X"00",X"00",
		X"00",X"00",X"03",X"07",X"05",X"0F",X"0E",X"0F",X"0B",X"0F",X"0E",X"0F",X"0B",X"0E",X"0F",X"0B",
		X"0B",X"0F",X"0E",X"0B",X"0F",X"0E",X"0F",X"0B",X"0F",X"0E",X"0F",X"05",X"07",X"03",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"0A",X"1F",X"1D",X"1F",X"16",X"1F",X"1D",X"1F",X"17",X"1D",X"1F",X"16",
		X"16",X"1F",X"1D",X"17",X"1F",X"1D",X"1F",X"16",X"1F",X"1D",X"1F",X"0A",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"0E",X"1F",X"15",X"3F",X"3A",X"3F",X"2D",X"3F",X"3B",X"3F",X"2E",X"3B",X"3F",X"2D",
		X"2D",X"3F",X"3B",X"2E",X"3F",X"3B",X"3F",X"2D",X"3F",X"3A",X"3F",X"15",X"1F",X"0E",X"00",X"00",
		X"00",X"00",X"1C",X"3E",X"2A",X"7F",X"75",X"7F",X"5B",X"7F",X"77",X"7F",X"5D",X"77",X"7F",X"5B",
		X"5B",X"7F",X"77",X"5D",X"7F",X"77",X"7F",X"5B",X"7F",X"75",X"7F",X"2A",X"3E",X"1C",X"00",X"00",
		X"00",X"7C",X"04",X"04",X"0E",X"08",X"08",X"08",X"08",X"0C",X"08",X"0A",X"08",X"0C",X"0A",X"08",
		X"0C",X"08",X"08",X"08",X"0C",X"08",X"0A",X"08",X"0C",X"08",X"0A",X"0C",X"06",X"04",X"7C",X"00",
		X"00",X"F8",X"08",X"08",X"1C",X"10",X"10",X"10",X"10",X"18",X"10",X"14",X"10",X"18",X"14",X"10",
		X"18",X"10",X"10",X"10",X"18",X"10",X"14",X"10",X"18",X"10",X"14",X"18",X"0C",X"08",X"F8",X"00",
		X"00",X"F0",X"10",X"10",X"38",X"20",X"20",X"20",X"20",X"30",X"20",X"28",X"20",X"30",X"28",X"20",
		X"30",X"20",X"20",X"20",X"30",X"20",X"28",X"20",X"30",X"20",X"28",X"30",X"18",X"10",X"F0",X"00",
		X"00",X"E0",X"20",X"20",X"70",X"40",X"40",X"40",X"40",X"60",X"40",X"50",X"40",X"60",X"50",X"40",
		X"60",X"40",X"40",X"40",X"60",X"40",X"50",X"40",X"60",X"40",X"50",X"60",X"30",X"20",X"E0",X"00",
		X"00",X"C0",X"40",X"40",X"E0",X"80",X"80",X"80",X"80",X"C0",X"80",X"A0",X"80",X"C0",X"A0",X"80",
		X"C0",X"80",X"80",X"80",X"C0",X"80",X"A0",X"80",X"C0",X"80",X"A0",X"C0",X"60",X"40",X"C0",X"00",
		X"00",X"80",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"00",X"80",X"40",X"00",
		X"80",X"00",X"00",X"00",X"80",X"00",X"40",X"00",X"80",X"00",X"40",X"80",X"C0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"0F",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"0F",X"00",
		X"00",X"1F",X"01",X"01",X"03",X"02",X"02",X"02",X"02",X"03",X"02",X"02",X"02",X"03",X"02",X"02",
		X"03",X"02",X"02",X"02",X"03",X"02",X"02",X"02",X"03",X"02",X"02",X"03",X"01",X"01",X"1F",X"00",
		X"00",X"3E",X"02",X"02",X"07",X"04",X"04",X"04",X"04",X"06",X"04",X"05",X"04",X"06",X"05",X"04",
		X"06",X"04",X"04",X"04",X"06",X"04",X"05",X"04",X"06",X"04",X"05",X"06",X"03",X"02",X"3E",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
