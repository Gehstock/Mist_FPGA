library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"E2",X"82",X"FE",X"7E",X"02",
		X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"04",X"08",X"04",X"FE",X"FE",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7C",X"FE",X"C6",X"C6",X"FE",X"7C",X"00",X"00",X"FE",X"FE",X"38",X"7C",X"EE",X"C6",X"00",
		X"00",X"60",X"60",X"00",X"0C",X"0E",X"06",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",
		X"00",X"44",X"6C",X"38",X"38",X"6C",X"44",X"00",X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",
		X"00",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",
		X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",
		X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",
		X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",
		X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",
		X"00",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",
		X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",
		X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",
		X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",
		X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"16",X"0E",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",
		X"00",X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",
		X"00",X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",
		X"00",X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",
		X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",
		X"00",X"00",X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"3E",X"FE",X"70",X"38",X"70",X"FE",X"3E",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"06",X"1E",X"F0",X"F0",X"1E",X"06",
		X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",
		X"00",X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",
		X"00",X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",
		X"00",X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",
		X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",
		X"00",X"00",X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"3E",X"FE",X"70",X"38",X"70",X"FE",X"3E",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"06",X"1E",X"F0",X"F0",X"1E",X"06",
		X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"60",X"60",X"08",X"1C",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"50",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"7E",X"81",X"BD",X"BD",X"A5",X"A5",X"81",X"7E",
		X"00",X"FF",X"FF",X"C3",X"C3",X"E7",X"7E",X"7E",X"FF",X"DB",X"DB",X"DB",X"7E",X"FF",X"C3",X"C3",
		X"F7",X"76",X"7E",X"FF",X"C3",X"C3",X"FF",X"7E",X"00",X"76",X"81",X"81",X"81",X"81",X"81",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"70",X"89",X"89",X"89",X"89",X"89",X"06",
		X"00",X"00",X"81",X"89",X"89",X"89",X"89",X"76",X"00",X"06",X"08",X"08",X"08",X"08",X"F7",X"00",
		X"00",X"06",X"89",X"89",X"89",X"89",X"89",X"70",X"00",X"76",X"89",X"89",X"89",X"89",X"89",X"70",
		X"00",X"06",X"01",X"01",X"01",X"01",X"01",X"76",X"00",X"76",X"89",X"89",X"89",X"89",X"89",X"76",
		X"00",X"06",X"89",X"89",X"89",X"89",X"89",X"76",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"50",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"6C",X"82",X"6C",X"00",X"6C",X"82",X"6C",X"00",X"00",X"00",X"EE",X"00",X"6C",X"82",X"6C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"E2",X"92",X"8C",
		X"00",X"00",X"00",X"00",X"82",X"92",X"92",X"6C",X"00",X"00",X"00",X"00",X"0E",X"10",X"10",X"EC",
		X"00",X"00",X"00",X"00",X"8E",X"92",X"92",X"E2",X"00",X"00",X"00",X"00",X"7C",X"92",X"92",X"60",
		X"00",X"00",X"00",X"00",X"82",X"42",X"22",X"1E",X"00",X"00",X"00",X"00",X"6C",X"92",X"92",X"6C",
		X"00",X"00",X"00",X"00",X"4C",X"92",X"92",X"7C",X"00",X"6C",X"82",X"6C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"FC",X"FE",X"AA",X"AA",X"D6",X"D6",X"FE",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"60",X"6F",X"7C",X"7C",X"6C",X"6F",X"7F",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"40",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",X"7F",X"C0",X"8A",X"AA",X"AA",
		X"40",X"40",X"40",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D5",X"D5",X"94",X"C0",X"7F",X"3F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"BD",X"D1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"02",
		X"D1",X"BD",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"38",X"10",X"40",X"00",X"10",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FC",X"FE",X"06",X"7E",X"F6",X"C6",X"C6",X"16",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"3F",X"FF",X"FF",X"F0",X"8A",X"AA",X"BF",X"86",
		X"16",X"C6",X"C6",X"F6",X"7E",X"06",X"FE",X"FC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"86",X"BF",X"AA",X"8A",X"F0",X"FF",X"FF",X"3F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"19",X"11",X"35",X"B7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"08",X"00",X"01",X"01",X"81",X"19",X"61",
		X"B7",X"35",X"11",X"19",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"61",X"19",X"81",X"01",X"01",X"00",X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"87",X"F7",X"FF",X"F7",X"C6",X"C4",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"FF",X"E1",X"84",X"92",X"8A",X"AA",X"BF",X"90",
		X"00",X"C4",X"C6",X"F7",X"FF",X"F7",X"87",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"90",X"BF",X"AA",X"8A",X"92",X"84",X"E1",X"FF",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"03",
		X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"07",X"8F",X"FF",X"00",X"00",X"80",X"C2",X"FF",X"FB",
		X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"30",X"3B",X"1F",X"1E",X"1F",X"1B",X"1B",X"1D",X"1D",
		X"FB",X"FF",X"C2",X"80",X"00",X"00",X"FF",X"8F",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",
		X"1D",X"1D",X"1B",X"1B",X"1F",X"1E",X"1F",X"3B",X"30",X"00",X"00",X"00",X"00",X"00",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"D0",X"F0",X"D0",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1F",X"F8",X"C5",X"15",X"5F",X"70",
		X"10",X"D0",X"F0",X"D0",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"5F",X"15",X"C5",X"F8",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"FC",X"77",X"E1",X"C1",X"85",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1E",X"1C",X"19",X"19",X"1B",X"1A",
		X"F7",X"FF",X"85",X"C1",X"E1",X"77",X"FC",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"1B",X"19",X"19",X"1C",X"1E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"38",X"FC",X"02",X"56",X"56",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"02",X"FC",X"38",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"FC",X"87",X"1F",X"31",X"B7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"B7",X"31",X"1F",X"87",X"FC",X"70",X"00",X"00",X"00",X"02",X"08",X"00",X"44",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"7F",X"F0",X"0A",X"AB",X"FE",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"AB",X"0A",X"F0",X"7F",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"01",X"00",X"00",X"1C",X"3F",X"41",X"5F",X"79",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"00",X"61",
		X"79",X"5F",X"41",X"3F",X"1C",X"00",X"00",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"89",X"00",X"00",X"10",X"80",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"FC",X"06",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"56",X"56",X"06",X"FC",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"1C",X"3F",X"41",X"5F",X"79",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"79",X"5F",X"41",X"3F",X"1C",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"00",X"78",X"78",X"03",X"03",X"03",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"7F",X"21",X"2D",X"21",X"21",X"7F",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"00",X"0E",X"1C",X"00",X"00",X"1C",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"20",X"20",X"18",X"00",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"18",X"FC",X"76",X"43",X"FF",X"FF",X"73",X"06",X"FC",X"18",X"18",X"00",X"00",
		X"18",X"18",X"3C",X"7E",X"D7",X"D7",X"FE",X"FE",X"FE",X"FE",X"D7",X"D7",X"7E",X"3C",X"18",X"18",
		X"08",X"10",X"00",X"00",X"00",X"78",X"CD",X"FD",X"FD",X"CD",X"78",X"00",X"00",X"00",X"10",X"08",
		X"21",X"42",X"00",X"00",X"00",X"21",X"12",X"0D",X"0D",X"12",X"21",X"00",X"00",X"00",X"42",X"21",
		X"90",X"92",X"92",X"92",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"48",X"48",X"48",X"48",
		X"24",X"24",X"24",X"24",X"1F",X"00",X"03",X"07",X"07",X"03",X"00",X"1F",X"92",X"92",X"92",X"12",
		X"00",X"0F",X"18",X"08",X"D8",X"0F",X"58",X"48",X"58",X"4F",X"18",X"CF",X"18",X"0F",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"07",X"07",X"06",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"10",X"02",X"02",X"02",X"02",X"10",X"C0",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"02",X"02",X"00",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"10",X"02",X"02",X"02",X"02",X"10",X"C0",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"30",X"30",X"30",X"00",X"30",X"36",X"36",X"30",X"00",X"30",X"30",X"30",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"10",X"02",X"02",X"02",X"02",X"10",X"C0",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"60",X"60",X"60",X"00",X"60",X"6E",X"6E",X"60",X"00",X"60",X"60",X"60",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"90",X"78",X"C8",X"C8",X"78",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"3D",X"7B",X"16",X"10",X"78",X"3C",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"46",X"46",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"90",X"FA",X"FD",X"FE",X"FE",X"DE",X"FC",X"EC",X"F8",X"FC",X"FC",X"FC",X"F8",X"38",X"10",
		X"00",X"33",X"7B",X"3F",X"3F",X"7E",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"5F",X"1F",X"29",X"18",
		X"00",X"16",X"BF",X"FE",X"F7",X"FF",X"BE",X"FC",X"78",X"FC",X"FE",X"DC",X"9C",X"FC",X"EA",X"C0",
		X"10",X"3B",X"7F",X"7F",X"7F",X"3B",X"7F",X"EF",X"6F",X"3F",X"7F",X"7F",X"FE",X"7F",X"73",X"20",
		X"21",X"FB",X"FE",X"FE",X"4C",X"8C",X"76",X"FD",X"FE",X"DD",X"78",X"7C",X"BE",X"FC",X"F8",X"70",
		X"05",X"7E",X"3F",X"7F",X"77",X"FB",X"F5",X"F7",X"79",X"7E",X"7F",X"5E",X"37",X"07",X"03",X"01",
		X"E0",X"D8",X"EC",X"5C",X"D6",X"AE",X"FF",X"77",X"EE",X"8C",X"AE",X"54",X"48",X"F8",X"30",X"C0",
		X"12",X"3B",X"7F",X"7F",X"7F",X"28",X"DF",X"D2",X"4D",X"75",X"FB",X"65",X"FB",X"65",X"2F",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"BE",X"F8",X"69",X"F2",X"76",X"FC",X"DC",X"F0",
		X"00",X"30",X"40",X"80",X"00",X"00",X"80",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"BC",X"F0",X"D5",X"F6",X"6D",X"27",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"01",X"49",X"6E",X"39",X"1F",X"6B",X"2D",X"7D",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"3F",X"BD",X"F7",X"F9",X"F9",X"82",X"87",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"90",X"F0",X"FC",X"FC",X"FC",X"F8",X"F8",X"B0",X"58",X"80",X"10",X"80",X"C0",X"00",X"00",
		X"00",X"05",X"09",X"93",X"EF",X"EF",X"7F",X"FD",X"FF",X"FF",X"FF",X"FD",X"F7",X"F5",X"FB",X"FF",
		X"80",X"B0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"FB",X"79",X"DB",X"F7",X"FB",X"D6",X"7F",X"F9",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"07",X"0B",X"3F",X"FF",X"7F",X"D5",X"DF",X"FF",X"7B",X"3D",X"C7",X"6B",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"5F",X"26",X"01",X"00",
		X"FF",X"EF",X"6F",X"F7",X"ED",X"FD",X"F7",X"7F",X"EF",X"AF",X"41",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"03",X"05",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"D0",X"FA",X"7E",X"FC",X"DE",X"FC",X"58",X"BC",X"F8",X"F0",X"70",X"C0",X"C0",X"80",X"00",
		X"00",X"07",X"1F",X"DB",X"EB",X"EB",X"FE",X"BF",X"5D",X"25",X"4B",X"A1",X"0D",X"53",X"13",X"0A",
		X"90",X"F8",X"FC",X"FC",X"FC",X"FA",X"7E",X"BC",X"FE",X"E5",X"EE",X"F4",X"E4",X"F0",X"E0",X"00",
		X"43",X"23",X"41",X"12",X"2D",X"4B",X"9D",X"E1",X"8F",X"FF",X"FF",X"7F",X"5F",X"FF",X"76",X"60",
		X"10",X"D6",X"D4",X"FF",X"FF",X"BF",X"FF",X"6F",X"FF",X"FF",X"FE",X"FC",X"FE",X"EC",X"EB",X"F0",
		X"00",X"01",X"02",X"07",X"0F",X"07",X"05",X"03",X"0F",X"BF",X"FD",X"7F",X"7F",X"1F",X"3B",X"3E",
		X"F0",X"EA",X"FA",X"F4",X"EC",X"F2",X"DF",X"FF",X"FF",X"FF",X"A7",X"FB",X"B0",X"33",X"01",X"00",
		X"1F",X"37",X"1F",X"17",X"15",X"17",X"3D",X"7F",X"7F",X"3B",X"5F",X"BF",X"5B",X"00",X"00",X"00",
		X"80",X"00",X"00",X"10",X"48",X"94",X"0C",X"12",X"02",X"28",X"16",X"01",X"8C",X"A4",X"40",X"50",
		X"12",X"60",X"8E",X"25",X"20",X"40",X"09",X"16",X"68",X"4E",X"A0",X"40",X"00",X"01",X"04",X"04",
		X"A8",X"C0",X"12",X"B0",X"40",X"06",X"04",X"22",X"D0",X"18",X"E0",X"10",X"20",X"88",X"40",X"20",
		X"00",X"02",X"01",X"00",X"42",X"80",X"00",X"00",X"80",X"34",X"40",X"23",X"0B",X"08",X"05",X"03",
		X"10",X"04",X"10",X"11",X"01",X"02",X"80",X"08",X"86",X"25",X"01",X"80",X"10",X"00",X"20",X"D0",
		X"0A",X"00",X"00",X"04",X"00",X"04",X"02",X"01",X"0C",X"0A",X"05",X"00",X"00",X"0A",X"00",X"02",
		X"00",X"80",X"20",X"00",X"80",X"44",X"80",X"22",X"25",X"0A",X"90",X"44",X"60",X"10",X"D0",X"00",
		X"00",X"48",X"04",X"00",X"14",X"4A",X"00",X"04",X"12",X"20",X"10",X"82",X"46",X"09",X"14",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"74",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"20",X"20",X"80",X"00",X"40",
		X"00",X"00",X"00",X"04",X"20",X"04",X"00",X"93",X"40",X"09",X"60",X"7A",X"F5",X"FA",X"F4",X"F8",
		X"00",X"20",X"20",X"00",X"80",X"00",X"20",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"BC",X"11",X"28",X"58",X"30",X"10",X"00",X"22",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"56",X"2E",X"52",X"0C",X"0F",X"BF",X"37",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"06",X"02",X"01",X"05",X"08",X"02",
		X"07",X"25",X"8F",X"0F",X"2C",X"8A",X"49",X"04",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"20",X"40",X"20",X"10",X"00",X"00",X"C0",X"80",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"01",X"00",X"00",X"A0",X"12",X"14",X"02",X"01",X"20",X"40",X"01",X"80",X"40",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"22",X"01",X"81",X"40",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",X"00",X"08",X"10",X"00",X"80",X"48",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",
		X"80",X"80",X"C0",X"40",X"20",X"40",X"C0",X"A0",X"05",X"0A",X"04",X"04",X"14",X"08",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"40",X"A0",X"D0",X"E8",X"F4",X"0A",X"05",X"05",X"0A",X"F4",X"E8",X"D0",X"A0",X"40",X"80",
		X"01",X"02",X"05",X"0B",X"17",X"2F",X"57",X"A2",X"A2",X"57",X"2F",X"17",X"0B",X"05",X"02",X"01",
		X"00",X"A0",X"80",X"0A",X"82",X"19",X"8A",X"2C",X"40",X"90",X"04",X"10",X"54",X"4E",X"0A",X"00",
		X"00",X"80",X"92",X"12",X"41",X"40",X"02",X"00",X"01",X"00",X"84",X"80",X"2E",X"23",X"04",X"00",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"20",X"20",X"20",X"20",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"01",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"1F",X"10",X"38",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"E0",X"60",X"00",X"08",X"3E",X"77",X"63",X"C1",X"C1",X"63",X"77",X"3E",X"08",
		X"00",X"00",X"00",X"0C",X"E8",X"E8",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"46",X"40",X"40",X"46",X"40",X"42",X"02",X"02",X"02",X"1E",X"10",X"38",X"10",
		X"00",X"00",X"80",X"00",X"00",X"00",X"30",X"00",X"80",X"04",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"08",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"C0",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"38",X"78",X"10",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"63",X"77",X"00",X"00",X"00",X"00",X"00",X"19",X"16",X"38",X"10",
		X"00",X"02",X"17",X"7E",X"FC",X"D6",X"74",X"7C",X"74",X"D4",X"F8",X"70",X"00",X"00",X"80",X"00",
		X"01",X"02",X"9E",X"BE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"BE",X"9E",X"81",X"00",X"00",
		X"00",X"60",X"70",X"60",X"60",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"23",X"03",X"0B",X"0B",X"07",X"9F",X"03",X"02",X"02",X"02",X"02",X"0E",X"1C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"C1",X"FB",X"FF",X"FF",X"FF",X"BF",X"87",X"C1",X"C3",X"E7",X"FF",X"FF",X"7E",X"3C",
		X"F0",X"FE",X"FF",X"FF",X"FF",X"CF",X"C1",X"C0",X"E1",X"F3",X"FF",X"7F",X"3F",X"0E",X"00",X"00",
		X"00",X"00",X"C1",X"FB",X"FF",X"3F",X"07",X"00",X"00",X"00",X"C1",X"FF",X"FF",X"3F",X"07",X"00",
		X"F0",X"FE",X"FF",X"EF",X"C3",X"C0",X"C0",X"E0",X"F0",X"FE",X"7F",X"0F",X"01",X"00",X"00",X"00",
		X"00",X"01",X"C1",X"FB",X"FF",X"FF",X"FF",X"BF",X"87",X"C1",X"C3",X"E7",X"FF",X"FF",X"7E",X"3C",
		X"F0",X"FE",X"FF",X"FF",X"7F",X"0F",X"01",X"00",X"01",X"CF",X"FF",X"FF",X"FE",X"F0",X"F0",X"00",
		X"00",X"00",X"01",X"C1",X"FB",X"FF",X"3F",X"FF",X"FF",X"FE",X"00",X"C0",X"F8",X"FF",X"3F",X"07",
		X"00",X"F0",X"FE",X"7F",X"0F",X"01",X"00",X"03",X"1F",X"FF",X"FE",X"7F",X"0F",X"01",X"00",X"00",
		X"00",X"00",X"C1",X"FB",X"FF",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FE",X"FF",X"7F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C1",X"FB",X"FF",X"FF",X"FF",X"BF",X"87",X"83",X"03",X"03",X"03",X"03",X"03",X"00",
		X"F0",X"FE",X"FF",X"FF",X"FF",X"CF",X"C3",X"C1",X"C1",X"C1",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"37",X"3F",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C1",X"C1",X"C1",X"03",X"07",X"07",X"C7",X"FF",X"FF",X"FF",X"3F",X"07",X"03",X"00",
		X"1E",X"3F",X"7F",X"FF",X"F1",X"E0",X"E0",X"FE",X"7F",X"3F",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"C1",X"FB",X"FF",X"FF",X"FF",X"BF",X"87",X"C1",X"C3",X"E7",X"FF",X"FF",X"7E",X"3C",
		X"F0",X"FE",X"FF",X"FF",X"3F",X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"01",X"C1",X"FB",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"FD",X"FF",X"FF",X"FF",X"3F",
		X"F0",X"FE",X"FF",X"FF",X"0F",X"00",X"03",X"07",X"03",X"F0",X"FE",X"FF",X"FF",X"0F",X"01",X"00",
		X"00",X"00",X"08",X"08",X"F8",X"08",X"08",X"00",X"F8",X"10",X"20",X"10",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"81",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",
		X"00",X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
