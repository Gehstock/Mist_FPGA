library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity vec_rom_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of vec_rom_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"A0",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"90",X"FF",X"73",X"FF",X"92",X"00",X"70",
		X"00",X"90",X"FF",X"77",X"FF",X"96",X"00",X"70",X"FF",X"92",X"FF",X"72",X"00",X"86",X"00",X"72",
		X"FE",X"87",X"FE",X"77",X"00",X"92",X"00",X"76",X"FE",X"81",X"00",X"72",X"FF",X"96",X"FF",X"72",
		X"7F",X"A3",X"FF",X"03",X"00",X"70",X"00",X"00",X"FF",X"96",X"FF",X"76",X"FE",X"81",X"00",X"76",
		X"00",X"92",X"00",X"72",X"FE",X"87",X"FE",X"73",X"00",X"86",X"00",X"76",X"FF",X"92",X"FF",X"76",
		X"FC",X"A1",X"F4",X"01",X"00",X"70",X"00",X"00",X"DB",X"F0",X"00",X"F9",X"CF",X"F0",X"00",X"F9",
		X"BB",X"F0",X"00",X"F9",X"AF",X"F0",X"00",X"F9",X"9B",X"F0",X"00",X"F9",X"8F",X"F0",X"00",X"F9",
		X"7B",X"F0",X"00",X"F9",X"6F",X"F0",X"00",X"F9",X"5B",X"F0",X"00",X"F9",X"4F",X"F0",X"00",X"F9",
		X"3B",X"F0",X"00",X"F9",X"2F",X"F0",X"7C",X"D0",X"E4",X"A0",X"5E",X"11",X"00",X"70",X"00",X"00",
		X"80",X"CA",X"78",X"CA",X"D8",X"CA",X"C7",X"CA",X"2C",X"CB",X"9B",X"CA",X"F3",X"CA",X"F3",X"CA",
		X"DD",X"CA",X"F3",X"EA",X"80",X"A0",X"90",X"01",X"00",X"70",X"00",X"00",X"73",X"F5",X"73",X"F1",
		X"78",X"F1",X"77",X"F1",X"77",X"F5",X"78",X"F5",X"80",X"31",X"00",X"02",X"75",X"F8",X"70",X"FD",
		X"71",X"F8",X"02",X"FD",X"2E",X"CB",X"63",X"CB",X"56",X"CB",X"63",X"CB",X"2C",X"CB",X"78",X"CA",
		X"02",X"CB",X"78",X"CA",X"F3",X"CA",X"BA",X"CA",X"2C",X"CB",X"BA",X"CA",X"D8",X"CA",X"8D",X"EA",
		X"C6",X"FF",X"C1",X"FE",X"C3",X"F1",X"CD",X"F1",X"C7",X"F1",X"C1",X"FD",X"D8",X"1E",X"32",X"EC",
		X"00",X"C4",X"3C",X"14",X"0A",X"46",X"D8",X"D8",X"D0",X"C8",X"B5",X"C8",X"96",X"C8",X"80",X"C8",
		X"0D",X"F8",X"78",X"F8",X"0D",X"FD",X"78",X"F8",X"09",X"FD",X"78",X"F8",X"0B",X"F1",X"78",X"F8",
		X"0A",X"F5",X"78",X"F8",X"08",X"F9",X"78",X"F8",X"09",X"F3",X"78",X"F8",X"0D",X"F3",X"78",X"F8",
		X"80",X"54",X"00",X"06",X"78",X"F8",X"0F",X"F1",X"78",X"F8",X"00",X"D0",X"00",X"30",X"80",X"07",
		X"78",X"F8",X"80",X"37",X"80",X"07",X"78",X"F8",X"80",X"37",X"80",X"03",X"78",X"F8",X"E0",X"40",
		X"A0",X"02",X"78",X"F8",X"C0",X"35",X"80",X"03",X"78",X"F8",X"80",X"33",X"00",X"00",X"78",X"F8",
		X"A0",X"42",X"E0",X"00",X"78",X"F8",X"A0",X"42",X"E0",X"04",X"78",X"F8",X"E0",X"44",X"80",X"07",
		X"78",X"F8",X"E0",X"40",X"A0",X"06",X"78",X"F8",X"00",X"D0",X"07",X"F8",X"78",X"F8",X"07",X"FF",
		X"78",X"F8",X"03",X"FF",X"78",X"F8",X"C0",X"40",X"40",X"02",X"78",X"F8",X"80",X"35",X"00",X"03",
		X"78",X"F8",X"00",X"FB",X"78",X"F8",X"40",X"42",X"C0",X"00",X"78",X"F8",X"40",X"42",X"C0",X"04",
		X"78",X"F8",X"C0",X"44",X"00",X"07",X"78",X"F8",X"C0",X"40",X"40",X"06",X"78",X"F8",X"00",X"D0",
		X"00",X"30",X"80",X"06",X"78",X"F8",X"80",X"36",X"80",X"06",X"78",X"F8",X"80",X"36",X"80",X"02",
		X"78",X"F8",X"40",X"31",X"C0",X"03",X"78",X"F8",X"40",X"35",X"80",X"02",X"78",X"F8",X"80",X"32",
		X"00",X"00",X"78",X"F8",X"C0",X"33",X"40",X"01",X"78",X"F8",X"C0",X"33",X"40",X"05",X"78",X"F8",
		X"A0",X"44",X"80",X"06",X"78",X"F8",X"40",X"31",X"C0",X"07",X"78",X"F8",X"00",X"D0",X"F3",X"C8",
		X"FF",X"C8",X"0D",X"C9",X"1A",X"C9",X"08",X"F9",X"79",X"F9",X"79",X"FD",X"7D",X"F6",X"79",X"F6",
		X"8F",X"F6",X"8F",X"F0",X"7D",X"F9",X"78",X"FA",X"79",X"F9",X"79",X"FD",X"00",X"D0",X"0A",X"F1",
		X"7A",X"F1",X"7D",X"F9",X"7E",X"F5",X"7E",X"F1",X"7D",X"FD",X"79",X"F6",X"7D",X"F6",X"79",X"FD",
		X"79",X"F1",X"8B",X"F5",X"8A",X"F3",X"7D",X"F9",X"00",X"D0",X"0D",X"F8",X"7E",X"F5",X"7A",X"F7",
		X"7A",X"F3",X"78",X"F7",X"79",X"F8",X"7A",X"F3",X"78",X"F9",X"7E",X"F3",X"7F",X"F0",X"7F",X"F7",
		X"7A",X"F5",X"00",X"D0",X"09",X"F0",X"7B",X"F1",X"68",X"F1",X"7F",X"F2",X"7F",X"F0",X"69",X"F6",
		X"7F",X"F0",X"78",X"F7",X"7A",X"F7",X"7B",X"F1",X"69",X"F5",X"69",X"F9",X"7F",X"F2",X"00",X"D0",
		X"29",X"C9",X"0E",X"F1",X"CA",X"F8",X"0B",X"F6",X"00",X"60",X"80",X"D6",X"DB",X"F6",X"CA",X"F8",
		X"DB",X"F2",X"DF",X"F2",X"CD",X"F2",X"CD",X"F8",X"CD",X"F6",X"DF",X"F6",X"00",X"D0",X"90",X"52",
		X"A8",X"52",X"CC",X"52",X"F0",X"52",X"14",X"53",X"36",X"53",X"5A",X"53",X"7E",X"53",X"A2",X"53",
		X"C6",X"53",X"EA",X"53",X"0E",X"54",X"32",X"54",X"56",X"54",X"7A",X"54",X"9E",X"54",X"C2",X"54",
		X"0F",X"F6",X"C8",X"FA",X"BD",X"F9",X"00",X"65",X"00",X"C3",X"00",X"65",X"00",X"C7",X"B9",X"F9",
		X"00",X"D0",X"CE",X"F9",X"CA",X"F9",X"00",X"D0",X"40",X"46",X"C0",X"06",X"00",X"52",X"30",X"C4",
		X"C0",X"41",X"20",X"C6",X"B0",X"64",X"18",X"C3",X"48",X"65",X"E0",X"C6",X"20",X"42",X"C0",X"C1",
		X"00",X"D0",X"D0",X"50",X"10",X"C6",X"60",X"42",X"C0",X"C3",X"00",X"D0",X"80",X"46",X"80",X"06",
		X"E0",X"43",X"C0",X"C4",X"A0",X"41",X"60",X"C6",X"68",X"64",X"20",X"C3",X"90",X"65",X"C0",X"C6",
		X"60",X"42",X"A0",X"C1",X"00",X"D0",X"90",X"50",X"30",X"C6",X"C0",X"42",X"80",X"C3",X"00",X"D0",
		X"C0",X"46",X"40",X"06",X"E0",X"43",X"20",X"C5",X"60",X"41",X"80",X"C6",X"18",X"64",X"28",X"C3",
		X"D0",X"65",X"98",X"C6",X"80",X"42",X"60",X"C1",X"00",X"D0",X"60",X"50",X"30",X"C6",X"20",X"43",
		X"40",X"C3",X"00",X"D0",X"0E",X"F7",X"C0",X"43",X"80",X"C5",X"20",X"41",X"A0",X"C6",X"38",X"60",
		X"28",X"C3",X"10",X"66",X"60",X"C6",X"A0",X"42",X"20",X"C1",X"00",X"D0",X"30",X"50",X"40",X"C6",
		X"60",X"43",X"E0",X"C2",X"00",X"D0",X"20",X"47",X"C0",X"05",X"80",X"43",X"E0",X"C5",X"E0",X"40",
		X"C0",X"C6",X"88",X"60",X"20",X"C3",X"48",X"66",X"30",X"C6",X"C0",X"42",X"E0",X"C0",X"00",X"D0",
		X"10",X"54",X"40",X"C6",X"A0",X"43",X"A0",X"C2",X"00",X"D0",X"60",X"47",X"60",X"05",X"60",X"43",
		X"40",X"C6",X"80",X"40",X"C0",X"C6",X"D8",X"60",X"10",X"C3",X"80",X"66",X"F0",X"C5",X"C0",X"42",
		X"80",X"C0",X"00",X"D0",X"40",X"54",X"30",X"C6",X"E0",X"43",X"40",X"C2",X"00",X"D0",X"80",X"47",
		X"00",X"05",X"20",X"43",X"80",X"C6",X"40",X"40",X"E0",X"C6",X"20",X"61",X"F8",X"C2",X"B0",X"66",
		X"B0",X"C5",X"E0",X"42",X"40",X"C0",X"00",X"D0",X"80",X"54",X"30",X"C6",X"10",X"52",X"F0",X"C0",
		X"00",X"D0",X"80",X"47",X"C0",X"04",X"E0",X"42",X"E0",X"C6",X"00",X"40",X"E0",X"C6",X"68",X"61",
		X"D8",X"C2",X"D8",X"66",X"68",X"C5",X"E0",X"42",X"00",X"C0",X"00",X"D0",X"B0",X"54",X"20",X"C6",
		X"20",X"52",X"B0",X"C0",X"00",X"D0",X"A0",X"47",X"60",X"04",X"80",X"42",X"20",X"C7",X"40",X"44",
		X"E0",X"C6",X"B0",X"61",X"B0",X"C2",X"F8",X"66",X"20",X"C5",X"E0",X"42",X"40",X"C4",X"00",X"D0",
		X"F0",X"54",X"10",X"C6",X"30",X"52",X"80",X"C0",X"00",X"D0",X"A0",X"47",X"00",X"00",X"40",X"42",
		X"60",X"C7",X"80",X"44",X"C0",X"C6",X"F0",X"61",X"80",X"C2",X"10",X"67",X"D8",X"C4",X"C0",X"42",
		X"80",X"C4",X"00",X"D0",X"40",X"46",X"E0",X"C7",X"30",X"52",X"40",X"C0",X"00",X"D0",X"A0",X"47",
		X"60",X"00",X"E0",X"41",X"80",X"C7",X"E0",X"44",X"C0",X"C6",X"30",X"62",X"48",X"C2",X"20",X"67",
		X"88",X"C4",X"C0",X"42",X"E0",X"C4",X"00",X"D0",X"A0",X"46",X"A0",X"C7",X"40",X"52",X"10",X"C0",
		X"00",X"D0",X"80",X"47",X"C0",X"00",X"80",X"41",X"C0",X"C7",X"20",X"45",X"A0",X"C6",X"60",X"62",
		X"10",X"C2",X"28",X"67",X"38",X"C4",X"A0",X"42",X"20",X"C5",X"00",X"D0",X"E0",X"46",X"60",X"C7",
		X"40",X"52",X"30",X"C4",X"00",X"D0",X"80",X"47",X"00",X"01",X"20",X"41",X"E0",X"C7",X"60",X"45",
		X"80",X"C6",X"98",X"62",X"D0",X"C1",X"28",X"67",X"18",X"C0",X"80",X"42",X"60",X"C5",X"00",X"D0",
		X"40",X"47",X"20",X"C7",X"30",X"52",X"60",X"C4",X"00",X"D0",X"60",X"47",X"60",X"01",X"C0",X"40",
		X"E0",X"C7",X"A0",X"45",X"60",X"C6",X"C0",X"62",X"90",X"C1",X"20",X"67",X"68",X"C0",X"60",X"42",
		X"A0",X"C5",X"00",X"D0",X"80",X"47",X"C0",X"C6",X"30",X"52",X"90",X"C4",X"00",X"D0",X"20",X"47",
		X"C0",X"01",X"30",X"50",X"00",X"C6",X"C0",X"45",X"20",X"C6",X"E0",X"62",X"48",X"C1",X"18",X"67",
		X"B0",X"C0",X"20",X"42",X"C0",X"C5",X"00",X"D0",X"C0",X"47",X"60",X"C6",X"10",X"52",X"D0",X"C4",
		X"00",X"D0",X"0A",X"F7",X"CE",X"F8",X"CD",X"FD",X"00",X"63",X"00",X"C1",X"00",X"67",X"00",X"C1",
		X"CD",X"F9",X"00",X"D0",X"CD",X"FE",X"CD",X"FA",X"00",X"D0",X"0E",X"F7",X"7A",X"F8",X"79",X"FD",
		X"00",X"63",X"00",X"75",X"00",X"67",X"00",X"75",X"79",X"F9",X"C0",X"60",X"80",X"02",X"9F",X"D0",
		X"70",X"FA",X"72",X"F2",X"72",X"F6",X"70",X"FE",X"06",X"F9",X"72",X"F8",X"02",X"F6",X"00",X"D0",
		X"70",X"FB",X"73",X"F0",X"71",X"F5",X"70",X"F5",X"75",X"F5",X"77",X"F0",X"03",X"F0",X"71",X"F5",
		X"70",X"F5",X"75",X"F5",X"77",X"F0",X"03",X"F8",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"06",X"FF",
		X"72",X"F8",X"02",X"F0",X"00",X"D0",X"70",X"FB",X"72",X"F0",X"72",X"F6",X"70",X"F6",X"76",X"F6",
		X"76",X"F0",X"03",X"F8",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"05",X"F7",X"77",X"F0",X"00",X"F7",
		X"72",X"F8",X"02",X"F0",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"05",X"F7",X"77",X"F0",X"00",X"F7",
		X"03",X"F8",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"70",X"F6",X"06",X"F6",X"72",X"F0",X"70",X"F6",
		X"76",X"F8",X"03",X"F8",X"00",X"D0",X"70",X"FB",X"00",X"F7",X"72",X"F8",X"00",X"F3",X"70",X"FF",
		X"02",X"F0",X"00",X"D0",X"72",X"F8",X"06",X"F0",X"70",X"FB",X"02",X"F0",X"76",X"F8",X"03",X"FF",
		X"00",X"D0",X"00",X"F2",X"72",X"F6",X"72",X"F0",X"70",X"FB",X"01",X"FF",X"00",X"D0",X"70",X"FB",
		X"03",X"F0",X"77",X"F7",X"73",X"F7",X"03",X"F0",X"00",X"D0",X"00",X"FB",X"70",X"FF",X"72",X"F8",
		X"02",X"F0",X"00",X"D0",X"70",X"FB",X"72",X"F6",X"72",X"F2",X"70",X"FF",X"02",X"F0",X"00",X"D0",
		X"70",X"FB",X"72",X"FF",X"70",X"FB",X"01",X"FF",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"70",X"FF",
		X"76",X"F8",X"03",X"F8",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"70",X"F7",X"76",X"F8",X"03",X"F7",
		X"03",X"F0",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"70",X"FE",X"76",X"F6",X"76",X"F0",X"02",X"F2",
		X"72",X"F6",X"02",X"F0",X"00",X"D0",X"70",X"FB",X"72",X"F8",X"70",X"F7",X"76",X"F8",X"01",X"F0",
		X"73",X"F7",X"02",X"F0",X"00",X"D0",X"72",X"F8",X"70",X"F3",X"76",X"F8",X"70",X"F3",X"72",X"F8",
		X"01",X"FF",X"00",X"D0",X"02",X"F0",X"70",X"FB",X"06",X"F0",X"72",X"F8",X"01",X"FF",X"00",X"D0",
		X"00",X"FB",X"70",X"FF",X"72",X"F8",X"70",X"FB",X"01",X"FF",X"00",X"D0",X"00",X"FB",X"71",X"FF",
		X"71",X"FB",X"01",X"FF",X"00",X"D0",X"00",X"FB",X"70",X"FF",X"72",X"F2",X"72",X"F6",X"70",X"FB",
		X"01",X"FF",X"00",X"D0",X"72",X"FB",X"06",X"F8",X"72",X"FF",X"02",X"F0",X"00",X"D0",X"02",X"F0",
		X"70",X"FA",X"76",X"F2",X"02",X"F8",X"76",X"F6",X"02",X"FE",X"00",X"D0",X"00",X"FB",X"72",X"F8",
		X"76",X"FF",X"72",X"F8",X"02",X"F0",X"00",X"D0",X"03",X"F8",X"00",X"D0",X"02",X"F0",X"70",X"FB",
		X"02",X"FF",X"00",X"D0",X"00",X"FB",X"72",X"F8",X"70",X"F7",X"76",X"F8",X"70",X"F7",X"72",X"F8",
		X"02",X"F0",X"00",X"D0",X"72",X"F8",X"70",X"FB",X"76",X"F8",X"00",X"F7",X"72",X"F8",X"02",X"F7",
		X"00",X"D0",X"00",X"FB",X"70",X"F7",X"72",X"F8",X"00",X"F3",X"70",X"FF",X"02",X"F0",X"00",X"D0",
		X"72",X"F8",X"70",X"F3",X"76",X"F8",X"70",X"F3",X"72",X"F8",X"01",X"FF",X"00",X"D0",X"00",X"F3",
		X"72",X"F8",X"70",X"F7",X"76",X"F8",X"70",X"FB",X"03",X"FF",X"00",X"D0",X"00",X"FB",X"72",X"F8",
		X"70",X"FF",X"02",X"F0",X"00",X"D0",X"72",X"F8",X"70",X"FB",X"76",X"F8",X"70",X"FF",X"00",X"F3",
		X"72",X"F8",X"02",X"F7",X"00",X"D0",X"02",X"F8",X"70",X"FB",X"76",X"F8",X"70",X"F7",X"72",X"F8",
		X"02",X"F7",X"00",X"D0",X"2C",X"CB",X"DD",X"CA",X"2E",X"CB",X"32",X"CB",X"3A",X"CB",X"41",X"CB",
		X"48",X"CB",X"4F",X"CB",X"56",X"CB",X"5B",X"CB",X"63",X"CB",X"78",X"CA",X"80",X"CA",X"8D",X"CA",
		X"93",X"CA",X"9B",X"CA",X"A3",X"CA",X"AA",X"CA",X"B3",X"CA",X"BA",X"CA",X"C1",X"CA",X"C7",X"CA",
		X"CD",X"CA",X"D2",X"CA",X"D8",X"CA",X"DD",X"CA",X"E3",X"CA",X"EA",X"CA",X"F3",X"CA",X"FB",X"CA",
		X"02",X"CB",X"08",X"CB",X"0E",X"CB",X"13",X"CB",X"1A",X"CB",X"1F",X"CB",X"26",X"CB",X"0B",X"13",
		X"19",X"2F",X"41",X"55",X"6F",X"77",X"7D",X"87",X"91",X"63",X"56",X"60",X"6E",X"3C",X"EC",X"4D",
		X"C0",X"A4",X"0A",X"EA",X"6C",X"08",X"00",X"EC",X"F2",X"B0",X"6E",X"3C",X"EC",X"48",X"5A",X"B8",
		X"66",X"92",X"42",X"9A",X"82",X"C3",X"12",X"0E",X"12",X"90",X"4C",X"4D",X"F1",X"A4",X"12",X"2D",
		X"D2",X"0A",X"64",X"C2",X"6C",X"0F",X"66",X"CD",X"82",X"6C",X"9A",X"C3",X"4A",X"85",X"C0",X"A6",
		X"6E",X"60",X"6C",X"9E",X"0A",X"C2",X"42",X"C4",X"C2",X"BA",X"60",X"49",X"F0",X"0C",X"12",X"C6",
		X"12",X"B0",X"00",X"A6",X"6E",X"60",X"58",X"ED",X"12",X"B5",X"E8",X"29",X"D2",X"0E",X"D8",X"4C",
		X"82",X"82",X"70",X"C2",X"6C",X"0B",X"6E",X"09",X"E6",X"B5",X"92",X"3E",X"00",X"A6",X"6E",X"60",
		X"6E",X"C1",X"6C",X"C0",X"00",X"59",X"62",X"48",X"66",X"D2",X"6D",X"18",X"4E",X"9B",X"64",X"09",
		X"02",X"A4",X"0A",X"ED",X"C0",X"18",X"4E",X"9B",X"64",X"08",X"C2",X"A4",X"0A",X"E8",X"00",X"20",
		X"4E",X"9B",X"64",X"B8",X"46",X"0D",X"20",X"2F",X"40",X"00",X"03",X"06",X"09",X"0C",X"10",X"13",
		X"16",X"19",X"1C",X"1F",X"22",X"25",X"28",X"2B",X"2E",X"31",X"33",X"36",X"39",X"3C",X"3F",X"41",
		X"44",X"47",X"49",X"4C",X"4E",X"51",X"53",X"55",X"58",X"5A",X"5C",X"5E",X"60",X"62",X"64",X"66",
		X"68",X"6A",X"6B",X"6D",X"6F",X"70",X"71",X"73",X"74",X"75",X"76",X"78",X"79",X"7A",X"7A",X"7B",
		X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
