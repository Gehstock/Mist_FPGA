library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"A2",X"AA",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A2",X"AA",X"A2",X"AA",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"3F",X"FF",X"30",X"0F",X"30",X"03",X"30",X"03",X"30",X"03",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"FF",X"3C",X"FF",X"00",X"00",
		X"00",X"00",X"03",X"FF",X"3F",X"FF",X"33",X"03",X"30",X"03",X"30",X"03",X"30",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"30",X"3F",X"FF",X"30",X"3F",X"30",X"30",X"30",X"30",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"30",X"FF",X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"CF",X"00",X"00",
		X"00",X"00",X"3C",X"FF",X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"30",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"3F",X"FF",X"30",X"C3",X"30",X"C3",X"3F",X"C3",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"30",X"FF",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"3F",X"C0",X"00",X"00",
		X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"8A",X"AA",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"8A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",
		X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"8A",X"AA",X"8A",X"AA",
		X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"FF",X"3F",X"C0",X"30",X"C0",X"30",X"C0",X"3F",X"FF",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"3F",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3C",X"0F",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3C",X"FF",X"30",X"C3",X"30",X"03",X"30",X"03",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"3F",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"3F",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"30",X"00",X"3F",X"FF",X"30",X"00",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"3F",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"30",X"3F",X"30",X"03",X"30",X"03",X"30",X"03",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"3F",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3C",X"FF",X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"CF",X"00",X"00",
		X"00",X"00",X"30",X"00",X"30",X"00",X"30",X"FF",X"3F",X"FF",X"30",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"00",X"00",X"FF",X"00",X"03",X"00",X"03",X"3F",X"FF",X"3F",X"C0",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"00",X"03",X"3F",X"FF",X"00",X"03",X"00",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"3F",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"00",X"00",X"C0",X"00",X"FF",X"00",X"FF",X"00",X"C0",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"0F",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"FF",X"3C",X"FF",X"00",X"00",
		X"AA",X"AA",X"A8",X"00",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"2A",X"AA",X"8A",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A2",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A8",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"A2",X"AA",X"A8",X"2A",X"AA",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"82",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"0F",X"00",X"03",
		X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FC",X"FF",X"3C",X"FF",X"0C",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"0F",X"00",X"03",
		X"00",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"00",
		X"FF",X"CF",X"FF",X"CF",X"FF",X"CF",X"FF",X"CF",X"FF",X"CF",X"FF",X"C0",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"00",X"0F",X"3F",X"CF",X"FF",X"CF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"3F",X"FF",X"3C",X"FF",X"30",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"C0",X"00",
		X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"00",X"3F",
		X"FF",X"F3",X"FF",X"F3",X"FF",X"F0",X"FF",X"F3",X"FF",X"F3",X"00",X"03",X"FF",X"3F",X"FF",X"3F",
		X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F3",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F3",X"FF",X"F3",X"FC",X"F3",X"F0",X"F0",X"00",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"C0",X"00",
		X"C0",X"00",X"F0",X"00",X"3C",X"00",X"3F",X"00",X"3F",X"C0",X"03",X"F0",X"F3",X"FC",X"F3",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"FF",X"FF",X"FF",X"FF",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",
		X"00",X"00",X"40",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"55",X"50",
		X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FD",X"7F",X"FD",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FD",X"7F",X"FD",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"AA",
		X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",
		X"03",X"FF",X"C0",X"3F",X"F0",X"03",X"FF",X"00",X"FF",X"C0",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"3F",X"FF",
		X"A0",X"00",X"AA",X"C0",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",
		X"FF",X"FF",X"3F",X"FD",X"0F",X"F5",X"C3",X"D5",X"F0",X"55",X"F1",X"55",X"F5",X"55",X"D5",X"55",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"AA",X"A8",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"80",X"AA",X"A8",X"0A",X"AA",X"00",X"AA",X"A0",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"F0",X"AF",X"FC",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"AA",X"80",X"AA",X"A0",X"2A",X"A8",X"0A",X"AA",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"54",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"55",X"00",
		X"0F",X"FF",X"C3",X"FD",X"F0",X"F5",X"FC",X"15",X"FC",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"55",X"55",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"00",X"00",X"00",X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"2A",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"40",X"55",X"40",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"80",X"02",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"40",X"00",X"00",X"00",
		X"55",X"50",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"55",X"50",
		X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"40",X"55",X"00",
		X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"02",X"55",X"0A",X"55",X"42",X"55",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"50",X"00",X"40",X"00",X"40",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"05",X"01",X"5F",X"07",X"F5",X"1D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"05",X"01",X"5F",X"07",X"FF",X"1F",X"FF",X"7F",X"FF",X"7F",X"FD",X"55",X"55",X"55",X"55",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"D5",X"55",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"55",X"55",X"00",X"00",X"00",X"00",
		X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"55",X"55",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"EA",X"A9",X"EA",X"A9",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",
		X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"55",X"55",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"FD",X"FF",X"FD",
		X"F0",X"40",X"F1",X"00",X"F4",X"00",X"D0",X"00",X"50",X"00",X"55",X"55",X"70",X"5B",X"70",X"5B",
		X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"59",X"F0",X"55",X"F0",X"54",X"F0",X"50",X"F0",X"40",
		X"D4",X"00",X"D0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"D0",X"FF",X"40",X"FD",X"00",X"FD",X"00",X"F4",X"00",
		X"00",X"7D",X"01",X"7D",X"01",X"FD",X"07",X"FD",X"1F",X"FD",X"5F",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"FF",X"40",X"FD",X"00",X"F4",X"00",X"D0",X"00",X"40",X"00",X"00",X"01",X"00",X"05",X"00",X"1D",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"D5",X"FD",X"50",X"F5",X"00",X"D4",X"00",X"50",X"00",X"40",X"00",
		X"03",X"AA",X"00",X"EA",X"00",X"3A",X"00",X"0E",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"15",X"AA",X"01",X"55",
		X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"55",X"F0",X"54",X"55",X"40",
		X"F0",X"5B",X"F0",X"5B",X"FC",X"5B",X"03",X"DB",X"00",X"FB",X"00",X"3B",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"3B",X"00",X"FB",X"01",X"DB",X"54",X"5B",X"F0",X"5B",X"F0",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"D0",X"00",X"F4",X"00",X"FD",X"00",X"FF",X"40",
		X"FF",X"40",X"FF",X"D0",X"FF",X"D0",X"FF",X"F4",X"FF",X"F4",X"FF",X"F4",X"FF",X"FD",X"FF",X"FD",
		X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"55",X"55",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"A9",X"EA",X"AA",X"EA",X"AA",
		X"EA",X"AA",X"EA",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"0E",X"AA",X"0E",X"AA",X"03",X"AA",
		X"01",X"AA",X"06",X"AA",X"06",X"AA",X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"03",X"AA",X"00",X"EA",X"00",X"3A",X"00",X"0E",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"06",X"00",X"1A",X"00",X"6A",X"01",X"AA",
		X"00",X"3A",X"00",X"3A",X"00",X"EA",X"03",X"AA",X"0E",X"AA",X"3A",X"AA",X"FA",X"AA",X"F5",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0E",
		X"EA",X"AA",X"EA",X"AA",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",X"F0",X"5B",
		X"F0",X"5B",X"F0",X"5B",X"70",X"59",X"F0",X"54",X"F0",X"54",X"F0",X"50",X"F0",X"40",X"F1",X"00",
		X"D0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"00",X"F4",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0D",X"00",X"39",X"00",X"39",
		X"00",X"E9",X"03",X"A9",X"0E",X"A9",X"3A",X"A9",X"3A",X"A9",X"EA",X"A9",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"F0",X"5B",X"F0",X"5B",
		X"55",X"55",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"FF",X"F5",X"FF",X"F4",X"FF",X"D0",X"FF",X"40",X"FD",X"00",X"F4",X"00",X"F4",X"00",
		X"55",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"40",X"00",X"10",X"00",X"04",X"00",X"01",X"00",X"00",X"40",X"00",X"10",X"00",X"04",X"00",X"01",
		X"01",X"55",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"AA",X"AA",
		X"80",X"00",X"20",X"00",X"08",X"00",X"02",X"00",X"00",X"80",X"00",X"20",X"00",X"08",X"00",X"02",
		X"80",X"02",X"20",X"08",X"08",X"20",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"FF",X"00",X"C3",X"00",X"C3",X"00",X"C3",X"00",X"C3",X"00",X"C3",X"00",X"C3",X"00",X"C3",X"00",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"30",X"00",X"0C",X"00",X"03",X"FF",
		X"C3",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"00",X"40",X"00",X"40",X"00",X"40",X"01",X"00",X"01",X"00",X"01",X"00",X"04",X"00",X"04",X"00",
		X"C0",X"00",X"30",X"00",X"0C",X"00",X"03",X"00",X"00",X"C0",X"00",X"30",X"00",X"0C",X"00",X"03",
		X"00",X"03",X"00",X"0F",X"00",X"33",X"00",X"C3",X"03",X"03",X"0C",X"03",X"30",X"03",X"C0",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"55",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"40",X"00",X"10",X"00",X"04",X"00",X"01",X"00",X"00",X"40",X"00",X"10",X"00",X"04",X"00",X"01",
		X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"1B",X"00",X"5B",X"01",X"5B",X"01",X"5B",X"04",X"5B",X"10",X"5B",X"50",X"5B",
		X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FD",X"50",X"F5",X"00",X"D4",X"00",X"D0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"F0",X"5B",X"F0",X"5B",
		X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"55",X"55",X"55",X"55",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"55",X"55",X"55",X"55",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7F",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7F",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"03",X"0C",X"3F",X"FF",X"F0",X"FF",X"F0",X"0C",X"3F",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"28",X"00",X"28",X"00",X"A8",X"02",X"A8",X"0A",X"A8",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"A8",X"00",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"14",X"00",X"01",X"55",
		X"10",X"00",X"10",X"00",X"10",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"01",X"00",X"01",X"00",
		X"01",X"40",X"00",X"40",X"00",X"10",X"00",X"14",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"10",X"00",X"10",X"55",X"55",X"00",X"10",X"55",X"55",X"00",X"10",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"14",X"00",X"55",X"05",X"00",X"50",X"00",
		X"01",X"10",X"01",X"10",X"01",X"10",X"04",X"10",X"04",X"10",X"04",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",
		X"80",X"00",X"20",X"00",X"08",X"00",X"02",X"00",X"00",X"80",X"00",X"20",X"00",X"08",X"00",X"02",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"C0",X"00",X"30",X"00",X"0C",X"00",X"03",X"00",X"00",X"C0",X"00",X"30",X"00",X"0C",X"00",X"03",
		X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",
		X"50",X"10",X"40",X"10",X"00",X"10",X"55",X"55",X"00",X"10",X"55",X"55",X"00",X"10",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"C0",X"03",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"C3",X"C3",X"C0",X"03",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"15",X"55",X"15",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"15",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",X"05",X"55",X"00",X"15",X"00",X"15",
		X"00",X"01",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"15",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"30",X"0C",X"30",X"00",X"00",
		X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"05",X"50",X"05",X"55",X"55",X"55",X"55",
		X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",
		X"55",X"55",X"55",X"55",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",
		X"50",X"50",X"50",X"50",X"50",X"55",X"50",X"55",X"50",X"05",X"50",X"05",X"55",X"55",X"55",X"55",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"00",X"55",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",X"50",X"50",X"50",X"50",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"55",X"50",
		X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"00",X"50",X"00",X"55",X"55",X"55",X"55",
		X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"00",X"55",X"00",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"55",
		X"55",X"55",X"55",X"55",X"50",X"55",X"50",X"55",X"00",X"00",X"00",X"00",X"50",X"00",X"50",X"00",
		X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"00",X"05",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"05",X"50",
		X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"50",X"55",X"50",X"55",X"50",X"00",X"50",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"55",X"50",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"55",X"50",
		X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FD",X"7F",X"FD",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FD",X"7F",X"FD",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"AA",
		X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",
		X"03",X"FF",X"C0",X"3F",X"F0",X"03",X"FF",X"00",X"FF",X"C0",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"3F",X"FF",
		X"A0",X"00",X"AA",X"C0",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",
		X"FF",X"FF",X"3F",X"FD",X"0F",X"F5",X"C3",X"D5",X"F0",X"55",X"F1",X"55",X"F5",X"55",X"D5",X"55",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"AA",X"A8",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"80",X"AA",X"A8",X"0A",X"AA",X"00",X"AA",X"A0",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"F0",X"AF",X"FC",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"AA",X"80",X"AA",X"A0",X"2A",X"A8",X"0A",X"AA",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"54",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"55",X"00",
		X"0F",X"FF",X"C3",X"FD",X"F0",X"F5",X"FC",X"15",X"FC",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"55",X"55",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"00",X"00",X"00",X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"2A",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"40",X"55",X"40",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"80",X"02",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"40",X"00",X"00",X"00",
		X"55",X"50",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"55",X"50",
		X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"40",X"55",X"00",
		X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"02",X"55",X"0A",X"55",X"42",X"55",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"50",X"00",X"40",X"00",X"40",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"05",X"01",X"5F",X"07",X"F5",X"1D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"05",X"01",X"5F",X"07",X"FF",X"1F",X"FF",X"7F",X"FF",X"7F",X"FD",X"55",X"55",X"55",X"55",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
