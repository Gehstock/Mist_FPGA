library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity F7 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of F7 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"3C",X"18",X"18",X"FF",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"18",X"18",X"7E",X"7E",X"BD",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"18",X"18",X"FF",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"99",X"18",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"4C",X"3E",X"3E",X"FE",X"7C",X"B8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"4C",X"3E",X"3E",X"FE",X"7C",X"B8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"18",X"9C",X"FE",X"FE",X"9C",X"18",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"18",X"9C",X"FE",X"FE",X"9C",X"18",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"30",X"F2",X"FF",X"F2",X"30",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"22",X"11",X"22",X"44",X"68",X"A0",X"3C",X"A0",X"68",X"44",X"22",X"11",X"22",X"44",X"00",
		X"90",X"48",X"24",X"24",X"44",X"68",X"E0",X"3C",X"A0",X"68",X"44",X"24",X"24",X"48",X"90",X"00",
		X"90",X"48",X"24",X"24",X"44",X"68",X"A0",X"3C",X"A0",X"68",X"44",X"24",X"24",X"48",X"90",X"00",
		X"10",X"88",X"44",X"33",X"44",X"68",X"E0",X"3C",X"A0",X"68",X"44",X"33",X"44",X"88",X"10",X"00",
		X"00",X"00",X"00",X"18",X"18",X"98",X"7F",X"8F",X"7F",X"1E",X"7C",X"B8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"18",X"18",X"6F",X"9F",X"2F",X"5E",X"BC",X"78",X"00",X"00",X"00",X"00",
		X"22",X"55",X"BE",X"74",X"02",X"61",X"C2",X"74",X"36",X"43",X"E0",X"40",X"36",X"7D",X"AE",X"44",
		X"14",X"94",X"42",X"F1",X"42",X"94",X"34",X"3C",X"3C",X"34",X"94",X"42",X"F1",X"42",X"94",X"14",
		X"00",X"24",X"4A",X"34",X"34",X"0C",X"3E",X"75",X"6D",X"2A",X"1C",X"34",X"34",X"4A",X"24",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"3C",X"1C",X"1C",X"1E",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"98",X"50",X"34",X"3C",X"3C",X"3C",X"3F",X"3E",X"3C",X"7C",X"BC",X"3C",X"7C",X"B8",X"98",
		X"00",X"86",X"FC",X"05",X"0F",X"0F",X"0F",X"7F",X"8F",X"8F",X"0F",X"1F",X"EF",X"8F",X"0E",X"06",
		X"01",X"06",X"0D",X"08",X"08",X"7C",X"FF",X"FC",X"F8",X"C8",X"CD",X"C6",X"C1",X"CC",X"E4",X"7C",
		X"01",X"06",X"0D",X"08",X"7C",X"FF",X"FC",X"C8",X"CD",X"C6",X"E1",X"60",X"30",X"18",X"44",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"A8",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"E8",X"A8",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"B1",X"42",X"81",X"02",X"00",X"29",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"59",X"96",X"01",X"83",X"82",X"84",X"EA",X"31",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7C",X"FE",X"7F",X"3E",X"7F",X"FE",X"7C",X"7E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"42",X"81",X"81",X"81",X"81",X"42",X"3C",
		X"3C",X"42",X"81",X"81",X"81",X"81",X"42",X"3C",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"30",X"F2",X"FF",X"F2",X"30",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"06",X"0F",X"03",X"0F",X"07",X"0E",X"0C",X"1C",X"0E",X"3F",X"0F",X"1F",X"0F",X"1E",X"0C",
		X"1C",X"0E",X"3F",X"7F",X"3F",X"3F",X"1E",X"1C",X"1C",X"1E",X"FF",X"FF",X"FF",X"FF",X"1E",X"1C",
		X"00",X"04",X"0E",X"02",X"0E",X"06",X"0C",X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0E",X"0C",X"00",
		X"00",X"0C",X"0E",X"6E",X"2E",X"0E",X"0C",X"00",X"00",X"0C",X"0E",X"6E",X"6E",X"0E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"18",X"18",X"7E",X"FF",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"18",X"18",X"7E",X"FF",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"18",X"99",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"18",X"99",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"4D",X"3E",X"3E",X"FE",X"7C",X"38",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"4D",X"3E",X"3E",X"FE",X"7C",X"38",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"18",X"9C",X"FE",X"FE",X"9C",X"18",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"18",X"9C",X"FE",X"FE",X"9C",X"18",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"22",X"22",X"22",X"44",X"68",X"A0",X"3C",X"E0",X"68",X"44",X"22",X"22",X"22",X"44",X"00",
		X"40",X"20",X"90",X"88",X"68",X"68",X"E0",X"3C",X"E0",X"68",X"68",X"88",X"90",X"20",X"40",X"00",
		X"44",X"22",X"22",X"22",X"44",X"68",X"A0",X"3C",X"E0",X"68",X"44",X"22",X"22",X"22",X"44",X"00",
		X"20",X"10",X"88",X"64",X"47",X"68",X"E0",X"3C",X"E0",X"68",X"47",X"64",X"88",X"10",X"20",X"00",
		X"00",X"00",X"00",X"18",X"18",X"D8",X"2F",X"9F",X"4F",X"3E",X"BC",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"18",X"18",X"7F",X"8F",X"3F",X"DE",X"3C",X"F8",X"00",X"00",X"00",X"00",
		X"34",X"42",X"E9",X"42",X"34",X"1C",X"36",X"43",X"E9",X"42",X"34",X"34",X"42",X"E9",X"42",X"34",
		X"28",X"66",X"DA",X"5D",X"BE",X"4C",X"7B",X"36",X"36",X"7B",X"4E",X"BE",X"1D",X"DA",X"66",X"14",
		X"00",X"00",X"08",X"10",X"1C",X"3E",X"31",X"74",X"2E",X"1C",X"7C",X"38",X"08",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"30",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"8C",X"68",X"1A",X"1E",X"1E",X"1E",X"1F",X"7E",X"9E",X"9E",X"1E",X"FE",X"9E",X"9C",X"8C",
		X"80",X"B0",X"A0",X"68",X"78",X"78",X"78",X"7E",X"7A",X"7A",X"FC",X"78",X"78",X"F8",X"F8",X"B0",
		X"01",X"06",X"0D",X"18",X"10",X"7C",X"FF",X"FC",X"D0",X"D8",X"CD",X"C6",X"E1",X"7C",X"04",X"0C",
		X"01",X"06",X"0D",X"08",X"7C",X"FF",X"FC",X"C8",X"CD",X"C6",X"C1",X"CC",X"D2",X"C4",X"CC",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"A8",X"B8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"E5",X"02",X"A2",X"85",X"20",X"63",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"36",X"DD",X"CF",X"67",X"46",X"FF",X"6E",X"A8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"7E",X"FE",X"6C",X"3E",X"7C",X"78",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
