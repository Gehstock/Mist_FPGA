library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bgscrn_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bgscrn_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"10",X"11",X"10",X"11",
		X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"13",X"12",X"13",
		X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"01",X"01",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"44",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"34",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"34",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"44",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"44",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"44",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"44",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"44",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"35",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"47",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"26",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"47",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"46",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"25",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"36",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"45",X"47",X"47",X"47",X"47",X"47",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",
		X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",
		X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",
		X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",X"56",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",
		X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",
		X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",X"57",X"54",
		X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",
		X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"65",X"04",X"27",X"75",X"27",X"2F",X"85",X"2F",X"37",X"95",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"51",X"53",X"04",X"64",X"04",X"27",X"74",X"27",X"2F",X"84",X"2F",X"37",X"94",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"50",X"52",X"04",X"63",X"04",X"27",X"73",X"27",X"2F",X"83",X"2F",X"37",X"93",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"49",X"48",X"04",X"62",X"04",X"27",X"72",X"27",X"2F",X"82",X"2F",X"37",X"92",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"4B",X"4A",X"04",X"62",X"04",X"27",X"72",X"27",X"2F",X"82",X"2F",X"37",X"92",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6F",X"01",X"01",X"01",X"01",
		X"01",X"14",X"16",X"04",X"61",X"04",X"27",X"71",X"27",X"2F",X"81",X"2F",X"37",X"92",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6E",X"01",X"01",X"01",X"01",
		X"01",X"15",X"17",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"91",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6D",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6C",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6B",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6A",X"01",X"1B",X"1A",X"44",
		X"45",X"51",X"53",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"01",X"19",X"18",X"46",
		X"47",X"50",X"52",X"04",X"65",X"04",X"27",X"75",X"27",X"2F",X"85",X"2F",X"37",X"95",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"68",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"64",X"04",X"27",X"74",X"27",X"2F",X"84",X"2F",X"37",X"94",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"67",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"04",X"63",X"04",X"27",X"73",X"27",X"2F",X"83",X"2F",X"37",X"93",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"66",X"01",X"01",X"01",X"01",
		X"01",X"41",X"43",X"04",X"62",X"04",X"27",X"72",X"27",X"2F",X"82",X"2F",X"37",X"92",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"40",X"42",X"04",X"62",X"04",X"27",X"72",X"27",X"2F",X"82",X"2F",X"37",X"92",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"49",X"48",X"04",X"60",X"04",X"27",X"70",X"27",X"2F",X"80",X"2F",X"37",X"90",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"4B",X"4A",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"14",X"16",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"15",X"17",X"04",X"04",X"04",X"27",X"27",X"27",X"2F",X"2F",X"2F",X"37",X"37",X"37",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"52",X"52",X"52",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
