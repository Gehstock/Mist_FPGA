library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_spr_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_spr_bit2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"7A",X"F2",X"00",X"10",X"1E",X"3F",X"71",X"EF",X"DF",X"5F",
		X"E2",X"72",X"04",X"00",X"00",X"00",X"00",X"00",X"5F",X"DF",X"EF",X"71",X"3F",X"1E",X"10",X"00",
		X"00",X"00",X"00",X"90",X"DA",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"7F",X"FC",X"DA",X"90",X"00",X"00",X"00",X"C2",X"98",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"7E",X"F8",X"F2",X"00",X"00",X"10",X"1F",X"3F",X"7F",X"EF",X"DF",
		X"62",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"5F",X"DF",X"7F",X"39",X"1F",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"96",X"DA",X"FD",X"FF",X"00",X"00",X"00",X"00",X"1E",X"1C",X"A2",X"C2",
		X"FF",X"FF",X"7F",X"FD",X"DA",X"90",X"00",X"00",X"C0",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"7D",X"CF",X"FC",X"F8",X"00",X"00",X"00",X"1F",X"AC",X"1F",X"77",X"63",
		X"70",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"DF",X"FF",X"7F",X"7F",X"FE",X"7F",X"1E",X"00",
		X"00",X"00",X"05",X"DF",X"26",X"37",X"98",X"FF",X"00",X"00",X"F0",X"FC",X"FE",X"6E",X"7A",X"B8",
		X"FF",X"FF",X"FF",X"FC",X"F0",X"80",X"00",X"00",X"C2",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"71",X"44",X"CE",X"C7",X"F0",X"7E",X"00",X"00",X"C0",X"5F",X"E0",X"0E",X"7F",X"3F",
		X"78",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"7B",X"E3",X"5F",X"FF",X"7F",X"3F",X"3F",X"1E",
		X"01",X"0F",X"0C",X"FF",X"1C",X"2F",X"17",X"FA",X"F0",X"1C",X"44",X"3E",X"5E",X"9E",X"F4",X"78",
		X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"00",X"00",X"A8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"71",X"44",X"CE",X"C7",X"F0",X"7E",X"00",X"00",X"C0",X"5F",X"E0",X"0E",X"7F",X"3F",
		X"78",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"7B",X"E3",X"5F",X"FF",X"7F",X"3F",X"3F",X"1E",
		X"01",X"0F",X"0C",X"FF",X"1C",X"2F",X"17",X"FA",X"F0",X"1C",X"44",X"3E",X"5E",X"9E",X"F4",X"78",
		X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"00",X"00",X"A8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"08",X"1C",X"38",X"4F",X"67",X"63",X"70",X"3F",X"9D",X"C0",X"00",
		X"3E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"7A",X"F2",X"00",X"13",X"1F",X"3D",X"70",X"E7",X"CF",X"4F",
		X"E2",X"72",X"04",X"00",X"00",X"00",X"00",X"00",X"4F",X"CF",X"E7",X"70",X"3D",X"1F",X"13",X"00",
		X"00",X"00",X"80",X"F0",X"FA",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"DF",X"FD",X"FA",X"F0",X"80",X"00",X"00",X"C2",X"88",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"7A",X"F2",X"00",X"13",X"1F",X"3D",X"70",X"E7",X"CF",X"4F",
		X"E2",X"72",X"04",X"00",X"00",X"00",X"00",X"00",X"4F",X"CF",X"E7",X"70",X"3D",X"1F",X"13",X"00",
		X"00",X"00",X"80",X"F0",X"FA",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"DF",X"FD",X"FA",X"F0",X"80",X"00",X"00",X"C2",X"88",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"7A",X"F2",X"00",X"13",X"1F",X"3F",X"70",X"EF",X"DF",X"5F",
		X"E2",X"72",X"04",X"00",X"00",X"00",X"00",X"00",X"5F",X"DF",X"EF",X"70",X"3F",X"1F",X"13",X"00",
		X"00",X"00",X"80",X"D0",X"DA",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"BF",X"FD",X"DA",X"D0",X"80",X"00",X"00",X"C2",X"88",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"7A",X"00",X"13",X"1F",X"3F",X"70",X"EF",X"DF",X"5F",
		X"72",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"DF",X"EF",X"70",X"3F",X"1F",X"13",X"00",
		X"00",X"00",X"80",X"D0",X"DA",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"BF",X"FD",X"DA",X"D0",X"80",X"00",X"00",X"C2",X"88",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"7A",X"F2",X"00",X"13",X"1F",X"3D",X"70",X"E7",X"CF",X"4F",
		X"E2",X"72",X"04",X"00",X"00",X"00",X"00",X"00",X"4F",X"CF",X"E7",X"70",X"3D",X"1F",X"13",X"00",
		X"00",X"00",X"80",X"F0",X"FA",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"DF",X"FD",X"FA",X"F0",X"80",X"00",X"00",X"C2",X"88",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"4E",X"3F",X"73",X"71",X"E7",X"CF",
		X"1A",X"72",X"E2",X"E0",X"70",X"00",X"00",X"00",X"4F",X"4F",X"CF",X"E7",X"70",X"39",X"1F",X"17",
		X"00",X"00",X"00",X"90",X"DA",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"FF",X"DF",X"F7",X"EC",X"C8",X"80",X"00",X"C2",X"88",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"01",X"08",X"3A",X"7B",X"5F",X"7B",X"E7",X"CF",X"CF",X"EF",X"6F",X"76",
		X"00",X"00",X"00",X"00",X"00",X"08",X"5F",X"FB",X"00",X"00",X"00",X"00",X"30",X"D8",X"0C",X"C4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DE",X"FB",X"F2",X"C4",X"C8",X"80",X"C0",X"00",X"00",X"00",X"00",
		X"71",X"79",X"30",X"00",X"00",X"00",X"00",X"00",X"78",X"3F",X"07",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"37",X"27",X"2F",
		X"00",X"00",X"00",X"01",X"02",X"00",X"09",X"37",X"00",X"40",X"B8",X"18",X"08",X"84",X"08",X"90",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"C0",X"80",X"80",X"80",X"80",X"80",X"00",X"80",
		X"00",X"00",X"00",X"00",X"05",X"08",X"1C",X"38",X"6F",X"67",X"63",X"70",X"3F",X"9D",X"C0",X"00",
		X"3E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F0",X"60",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"7A",X"00",X"10",X"1E",X"3F",X"71",X"EF",X"DF",X"5F",
		X"72",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"DF",X"EF",X"71",X"3F",X"1E",X"10",X"00",
		X"00",X"00",X"00",X"90",X"DA",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E8",X"C2",
		X"FF",X"7F",X"FC",X"DA",X"90",X"00",X"00",X"00",X"C2",X"98",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"7D",X"7F",X"7F",X"3E",X"0F",X"3F",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"80",
		X"7F",X"67",X"03",X"2E",X"36",X"08",X"1C",X"0E",X"60",X"F0",X"78",X"78",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"08",X"1C",X"38",X"4F",X"67",X"63",X"70",X"3F",X"9D",X"C0",X"00",
		X"3E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"3F",X"3F",X"3F",X"38",X"3F",X"3F",X"00",X"F8",X"FC",X"FC",X"FC",X"1C",X"FC",X"FC",
		X"3F",X"3F",X"38",X"3F",X"3F",X"3F",X"3F",X"38",X"FC",X"FC",X"1C",X"FC",X"FC",X"FC",X"FC",X"1C",
		X"3F",X"3F",X"3F",X"3F",X"38",X"3F",X"3F",X"3F",X"FC",X"FC",X"FC",X"FC",X"1C",X"FC",X"FC",X"FC",
		X"3F",X"38",X"7F",X"7F",X"7F",X"7F",X"7F",X"38",X"FC",X"1C",X"FC",X"FC",X"FC",X"FC",X"FC",X"1C",
		X"3F",X"3F",X"3F",X"3F",X"38",X"3F",X"3F",X"3F",X"FC",X"FC",X"FC",X"FC",X"1C",X"FC",X"FC",X"FC",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"FC",X"FC",X"9C",X"9C",X"9C",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"38",X"3F",X"3F",X"3F",X"FC",X"FC",X"FC",X"FC",X"1C",X"FC",X"FC",X"FC",
		X"3F",X"3F",X"3B",X"3B",X"39",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",
		X"00",X"03",X"47",X"BF",X"FA",X"B3",X"E7",X"AF",X"00",X"FE",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"87",X"B8",X"E0",X"E7",X"EF",X"CF",X"FE",X"FD",X"CF",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"F8",X"CF",X"83",X"B3",X"AB",X"00",X"00",X"FF",X"18",X"FF",X"FF",X"FF",X"FF",
		X"A3",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"0F",X"FF",X"F9",X"E1",X"EB",X"00",X"80",X"FE",X"D9",X"C7",X"3F",X"FF",X"FF",
		X"E3",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FD",
		X"00",X"03",X"07",X"7F",X"1E",X"01",X"3F",X"3F",X"00",X"FE",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",
		X"7F",X"31",X"0C",X"41",X"4F",X"5F",X"7F",X"5F",X"C0",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FE",X"CF",X"82",X"B2",X"AA",X"00",X"00",X"FF",X"B8",X"DF",X"1F",X"DE",X"9F",
		X"A2",X"82",X"82",X"82",X"82",X"83",X"83",X"83",X"1F",X"1F",X"1F",X"1D",X"1F",X"FF",X"FE",X"FD",
		X"00",X"FF",X"FF",X"1F",X"FF",X"F9",X"20",X"AA",X"00",X"80",X"FE",X"DD",X"C7",X"3F",X"FF",X"FF",
		X"E2",X"E0",X"E0",X"E0",X"E0",X"E0",X"60",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"87",X"87",X"87",X"85",X"86",X"85",X"86",X"A5",X"FD",X"FE",X"FF",X"F7",X"4D",X"17",X"0F",X"17",
		X"AE",X"B5",X"86",X"CD",X"FE",X"FF",X"00",X"00",X"8F",X"F6",X"AF",X"57",X"B8",X"FF",X"00",X"00",
		X"A0",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E2",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"20",X"F9",X"FF",X"1F",X"FF",X"FF",X"00",X"FF",X"FF",X"3F",X"C7",X"DD",X"FE",X"80",X"00",
		X"5F",X"7F",X"5F",X"4F",X"41",X"0C",X"31",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"C0",
		X"3F",X"3F",X"01",X"1E",X"7F",X"07",X"03",X"00",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FE",X"00",
		X"00",X"00",X"00",X"03",X"07",X"1F",X"39",X"3B",X"00",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"79",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"40",X"FF",X"E4",X"F4",X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"21",X"2F",
		X"FF",X"7F",X"9F",X"DF",X"3F",X"1F",X"1F",X"1F",X"FF",X"FF",X"F5",X"F9",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"F0",X"F8",X"FE",X"FD",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"6F",X"47",X"C7",
		X"00",X"00",X"01",X"03",X"01",X"01",X"01",X"01",X"88",X"87",X"8F",X"9F",X"1F",X"0F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"F1",X"FF",
		X"FF",X"F9",X"ED",X"EF",X"ED",X"FD",X"FD",X"FD",X"27",X"FF",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"E2",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"F0",X"3C",X"5C",X"FE",X"F6",X"F2",X"F2",X"80",X"80",X"C0",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"DF",X"BF",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"DF",X"DF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"A8",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"F2",X"F3",X"F3",X"F2",X"F2",X"F3",X"F3",X"F1",X"F9",X"F9",X"F9",X"F9",X"F1",X"FB",X"FF",
		X"00",X"00",X"00",X"D5",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"90",X"50",X"50",X"D0",
		X"BF",X"BF",X"DF",X"BF",X"BF",X"DF",X"BF",X"BF",X"F0",X"F0",X"F0",X"F0",X"F0",X"D0",X"50",X"50",
		X"00",X"03",X"47",X"BF",X"FA",X"B3",X"E7",X"AF",X"00",X"FE",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"87",X"B8",X"E0",X"E7",X"EF",X"EF",X"FE",X"FD",X"CF",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"F8",X"CF",X"83",X"B3",X"AB",X"00",X"00",X"FF",X"18",X"FF",X"FF",X"FF",X"FF",
		X"A3",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"0F",X"FF",X"F9",X"E1",X"EB",X"00",X"80",X"FE",X"D9",X"C7",X"3F",X"FF",X"FF",
		X"E3",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FD",
		X"00",X"03",X"07",X"7F",X"1E",X"01",X"3F",X"3F",X"00",X"FE",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",
		X"7F",X"31",X"0C",X"41",X"4F",X"5F",X"7F",X"5F",X"C0",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FE",X"CF",X"82",X"B2",X"AB",X"00",X"00",X"FF",X"B8",X"FF",X"4F",X"EE",X"FF",
		X"A2",X"83",X"82",X"83",X"82",X"83",X"83",X"83",X"EF",X"FF",X"EF",X"BD",X"0F",X"FF",X"FE",X"FD",
		X"00",X"FF",X"FF",X"1F",X"FF",X"F9",X"20",X"AA",X"00",X"80",X"FE",X"DD",X"C7",X"3F",X"FF",X"FF",
		X"E2",X"E0",X"E0",X"E0",X"E0",X"E0",X"60",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"A3",X"FD",X"FE",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",
		X"AB",X"B3",X"83",X"CF",X"FE",X"FF",X"00",X"00",X"7F",X"3E",X"FF",X"FF",X"B8",X"FF",X"00",X"00",
		X"A0",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E2",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"20",X"F9",X"FF",X"1F",X"FF",X"FF",X"00",X"FF",X"FF",X"3F",X"C7",X"DD",X"FE",X"80",X"00",
		X"5F",X"7F",X"5F",X"4F",X"41",X"0C",X"31",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"C0",
		X"3F",X"3F",X"01",X"1E",X"7F",X"07",X"03",X"00",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FE",X"00",
		X"00",X"00",X"00",X"03",X"07",X"1F",X"39",X"3B",X"00",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"79",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"40",X"FF",X"E4",X"F4",X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"21",X"2F",
		X"FF",X"7F",X"9F",X"DF",X"3F",X"1F",X"1F",X"1F",X"FF",X"FF",X"F5",X"F9",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"F0",X"F8",X"FE",X"FD",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"6F",X"47",X"C7",
		X"00",X"00",X"01",X"03",X"01",X"01",X"01",X"01",X"88",X"87",X"8F",X"9F",X"1F",X"0F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"F1",X"FF",
		X"FF",X"F9",X"ED",X"EF",X"ED",X"FD",X"FD",X"FD",X"27",X"FF",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"60",X"E0",X"E2",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"F0",X"3C",X"5C",X"FE",X"F6",X"F2",X"F2",X"80",X"80",X"C0",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"DF",X"BF",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"EF",X"EF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"48",X"FF",X"FF",X"FF",X"F3",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"F2",X"F3",X"F3",X"F2",X"F2",X"F3",X"F3",X"F1",X"F9",X"F9",X"F9",X"F9",X"F1",X"FB",X"FF",
		X"00",X"00",X"00",X"EA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"90",X"50",X"50",X"D0",
		X"BF",X"BF",X"DF",X"BF",X"BF",X"DF",X"BF",X"BF",X"F0",X"F0",X"F0",X"F0",X"F0",X"D0",X"50",X"50",
		X"00",X"01",X"03",X"10",X"26",X"37",X"27",X"27",X"00",X"FF",X"40",X"00",X"FB",X"00",X"40",X"67",
		X"37",X"27",X"27",X"27",X"27",X"27",X"37",X"37",X"0F",X"4F",X"6F",X"0F",X"4F",X"6F",X"0F",X"0F",
		X"10",X"8F",X"F0",X"60",X"61",X"63",X"66",X"E4",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"E4",X"E4",X"E4",X"E4",X"E4",X"E4",X"E4",X"E6",X"3E",X"63",X"40",X"40",X"60",X"3C",X"07",X"00",
		X"37",X"37",X"27",X"27",X"27",X"27",X"37",X"27",X"0F",X"0F",X"6F",X"4F",X"0F",X"6F",X"4F",X"0F",
		X"27",X"37",X"27",X"26",X"10",X"03",X"01",X"00",X"67",X"40",X"00",X"FB",X"00",X"00",X"FF",X"00",
		X"E3",X"E1",X"E0",X"E0",X"E7",X"E4",X"E4",X"E4",X"00",X"F0",X"1E",X"03",X"C1",X"41",X"63",X"3E",
		X"E4",X"E2",X"63",X"60",X"60",X"F0",X"9F",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",
		X"80",X"7F",X"00",X"00",X"C0",X"60",X"30",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"F0",X"01",X"03",X"C2",X"66",X"00",X"00",X"3F",X"E0",X"80",X"00",X"0E",X"1E",
		X"86",X"7F",X"00",X"00",X"03",X"03",X"03",X"03",X"01",X"FF",X"00",X"00",X"FF",X"F1",X"F1",X"F1",
		X"03",X"03",X"83",X"E3",X"63",X"33",X"13",X"13",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0E",X"3C",X"78",X"70",X"60",X"41",X"03",X"07",X"0E",
		X"1B",X"11",X"30",X"E0",X"80",X"00",X"FF",X"00",X"00",X"80",X"E0",X"3F",X"00",X"00",X"FF",X"00",
		X"1F",X"37",X"67",X"C7",X"C7",X"87",X"0F",X"0B",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"1B",X"33",X"E3",X"83",X"00",X"00",X"FF",X"06",X"F0",X"F0",X"F1",X"FF",X"00",X"00",X"FF",X"01",
		X"A3",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"FF",X"00",X"00",X"1F",X"11",X"11",X"11",
		X"00",X"00",X"FF",X"81",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"91",X"D1",X"51",X"71",X"31",
		X"A0",X"7F",X"00",X"00",X"01",X"01",X"01",X"01",X"34",X"FA",X"02",X"00",X"F0",X"12",X"10",X"10",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"10",X"10",X"12",X"10",X"10",X"12",X"10",
		X"7C",X"C6",X"82",X"82",X"82",X"82",X"86",X"FC",X"31",X"31",X"31",X"31",X"31",X"30",X"38",X"28",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"23",X"2C",X"66",X"C3",X"80",X"00",X"00",X"FF",X"61",
		X"01",X"01",X"01",X"01",X"81",X"81",X"E1",X"3F",X"10",X"12",X"10",X"10",X"12",X"10",X"10",X"12",
		X"00",X"00",X"80",X"FF",X"00",X"00",X"FF",X"20",X"10",X"10",X"12",X"F0",X"00",X"02",X"FE",X"30",
		X"00",X"01",X"03",X"10",X"26",X"37",X"27",X"27",X"00",X"FF",X"40",X"00",X"FB",X"00",X"00",X"27",
		X"37",X"27",X"27",X"27",X"27",X"27",X"37",X"37",X"0F",X"0F",X"2F",X"0F",X"0F",X"2F",X"0F",X"0F",
		X"37",X"37",X"27",X"27",X"27",X"27",X"37",X"27",X"0F",X"0F",X"2F",X"0F",X"0F",X"2F",X"0F",X"0F",
		X"27",X"37",X"27",X"26",X"10",X"03",X"01",X"00",X"27",X"00",X"00",X"FB",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"3C",X"7A",X"00",X"00",X"2F",X"3F",X"31",X"70",X"EF",X"DF",
		X"F2",X"E2",X"72",X"00",X"00",X"00",X"00",X"00",X"5F",X"5F",X"DF",X"EF",X"71",X"3F",X"1F",X"00",
		X"00",X"00",X"00",X"9E",X"E7",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"3E",X"04",X"E2",X"C2",
		X"FF",X"FF",X"BF",X"EE",X"CC",X"98",X"10",X"00",X"C0",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"BF",X"E3",
		X"00",X"01",X"3D",X"74",X"F4",X"E2",X"70",X"00",X"CF",X"9F",X"9F",X"9F",X"DF",X"EF",X"3F",X"1F",
		X"00",X"00",X"00",X"03",X"2F",X"F7",X"FF",X"FF",X"00",X"00",X"38",X"C6",X"82",X"C2",X"E0",X"C4",
		X"FF",X"FF",X"FF",X"FF",X"B4",X"E6",X"C4",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"06",X"18",X"70",X"41",X"E5",X"0C",X"6F",X"F7",X"31",X"4F",X"EF",X"9F",X"9F",
		X"00",X"01",X"03",X"07",X"3F",X"FE",X"B1",X"EF",X"38",X"FC",X"FC",X"E8",X"80",X"80",X"08",X"80",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FA",X"F0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E5",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"EF",X"43",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"06",X"18",X"70",X"41",X"E5",X"0C",X"6F",X"F7",X"31",X"4F",X"EF",X"9F",X"9F",
		X"E5",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"EF",X"43",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"7C",X"C6",X"86",X"93",X"39",X"79",X"9E",X"86",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"7E",X"02",X"02",X"00",X"00",X"08",X"08",
		X"00",X"00",X"00",X"00",X"1F",X"9F",X"80",X"80",X"00",X"01",X"03",X"09",X"C3",X"E6",X"7A",X"64",
		X"00",X"00",X"80",X"C0",X"61",X"33",X"1B",X"71",X"47",X"43",X"60",X"F8",X"FF",X"FF",X"E1",X"00",
		X"F8",X"CC",X"04",X"26",X"F6",X"F2",X"3E",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"BC",X"C4",X"6C",X"38",X"98",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"60",X"40",X"00",X"80",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"D8",X"98",X"38",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"20",X"67",X"4E",X"5E",X"64",X"20",X"33",X"A0",X"F0",X"80",X"40",X"47",X"80",X"80",X"80",
		X"1F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"0B",X"0B",X"0F",X"0F",X"0C",X"0C",X"0C",X"1C",X"1C",X"3E",X"3E",X"FE",X"0E",X"07",X"06",
		X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"04",X"1E",X"04",X"00",X"02",X"07",X"1D",X"39",X"21",X"00",
		X"00",X"00",X"00",X"00",X"04",X"1F",X"31",X"23",X"00",X"00",X"00",X"00",X"00",X"B8",X"90",X"96",
		X"67",X"4E",X"5E",X"6C",X"28",X"3A",X"1E",X"06",X"CD",X"59",X"33",X"67",X"6E",X"CE",X"CC",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"7C",X"E6",X"82",X"92",X"38",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"94",X"C3",X"C5",X"78",X"00",X"00",X"01",
		X"03",X"07",X"0D",X"18",X"30",X"20",X"00",X"00",X"30",X"FF",X"CF",X"80",X"81",X"7F",X"7E",X"7C",
		X"00",X"70",X"7C",X"99",X"82",X"06",X"0C",X"8C",X"F8",X"F0",X"E0",X"20",X"00",X"00",X"00",X"00",
		X"03",X"06",X"04",X"0C",X"09",X"0F",X"2E",X"74",X"E0",X"30",X"30",X"98",X"C8",X"F8",X"FC",X"10",
		X"CC",X"FF",X"73",X"20",X"20",X"1F",X"1F",X"1F",X"74",X"CC",X"FC",X"3C",X"40",X"FC",X"B8",X"00",
		X"88",X"80",X"3A",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"31",X"20",X"65",X"6F",X"4F",X"7C",X"70",X"00",X"80",X"C0",X"D0",X"D8",X"50",X"C4",X"9C",
		X"30",X"21",X"B7",X"AE",X"A8",X"F1",X"E3",X"E3",X"78",X"E6",X"9C",X"78",X"F0",X"C0",X"80",X"00",
		X"00",X"00",X"02",X"02",X"02",X"03",X"07",X"07",X"C1",X"87",X"DE",X"B9",X"A3",X"C7",X"8E",X"8C",
		X"0C",X"0C",X"18",X"18",X"30",X"30",X"00",X"00",X"5E",X"3E",X"1E",X"0C",X"0C",X"1C",X"10",X"00",
		X"03",X"03",X"07",X"04",X"00",X"C4",X"EC",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"08",X"04",X"01",X"07",X"C7",X"60",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"06",X"04",X"0C",X"06",X"0C",X"0C",X"80",X"E0",X"33",X"11",X"90",
		X"09",X"0D",X"0C",X"04",X"06",X"03",X"00",X"00",X"FC",X"FF",X"93",X"00",X"60",X"C0",X"80",X"00",
		X"FD",X"B4",X"BE",X"9A",X"1E",X"38",X"18",X"0C",X"E0",X"F8",X"FC",X"78",X"08",X"04",X"03",X"03",
		X"0C",X"06",X"06",X"00",X"00",X"00",X"01",X"01",X"06",X"1E",X"18",X"00",X"06",X"FC",X"88",X"18",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"C6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"0C",X"08",X"00",X"70",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"03",X"03",X"01",X"01",X"00",X"00",X"24",X"72",X"72",X"26",X"04",X"9C",X"F8",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"3E",X"77",X"47",X"CF",X"9C",X"00",X"00",X"88",X"6C",X"6C",X"6C",X"6C",X"6C",
		X"9C",X"CD",X"67",X"66",X"3F",X"0A",X"02",X"02",X"6C",X"36",X"B6",X"B7",X"F7",X"D3",X"FB",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"0B",X"0D",X"35",X"06",X"F2",X"CB",
		X"02",X"06",X"04",X"06",X"06",X"02",X"03",X"01",X"CB",X"69",X"E5",X"F4",X"59",X"0A",X"3F",X"F1",
		X"2C",X"BF",X"B7",X"BB",X"78",X"5C",X"9D",X"AF",X"00",X"80",X"F8",X"FC",X"C5",X"81",X"01",X"01",
		X"C6",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"C0",X"E0",X"30",X"11",X"03",X"02",
		X"00",X"0C",X"06",X"06",X"56",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"02",X"22",X"60",X"60",X"E0",X"D0",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D9",X"9C",X"9D",X"C9",X"61",X"63",X"3E",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"07",X"DF",X"DF",X"07",X"00",X"03",X"02",X"C0",X"F3",X"FC",X"FC",X"F3",X"C0",X"80",X"00",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"1F",X"7F",X"7F",X"7F",X"7F",X"3F",X"0F",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"F8",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FC",X"FF",X"FF",X"FF",X"FF",X"9F",X"8F",X"8E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"1F",X"7F",X"CB",X"FF",X"FE",X"0A",X"48",X"FD",X"D8",X"AE",X"E3",X"B3",X"2B",
		X"7C",X"38",X"34",X"1F",X"07",X"00",X"00",X"00",X"70",X"AA",X"17",X"97",X"DF",X"EF",X"77",X"3B",
		X"80",X"71",X"B9",X"89",X"53",X"FF",X"3F",X"15",X"C0",X"10",X"F0",X"F4",X"3F",X"7F",X"AB",X"5E",
		X"CA",X"F7",X"FF",X"F6",X"F7",X"F0",X"E5",X"E0",X"F5",X"C0",X"BA",X"EA",X"C0",X"20",X"00",X"10",
		X"04",X"00",X"00",X"1F",X"7D",X"CB",X"FF",X"FC",X"1C",X"58",X"91",X"53",X"FF",X"AE",X"75",X"3F",
		X"79",X"27",X"33",X"1F",X"06",X"01",X"00",X"00",X"5D",X"98",X"FF",X"3F",X"8F",X"E7",X"DF",X"3F",
		X"00",X"07",X"3F",X"F1",X"C7",X"7C",X"E1",X"DF",X"20",X"D8",X"F0",X"FC",X"7F",X"F7",X"FD",X"EA",
		X"9E",X"F6",X"FA",X"F3",X"F6",X"E5",X"FA",X"D4",X"F4",X"A0",X"31",X"90",X"EA",X"80",X"80",X"00",
		X"1F",X"3F",X"3F",X"3F",X"7F",X"FD",X"FF",X"FB",X"88",X"C0",X"C8",X"F3",X"F7",X"FF",X"EC",X"54",
		X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"7E",X"81",X"4B",X"3C",X"BA",X"D4",X"81",X"16",X"1E",
		X"1F",X"3F",X"3F",X"DE",X"FF",X"FE",X"B5",X"3B",X"00",X"80",X"80",X"20",X"D0",X"FE",X"BA",X"7C",
		X"7A",X"CB",X"BD",X"7F",X"E6",X"0D",X"1D",X"7F",X"FA",X"FA",X"FC",X"BC",X"FE",X"FE",X"BE",X"2E",
		X"7E",X"FF",X"FC",X"FF",X"FA",X"FE",X"FF",X"FF",X"DE",X"FE",X"27",X"AC",X"DA",X"FE",X"77",X"CB",
		X"FB",X"FF",X"FD",X"7F",X"3F",X"3F",X"3F",X"1F",X"EF",X"FE",X"FF",X"F7",X"F3",X"C0",X"C0",X"80",
		X"76",X"C5",X"2D",X"13",X"6F",X"85",X"41",X"38",X"2E",X"9E",X"EE",X"FA",X"FD",X"FD",X"FC",X"FE",
		X"9F",X"B7",X"EE",X"FF",X"5E",X"3F",X"3F",X"1F",X"6D",X"90",X"FC",X"F4",X"A0",X"80",X"80",X"00",
		X"1F",X"3F",X"3F",X"3F",X"7E",X"FD",X"FF",X"FB",X"98",X"C0",X"CB",X"DF",X"BA",X"B5",X"C2",X"DE",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FE",X"7D",X"BD",X"7F",X"BE",X"B8",X"DA",X"E7",X"EF",X"FF",
		X"1F",X"3F",X"3B",X"D6",X"BE",X"FF",X"A5",X"9B",X"00",X"80",X"80",X"30",X"E0",X"C6",X"88",X"5C",
		X"5A",X"3F",X"BD",X"7E",X"E5",X"0C",X"1B",X"7F",X"38",X"F8",X"2F",X"6E",X"D6",X"6E",X"DE",X"EA",
		X"71",X"F9",X"FF",X"FD",X"FC",X"F6",X"FF",X"FF",X"EF",X"DE",X"EF",X"FC",X"33",X"D2",X"40",X"B9",
		X"FA",X"FF",X"FC",X"7F",X"3F",X"3F",X"3F",X"1F",X"E4",X"76",X"FB",X"C5",X"E2",X"C0",X"C0",X"80",
		X"F8",X"FD",X"BF",X"FF",X"6D",X"91",X"D1",X"78",X"2E",X"96",X"CA",X"E0",X"FD",X"F8",X"FC",X"BC",
		X"EE",X"B7",X"FB",X"FD",X"5E",X"3F",X"3F",X"1F",X"4C",X"50",X"DC",X"C4",X"3A",X"88",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"3D",X"79",X"00",X"10",X"19",X"3C",X"B0",X"AF",X"FF",X"FF",
		X"71",X"39",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"AF",X"B0",X"33",X"1F",X"10",X"00",
		X"00",X"00",X"00",X"D8",X"6E",X"A7",X"DD",X"EB",X"00",X"00",X"00",X"00",X"1C",X"70",X"B8",X"C6",
		X"EB",X"DD",X"A7",X"6E",X"D8",X"00",X"00",X"00",X"C6",X"98",X"70",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"7C",X"FB",X"F1",X"00",X"00",X"10",X"1F",X"31",X"FE",X"AF",X"FF",
		X"61",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"AF",X"30",X"1B",X"17",X"00",
		X"00",X"00",X"00",X"18",X"9E",X"4E",X"B7",X"D9",X"00",X"00",X"00",X"00",X"7C",X"E0",X"BA",X"C6",
		X"EB",X"EB",X"D8",X"B6",X"5C",X"88",X"18",X"00",X"C4",X"90",X"1C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"7D",X"CB",X"FD",X"F8",X"00",X"00",X"00",X"00",X"D0",X"5F",X"31",X"BE",
		X"73",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"BF",X"FF",X"FF",X"FF",X"BF",X"1F",X"17",X"00",
		X"00",X"00",X"09",X"1F",X"7B",X"5B",X"CC",X"7D",X"00",X"00",X"F0",X"BC",X"BE",X"EE",X"7A",X"A4",
		X"BB",X"CB",X"E8",X"EA",X"94",X"44",X"00",X"00",X"C4",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"71",X"CE",X"C8",X"F1",X"7E",X"38",X"00",X"00",X"C0",X"60",X"43",X"0F",X"30",X"F6",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FF",X"BF",X"3F",X"1F",X"1F",X"0F",
		X"01",X"17",X"1F",X"7A",X"EC",X"3B",X"9C",X"FD",X"F0",X"1C",X"E6",X"66",X"1E",X"7C",X"C4",X"30",
		X"7B",X"9B",X"E8",X"EC",X"E8",X"80",X"00",X"00",X"C4",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"71",X"CE",X"C8",X"F1",X"7E",X"38",X"00",X"00",X"C0",X"60",X"43",X"0F",X"30",X"F6",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FF",X"BF",X"3F",X"1F",X"1F",X"0F",
		X"01",X"17",X"1F",X"7A",X"EC",X"3B",X"9C",X"FD",X"F0",X"1C",X"E6",X"66",X"1E",X"7C",X"C4",X"30",
		X"7B",X"9B",X"E8",X"EC",X"E8",X"80",X"00",X"00",X"C4",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"3D",X"79",X"00",X"10",X"19",X"3C",X"B0",X"AF",X"FF",X"FF",
		X"71",X"39",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"AF",X"B0",X"33",X"1F",X"10",X"00",
		X"00",X"00",X"00",X"D8",X"6E",X"A7",X"DD",X"EB",X"00",X"00",X"00",X"00",X"1C",X"70",X"98",X"C6",
		X"EB",X"DD",X"A7",X"6E",X"D8",X"00",X"00",X"00",X"C6",X"98",X"70",X"1C",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"1F",X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"1E",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"7F",X"7F",X"7F",X"7F",X"73",X"73",X"71",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"22",X"22",
		X"00",X"7F",X"74",X"00",X"00",X"E0",X"20",X"3F",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"09",X"09",X"09",X"09",X"09",
		X"00",X"00",X"FF",X"80",X"C0",X"F4",X"FF",X"00",X"09",X"09",X"F9",X"01",X"01",X"01",X"FF",X"00",
		X"74",X"40",X"40",X"00",X"00",X"7F",X"50",X"00",X"02",X"02",X"00",X"00",X"00",X"FE",X"02",X"02",
		X"18",X"71",X"74",X"00",X"00",X"7F",X"74",X"00",X"00",X"FE",X"02",X"02",X"00",X"FE",X"02",X"02",
		X"00",X"00",X"00",X"03",X"1E",X"F0",X"86",X"C3",X"00",X"0F",X"79",X"C1",X"01",X"07",X"1C",X"90",
		X"C3",X"F8",X"FA",X"1E",X"03",X"00",X"00",X"00",X"90",X"1C",X"07",X"01",X"C1",X"79",X"0F",X"00",
		X"00",X"3F",X"20",X"00",X"00",X"5F",X"34",X"00",X"00",X"FC",X"06",X"0A",X"0A",X"FA",X"02",X"00",
		X"00",X"3F",X"01",X"02",X"02",X"5E",X"74",X"00",X"00",X"00",X"80",X"80",X"80",X"FE",X"02",X"02",
		X"00",X"7F",X"C0",X"80",X"B0",X"BF",X"90",X"90",X"00",X"FE",X"03",X"01",X"01",X"F9",X"09",X"09",
		X"90",X"D0",X"9F",X"C0",X"E0",X"FA",X"7F",X"00",X"09",X"09",X"F9",X"01",X"01",X"03",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"78",X"1F",X"03",X"00",X"7F",X"74",X"00",X"1E",X"72",X"C2",X"00",X"00",X"7E",X"02",X"02",
		X"00",X"7F",X"C6",X"8E",X"9F",X"9E",X"93",X"93",X"00",X"FE",X"03",X"01",X"01",X"79",X"49",X"C9",
		X"93",X"D0",X"9F",X"C0",X"E0",X"FA",X"7F",X"00",X"C9",X"09",X"F9",X"01",X"01",X"03",X"FE",X"00",
		X"00",X"38",X"08",X"08",X"00",X"5F",X"34",X"00",X"00",X"1C",X"06",X"02",X"02",X"FA",X"02",X"00",
		X"00",X"60",X"21",X"20",X"20",X"60",X"74",X"00",X"00",X"06",X"82",X"82",X"82",X"82",X"02",X"02",
		X"00",X"7F",X"50",X"00",X"00",X"7E",X"74",X"00",X"00",X"FE",X"02",X"02",X"00",X"7E",X"02",X"02",
		X"00",X"38",X"08",X"08",X"00",X"5F",X"34",X"00",X"00",X"1C",X"06",X"02",X"02",X"FA",X"02",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"21",X"18",X"01",
		X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"07",X"1A",X"39",X"19",X"B3",X"F6",X"18",X"00",
		X"00",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"68",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"10",X"40",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"03",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"DF",X"06",X"23",X"13",X"B7",X"F6",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"68",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"08",X"03",X"04",X"0B",X"13",X"A0",X"40",X"0F",X"16",X"7F",X"1F",X"CF",X"E6",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"04",X"01",X"03",X"01",X"03",X"02",X"17",X"7F",X"1F",X"8F",X"C6",X"1C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"68",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"04",X"01",X"03",X"01",X"00",X"02",X"17",X"7F",X"1F",X"8F",X"C6",X"1C",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"0B",X"1B",X"10",X"32",X"24",X"17",X"7F",X"1F",X"CF",X"E6",X"18",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"0F",X"00",X"08",X"04",X"00",X"00",X"00",X"E0",X"E0",X"08",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",
		X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"34",X"18",X"B1",X"F3",X"F6",X"18",X"00",X"00",
		X"08",X"18",X"30",X"60",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"0F",X"00",X"00",X"04",X"00",X"00",X"00",X"E0",X"E0",X"08",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"36",X"1C",X"B0",X"F1",X"F6",X"18",X"00",X"00",
		X"00",X"00",X"0C",X"0C",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"0F",X"00",X"00",X"04",X"00",X"00",X"00",X"E0",X"E0",X"08",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",
		X"07",X"07",X"03",X"03",X"03",X"01",X"01",X"00",X"E0",X"E0",X"F0",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"F9",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",
		X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"C0",X"C0",
		X"1F",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"C0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"FF",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"7F",X"7E",X"7C",X"7E",X"3E",X"3F",X"3F",X"1F",
		X"FC",X"FF",X"FF",X"7F",X"3F",X"1F",X"07",X"00",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"1F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"8F",X"80",X"C0",X"C0",X"C0",X"F0",X"FF",X"FF",
		X"FF",X"0F",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"3F",X"00",X"0F",X"3F",X"3F",X"7F",
		X"07",X"00",X"00",X"80",X"FE",X"FF",X"FF",X"FF",X"F8",X"FC",X"FC",X"7E",X"7E",X"FE",X"FE",X"FE",
		X"FF",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FE",X"FC",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"80",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"FE",X"FE",X"7E",X"7E",X"3E",X"3C",X"10",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"FE",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"FC",X"FE",X"FF",X"22",X"23",X"A3",X"A1",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"38",X"28",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"20",X"20",X"22",X"23",X"23",X"23",X"23",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"21",X"21",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"21",X"3F",X"3F",X"3F",X"2F",X"23",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"22",X"23",X"23",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"38",X"38",X"28",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"21",X"21",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"21",X"21",X"21",X"23",X"23",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"21",X"21",X"21",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"2F",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"22",X"23",X"23",X"23",X"23",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"38",X"38",X"28",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"C0",X"81",X"01",X"22",X"00",X"20",X"00",X"40",X"00",X"80",X"00",X"00",
		X"36",X"3C",X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"60",X"C0",X"80",X"80",X"80",X"F0",X"FF",X"FF",X"70",X"18",X"0C",X"06",X"03",X"01",X"C1",X"FF",
		X"00",X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0F",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"1F",X"03",X"00",
		X"FE",X"03",X"00",X"00",X"00",X"80",X"F0",X"FF",X"00",X"F8",X"0F",X"00",X"00",X"00",X"00",X"C0",
		X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"80",X"F0",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"38",X"60",X"00",X"00",X"00",X"00",X"F8",X"0F",X"00",X"00",
		X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0F",X"00",X"00",X"00",
		X"FF",X"FC",X"F0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"07",X"07",X"05",X"04",X"04",X"04",X"07",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",
		X"00",X"C0",X"7E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0F",X"00",X"00",X"00",
		X"F0",X"FF",X"FF",X"3F",X"01",X"01",X"0F",X"3F",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"60",X"C0",X"80",X"80",X"80",X"F0",X"FF",X"FF",X"70",X"18",X"0C",X"06",X"03",X"01",X"C1",X"FF",
		X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"1F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E1",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",
		X"78",X"38",X"3C",X"1C",X"1C",X"0E",X"0E",X"0E",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",
		X"07",X"07",X"07",X"07",X"06",X"04",X"80",X"80",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"E0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",X"00",X"00",
		X"00",X"FC",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"F0",X"1E",X"03",X"00",X"00",X"00",X"00",X"F0",
		X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FC",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"E0",X"FE",X"FF",X"7F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"7C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C6",X"C7",X"E7",X"07",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",
		X"00",X"FC",X"FF",X"FF",X"0F",X"00",X"01",X"03",X"01",X"01",X"E1",X"E1",X"E1",X"60",X"E0",X"E0",
		X"83",X"87",X"C7",X"47",X"46",X"46",X"46",X"46",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"07",X"07",X"07",X"07",X"06",X"04",X"80",X"80",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E1",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"78",X"38",X"3C",X"1C",X"1C",X"0E",X"0E",X"0E",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"8C",X"84",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"30",X"FC",X"FC",X"BC",X"8C",X"CC",X"8C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"40",X"00",X"00",X"00",X"04",X"8E",X"FF",X"FF",X"78",X"3C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",
		X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"F8",X"0F",X"01",X"7F",X"FF",X"FF",X"E1",X"0C",X"0C",X"0C",X"8C",X"84",X"FC",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"0F",X"01",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"8C",
		X"00",X"00",X"00",X"C0",X"FF",X"FF",X"FF",X"03",X"84",X"FC",X"FC",X"FC",X"BC",X"8C",X"CC",X"8C",
		X"00",X"00",X"80",X"E0",X"30",X"18",X"0C",X"04",X"70",X"38",X"38",X"38",X"18",X"1C",X"1C",X"1C",
		X"C6",X"FE",X"FE",X"FF",X"03",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"8C",X"0C",X"0C",X"0C",
		X"0F",X"01",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"0C",X"8C",X"84",X"FC",X"00",X"00",X"00",X"00",
		X"3F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"70",
		X"00",X"00",X"C0",X"FF",X"FF",X"FF",X"03",X"00",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"CC",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"7F",X"03",X"00",X"00",X"E0",X"38",X"0C",X"06",X"FC",X"FC",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"02",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"8C",X"8C",X"8C",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0C",X"8C",X"84",X"FC",X"00",X"00",X"00",X"FC",
		X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"18",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"30",X"FC",X"FC",X"BC",X"8C",X"CC",X"8C",X"0C",
		X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"61",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",
		X"40",X"00",X"00",X"00",X"04",X"8E",X"FF",X"FF",X"78",X"3C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",
		X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F9",X"F0",X"E9",X"EF",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"1F",
		X"00",X"1E",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FF",X"F3",X"FA",X"00",
		X"FF",X"E1",X"EA",X"FA",X"F9",X"FF",X"FF",X"FF",X"9F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"00",X"FA",X"F3",X"FF",X"07",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F9",X"F0",X"E9",X"EF",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"1F",
		X"00",X"1C",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FC",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"03",X"FF",X"F3",X"FA",X"00",
		X"FF",X"E1",X"EA",X"FA",X"F9",X"FF",X"FF",X"FF",X"9F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",X"00",X"00",
		X"F8",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"00",X"FA",X"F3",X"FF",X"07",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"9F",X"1E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
