`define BUILD_DATE "190304"
`define BUILD_TIME "221722"
