`define BUILD_DATE "190415"
`define BUILD_TIME "175456"
