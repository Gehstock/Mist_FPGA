library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"3E",X"00",X"ED",X"47",X"C3",X"24",X"92",X"77",X"23",X"10",X"FC",X"C9",X"C3",X"18",X"04",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"78",X"87",X"D7",X"5F",X"23",X"56",X"EB",X"C9",
		X"E1",X"87",X"D7",X"5F",X"23",X"56",X"EB",X"E9",X"E1",X"46",X"23",X"4E",X"23",X"E5",X"18",X"12",
		X"11",X"90",X"4C",X"06",X"10",X"C3",X"51",X"00",X"F5",X"ED",X"57",X"B7",X"20",X"27",X"F1",X"C3",
		X"4F",X"9F",X"2A",X"80",X"4C",X"70",X"2C",X"71",X"2C",X"20",X"02",X"2E",X"C0",X"22",X"80",X"4C",
		X"C9",X"1A",X"A7",X"28",X"06",X"1C",X"1C",X"1C",X"10",X"F7",X"C9",X"E1",X"06",X"03",X"7E",X"12",
		X"23",X"1C",X"10",X"FA",X"E9",X"32",X"C0",X"50",X"AF",X"32",X"00",X"50",X"F3",X"C5",X"D5",X"E5",
		X"DD",X"E5",X"FD",X"E5",X"21",X"8C",X"4E",X"11",X"50",X"50",X"01",X"10",X"00",X"ED",X"B0",X"3A",
		X"9C",X"4E",X"A7",X"3A",X"CF",X"4E",X"28",X"03",X"3A",X"9F",X"4E",X"32",X"45",X"50",X"3A",X"AC",
		X"4E",X"A7",X"3A",X"DF",X"4E",X"28",X"03",X"3A",X"AF",X"4E",X"32",X"4A",X"50",X"3A",X"BC",X"4E",
		X"A7",X"3A",X"EF",X"4E",X"28",X"03",X"3A",X"BF",X"4E",X"32",X"4F",X"50",X"21",X"02",X"4C",X"11",
		X"22",X"4C",X"01",X"0A",X"06",X"7E",X"07",X"07",X"12",X"2C",X"1C",X"ED",X"A0",X"10",X"F6",X"09",
		X"EB",X"09",X"EB",X"0E",X"0C",X"ED",X"B0",X"21",X"22",X"4C",X"11",X"F2",X"4F",X"01",X"0C",X"00",
		X"ED",X"B0",X"21",X"32",X"4C",X"11",X"62",X"50",X"01",X"0C",X"00",X"ED",X"B0",X"CD",X"37",X"01",
		X"CD",X"8E",X"01",X"CD",X"00",X"B0",X"3A",X"00",X"4E",X"A7",X"28",X"0C",X"CD",X"13",X"88",X"CD",
		X"F8",X"01",X"CD",X"3E",X"02",X"CD",X"8E",X"02",X"3A",X"00",X"4E",X"3D",X"20",X"0F",X"32",X"AC",
		X"4E",X"32",X"BC",X"4E",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"32",X"EC",X"4E",X"CD",X"A3",X"9B",
		X"CD",X"58",X"9B",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3A",X"00",X"4E",X"A7",X"28",X"07",
		X"3A",X"80",X"50",X"07",X"D2",X"00",X"00",X"3E",X"01",X"32",X"00",X"50",X"FB",X"F1",X"C9",X"06",
		X"A0",X"0A",X"60",X"0A",X"60",X"0A",X"A0",X"21",X"84",X"4C",X"34",X"23",X"35",X"23",X"11",X"2F",
		X"01",X"01",X"01",X"04",X"34",X"7E",X"E6",X"0F",X"EB",X"BE",X"20",X"13",X"0C",X"1A",X"C6",X"10",
		X"E6",X"F0",X"12",X"23",X"BE",X"20",X"08",X"0C",X"EB",X"36",X"00",X"23",X"13",X"10",X"E5",X"21",
		X"8A",X"4C",X"71",X"21",X"8B",X"4C",X"7E",X"87",X"87",X"86",X"3C",X"77",X"21",X"8C",X"4C",X"7E",
		X"87",X"86",X"87",X"87",X"86",X"3C",X"77",X"2A",X"8D",X"4C",X"54",X"5D",X"29",X"29",X"19",X"EB",
		X"29",X"29",X"29",X"29",X"29",X"29",X"19",X"23",X"22",X"8D",X"4C",X"C9",X"FF",X"FF",X"21",X"90",
		X"4C",X"3A",X"8A",X"4C",X"4F",X"06",X"10",X"7E",X"A7",X"28",X"46",X"E6",X"C0",X"07",X"07",X"B9",
		X"30",X"3F",X"35",X"7E",X"E6",X"3F",X"20",X"39",X"77",X"C5",X"E5",X"2C",X"7E",X"2C",X"46",X"21",
		X"DF",X"01",X"E5",X"E7",X"81",X"B2",X"0D",X"B2",X"27",X"B1",X"68",X"86",X"15",X"83",X"20",X"83",
		X"E7",X"01",X"BB",X"91",X"C0",X"91",X"C5",X"91",X"D2",X"01",X"DA",X"01",X"EB",X"01",X"44",X"B0",
		X"44",X"B0",X"EF",X"1C",X"14",X"AF",X"32",X"39",X"4F",X"C9",X"21",X"22",X"4E",X"34",X"C9",X"E1",
		X"C1",X"2C",X"2C",X"2C",X"10",X"B1",X"C9",X"EF",X"1C",X"86",X"C9",X"78",X"A7",X"3E",X"00",X"20",
		X"03",X"32",X"27",X"4F",X"32",X"26",X"4F",X"C9",X"3A",X"6E",X"4E",X"FE",X"99",X"17",X"32",X"06",
		X"50",X"1F",X"D0",X"3A",X"00",X"50",X"47",X"CB",X"00",X"3A",X"66",X"4E",X"17",X"E6",X"0F",X"32",
		X"66",X"4E",X"D6",X"0C",X"CC",X"70",X"02",X"CB",X"00",X"3A",X"67",X"4E",X"17",X"E6",X"0F",X"32",
		X"67",X"4E",X"D6",X"0C",X"C2",X"2B",X"02",X"21",X"69",X"4E",X"34",X"CB",X"00",X"3A",X"68",X"4E",
		X"17",X"E6",X"0F",X"32",X"68",X"4E",X"D6",X"0C",X"C0",X"21",X"69",X"4E",X"34",X"C9",X"3A",X"69",
		X"4E",X"A7",X"C8",X"47",X"3A",X"6A",X"4E",X"5F",X"FE",X"00",X"C2",X"55",X"02",X"3E",X"01",X"32",
		X"07",X"50",X"CD",X"70",X"02",X"7B",X"FE",X"08",X"C2",X"5F",X"02",X"AF",X"32",X"07",X"50",X"1C",
		X"7B",X"32",X"6A",X"4E",X"D6",X"10",X"C0",X"32",X"6A",X"4E",X"05",X"78",X"32",X"69",X"4E",X"C9",
		X"3A",X"6B",X"4E",X"21",X"6C",X"4E",X"34",X"96",X"C0",X"77",X"3A",X"6D",X"4E",X"21",X"6E",X"4E",
		X"86",X"27",X"D2",X"87",X"02",X"3E",X"99",X"77",X"3E",X"01",X"32",X"9C",X"4E",X"C9",X"21",X"DA",
		X"4D",X"34",X"DD",X"21",X"D8",X"43",X"FD",X"21",X"C5",X"43",X"3A",X"00",X"4E",X"FE",X"03",X"CA",
		X"B1",X"02",X"3A",X"03",X"4E",X"FE",X"02",X"D2",X"B1",X"02",X"CD",X"D6",X"02",X"CD",X"E3",X"02",
		X"C9",X"3A",X"09",X"4E",X"A7",X"3A",X"DA",X"4D",X"C2",X"C6",X"02",X"CB",X"67",X"CC",X"D6",X"02",
		X"C4",X"F0",X"02",X"C3",X"CE",X"02",X"CB",X"67",X"CC",X"E3",X"02",X"C4",X"FD",X"02",X"3A",X"70",
		X"4E",X"A7",X"CC",X"FD",X"02",X"C9",X"DD",X"36",X"00",X"50",X"DD",X"36",X"01",X"55",X"DD",X"36",
		X"02",X"31",X"C9",X"FD",X"36",X"00",X"50",X"FD",X"36",X"01",X"55",X"FD",X"36",X"02",X"32",X"C9",
		X"DD",X"36",X"00",X"40",X"DD",X"36",X"01",X"40",X"DD",X"36",X"02",X"40",X"C9",X"FD",X"36",X"00",
		X"40",X"FD",X"36",X"01",X"40",X"FD",X"36",X"02",X"40",X"C9",X"00",X"FF",X"01",X"00",X"00",X"01",
		X"FF",X"00",X"78",X"A7",X"20",X"04",X"2A",X"0A",X"4E",X"7E",X"DD",X"21",X"9A",X"03",X"47",X"87",
		X"87",X"80",X"80",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"7E",X"00",X"87",X"47",X"87",X"87",X"4F",
		X"87",X"87",X"81",X"80",X"5F",X"16",X"00",X"21",X"8F",X"04",X"19",X"CD",X"18",X"04",X"DD",X"7E",
		X"01",X"32",X"BC",X"4D",X"DD",X"7E",X"02",X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"5F",X"04",
		X"19",X"CD",X"50",X"04",X"DD",X"7E",X"03",X"87",X"5F",X"16",X"00",X"FD",X"21",X"7D",X"04",X"FD",
		X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"C7",X"4D",X"DD",X"7E",X"04",X"87",X"5F",X"16",
		X"00",X"FD",X"21",X"6B",X"04",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"C9",X"4D",
		X"DD",X"7E",X"05",X"87",X"5F",X"16",X"00",X"FD",X"21",X"59",X"04",X"FD",X"19",X"FD",X"6E",X"00",
		X"FD",X"66",X"01",X"CD",X"CB",X"0B",X"CD",X"98",X"9A",X"C9",X"03",X"01",X"01",X"00",X"02",X"00",
		X"04",X"01",X"02",X"01",X"03",X"00",X"04",X"01",X"03",X"02",X"04",X"01",X"04",X"02",X"03",X"02",
		X"05",X"01",X"05",X"00",X"03",X"02",X"06",X"02",X"05",X"01",X"03",X"03",X"06",X"02",X"05",X"02",
		X"03",X"03",X"06",X"02",X"05",X"02",X"03",X"03",X"06",X"02",X"05",X"00",X"03",X"04",X"06",X"02",
		X"05",X"01",X"03",X"04",X"07",X"02",X"05",X"02",X"03",X"04",X"07",X"02",X"05",X"02",X"03",X"05",
		X"07",X"02",X"05",X"00",X"03",X"05",X"07",X"02",X"05",X"02",X"03",X"05",X"07",X"02",X"05",X"01",
		X"03",X"06",X"07",X"02",X"05",X"02",X"03",X"06",X"07",X"02",X"05",X"02",X"03",X"06",X"08",X"02",
		X"05",X"02",X"03",X"06",X"08",X"02",X"05",X"02",X"03",X"07",X"08",X"02",X"05",X"02",X"03",X"07",
		X"08",X"02",X"06",X"02",X"03",X"07",X"08",X"02",X"11",X"52",X"4D",X"01",X"08",X"00",X"ED",X"B0",
		X"E5",X"11",X"00",X"4F",X"01",X"0C",X"00",X"ED",X"B0",X"E1",X"11",X"5A",X"4D",X"01",X"14",X"00",
		X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",X"42",X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",X"42",
		X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",X"42",X"ED",X"B0",X"01",X"0E",X"00",X"ED",X"B0",X"C9",
		X"11",X"C4",X"4D",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"F0",X"00",X"F0",X"00",X"B4",X"00",X"14",
		X"1E",X"46",X"00",X"1E",X"3C",X"00",X"00",X"32",X"00",X"00",X"00",X"40",X"00",X"38",X"00",X"30",
		X"00",X"28",X"00",X"20",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"14",X"0A",X"1E",
		X"0F",X"28",X"14",X"32",X"19",X"3C",X"1E",X"50",X"28",X"64",X"32",X"78",X"3C",X"8C",X"46",X"55",
		X"2A",X"55",X"2A",X"55",X"55",X"55",X"55",X"55",X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"25",
		X"25",X"25",X"25",X"22",X"22",X"22",X"22",X"01",X"01",X"01",X"01",X"58",X"02",X"08",X"07",X"60",
		X"09",X"10",X"0E",X"68",X"10",X"70",X"17",X"14",X"19",X"52",X"4A",X"A5",X"94",X"AA",X"2A",X"55",
		X"55",X"55",X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"92",X"24",X"25",X"49",X"48",X"24",X"22",
		X"91",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"2A",X"55",X"2A",X"55",X"55",X"55",X"55",X"AA",X"2A",X"55",X"55",X"55",
		X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"48",X"24",X"22",X"91",X"21",X"44",X"44",X"08",X"58",
		X"02",X"34",X"08",X"D8",X"09",X"B4",X"0F",X"58",X"11",X"08",X"16",X"34",X"17",X"55",X"55",X"55",
		X"55",X"D5",X"6A",X"D5",X"6A",X"AA",X"6A",X"55",X"D5",X"55",X"55",X"55",X"55",X"AA",X"2A",X"55",
		X"55",X"92",X"24",X"92",X"24",X"22",X"22",X"22",X"22",X"A4",X"01",X"54",X"06",X"F8",X"07",X"A8",
		X"0C",X"D4",X"0D",X"84",X"12",X"B0",X"13",X"D5",X"6A",X"D5",X"6A",X"D6",X"5A",X"AD",X"B5",X"D6",
		X"5A",X"AD",X"B5",X"D5",X"6A",X"D5",X"6A",X"AA",X"6A",X"55",X"D5",X"92",X"24",X"25",X"49",X"48",
		X"24",X"22",X"91",X"A4",X"01",X"54",X"06",X"F8",X"07",X"A8",X"0C",X"D4",X"0D",X"FE",X"FF",X"FF",
		X"FF",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"B6",X"6D",X"6D",X"DB",X"6D",X"6D",X"6D",
		X"6D",X"D6",X"5A",X"AD",X"B5",X"25",X"25",X"25",X"25",X"92",X"24",X"92",X"24",X"2C",X"01",X"DC",
		X"05",X"08",X"07",X"B8",X"0B",X"E4",X"0C",X"FE",X"FF",X"FF",X"FF",X"D5",X"6A",X"D5",X"6A",X"D5",
		X"6A",X"D5",X"6A",X"B6",X"6D",X"6D",X"DB",X"6D",X"6D",X"6D",X"6D",X"D6",X"5A",X"AD",X"B5",X"48",
		X"24",X"22",X"91",X"92",X"24",X"92",X"24",X"2C",X"01",X"DC",X"05",X"08",X"07",X"B8",X"0B",X"E4",
		X"0C",X"FE",X"FF",X"FF",X"FF",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",
		X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"CD",X"8B",X"85",
		X"C8",X"2A",X"B0",X"4D",X"7C",X"B5",X"C0",X"21",X"CC",X"4E",X"CB",X"C6",X"C9",X"06",X"1E",X"DD",
		X"21",X"0A",X"4E",X"FD",X"21",X"38",X"4E",X"DD",X"56",X"00",X"FD",X"5E",X"00",X"FD",X"72",X"00",
		X"DD",X"73",X"00",X"DD",X"23",X"FD",X"23",X"10",X"EE",X"C9",X"CD",X"34",X"0B",X"C0",X"21",X"0B",
		X"4C",X"3A",X"B1",X"4D",X"A7",X"20",X"06",X"3A",X"33",X"4E",X"A7",X"20",X"06",X"3E",X"1C",X"BE",
		X"C8",X"77",X"C9",X"CD",X"46",X"0B",X"3A",X"BC",X"4E",X"A7",X"20",X"05",X"3E",X"02",X"32",X"EC",
		X"4E",X"3A",X"CC",X"4D",X"0F",X"7E",X"30",X"06",X"FE",X"0C",X"C8",X"36",X"0C",X"C9",X"FE",X"1C",
		X"C8",X"36",X"1C",X"C9",X"C8",X"36",X"0C",X"C9",X"FE",X"1C",X"C8",X"36",X"1C",X"C9",X"AF",X"32",
		X"33",X"4E",X"18",X"CD",X"21",X"D0",X"4D",X"34",X"3E",X"08",X"BE",X"C0",X"36",X"00",X"3A",X"CC",
		X"4D",X"EE",X"01",X"32",X"CC",X"4D",X"21",X"33",X"4F",X"06",X"06",X"34",X"23",X"10",X"FC",X"C9",
		X"3A",X"B2",X"4D",X"A7",X"C0",X"3A",X"CD",X"4D",X"FE",X"07",X"C8",X"87",X"2A",X"CE",X"4D",X"23",
		X"22",X"CE",X"4D",X"5F",X"16",X"00",X"DD",X"21",X"92",X"4D",X"DD",X"19",X"DD",X"5E",X"00",X"DD",
		X"56",X"01",X"A7",X"ED",X"52",X"C0",X"CB",X"3F",X"3C",X"32",X"CD",X"4D",X"21",X"01",X"01",X"22",
		X"BD",X"4D",X"22",X"BF",X"4D",X"C9",X"2A",X"B0",X"4D",X"7C",X"B5",X"C0",X"21",X"28",X"4E",X"7E",
		X"3C",X"77",X"D6",X"28",X"D8",X"E7",X"44",X"B0",X"44",X"B0",X"9A",X"07",X"49",X"07",X"B0",X"06",
		X"21",X"28",X"4E",X"36",X"00",X"23",X"3E",X"99",X"86",X"27",X"77",X"38",X"33",X"23",X"3E",X"99",
		X"86",X"27",X"77",X"38",X"0B",X"21",X"00",X"00",X"22",X"29",X"4E",X"3E",X"0D",X"32",X"B1",X"4D",
		X"21",X"2C",X"4E",X"AF",X"77",X"3A",X"29",X"4E",X"ED",X"67",X"23",X"77",X"3A",X"2A",X"4E",X"ED",
		X"67",X"CD",X"FF",X"90",X"11",X"2D",X"4E",X"21",X"61",X"43",X"01",X"03",X"02",X"C3",X"CD",X"90",
		X"A7",X"20",X"DD",X"23",X"86",X"20",X"D9",X"18",X"D2",X"74",X"E1",X"73",X"75",X"72",X"E0",X"67",
		X"6A",X"65",X"10",X"64",X"66",X"67",X"6A",X"68",X"10",X"64",X"66",X"6C",X"77",X"69",X"11",X"6B",
		X"6E",X"6C",X"77",X"6D",X"12",X"6B",X"6E",X"78",X"71",X"76",X"13",X"6F",X"70",X"78",X"71",X"79",
		X"13",X"6F",X"70",X"63",X"40",X"46",X"43",X"6D",X"40",X"52",X"43",X"7B",X"40",X"69",X"40",X"4D",
		X"43",X"72",X"40",X"5B",X"43",X"E3",X"42",X"0F",X"01",X"07",X"08",X"02",X"0F",X"03",X"05",X"04",
		X"06",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"21",X"2A",X"4E",X"3E",X"0F",X"A6",X"28",
		X"08",X"47",X"3E",X"00",X"0E",X"0A",X"81",X"10",X"FD",X"47",X"2B",X"7E",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"80",X"E7",X"44",X"B0",X"44",X"B0",X"8D",X"08",X"44",X"B0",X"44",X"B0",X"89",X"08",
		X"44",X"B0",X"44",X"B0",X"85",X"08",X"44",X"B0",X"44",X"B0",X"00",X"02",X"10",X"00",X"00",X"21",
		X"00",X"00",X"32",X"10",X"00",X"43",X"01",X"00",X"14",X"00",X"00",X"31",X"00",X"00",X"23",X"00",
		X"40",X"02",X"10",X"04",X"40",X"01",X"30",X"04",X"20",X"03",X"21",X"2B",X"4E",X"34",X"3E",X"1F",
		X"A6",X"21",X"7A",X"07",X"D7",X"A7",X"C8",X"F5",X"E6",X"0F",X"CD",X"3A",X"08",X"F1",X"0F",X"0F",
		X"0F",X"0F",X"E6",X"0F",X"C3",X"D1",X"07",X"40",X"C4",X"C5",X"40",X"C2",X"C0",X"40",X"C4",X"C5",
		X"40",X"C2",X"C0",X"40",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"40",X"C2",X"C0",X"40",X"C4",X"C5",
		X"40",X"E7",X"44",X"B0",X"DE",X"07",X"E7",X"07",X"06",X"08",X"0F",X"08",X"2E",X"08",X"21",X"C4",
		X"40",X"11",X"C5",X"07",X"C3",X"56",X"09",X"21",X"C7",X"42",X"11",X"B8",X"07",X"CD",X"56",X"09",
		X"3A",X"1E",X"4E",X"A7",X"C8",X"3A",X"0A",X"47",X"32",X"20",X"4E",X"3E",X"1A",X"32",X"0A",X"43",
		X"3E",X"0C",X"32",X"0A",X"47",X"C9",X"21",X"CE",X"40",X"11",X"C5",X"07",X"C3",X"56",X"09",X"21",
		X"D3",X"42",X"11",X"C5",X"07",X"CD",X"56",X"09",X"3A",X"1F",X"4E",X"A7",X"C8",X"3A",X"16",X"47",
		X"32",X"21",X"4E",X"3E",X"1A",X"32",X"16",X"43",X"3E",X"0C",X"32",X"16",X"47",X"C9",X"CD",X"DE",
		X"07",X"CD",X"E7",X"07",X"CD",X"06",X"08",X"C3",X"0F",X"08",X"E7",X"44",X"B0",X"47",X"08",X"50",
		X"08",X"60",X"08",X"69",X"08",X"79",X"08",X"21",X"C4",X"40",X"11",X"C4",X"07",X"C3",X"56",X"09",
		X"21",X"C7",X"42",X"11",X"B7",X"07",X"CD",X"56",X"09",X"3A",X"20",X"4E",X"C3",X"B0",X"0A",X"C9",
		X"21",X"CE",X"40",X"11",X"C4",X"07",X"C3",X"56",X"09",X"21",X"D3",X"42",X"11",X"C4",X"07",X"CD",
		X"56",X"09",X"3A",X"21",X"4E",X"C3",X"B9",X"0A",X"C9",X"CD",X"47",X"08",X"CD",X"50",X"08",X"CD",
		X"60",X"08",X"C3",X"69",X"08",X"0E",X"01",X"18",X"0A",X"0E",X"02",X"18",X"06",X"0E",X"03",X"18",
		X"02",X"0E",X"04",X"3A",X"29",X"4E",X"E6",X"0F",X"21",X"37",X"07",X"D7",X"FE",X"0F",X"C8",X"3D",
		X"47",X"21",X"16",X"4E",X"D7",X"B9",X"C0",X"3C",X"77",X"87",X"86",X"87",X"4F",X"7E",X"FE",X"05",
		X"30",X"13",X"FE",X"01",X"20",X"07",X"3E",X"01",X"32",X"AC",X"4E",X"18",X"08",X"21",X"41",X"07",
		X"78",X"D7",X"32",X"BC",X"4E",X"21",X"F9",X"06",X"7D",X"81",X"6F",X"3E",X"00",X"8C",X"67",X"E5",
		X"21",X"23",X"07",X"3E",X"07",X"B8",X"20",X"05",X"3A",X"0D",X"4E",X"80",X"47",X"DF",X"D1",X"CD",
		X"3D",X"09",X"C9",X"78",X"21",X"16",X"4E",X"D7",X"36",X"00",X"21",X"F9",X"06",X"18",X"E0",X"78",
		X"21",X"16",X"4E",X"D7",X"18",X"B1",X"78",X"21",X"16",X"4E",X"D7",X"18",X"AC",X"78",X"21",X"16",
		X"4E",X"D7",X"A7",X"C8",X"18",X"A1",X"06",X"08",X"C5",X"05",X"CD",X"FD",X"08",X"C1",X"10",X"F8",
		X"C9",X"06",X"08",X"C5",X"05",X"CD",X"EF",X"08",X"C1",X"10",X"F8",X"C9",X"06",X"08",X"C5",X"05",
		X"CD",X"F6",X"08",X"C1",X"10",X"F8",X"C9",X"06",X"08",X"C5",X"05",X"CD",X"E3",X"08",X"C1",X"10",
		X"F8",X"3A",X"0D",X"4E",X"EE",X"01",X"C6",X"07",X"47",X"CD",X"E3",X"08",X"C9",X"06",X"03",X"D5",
		X"DD",X"E1",X"11",X"1F",X"00",X"DD",X"7E",X"00",X"77",X"23",X"DD",X"23",X"DD",X"7E",X"00",X"77",
		X"DD",X"23",X"19",X"10",X"F0",X"C9",X"06",X"04",X"C5",X"1A",X"77",X"23",X"13",X"1A",X"77",X"23",
		X"13",X"1A",X"77",X"13",X"01",X"1E",X"00",X"09",X"C1",X"10",X"ED",X"C9",X"03",X"02",X"9C",X"43",
		X"E0",X"D1",X"C3",X"D0",X"D0",X"D0",X"03",X"02",X"53",X"40",X"D0",X"D0",X"D0",X"6A",X"D6",X"C7",
		X"03",X"02",X"9C",X"43",X"66",X"D1",X"C3",X"D0",X"D0",X"D0",X"03",X"02",X"53",X"40",X"D0",X"D0",
		X"D0",X"E1",X"D6",X"C7",X"03",X"06",X"3C",X"41",X"CE",X"D8",X"C3",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"CF",X"D7",X"C7",X"03",X"03",X"96",X"41",X"40",X"D9",
		X"DA",X"D0",X"D0",X"D0",X"CF",X"F9",X"DE",X"03",X"04",X"19",X"42",X"CE",X"F8",X"DA",X"D0",X"D0",
		X"D0",X"D0",X"D0",X"D0",X"40",X"DB",X"DE",X"03",X"03",X"0E",X"42",X"CE",X"F8",X"DA",X"D0",X"D0",
		X"D0",X"CF",X"D7",X"C7",X"03",X"03",X"8A",X"41",X"40",X"D9",X"DA",X"D0",X"D0",X"D0",X"63",X"F9",
		X"DE",X"03",X"04",X"07",X"42",X"CE",X"F8",X"DA",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"CF",X"D7",
		X"C7",X"03",X"03",X"84",X"41",X"40",X"D9",X"DA",X"D0",X"D0",X"D0",X"40",X"DB",X"DE",X"02",X"01",
		X"FA",X"41",X"1C",X"1D",X"02",X"01",X"77",X"41",X"1C",X"1D",X"04",X"01",X"F2",X"41",X"1C",X"1D",
		X"1D",X"1D",X"03",X"01",X"EB",X"41",X"1C",X"1D",X"1D",X"03",X"01",X"EB",X"42",X"1C",X"1D",X"1D",
		X"02",X"01",X"E5",X"41",X"1C",X"1D",X"E4",X"78",X"94",X"09",X"1C",X"80",X"B4",X"80",X"AA",X"09",
		X"1C",X"80",X"CC",X"80",X"B7",X"09",X"1C",X"00",X"74",X"78",X"C7",X"09",X"1C",X"00",X"54",X"58",
		X"D4",X"09",X"1C",X"00",X"3C",X"80",X"E1",X"09",X"1C",X"00",X"24",X"58",X"F1",X"09",X"1C",X"00",
		X"20",X"20",X"1C",X"00",X"38",X"E0",X"1C",X"80",X"70",X"20",X"1C",X"00",X"98",X"E0",X"1C",X"80",
		X"E0",X"20",X"1C",X"00",X"50",X"20",X"1C",X"00",X"70",X"E0",X"1C",X"80",X"98",X"20",X"1C",X"00",
		X"24",X"02",X"02",X"02",X"02",X"10",X"FF",X"FF",X"28",X"16",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"01",X"BC",X"38",X"1A",X"20",X"0C",X"3E",X"00",X"BD",X"20",X"13",X"21",X"00",X"15",X"22",
		X"30",X"4E",X"C9",X"3E",X"50",X"BD",X"38",X"F4",X"21",X"00",X"20",X"22",X"30",X"4E",X"C9",X"22",
		X"30",X"4E",X"C9",X"30",X"4E",X"AF",X"96",X"27",X"77",X"23",X"3E",X"10",X"9E",X"27",X"77",X"C9",
		X"32",X"0A",X"47",X"3E",X"40",X"32",X"0A",X"43",X"C9",X"32",X"16",X"47",X"3E",X"40",X"32",X"16",
		X"43",X"C9",X"21",X"22",X"0F",X"DD",X"21",X"2A",X"0F",X"18",X"07",X"21",X"8C",X"0F",X"DD",X"21",
		X"94",X"0F",X"06",X"00",X"DD",X"09",X"79",X"3D",X"0F",X"E6",X"06",X"4F",X"09",X"5E",X"23",X"56",
		X"DD",X"7E",X"00",X"12",X"C9",X"21",X"00",X"0F",X"18",X"03",X"21",X"6A",X"0F",X"06",X"00",X"5E",
		X"23",X"56",X"D5",X"DD",X"E1",X"79",X"0F",X"30",X"05",X"11",X"00",X"04",X"DD",X"19",X"23",X"79",
		X"87",X"87",X"4F",X"09",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"20",X"23",X"7E",X"DD",
		X"77",X"40",X"23",X"7E",X"DD",X"77",X"60",X"C9",X"22",X"D7",X"4D",X"0E",X"04",X"CD",X"EA",X"0A",
		X"0E",X"05",X"CD",X"EA",X"0A",X"C9",X"22",X"D7",X"4D",X"0E",X"02",X"CD",X"EA",X"0A",X"0E",X"03",
		X"CD",X"EA",X"0A",X"C9",X"CD",X"82",X"85",X"47",X"3A",X"1A",X"4F",X"D6",X"09",X"0E",X"00",X"38",
		X"02",X"0E",X"0F",X"78",X"B1",X"C9",X"E5",X"2A",X"D7",X"4D",X"2D",X"20",X"10",X"3A",X"C9",X"4D",
		X"6F",X"24",X"3E",X"0F",X"A4",X"28",X"0B",X"E5",X"4F",X"CD",X"CB",X"0A",X"E1",X"22",X"D7",X"4D",
		X"E1",X"C9",X"CD",X"6E",X"0B",X"AF",X"32",X"33",X"4E",X"E1",X"36",X"1C",X"E1",X"C9",X"3A",X"1E",
		X"4E",X"4F",X"3A",X"1F",X"4E",X"B1",X"21",X"01",X"0F",X"28",X"0E",X"22",X"D7",X"4D",X"0E",X"00",
		X"CD",X"EA",X"0A",X"0E",X"01",X"CD",X"EA",X"0A",X"C9",X"CD",X"18",X"0B",X"C9",X"3A",X"3F",X"4F",
		X"B7",X"20",X"04",X"3A",X"40",X"50",X"C9",X"2A",X"3D",X"4F",X"2D",X"20",X"13",X"3A",X"3B",X"4F",
		X"6F",X"24",X"3E",X"0F",X"A4",X"28",X"0E",X"22",X"3D",X"4F",X"4F",X"CD",X"C2",X"0A",X"E1",X"C9",
		X"22",X"3D",X"4F",X"E1",X"C9",X"21",X"01",X"0F",X"22",X"3D",X"4F",X"0E",X"02",X"CD",X"E5",X"0A",
		X"0E",X"03",X"CD",X"E5",X"0A",X"AF",X"32",X"3F",X"4F",X"E1",X"C9",X"22",X"A1",X"4D",X"3A",X"13",
		X"4E",X"87",X"4F",X"06",X"00",X"21",X"3A",X"0F",X"09",X"5E",X"23",X"56",X"EB",X"22",X"3B",X"4F",
		X"AF",X"32",X"3F",X"4F",X"C9",X"CD",X"40",X"93",X"0E",X"00",X"CD",X"E5",X"0A",X"0E",X"00",X"CD",
		X"EA",X"0A",X"C9",X"CD",X"0F",X"91",X"0E",X"01",X"CD",X"E5",X"0A",X"0E",X"01",X"CD",X"EA",X"0A",
		X"C9",X"47",X"2F",X"E6",X"0F",X"CA",X"B0",X"8B",X"2A",X"41",X"4F",X"7D",X"B4",X"28",X"19",X"3A",
		X"09",X"4D",X"FE",X"58",X"38",X"0C",X"FE",X"68",X"38",X"17",X"FE",X"90",X"38",X"04",X"FE",X"A0",
		X"38",X"0F",X"21",X"00",X"00",X"22",X"41",X"4F",X"78",X"CB",X"4F",X"CA",X"FF",X"8C",X"C3",X"A1",
		X"8B",X"78",X"2A",X"41",X"4F",X"E9",X"0F",X"D2",X"0D",X"8D",X"0F",X"D2",X"0D",X"8D",X"0F",X"D2",
		X"06",X"8D",X"C3",X"06",X"8D",X"0F",X"D2",X"FF",X"8C",X"0F",X"D2",X"FF",X"8C",X"0F",X"D2",X"14",
		X"8D",X"C3",X"14",X"8D",X"0F",X"D2",X"0D",X"8D",X"0F",X"D2",X"FF",X"8C",X"0F",X"D2",X"0D",X"8D",
		X"C3",X"FF",X"8C",X"0F",X"D2",X"06",X"8D",X"0F",X"D2",X"14",X"8D",X"0F",X"D2",X"06",X"8D",X"C3",
		X"14",X"8D",X"E6",X"07",X"FE",X"04",X"C0",X"D1",X"ED",X"5B",X"08",X"4D",X"21",X"CC",X"0F",X"06",
		X"08",X"7B",X"BE",X"23",X"20",X"18",X"7A",X"BE",X"20",X"14",X"21",X"DC",X"0F",X"3E",X"08",X"90",
		X"E6",X"06",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"ED",X"53",X"41",X"4F",X"C9",X"23",X"10",
		X"E0",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D1",X"42",X"FC",X"05",X"05",X"EC",X"1D",X"1D",X"1D",X"1D",X"FC",X"05",X"05",X"EC",X"1D",X"1D",
		X"1D",X"1D",X"FC",X"05",X"05",X"EC",X"1B",X"1B",X"1B",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"31",X"43",X"11",X"43",X"F1",X"42",X"D1",X"42",X"EC",X"ED",X"EE",X"EF",X"FA",X"08",
		X"07",X"06",X"01",X"08",X"07",X"06",X"01",X"FF",X"FE",X"FD",X"12",X"00",X"16",X"00",X"1A",X"00",
		X"1E",X"00",X"25",X"00",X"2D",X"00",X"34",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",
		X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",
		X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"D1",X"40",X"FB",X"01",X"01",X"FA",
		X"1D",X"1D",X"1D",X"1D",X"FC",X"05",X"05",X"EC",X"1D",X"1D",X"1D",X"1D",X"FC",X"05",X"05",X"EC",
		X"1B",X"1B",X"1B",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"31",X"41",X"11",X"41",
		X"F1",X"40",X"D1",X"40",X"EC",X"ED",X"EE",X"EF",X"FA",X"08",X"07",X"06",X"01",X"08",X"07",X"06",
		X"01",X"FF",X"FE",X"FD",X"08",X"1A",X"0C",X"00",X"09",X"1D",X"0D",X"00",X"0A",X"1F",X"0E",X"00",
		X"0B",X"1B",X"0F",X"00",X"0C",X"1E",X"08",X"00",X"0D",X"13",X"09",X"00",X"0E",X"1B",X"0A",X"00",
		X"0F",X"0C",X"0B",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"9C",X"5C",X"94",X"64",
		X"94",X"5C",X"8C",X"64",X"9C",X"9C",X"94",X"94",X"94",X"9C",X"8C",X"94",X"36",X"0C",X"45",X"0C",
		X"54",X"0C",X"63",X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr(11 downto 0))));
	end if;
end process;
end architecture;
