library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity char_rom2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of char_rom2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"DE",X"9E",X"2F",X"4B",X"4B",X"9F",X"5F",X"0F",X"E0",X"F0",X"A4",X"5A",X"3C",X"9E",X"0F",X"2F",
		X"1E",X"3C",X"68",X"5A",X"69",X"2D",X"3C",X"3C",X"E0",X"C1",X"D0",X"50",X"E0",X"A4",X"E0",X"30",
		X"0F",X"0F",X"1E",X"2D",X"0F",X"5B",X"0F",X"0F",X"4B",X"3F",X"0F",X"0F",X"87",X"1E",X"3C",X"94",
		X"0F",X"3F",X"0F",X"0F",X"0F",X"3F",X"2F",X"0F",X"87",X"96",X"AF",X"2F",X"87",X"0F",X"0F",X"4B",
		X"0F",X"38",X"33",X"33",X"2A",X"19",X"0C",X"0F",X"E1",X"ED",X"FE",X"76",X"ED",X"21",X"03",X"0F",
		X"4F",X"4F",X"0F",X"0F",X"6F",X"2F",X"8F",X"0F",X"B4",X"5A",X"B4",X"3C",X"1E",X"8F",X"4F",X"0F",
		X"2D",X"1E",X"3C",X"2D",X"1E",X"2D",X"1E",X"0F",X"B0",X"78",X"78",X"F0",X"E1",X"E1",X"F0",X"B4",
		X"0F",X"1E",X"3C",X"2D",X"78",X"5A",X"3C",X"78",X"C3",X"5A",X"F0",X"E1",X"B0",X"D2",X"B4",X"70",
		X"1E",X"0F",X"2D",X"0F",X"0F",X"1F",X"4B",X"0F",X"1E",X"2F",X"0F",X"0F",X"4B",X"0F",X"87",X"3C",
		X"0F",X"CF",X"5F",X"4F",X"0F",X"3F",X"2F",X"0F",X"0F",X"87",X"4B",X"8F",X"87",X"1F",X"0F",X"0F",
		X"3E",X"33",X"33",X"7F",X"2A",X"08",X"09",X"0F",X"78",X"D4",X"FE",X"BB",X"FE",X"30",X"21",X"0F",
		X"C7",X"73",X"31",X"10",X"10",X"00",X"00",X"70",X"0F",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"F0",
		X"2D",X"5E",X"6F",X"2F",X"2D",X"4F",X"1F",X"3F",X"6F",X"9F",X"6B",X"9E",X"4F",X"B4",X"69",X"4B",
		X"8F",X"69",X"0F",X"6F",X"0F",X"BF",X"2F",X"0F",X"6F",X"3F",X"4F",X"2F",X"87",X"4B",X"9E",X"2D",
		X"3C",X"2F",X"6F",X"1E",X"AD",X"4F",X"1F",X"7F",X"6F",X"4F",X"0F",X"4F",X"DB",X"0F",X"5A",X"69",
		X"2D",X"4F",X"5E",X"96",X"1F",X"4F",X"97",X"2F",X"8F",X"CF",X"2F",X"C7",X"0F",X"4F",X"1E",X"2D",
		X"40",X"E0",X"B0",X"58",X"B4",X"F0",X"3C",X"0F",X"58",X"A0",X"D0",X"78",X"F0",X"F0",X"C3",X"0F",
		X"AF",X"FF",X"BB",X"99",X"CC",X"6E",X"B7",X"D3",X"9E",X"EF",X"BF",X"CF",X"EF",X"77",X"55",X"3B",
		X"97",X"2D",X"1E",X"69",X"C3",X"97",X"6F",X"BF",X"FF",X"7F",X"F0",X"3C",X"EF",X"0F",X"2F",X"6D",
		X"0F",X"1E",X"6F",X"4F",X"1F",X"0C",X"7F",X"3F",X"ED",X"0F",X"2E",X"CC",X"00",X"FF",X"DF",X"66",
		X"1E",X"0F",X"4B",X"8F",X"2F",X"2D",X"4F",X"0F",X"69",X"B4",X"69",X"96",X"0F",X"4F",X"8F",X"0F",
		X"F0",X"B0",X"F0",X"F0",X"B4",X"B4",X"5A",X"3C",X"F0",X"F0",X"78",X"F0",X"E0",X"F0",X"B4",X"F0",
		X"E0",X"E0",X"F0",X"B0",X"B0",X"F0",X"F0",X"F0",X"B7",X"37",X"53",X"13",X"A1",X"90",X"C0",X"E0",
		X"58",X"D0",X"D0",X"D0",X"E0",X"E1",X"C0",X"E0",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"B7",
		X"0F",X"4B",X"1E",X"9E",X"3D",X"2D",X"2C",X"48",X"2D",X"4B",X"43",X"47",X"1F",X"C7",X"6F",X"5F",
		X"0F",X"0F",X"0F",X"87",X"4B",X"0F",X"8F",X"0F",X"0F",X"3C",X"0F",X"6F",X"2F",X"0F",X"1E",X"3C",
		X"4F",X"4F",X"1E",X"2D",X"AF",X"4F",X"0F",X"0F",X"0F",X"3C",X"4F",X"6F",X"0F",X"0F",X"4B",X"8F",
		X"0F",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"F0",X"0F",X"CF",X"8F",X"8F",X"8F",X"C7",X"63",X"F1",
		X"2D",X"4F",X"1F",X"4B",X"1E",X"6F",X"3F",X"8F",X"4B",X"3C",X"CF",X"2F",X"87",X"D3",X"0F",X"4F",
		X"2F",X"69",X"1F",X"4F",X"1E",X"69",X"97",X"87",X"A7",X"0F",X"DA",X"AD",X"4F",X"5F",X"0F",X"2F",
		X"0F",X"2F",X"BF",X"2D",X"5B",X"4F",X"1F",X"A5",X"C3",X"D7",X"0F",X"2F",X"5E",X"2D",X"9E",X"CF",
		X"0F",X"2F",X"5B",X"0F",X"6D",X"C7",X"1F",X"0F",X"5E",X"0F",X"3F",X"4B",X"AF",X"B4",X"2F",X"8F",
		X"C3",X"0F",X"0B",X"96",X"2F",X"0F",X"4B",X"0F",X"6F",X"1E",X"2F",X"0F",X"2D",X"87",X"0F",X"0F",
		X"0F",X"1F",X"1F",X"0F",X"4F",X"BE",X"FC",X"F7",X"EA",X"7B",X"7B",X"E2",X"C7",X"C7",X"AD",X"0F",
		X"00",X"08",X"86",X"69",X"F4",X"5A",X"3D",X"0F",X"00",X"00",X"00",X"00",X"08",X"80",X"84",X"C0",
		X"0F",X"DD",X"00",X"00",X"00",X"CC",X"AA",X"00",X"0F",X"AB",X"11",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"78",X"B4",X"69",X"1E",X"0F",X"0F",X"0F",X"F0",X"78",X"E1",X"B4",X"E1",X"0F",X"0F",X"0F",
		X"21",X"90",X"C0",X"E0",X"F0",X"E1",X"B0",X"B0",X"FF",X"7F",X"97",X"21",X"80",X"78",X"F0",X"B0",
		X"99",X"AA",X"88",X"DD",X"CC",X"CC",X"FF",X"D5",X"FF",X"FF",X"77",X"BB",X"55",X"00",X"00",X"FF",
		X"33",X"33",X"67",X"33",X"77",X"33",X"BB",X"99",X"FF",X"FF",X"FF",X"BB",X"BF",X"77",X"FF",X"FF",
		X"4F",X"4F",X"9F",X"3F",X"5D",X"5D",X"BB",X"BB",X"7F",X"AF",X"AF",X"77",X"DF",X"BB",X"EF",X"57",
		X"0F",X"97",X"97",X"3F",X"4B",X"1E",X"69",X"87",X"0F",X"78",X"C7",X"87",X"4F",X"1F",X"4F",X"8F",
		X"CC",X"AD",X"1F",X"0F",X"1E",X"2F",X"2F",X"0F",X"17",X"B7",X"4F",X"3F",X"6E",X"5F",X"AF",X"5F",
		X"0F",X"CB",X"1F",X"4F",X"0F",X"6F",X"2F",X"0F",X"0F",X"87",X"4B",X"8F",X"0F",X"1F",X"2E",X"88",
		X"90",X"90",X"90",X"90",X"90",X"80",X"80",X"00",X"E7",X"E7",X"E7",X"E7",X"E7",X"63",X"31",X"10",
		X"0F",X"87",X"C3",X"B1",X"90",X"90",X"90",X"90",X"0F",X"0F",X"2F",X"EF",X"E7",X"E7",X"E7",X"E7",
		X"F0",X"F0",X"F0",X"E0",X"E1",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",X"00",X"00",X"78",X"3C",X"1E",
		X"2F",X"8F",X"1F",X"4E",X"2D",X"4F",X"8F",X"0E",X"5B",X"6D",X"ED",X"76",X"77",X"77",X"77",X"77",
		X"0F",X"4F",X"0F",X"1E",X"1E",X"2F",X"6F",X"0F",X"1E",X"2F",X"5E",X"2F",X"2D",X"CF",X"4F",X"0F",
		X"66",X"CE",X"7F",X"DF",X"77",X"AE",X"2F",X"07",X"03",X"03",X"47",X"07",X"16",X"2F",X"6F",X"0F",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"22",X"47",X"23",X"01",X"23",X"23",X"01",X"23",X"23",
		X"2F",X"3F",X"8F",X"47",X"11",X"00",X"00",X"00",X"1E",X"5E",X"2F",X"4F",X"0F",X"AF",X"47",X"23",
		X"F0",X"F0",X"90",X"78",X"E1",X"78",X"2D",X"0F",X"E1",X"A5",X"D2",X"70",X"A5",X"C3",X"0F",X"0F",
		X"FF",X"FF",X"EF",X"0F",X"70",X"00",X"F0",X"D2",X"FF",X"FF",X"3F",X"C3",X"30",X"CC",X"3C",X"F0",
		X"FF",X"FF",X"EE",X"FF",X"FF",X"EF",X"11",X"CC",X"FF",X"7F",X"FF",X"FF",X"EF",X"DD",X"FF",X"00",
		X"4F",X"EF",X"CF",X"AB",X"DF",X"FF",X"EF",X"FF",X"0F",X"0F",X"0F",X"8F",X"CF",X"5F",X"FF",X"BB",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"2D",X"CF",X"0F",X"0F",X"0F",X"4B",X"8F",X"0F",
		X"78",X"C3",X"0F",X"3D",X"4F",X"0F",X"3F",X"4F",X"F0",X"1E",X"2D",X"CF",X"2F",X"0F",X"1E",X"0F",
		X"FF",X"7F",X"CC",X"FF",X"EF",X"77",X"FF",X"8F",X"FF",X"9F",X"FF",X"FF",X"EF",X"BB",X"FF",X"0F",
		X"0F",X"6F",X"5E",X"0F",X"DD",X"00",X"00",X"77",X"AD",X"8F",X"0F",X"6E",X"88",X"00",X"00",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"D0",X"B0",X"F0",X"70",X"70",X"70",X"00",X"00",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"00",X"10",X"E0",X"E0",X"E8",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",
		X"FF",X"BB",X"FF",X"FF",X"EE",X"88",X"03",X"1F",X"ED",X"ED",X"ED",X"25",X"4F",X"1E",X"A7",X"0F",
		X"0F",X"3F",X"1F",X"0F",X"0F",X"7D",X"2F",X"0F",X"4A",X"A5",X"1E",X"0F",X"7E",X"1F",X"0F",X"0F",
		X"0F",X"1E",X"1E",X"0F",X"1E",X"0F",X"0F",X"0F",X"78",X"A0",X"58",X"A0",X"68",X"D2",X"B4",X"F0",
		X"8F",X"1F",X"4F",X"0F",X"0F",X"2D",X"1E",X"0F",X"0F",X"0F",X"0F",X"5A",X"E7",X"0F",X"3C",X"68",
		X"3C",X"3B",X"33",X"77",X"11",X"00",X"0C",X"0E",X"C3",X"E9",X"FC",X"76",X"FE",X"FE",X"65",X"43",
		X"87",X"2F",X"87",X"4B",X"0F",X"4B",X"87",X"0F",X"1E",X"1E",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"EF",X"CF",X"DF",X"2F",X"00",X"70",X"87",X"0F",X"8F",X"9E",X"0F",X"70",X"43",X"87",X"2F",X"2F",
		X"DF",X"FF",X"BB",X"FF",X"EF",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"CF",X"0F",X"0F",
		X"0F",X"0F",X"1E",X"AF",X"5F",X"2F",X"CF",X"FF",X"0F",X"0F",X"0F",X"87",X"0F",X"4F",X"8F",X"4F",
		X"0F",X"2D",X"4F",X"0F",X"0F",X"1E",X"3F",X"0F",X"5A",X"1E",X"5A",X"0F",X"2D",X"87",X"0F",X"0F",
		X"0F",X"F0",X"1E",X"4B",X"1E",X"0F",X"D2",X"1E",X"CC",X"3F",X"C3",X"78",X"3C",X"D2",X"B4",X"69",
		X"EE",X"55",X"EE",X"CC",X"AA",X"CC",X"DD",X"66",X"CC",X"26",X"88",X"44",X"9B",X"00",X"44",X"00",
		X"0F",X"0F",X"08",X"00",X"00",X"00",X"00",X"08",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"8E",X"2D",X"6F",X"2F",X"CB",X"5F",X"0F",X"FF",X"77",X"33",X"00",X"08",X"0C",X"4B",X"8F",
		X"87",X"1F",X"0F",X"6B",X"8F",X"5F",X"0E",X"0E",X"0F",X"3C",X"79",X"FF",X"FF",X"EE",X"DD",X"FF",
		X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",
		X"8F",X"0F",X"F0",X"F7",X"FF",X"FF",X"FF",X"FF",X"1F",X"E1",X"ED",X"FC",X"FE",X"FE",X"CF",X"CF",
		X"F0",X"48",X"D2",X"E1",X"1E",X"0F",X"4F",X"1F",X"10",X"E1",X"B0",X"D2",X"F0",X"0F",X"2F",X"0F",
		X"3B",X"3B",X"3B",X"1D",X"95",X"A6",X"C3",X"69",X"1E",X"0F",X"AF",X"8F",X"EF",X"77",X"08",X"0F",
		X"1F",X"0F",X"4B",X"1E",X"3C",X"4B",X"B7",X"6F",X"AA",X"7F",X"0F",X"F0",X"0F",X"9E",X"4F",X"3F",
		X"0F",X"4F",X"0F",X"1E",X"6F",X"4F",X"0F",X"0E",X"1E",X"7E",X"8F",X"87",X"0F",X"0F",X"CC",X"DF",
		X"2F",X"0F",X"1E",X"6F",X"2F",X"0F",X"6F",X"1F",X"87",X"0F",X"3C",X"4F",X"2F",X"4F",X"0F",X"0F",
		X"5E",X"BD",X"D2",X"C7",X"2F",X"0F",X"0F",X"0F",X"2F",X"0F",X"0F",X"87",X"2F",X"2F",X"0F",X"0F",
		X"8F",X"0F",X"1F",X"1F",X"3E",X"8F",X"0F",X"3C",X"3D",X"6D",X"79",X"1F",X"7B",X"2D",X"69",X"A7",
		X"0F",X"2D",X"1E",X"2D",X"2D",X"2D",X"1E",X"8F",X"B4",X"5A",X"1E",X"0F",X"87",X"0F",X"3C",X"2D",
		X"5A",X"87",X"A5",X"4B",X"D2",X"A5",X"4B",X"69",X"E6",X"E2",X"FD",X"7D",X"7F",X"2D",X"B4",X"5A",
		X"00",X"00",X"88",X"6E",X"B7",X"D3",X"69",X"3C",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"4C",
		X"0F",X"BF",X"0F",X"1E",X"6F",X"2F",X"0F",X"0F",X"AD",X"0F",X"0F",X"3C",X"3F",X"7F",X"77",X"33",
		X"0F",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"77",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"BB",X"FF",X"FF",X"22",X"01",X"17",X"0F",X"ED",X"CB",X"ED",X"CF",X"8F",X"3F",X"2F",X"9E",
		X"0F",X"E1",X"FC",X"FE",X"BB",X"FF",X"77",X"EE",X"BE",X"0F",X"3F",X"1F",X"D2",X"CB",X"ED",X"ED",
		X"E1",X"E1",X"E1",X"10",X"00",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",X"E1",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"A7",X"97",X"C3",X"0F",X"0F",X"0F",X"0F",X"0F",X"84",X"2F",X"4F",X"9F",X"1E",X"6F",X"7C",X"0F",
		X"9F",X"CF",X"0F",X"3F",X"FF",X"FE",X"ED",X"DA",X"EA",X"FB",X"FB",X"95",X"B7",X"2F",X"0F",X"0F",
		X"22",X"88",X"08",X"B7",X"5B",X"6D",X"1E",X"5B",X"00",X"00",X"00",X"00",X"00",X"88",X"19",X"A6",
		X"9E",X"3F",X"2F",X"0F",X"0F",X"88",X"00",X"CC",X"97",X"1E",X"6F",X"4F",X"0F",X"67",X"11",X"00",
		X"2D",X"6F",X"2F",X"1E",X"6F",X"4F",X"2F",X"0F",X"3B",X"19",X"08",X"08",X"84",X"0E",X"8F",X"2D",
		X"2D",X"4F",X"1D",X"4E",X"A6",X"0D",X"0B",X"07",X"88",X"99",X"23",X"47",X"0F",X"0F",X"0F",X"0F",
		X"EF",X"FF",X"AB",X"BB",X"7F",X"DF",X"3F",X"87",X"FF",X"FF",X"AA",X"EE",X"4C",X"AA",X"4C",X"08",
		X"7F",X"6E",X"5D",X"7F",X"7F",X"6E",X"7F",X"EF",X"55",X"BB",X"9D",X"EF",X"46",X"FF",X"55",X"FF",
		X"00",X"00",X"00",X"44",X"00",X"00",X"22",X"99",X"00",X"00",X"00",X"22",X"00",X"CC",X"55",X"BB",
		X"1D",X"19",X"3B",X"2A",X"80",X"8C",X"2D",X"4F",X"FF",X"DD",X"77",X"FF",X"11",X"1D",X"8C",X"4F",
		X"3F",X"1F",X"0F",X"C3",X"F8",X"55",X"EE",X"BB",X"4B",X"1E",X"6F",X"1F",X"87",X"C3",X"FB",X"C3",
		X"3F",X"5F",X"0F",X"47",X"11",X"00",X"00",X"00",X"0F",X"2D",X"5F",X"2F",X"0F",X"8F",X"67",X"00",
		X"0E",X"0C",X"0C",X"0C",X"0C",X"0E",X"0F",X"0F",X"77",X"77",X"77",X"33",X"22",X"00",X"00",X"0F",
		X"4F",X"A7",X"1E",X"7F",X"3E",X"DA",X"4F",X"0F",X"4F",X"78",X"FF",X"55",X"FF",X"B3",X"19",X"22",
		X"6B",X"8F",X"0F",X"0E",X"0F",X"0F",X"0F",X"8F",X"77",X"33",X"11",X"33",X"11",X"2A",X"0F",X"1F",
		X"0F",X"0F",X"8F",X"BE",X"0F",X"2D",X"4F",X"0F",X"4B",X"8F",X"1E",X"79",X"3B",X"3B",X"3B",X"33",
		X"1E",X"39",X"77",X"77",X"22",X"19",X"08",X"0E",X"87",X"C3",X"F8",X"FE",X"DC",X"BA",X"ED",X"47",
		X"88",X"88",X"00",X"88",X"99",X"01",X"23",X"47",X"27",X"9E",X"8F",X"3F",X"3D",X"4F",X"CF",X"0F",
		X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"5E",X"2F",X"8F",X"AF",X"37",X"07",X"07",
		X"1F",X"0F",X"1E",X"2F",X"6F",X"0F",X"0F",X"03",X"1E",X"3E",X"7F",X"0F",X"2D",X"AD",X"8F",X"0F",
		X"DD",X"BB",X"EE",X"33",X"00",X"00",X"0B",X"0F",X"87",X"CB",X"ED",X"FE",X"65",X"4B",X"0F",X"0F",
		X"07",X"4F",X"5F",X"0F",X"1E",X"6F",X"4F",X"0F",X"4B",X"CB",X"0F",X"8F",X"1E",X"6F",X"CF",X"0F",
		X"00",X"00",X"11",X"00",X"11",X"23",X"03",X"47",X"07",X"8F",X"2F",X"7F",X"0F",X"4B",X"AD",X"4F",
		X"44",X"88",X"88",X"88",X"44",X"88",X"88",X"00",X"23",X"23",X"23",X"23",X"47",X"47",X"47",X"47",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"01",X"11",X"11",X"11",X"11",X"01",X"23",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"23",X"23",X"23",X"23",X"23",X"11",X"11",
		X"47",X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"CF",X"2D",X"7E",X"AF",X"8F",X"57",X"47",X"23",
		X"0F",X"87",X"C2",X"D3",X"D3",X"C3",X"80",X"00",X"0F",X"1E",X"30",X"B8",X"B8",X"3C",X"10",X"00",
		X"BB",X"FF",X"FF",X"EE",X"89",X"16",X"2F",X"0F",X"ED",X"E9",X"07",X"1E",X"3F",X"6B",X"8F",X"8F",
		X"0F",X"87",X"F0",X"FE",X"BB",X"DD",X"FF",X"FF",X"CB",X"3F",X"2F",X"87",X"D3",X"CB",X"ED",X"ED",
		X"FF",X"FF",X"FF",X"FF",X"11",X"0C",X"0F",X"4F",X"FE",X"ED",X"8F",X"8F",X"CB",X"0F",X"2F",X"6D",
		X"BC",X"3D",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"D3",X"E9",X"FC",X"FE",X"FC",X"FE",X"FE",
		X"E0",X"E0",X"E0",X"C1",X"C1",X"C1",X"D1",X"E0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"9F",X"EF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"81",X"03",X"07",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"01",X"01",X"81",X"91",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"4F",X"1F",X"0F",X"0F",X"1F",X"FF",X"FF",X"0F",X"0F",X"8F",X"0F",X"69",X"9E",X"CF",X"AF",
		X"DF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"00",X"70",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"2F",X"6F",X"0F",X"1E",X"2F",X"EF",X"EF",X"87",X"0F",X"0F",X"0F",X"97",X"F7",X"7F",X"FF",
		X"FF",X"EF",X"EF",X"00",X"C0",X"F0",X"F0",X"F0",X"0F",X"8F",X"8F",X"CF",X"03",X"80",X"F0",X"F0",
		X"0F",X"0F",X"2F",X"1F",X"0F",X"1E",X"EF",X"FF",X"2D",X"0F",X"AD",X"8F",X"0F",X"87",X"69",X"1E",
		X"0C",X"9D",X"1D",X"08",X"0C",X"0E",X"4E",X"2F",X"FF",X"FF",X"77",X"DD",X"FF",X"44",X"01",X"0F",
		X"FF",X"FF",X"FF",X"00",X"10",X"F0",X"F0",X"F0",X"EF",X"DF",X"11",X"00",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"2F",X"6F",X"0F",X"1F",X"3F",X"FF",X"FF",X"0F",X"8F",X"0F",X"3C",X"CF",X"EF",X"EF",X"FF",
		X"0F",X"0F",X"0F",X"1F",X"2F",X"0F",X"0F",X"1F",X"0F",X"2F",X"6F",X"0F",X"0F",X"4F",X"1F",X"3F",
		X"EF",X"DF",X"AE",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"2F",X"6F",X"0F",X"0F",X"3C",X"CF",X"EF",X"0F",X"0F",X"0F",X"2F",X"0F",X"C3",X"4B",X"3C",
		X"FF",X"FF",X"FF",X"EF",X"00",X"F0",X"F0",X"F0",X"8F",X"4F",X"4F",X"EF",X"01",X"E0",X"F0",X"F0",
		X"0F",X"0F",X"4F",X"0F",X"3F",X"0F",X"FE",X"FF",X"0F",X"2D",X"0F",X"8F",X"0F",X"0F",X"F0",X"0F",
		X"1E",X"0F",X"0F",X"4B",X"87",X"97",X"87",X"0F",X"0F",X"0F",X"2D",X"0F",X"8F",X"2F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"1E",X"1E",X"0F",X"0F",X"1E",X"4F",X"4F",X"0F",X"1E",X"2F",X"87",X"87",X"0F",
		X"0F",X"2F",X"CF",X"8F",X"1E",X"1E",X"1E",X"1E",X"87",X"87",X"87",X"87",X"1E",X"2F",X"6F",X"0F",
		X"C3",X"3C",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",X"4F",X"0F",X"C3",X"4B",X"4B",X"87",
		X"EF",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"4F",X"47",X"03",X"03",X"81",X"C1",X"C1",X"E0",
		X"0F",X"0F",X"4B",X"3C",X"8F",X"CF",X"CF",X"DF",X"0F",X"4F",X"2F",X"87",X"87",X"78",X"0F",X"CF",
		X"1F",X"2F",X"5F",X"6E",X"08",X"70",X"F0",X"F0",X"FF",X"FF",X"CC",X"10",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"2F",X"6F",X"0F",X"0F",X"97",X"0F",X"87",X"87",X"0F",X"0F",X"1F",X"3F",X"FF",
		X"2F",X"8F",X"0F",X"0C",X"3B",X"19",X"1D",X"95",X"0F",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"BB",
		X"8F",X"8F",X"8F",X"01",X"00",X"F0",X"F0",X"F0",X"6F",X"6F",X"FF",X"EE",X"00",X"F0",X"F0",X"F0",
		X"0F",X"4F",X"1F",X"0F",X"87",X"69",X"1E",X"1E",X"0F",X"8F",X"0F",X"4F",X"0F",X"0F",X"87",X"7F",
		X"0F",X"0F",X"0F",X"2F",X"0F",X"87",X"78",X"8F",X"0F",X"C3",X"0F",X"0F",X"4F",X"0F",X"1F",X"F7",
		X"7F",X"FF",X"33",X"91",X"E0",X"F0",X"F0",X"F0",X"AF",X"AF",X"FF",X"CF",X"23",X"C0",X"F0",X"F0",
		X"0F",X"2D",X"8F",X"4F",X"0F",X"1F",X"3F",X"7F",X"0F",X"0F",X"0F",X"1F",X"C3",X"4B",X"3C",X"8F",
		X"3F",X"3F",X"3F",X"5F",X"6F",X"23",X"C0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"10",X"F0",
		X"0F",X"4F",X"0F",X"2F",X"4F",X"0F",X"87",X"F3",X"0F",X"4B",X"87",X"0F",X"0F",X"1F",X"FF",X"FF",
		X"1E",X"1F",X"1D",X"3B",X"19",X"0C",X"0F",X"0F",X"0F",X"C3",X"ED",X"FE",X"FE",X"8B",X"07",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"10",X"EE",X"6E",X"DC",X"B8",X"30",X"70",X"F0",X"F0",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"70",X"70",X"70",X"30",X"30",X"98",X"98",X"8C",
		X"77",X"33",X"D1",X"E0",X"F0",X"F0",X"F0",X"F0",X"EE",X"DC",X"B8",X"30",X"F0",X"F0",X"F0",X"F0",
		X"4B",X"2D",X"2D",X"2D",X"1E",X"1E",X"1F",X"3F",X"0F",X"0F",X"0F",X"1F",X"B7",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"2F",X"7F",X"2F",X"0F",X"C3",X"4B",X"2D",X"4B",X"0F",X"0F",X"0F",X"2F",X"0F",X"0F",
		X"FF",X"FF",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"03",X"C0",X"F0",X"F0",X"F0",
		X"0F",X"8F",X"0F",X"2D",X"DE",X"CF",X"EF",X"EF",X"4F",X"AF",X"4F",X"0F",X"87",X"F0",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"00",X"70",X"F0",X"F0",X"F0",X"CC",X"98",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"2D",X"4F",X"4F",X"0F",X"7F",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"BF",
		X"0F",X"2F",X"4F",X"0F",X"0F",X"EF",X"EF",X"FF",X"0F",X"2D",X"0F",X"0F",X"D3",X"5B",X"7B",X"3F",
		X"0F",X"0F",X"0F",X"1F",X"1F",X"37",X"80",X"F0",X"FF",X"FF",X"FF",X"FF",X"7F",X"4C",X"10",X"F0",
		X"4B",X"0F",X"0F",X"8F",X"9F",X"0F",X"87",X"78",X"0F",X"0F",X"2D",X"8F",X"0F",X"8F",X"0F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"FF",X"FF",X"EE",X"CC",X"98",X"70",X"F0",X"F0",
		X"0F",X"8F",X"4F",X"0F",X"0F",X"FF",X"FF",X"FF",X"1E",X"4F",X"CF",X"0F",X"7F",X"FF",X"FF",X"FF",
		X"4F",X"0F",X"0F",X"0F",X"2F",X"4F",X"3F",X"0F",X"3F",X"1F",X"5B",X"87",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"1F",X"0F",X"0F",X"2F",X"6F",X"0F",X"0F",X"2F",X"0F",X"8F",X"0F",X"1F",X"1F",X"3F",X"3F",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"AF",X"47",X"07",X"07",X"07",X"83",X"C1",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"7F",X"FF",X"FF",X"AE",X"AE",X"88",X"70",X"EF",X"DF",X"CC",X"00",X"00",X"30",X"70",X"F0",
		X"0F",X"1F",X"4F",X"6F",X"2F",X"0F",X"0F",X"0F",X"4B",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"6F",
		X"7F",X"9F",X"FF",X"8C",X"10",X"F0",X"F0",X"F0",X"EE",X"DC",X"98",X"70",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"1E",X"6F",X"4F",X"0F",X"97",X"F7",X"7F",X"0F",X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"1F",X"87",X"69",X"3C",X"8F",X"CF",
		X"9F",X"7F",X"3F",X"DF",X"8C",X"98",X"70",X"70",X"FF",X"FF",X"CC",X"00",X"10",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"2F",X"0F",X"0F",X"0F",X"C3",X"0F",X"2D",X"8F",X"0F",X"6F",X"0F",X"ED",X"FF",
		X"BF",X"FF",X"7F",X"CC",X"00",X"30",X"F0",X"F0",X"FF",X"CC",X"00",X"10",X"70",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"2F",X"4F",X"0F",X"1F",X"BF",X"1E",X"4F",X"0F",X"0F",X"0F",X"7F",X"FF",X"FF",
		X"FF",X"EE",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"6F",X"00",X"00",X"80",X"C0",X"F0",X"F0",X"F0",
		X"0F",X"2F",X"0F",X"6F",X"FF",X"FF",X"EF",X"FF",X"3F",X"1F",X"0F",X"C3",X"3C",X"8F",X"CF",X"AF",
		X"CC",X"CC",X"CC",X"CC",X"EE",X"EE",X"6E",X"6E",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",
		X"07",X"91",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"2F",X"CF",X"0F",X"07",X"03",X"01",X"C1",X"E0",
		X"0F",X"0F",X"5B",X"4B",X"2D",X"3C",X"0F",X"0F",X"0F",X"8F",X"0F",X"4F",X"0F",X"0F",X"E1",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"03",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"07",X"03",X"81",X"C1",X"E0",
		X"1E",X"2F",X"6F",X"0F",X"78",X"1E",X"8F",X"8F",X"1E",X"0F",X"0F",X"4F",X"0F",X"C3",X"78",X"1E",
		X"1F",X"8F",X"2F",X"4F",X"0F",X"1F",X"1F",X"3F",X"1F",X"EF",X"7F",X"DF",X"DF",X"FF",X"FF",X"CC",
		X"3F",X"3F",X"DF",X"AF",X"EE",X"CC",X"98",X"70",X"FF",X"EE",X"CC",X"88",X"10",X"70",X"F0",X"F0",
		X"0F",X"0F",X"3F",X"4F",X"0F",X"0F",X"3F",X"3F",X"4B",X"0F",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"8F",X"4F",X"0F",X"C3",X"3F",X"3F",X"0F",X"87",X"4B",X"0F",X"0F",X"0F",X"FF",X"FF",
		X"7F",X"88",X"00",X"30",X"F0",X"F0",X"F0",X"F0",X"BF",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"2F",X"4F",X"4F",X"1F",X"3F",X"FF",X"FF",X"87",X"2F",X"0F",X"3E",X"EF",X"EF",X"DF",X"BF",
		X"00",X"10",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"2F",X"6F",X"0F",X"3F",X"CF",X"FF",X"FF",X"FF",X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"EE",X"18",
		X"0F",X"33",X"01",X"00",X"00",X"00",X"80",X"E0",X"4F",X"8F",X"0F",X"0F",X"07",X"07",X"03",X"03",
		X"0F",X"0F",X"1F",X"2F",X"0F",X"C3",X"0F",X"0F",X"2D",X"4B",X"0F",X"4F",X"0F",X"2F",X"7E",X"9E",
		X"07",X"80",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"1F",X"33",X"C0",X"F0",X"F0",X"F0",X"F0",
		X"4B",X"2D",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"4F",X"CF",X"0F",X"87",X"69",X"3C",X"0F",X"0F",
		X"3F",X"0F",X"0F",X"1F",X"2F",X"0F",X"8F",X"CB",X"0F",X"2D",X"4B",X"0F",X"0F",X"2F",X"6F",X"0F",
		X"67",X"81",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"07",X"03",X"83",X"81",X"E0",
		X"E1",X"3C",X"0F",X"0F",X"0F",X"0F",X"3F",X"2F",X"0F",X"87",X"D3",X"4B",X"69",X"AD",X"1E",X"0F",
		X"FF",X"88",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"EF",X"33",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"8F",X"CF",X"EF",X"FF",X"FF",X"CC",X"B8",X"70",X"3F",X"0F",X"1F",X"0E",X"10",X"F0",X"F0",X"F0",
		X"88",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"67",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"1F",X"87",X"69",X"3C",X"0F",X"8F",X"8F",X"9E",X"8F",X"8F",X"0F",X"D3",X"B7",X"7F",X"5F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"8F",X"01",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"81",X"C1",
		X"0F",X"0F",X"0F",X"E1",X"1E",X"0F",X"0F",X"8F",X"1E",X"4F",X"AF",X"0F",X"0F",X"C3",X"3C",X"1E",
		X"FF",X"FF",X"CC",X"10",X"F0",X"F0",X"F0",X"F0",X"BF",X"19",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"98",X"70",X"F0",X"88",X"10",X"10",X"30",X"70",X"F0",X"F0",X"F0",
		X"9F",X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"CC",X"88",
		X"0F",X"4F",X"0F",X"1F",X"2F",X"4F",X"2F",X"0F",X"2D",X"4B",X"0F",X"0F",X"0F",X"1F",X"3F",X"7F",
		X"3F",X"BF",X"DF",X"37",X"80",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"88",X"70",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"2F",X"5F",X"0F",X"87",X"F1",X"1F",X"0F",X"C3",X"0F",X"0F",X"2F",X"0F",X"3F",X"FF",
		X"07",X"03",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"3F",X"DF",X"57",X"00",X"F0",X"F0",X"F0",X"F0",
		X"4B",X"2D",X"1E",X"0F",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"97",X"1F",X"C3",X"4B",X"3C",
		X"4B",X"0F",X"8F",X"1F",X"1F",X"0F",X"87",X"4B",X"0F",X"0F",X"4B",X"8F",X"0F",X"1E",X"2F",X"0F",
		X"6F",X"7F",X"4C",X"00",X"F0",X"F0",X"F0",X"F0",X"FF",X"7F",X"7F",X"00",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"7F",X"BF",X"00",X"F0",X"F0",X"F0",X"F0",X"3F",X"9F",X"88",X"70",X"F0",X"F0",X"F0",X"F0",
		X"EF",X"77",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"8F",X"4F",X"4F",X"47",X"23",X"C1",X"E0",X"E0",
		X"0F",X"5E",X"4F",X"0F",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"C3",X"78",X"0F",X"8F",
		X"0F",X"07",X"33",X"91",X"C0",X"F0",X"F0",X"F0",X"7F",X"FF",X"FF",X"BF",X"57",X"80",X"F0",X"F0",
		X"87",X"4B",X"2D",X"2D",X"1E",X"0F",X"0F",X"0F",X"0F",X"2F",X"4F",X"2F",X"87",X"87",X"4B",X"3D",
		X"3C",X"3F",X"3B",X"11",X"1D",X"0E",X"4E",X"2F",X"4B",X"E5",X"FE",X"FE",X"CD",X"8B",X"17",X"0F",
		X"0F",X"0F",X"07",X"00",X"E0",X"F0",X"F0",X"F0",X"1F",X"1F",X"0F",X"07",X"01",X"80",X"F0",X"F0",
		X"0F",X"0F",X"1F",X"2F",X"1F",X"87",X"69",X"1E",X"1E",X"2D",X"8F",X"0F",X"0F",X"0F",X"0F",X"F1",
		X"EF",X"4C",X"88",X"00",X"00",X"00",X"30",X"70",X"0F",X"01",X"00",X"00",X"10",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"78",X"3F",X"DF",X"CF",X"EF",X"0F",X"2F",X"0F",X"C3",X"F8",X"8F",X"CF",X"8F",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"CC",X"CC",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"7F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"EE",X"B8",X"B8",X"70",X"70",X"70",X"70",X"70",X"70",
		X"FF",X"FF",X"7F",X"37",X"00",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"00",X"70",X"F0",X"F0",X"F0",
		X"0F",X"2D",X"0F",X"8F",X"0F",X"0F",X"1F",X"FF",X"0F",X"0F",X"0F",X"8F",X"0F",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"18",X"0F",X"DB",X"ED",X"ED",X"ED",X"DB",X"CB",X"A7",X"0F",
		X"C3",X"CB",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"0F",X"9F",X"0F",X"2F",X"87",X"87",X"DB",X"CB",
		X"33",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"BF",X"DF",X"33",X"80",X"F0",X"F0",X"F0",X"F0",
		X"2D",X"2D",X"4B",X"3C",X"1E",X"0F",X"3F",X"3F",X"4F",X"0F",X"0F",X"2F",X"0F",X"0F",X"EF",X"DF",
		X"0F",X"0F",X"3F",X"6F",X"0F",X"87",X"4B",X"2D",X"2D",X"4B",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",
		X"FF",X"FF",X"FF",X"88",X"00",X"30",X"F0",X"F0",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",
		X"87",X"0F",X"1F",X"2F",X"8F",X"0F",X"0F",X"FF",X"0F",X"69",X"0F",X"CF",X"0F",X"0F",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"7F",X"9F",X"CC",X"10",X"F0",X"F0",X"EE",X"EE",X"98",X"30",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"2F",X"4F",X"2F",X"0F",X"1F",X"FF",X"5B",X"B7",X"3F",X"3F",X"7F",X"5F",X"EF",X"FF",
		X"0F",X"1F",X"11",X"00",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"2F",X"6F",X"0F",X"C3",X"69",X"1E",X"0F",X"4B",X"0F",X"0F",X"2F",X"4F",X"0F",X"F7",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E0",X"00",X"00",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"0D",X"89",X"89",X"CD",X"CD",X"EF",X"EF",
		X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",X"EF",X"EE",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"7C",X"7C",X"7C",X"F0",X"F0",X"1F",X"1F",X"1F",
		X"EF",X"EF",X"CF",X"CF",X"8F",X"8F",X"0F",X"0F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"BC",X"FC",X"7C",X"7C",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",
		X"3F",X"0F",X"3C",X"3C",X"0C",X"0C",X"3C",X"3F",X"FF",X"0F",X"F0",X"F0",X"00",X"00",X"F0",X"FF",
		X"3F",X"3F",X"0F",X"3C",X"3C",X"0F",X"3F",X"3F",X"FF",X"FF",X"0F",X"F0",X"F0",X"0F",X"FF",X"FF",
		X"00",X"08",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"6D",X"6D",X"4F",X"0F",X"87",X"87",X"87",X"87",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"87",X"87",X"4B",X"2D",X"6D",X"6D",X"6D",X"6D",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"0F",X"2F",X"6E",X"0E",X"4C",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"4F",X"4F",X"1F",X"3F",X"4F",X"1F",X"2F",X"8F",X"CF",X"0E",X"4E",X"0C",X"0C",X"08",X"08",
		X"3D",X"4F",X"1F",X"4B",X"1E",X"6F",X"3F",X"8F",X"6B",X"1E",X"CF",X"2F",X"8F",X"D3",X"0F",X"4F",
		X"2F",X"2D",X"1F",X"4F",X"1E",X"3D",X"1F",X"87",X"A7",X"0F",X"FA",X"8F",X"4F",X"5F",X"0F",X"2F",
		X"0F",X"2F",X"BF",X"0F",X"2F",X"4F",X"1F",X"0F",X"08",X"08",X"0C",X"0C",X"CE",X"0E",X"8F",X"CF",
		X"08",X"08",X"0C",X"0C",X"4E",X"4E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"0F",X"0F",X"D3",X"D3",X"D3",X"D3",X"D3",X"D3",X"0F",X"0F",
		X"FF",X"0F",X"F0",X"F0",X"00",X"00",X"F0",X"FF",X"FF",X"0F",X"F0",X"F0",X"00",X"00",X"F0",X"FF",
		X"C8",X"C8",X"48",X"C0",X"C0",X"48",X"C8",X"C8",X"D3",X"D3",X"C3",X"D2",X"D2",X"C3",X"D3",X"D3",
		X"00",X"00",X"BC",X"C8",X"C8",X"C8",X"C8",X"C8",X"00",X"00",X"1F",X"D3",X"D3",X"D3",X"D3",X"D3",
		X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"D3",X"D3",X"D3",X"D3",X"D3",X"D3",X"D3",X"D3",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"62",X"62",X"62",X"06",X"02",X"10",X"10",X"10",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"10",X"10",X"20",X"60",X"62",X"62",X"62",X"62",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"BF",X"FF",X"F7",X"D7",X"F3",X"F3",X"F1",X"F1",
		X"DF",X"FF",X"E7",X"F7",X"F3",X"F3",X"F1",X"F1",X"FF",X"DF",X"FF",X"6F",X"FF",X"EF",X"EF",X"FF",
		X"DF",X"BB",X"EE",X"BF",X"EF",X"BB",X"DD",X"FF",X"BF",X"EF",X"77",X"DD",X"57",X"BF",X"FF",X"BB",
		X"FF",X"DD",X"44",X"DF",X"BF",X"EE",X"FF",X"5F",X"BF",X"7F",X"FF",X"BB",X"EF",X"FF",X"6F",X"BB",
		X"F1",X"F1",X"F3",X"D3",X"F7",X"F7",X"FF",X"DF",X"BF",X"EF",X"FF",X"3F",X"EF",X"DF",X"FF",X"EF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F3",X"F3",X"F7",X"C7",X"FF",X"FF",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"0F",X"0F",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"0F",X"0F",
		X"DE",X"DE",X"0F",X"F0",X"F0",X"0F",X"DE",X"DE",X"B7",X"B7",X"0F",X"F0",X"F0",X"0F",X"B7",X"B7",
		X"CF",X"0F",X"F0",X"F0",X"00",X"00",X"F0",X"CF",X"3F",X"0F",X"F0",X"F0",X"00",X"00",X"F0",X"3F",
		X"00",X"00",X"CF",X"DE",X"DE",X"DE",X"DE",X"DE",X"00",X"00",X"3F",X"B7",X"B7",X"B7",X"B7",X"B7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"9F",X"9F",X"DF",X"DF",X"FF",X"EF",
		X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",X"EF",X"EF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"EF",X"EF",X"CF",X"CF",X"8F",X"8F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"DF",X"DF",X"9F",X"9F",X"1F",X"1F",
		X"8B",X"B8",X"B8",X"B8",X"90",X"C0",X"E0",X"E0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"80",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"90",X"90",X"80",X"C3",X"90",X"90",X"90",X"90",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"90",X"90",X"90",X"90",X"80",X"C3",X"90",X"90",X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",
		X"C3",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"0E",X"BF",X"BC",X"B8",X"B8",X"B8",X"88",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"DE",X"9E",X"3C",X"F0",X"E1",X"0F",X"FF",X"FF",X"B7",X"B7",X"B7",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"DE",X"DE",X"1E",X"D2",X"D2",X"1E",X"DE",X"DE",X"B7",X"B7",X"87",X"96",X"96",X"87",X"B7",X"B7",
		X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"0F",X"0F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"0E",
		X"0F",X"0F",X"F0",X"F0",X"00",X"00",X"F0",X"0F",X"CC",X"0C",X"84",X"84",X"40",X"40",X"84",X"CC",
		X"FF",X"B8",X"A8",X"A8",X"08",X"C0",X"80",X"80",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0E",X"0E",X"0C",X"0C",X"08",X"08",
		X"80",X"08",X"CC",X"0C",X"A8",X"A8",X"B8",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"DD",X"5D",X"DD",X"DD",X"DD",X"2B",X"0F",X"8F",X"4F",X"1E",X"6F",X"0F",X"3E",X"4F",X"0F",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"C0",X"90",X"34",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"30",
		X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F3",X"F3",X"11",X"0F",X"F3",X"F3",X"F3",X"F3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F3",X"F3",X"F3",X"F3",X"11",X"0F",X"F3",X"F3",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"3C",X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"CC",X"0C",X"0C",X"84",X"84",X"0C",X"CC",X"CC",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"0F",X"8F",X"9F",X"FD",X"DF",X"FF",X"EF",
		X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",X"EF",X"EF",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EE",X"CC",X"CC",X"8E",X"8E",X"0E",X"F0",
		X"00",X"00",X"9F",X"69",X"69",X"69",X"69",X"69",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"7F",X"A6",X"A6",X"A6",X"86",X"70",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"10",X"F0",X"F0",X"F0",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"F0",X"F0",X"3F",X"3F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"F0",X"F0",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",
		X"F0",X"0F",X"FF",X"2F",X"A6",X"A6",X"A6",X"A6",X"F0",X"0F",X"FF",X"1F",X"E1",X"E1",X"E1",X"00",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"33",X"C0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"11",X"80",X"F0",X"F0",
		X"0F",X"0F",X"1F",X"2F",X"0F",X"0F",X"FF",X"FF",X"08",X"08",X"0C",X"0C",X"0E",X"EE",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"77",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"C0",X"80",X"80",
		X"F0",X"F0",X"0F",X"0F",X"FF",X"F0",X"F0",X"F0",X"80",X"80",X"0C",X"0C",X"EE",X"E0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"EF",X"CF",X"DE",X"DE",X"DE",X"FF",X"FF",X"0F",X"78",X"F0",X"C3",X"97",X"B7",
		X"F0",X"B7",X"93",X"81",X"80",X"90",X"B0",X"F0",X"F0",X"FE",X"DE",X"9E",X"1E",X"96",X"D2",X"F0",
		X"FF",X"B8",X"B8",X"B8",X"08",X"F0",X"F0",X"F0",X"FF",X"E1",X"E1",X"E1",X"10",X"F0",X"F0",X"F0",
		X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"0F",X"37",X"61",X"54",X"54",X"40",X"73",X"00",X"0F",X"CF",X"0F",X"A7",X"A7",X"61",X"CF",X"01",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",
		X"F0",X"0F",X"FF",X"0F",X"B8",X"B8",X"B8",X"88",X"F0",X"0F",X"FF",X"0F",X"E1",X"E1",X"E1",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"F0",X"F0",X"00",X"00",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"F0",X"F0",X"F0",X"FF",X"FF",X"EE",X"0E",X"0C",X"C0",X"80",X"80",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"4B",X"1E",X"BE",X"AF",X"8F",X"9E",X"AF",X"8F",
		X"0F",X"0F",X"8F",X"FF",X"FF",X"CF",X"EF",X"EF",X"7C",X"7C",X"7C",X"E8",X"FC",X"1F",X"1F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"EF",X"EF",X"CC",X"CC",X"88",X"8F",X"0F",X"0F",X"1F",X"1F",X"01",X"03",X"00",X"7C",X"7C",X"7C",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",
		X"FF",X"FF",X"0F",X"F0",X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"0F",X"F0",X"F0",X"0F",X"FF",X"FF",
		X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",
		X"CF",X"CF",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"F0",X"F0",
		X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"F0",X"F0",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"0F",X"87",X"C2",X"D3",X"D3",X"C3",X"80",X"00",X"0F",X"1E",X"30",X"B8",X"B8",X"3C",X"10",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7C",X"7C",X"E8",X"E8",X"DF",X"DF",X"FF",X"EF",
		X"00",X"00",X"88",X"88",X"CC",X"CF",X"EF",X"EF",X"00",X"00",X"00",X"03",X"03",X"7C",X"7C",X"7C",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"0F",X"1F",X"2F",X"8F",X"CF",X"67",X"23",X"33",X"4B",X"9E",X"4B",X"2D",X"CF",X"4F",X"1F",X"0F",
		X"10",X"20",X"20",X"02",X"40",X"84",X"0C",X"08",X"10",X"10",X"10",X"31",X"20",X"62",X"40",X"84",
		X"0C",X"0C",X"0C",X"0C",X"08",X"08",X"18",X"18",X"62",X"62",X"44",X"C4",X"80",X"88",X"88",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"08",X"00",X"00",X"10",X"10",X"11",X"31",X"20",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"3E",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",
		X"3C",X"3C",X"9E",X"0F",X"6D",X"1F",X"AD",X"3E",X"78",X"F0",X"F0",X"F0",X"78",X"B4",X"8F",X"2F",
		X"0F",X"5A",X"A5",X"1E",X"3C",X"E1",X"2D",X"78",X"68",X"E0",X"C0",X"C1",X"40",X"E0",X"E0",X"A1",
		X"0F",X"0F",X"2D",X"1F",X"6B",X"2F",X"87",X"5A",X"0F",X"5B",X"3F",X"87",X"DB",X"2D",X"4B",X"2C",
		X"0F",X"97",X"0F",X"2F",X"5A",X"0F",X"5F",X"87",X"DB",X"CB",X"87",X"6D",X"4F",X"87",X"3D",X"7B",
		X"C0",X"F0",X"D0",X"78",X"E0",X"D2",X"F0",X"3C",X"07",X"00",X"F0",X"E1",X"D0",X"E1",X"69",X"D2",
		X"2B",X"3B",X"23",X"3B",X"19",X"4C",X"A6",X"C3",X"0F",X"0F",X"AF",X"DF",X"FF",X"FF",X"00",X"4D",
		X"2D",X"4F",X"1F",X"4B",X"1E",X"6F",X"3F",X"00",X"4B",X"3C",X"CF",X"2F",X"87",X"D3",X"0F",X"00",
		X"2D",X"5E",X"6F",X"2F",X"2D",X"4F",X"1F",X"3F",X"6F",X"9F",X"2F",X"9E",X"4F",X"B4",X"69",X"4B",
		X"8F",X"69",X"0F",X"6F",X"0F",X"BF",X"2F",X"0F",X"6F",X"1F",X"2F",X"87",X"4B",X"0F",X"9E",X"2D",
		X"3C",X"2F",X"6F",X"1E",X"AD",X"4F",X"1F",X"7F",X"6F",X"4F",X"0F",X"4F",X"DB",X"0F",X"5A",X"69",
		X"2D",X"4F",X"5E",X"96",X"1F",X"4F",X"97",X"2F",X"8F",X"CF",X"2F",X"C7",X"0F",X"4F",X"1E",X"2D",
		X"8F",X"8F",X"0F",X"0F",X"0F",X"0E",X"0E",X"1D",X"0F",X"0F",X"0F",X"07",X"07",X"CF",X"CF",X"8F",
		X"0F",X"0E",X"0E",X"1D",X"1D",X"3B",X"0B",X"47",X"34",X"9E",X"1E",X"0F",X"0F",X"0F",X"0E",X"0E",
		X"56",X"56",X"DE",X"8F",X"8F",X"0F",X"0F",X"0F",X"2C",X"86",X"86",X"D1",X"C1",X"2B",X"29",X"74",
		X"2C",X"86",X"95",X"D1",X"D1",X"7B",X"2B",X"3A",X"FC",X"F8",X"F8",X"F0",X"F0",X"78",X"78",X"3C",
		X"78",X"78",X"78",X"F0",X"F0",X"F8",X"F8",X"FC",X"F7",X"F7",X"F3",X"F3",X"F1",X"F1",X"70",X"30",
		X"7F",X"7F",X"7B",X"3F",X"3D",X"3D",X"3C",X"78",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"70",X"70",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"2E",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"3F",X"35",X"35",X"34",
		X"1E",X"39",X"3B",X"3B",X"3B",X"08",X"86",X"2D",X"87",X"E9",X"FE",X"ED",X"FE",X"DC",X"03",X"0F",
		X"1E",X"19",X"1D",X"11",X"19",X"08",X"0C",X"0D",X"87",X"E9",X"FE",X"FE",X"ED",X"FE",X"32",X"09",
		X"3C",X"3F",X"33",X"77",X"33",X"3B",X"19",X"0C",X"A7",X"CB",X"ED",X"FE",X"FE",X"ED",X"03",X"17",
		X"2D",X"5E",X"6F",X"2F",X"2D",X"4F",X"1F",X"00",X"6F",X"9F",X"2F",X"9E",X"4F",X"B4",X"4B",X"00",
		X"2D",X"4F",X"1F",X"4B",X"1E",X"6F",X"3F",X"8F",X"4B",X"3C",X"CF",X"2F",X"87",X"D3",X"0F",X"4F",
		X"2F",X"69",X"1F",X"4F",X"1E",X"69",X"97",X"87",X"A7",X"0F",X"DA",X"AD",X"4F",X"5F",X"0F",X"2F",
		X"0F",X"2F",X"BF",X"0F",X"5B",X"4F",X"1F",X"A5",X"C3",X"D7",X"0F",X"2F",X"5E",X"2D",X"9E",X"CF",
		X"0F",X"2F",X"5B",X"0F",X"6D",X"C7",X"1F",X"0F",X"5E",X"0F",X"3F",X"4B",X"AF",X"B4",X"2F",X"8F",
		X"FE",X"DE",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"96",X"96",X"C3",X"C3",X"69",X"68",X"0C",
		X"2C",X"86",X"95",X"D1",X"B3",X"77",X"FF",X"EF",X"76",X"FF",X"FE",X"FC",X"F8",X"F8",X"78",X"3C",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"78",X"78",X"3C",X"87",X"87",X"C3",X"C3",X"E1",X"A1",X"B0",X"76",
		X"86",X"86",X"D1",X"D1",X"A3",X"A3",X"74",X"74",X"07",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"3B",X"19",X"1D",X"1D",X"0C",X"0E",X"0E",X"0F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"56",X"56",
		X"B3",X"B3",X"33",X"77",X"FF",X"77",X"77",X"3B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"86",X"86",X"C3",X"C2",X"C0",X"D1",X"91",X"FF",X"FF",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"87",X"C3",X"43",X"43",X"61",X"21",X"21",X"30",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"3F",X"5B",X"8F",X"3C",X"78",X"C3",X"C7",X"2F",X"FF",X"CF",X"78",X"F2",X"5A",X"AF",X"CF",X"8F",
		X"0F",X"CB",X"2F",X"2E",X"BB",X"6F",X"BF",X"FF",X"CB",X"1F",X"CC",X"00",X"EE",X"CC",X"8C",X"5D",
		X"21",X"87",X"A7",X"C3",X"A5",X"C3",X"96",X"69",X"69",X"1E",X"8F",X"BF",X"2F",X"0F",X"9E",X"2F",
		X"0F",X"2F",X"BF",X"2D",X"5B",X"4F",X"1F",X"00",X"C3",X"D7",X"0F",X"2F",X"5E",X"2D",X"9E",X"00",
		X"D8",X"D8",X"D8",X"D8",X"D9",X"C8",X"B8",X"FF",X"F1",X"F2",X"F4",X"F8",X"F0",X"00",X"F0",X"FF",
		X"D8",X"D8",X"D8",X"D8",X"D8",X"D8",X"D8",X"D8",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"0F",X"FF",X"F8",X"D8",X"C8",X"D8",X"D8",X"D8",X"0F",X"FF",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",
		X"0F",X"FF",X"F0",X"F0",X"F0",X"00",X"F0",X"FF",X"0F",X"FF",X"F0",X"F0",X"F0",X"00",X"F0",X"FF",
		X"F0",X"F0",X"E0",X"C0",X"91",X"33",X"67",X"CF",X"91",X"33",X"67",X"CF",X"8F",X"0F",X"0F",X"0F",
		X"87",X"87",X"C3",X"C3",X"E1",X"E1",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"91",X"D1",X"59",X"48",X"2C",X"2C",X"0E",X"0F",
		X"E0",X"E0",X"68",X"78",X"3C",X"3C",X"1E",X"1E",X"FF",X"FF",X"77",X"77",X"77",X"33",X"B3",X"B3",
		X"8F",X"CF",X"03",X"83",X"81",X"C1",X"C1",X"C0",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"8F",X"8F",X"8F",X"CF",X"CF",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"8F",X"2F",X"9F",X"6B",X"9F",X"FF",X"FE",X"FC",X"E2",X"6A",X"4A",X"5B",X"D3",X"97",X"87",X"2D",
		X"88",X"6E",X"2C",X"F3",X"A7",X"8F",X"7C",X"97",X"00",X"00",X"00",X"88",X"4C",X"CC",X"4C",X"6A",
		X"2F",X"FF",X"00",X"00",X"00",X"19",X"11",X"44",X"2F",X"EF",X"11",X"00",X"00",X"00",X"88",X"88",
		X"3C",X"2F",X"6F",X"1E",X"AD",X"4F",X"1F",X"00",X"6F",X"4F",X"0F",X"4F",X"DB",X"0F",X"5A",X"00",
		X"68",X"68",X"68",X"68",X"68",X"48",X"78",X"0F",X"B7",X"97",X"87",X"F0",X"00",X"00",X"F0",X"0F",
		X"78",X"0F",X"4B",X"69",X"68",X"68",X"68",X"68",X"F0",X"0F",X"0F",X"0F",X"F0",X"84",X"97",X"B7",
		X"DC",X"9C",X"1C",X"F0",X"00",X"00",X"F0",X"0F",X"1E",X"1E",X"1E",X"1E",X"1E",X"16",X"D2",X"0F",
		X"F0",X"0F",X"0F",X"0F",X"F0",X"10",X"9C",X"DC",X"F0",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F7",X"F7",X"F3",X"73",X"73",X"F3",X"F7",X"CF",X"FF",X"FF",X"FF",X"EF",X"CF",X"8F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",
		X"0F",X"8F",X"8F",X"8F",X"CF",X"CF",X"CF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"4F",X"5F",X"8F",X"0F",X"2D",X"1E",X"6F",X"0F",X"87",X"1F",X"0F",X"6D",X"CB",X"1E",X"3E",X"2F",
		X"44",X"55",X"33",X"7F",X"BF",X"FF",X"AA",X"EF",X"47",X"47",X"16",X"07",X"9F",X"9E",X"2F",X"4F",
		X"00",X"00",X"00",X"00",X"22",X"00",X"44",X"00",X"47",X"23",X"23",X"23",X"23",X"23",X"23",X"67",
		X"3E",X"2F",X"8F",X"67",X"11",X"00",X"00",X"00",X"0F",X"2D",X"AD",X"4F",X"1E",X"8F",X"57",X"47",
		X"0F",X"0F",X"2F",X"6D",X"5A",X"AF",X"0F",X"4B",X"C1",X"F0",X"68",X"3C",X"1E",X"6B",X"8F",X"0F",
		X"1E",X"3C",X"3C",X"2D",X"3C",X"3C",X"1E",X"1E",X"68",X"94",X"50",X"E0",X"B0",X"D2",X"E0",X"B4",
		X"4B",X"8F",X"2D",X"4F",X"1E",X"0F",X"2D",X"0F",X"4B",X"1F",X"0F",X"2D",X"4F",X"0F",X"5A",X"F0",
		X"D8",X"D8",X"D0",X"E0",X"F0",X"00",X"F0",X"FF",X"E3",X"E3",X"E3",X"E3",X"63",X"23",X"E3",X"EF",
		X"0F",X"FF",X"F0",X"F0",X"F0",X"10",X"D0",X"D0",X"0F",X"EF",X"E7",X"EB",X"E3",X"E3",X"E3",X"E3",
		X"2D",X"4F",X"1F",X"4B",X"1E",X"6F",X"3F",X"07",X"4B",X"3C",X"CF",X"0F",X"87",X"D3",X"0F",X"4F",
		X"25",X"56",X"67",X"27",X"25",X"47",X"17",X"37",X"6F",X"9F",X"2F",X"9E",X"4F",X"B4",X"69",X"4B",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"8F",X"0F",X"FF",X"FF",X"8F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"4F",X"FF",X"FF",X"8F",X"0F",X"0F",X"FF",
		X"0F",X"7F",X"7F",X"4F",X"0F",X"0F",X"0F",X"0F",X"1F",X"FF",X"FF",X"0F",X"0F",X"0F",X"7F",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"8F",X"0F",X"8F",X"8F",X"DF",X"AF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"7F",X"0F",X"0F",X"7F",X"FF",X"8F",X"4F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"EF",X"8F",X"0F",X"7F",X"FF",X"8F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"EF",X"1F",X"3F",X"EF",X"BF",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7F",X"FF",X"8F",X"4F",X"FF",X"FF",X"8F",
		X"2F",X"0F",X"0F",X"DF",X"DF",X"1F",X"0F",X"0F",X"1F",X"0F",X"1F",X"FF",X"FF",X"1F",X"0F",X"0F",
		X"0F",X"0F",X"1F",X"3F",X"2F",X"1F",X"3F",X"3F",X"0F",X"1F",X"FF",X"FF",X"0F",X"1F",X"FF",X"FF",
		X"1F",X"0F",X"0F",X"1F",X"1F",X"FF",X"7F",X"1F",X"EF",X"0F",X"0F",X"2F",X"1F",X"FF",X"EF",X"0F",
		X"0F",X"0F",X"0F",X"1F",X"3F",X"2F",X"2F",X"3F",X"0F",X"0F",X"0F",X"EF",X"FF",X"1F",X"1F",X"FF",
		X"F0",X"B0",X"F0",X"5A",X"F0",X"3C",X"4F",X"1F",X"00",X"B0",X"52",X"F0",X"A5",X"D2",X"4B",X"8F",
		X"07",X"61",X"07",X"67",X"07",X"36",X"27",X"07",X"6F",X"3F",X"4F",X"2F",X"87",X"4B",X"9E",X"2D",
		X"34",X"27",X"67",X"16",X"25",X"47",X"17",X"77",X"6F",X"4F",X"0F",X"4F",X"DB",X"0F",X"5A",X"69",
		X"25",X"47",X"56",X"16",X"17",X"47",X"17",X"27",X"8F",X"CF",X"2F",X"C7",X"0F",X"4F",X"1E",X"2D",
		X"8F",X"8F",X"4F",X"CF",X"8F",X"0F",X"0F",X"0F",X"3F",X"2F",X"0F",X"0F",X"3F",X"2F",X"0F",X"0F",
		X"0F",X"4F",X"CF",X"CF",X"4F",X"0F",X"4F",X"CF",X"2F",X"3F",X"1F",X"0F",X"2F",X"3F",X"0F",X"0F",
		X"4F",X"CF",X"CF",X"4F",X"0F",X"4F",X"CF",X"CF",X"0F",X"3F",X"3F",X"2F",X"0F",X"1F",X"3F",X"2F",
		X"CF",X"DF",X"5F",X"1F",X"4F",X"CF",X"8F",X"0F",X"0F",X"FF",X"FF",X"0F",X"0F",X"1F",X"3F",X"1F",
		X"DF",X"9F",X"1F",X"4F",X"CF",X"CF",X"0F",X"4F",X"FF",X"FF",X"1F",X"2F",X"2F",X"3F",X"1F",X"0F",
		X"8F",X"0F",X"0F",X"0F",X"8F",X"CF",X"4F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"CF",X"8F",X"0F",X"0F",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"4F",X"CF",X"CF",X"0F",X"4F",X"CF",X"CF",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"8F",X"0F",X"1F",X"0F",X"0F",X"FF",X"FF",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",
		X"3B",X"3B",X"19",X"19",X"4C",X"A6",X"D3",X"E1",X"0F",X"5F",X"AF",X"EF",X"FF",X"33",X"00",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"0F",X"0F",X"3F",X"1F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",
		X"4B",X"8F",X"1E",X"3D",X"6B",X"E7",X"E7",X"7F",X"0F",X"E1",X"96",X"0F",X"4B",X"2F",X"5E",X"0F",
		X"0F",X"3D",X"4F",X"0F",X"7F",X"CC",X"11",X"1F",X"5E",X"87",X"1F",X"FF",X"CC",X"00",X"DF",X"77",
		X"16",X"0F",X"A7",X"1F",X"0F",X"4B",X"87",X"1E",X"97",X"5B",X"2F",X"4F",X"0F",X"AD",X"6D",X"4F",
		X"8F",X"CF",X"3F",X"EF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1F",X"FF",X"EF",X"0F",X"0F",X"8F",X"7F",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"9F",X"FF",X"FF",X"1F",X"0F",X"EF",X"FF",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1F",X"FF",X"FF",X"1F",X"0F",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"2F",X"1F",X"1F",X"FF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"3F",X"3F",X"0F",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"2F",X"8F",X"4F",X"0F",X"9F",X"FE",X"FE",X"69",X"F3",X"E3",X"7B",X"FB",X"D5",X"3F",X"3F",X"2F",
		X"88",X"4C",X"F3",X"78",X"3C",X"9E",X"2F",X"4F",X"00",X"00",X"00",X"88",X"C4",X"C4",X"E2",X"6A",
		X"0F",X"0F",X"CF",X"8F",X"8F",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",X"CF",X"CF",X"4F",
		X"0F",X"FF",X"FF",X"8F",X"0F",X"FF",X"FF",X"8F",X"4F",X"CF",X"8F",X"8F",X"4F",X"CF",X"8F",X"0F",
		X"6F",X"EF",X"4F",X"2F",X"FF",X"FF",X"8F",X"0F",X"0F",X"0F",X"0F",X"4F",X"CF",X"CF",X"4F",X"0F",
		X"0F",X"0F",X"4F",X"4F",X"FF",X"FF",X"4F",X"0F",X"4F",X"0F",X"8F",X"4F",X"CF",X"8F",X"0F",X"0F",
		X"0F",X"0F",X"7F",X"FF",X"8F",X"4F",X"FF",X"FF",X"0F",X"4F",X"CF",X"CF",X"0F",X"4F",X"CF",X"CF",
		X"0F",X"6F",X"6F",X"AF",X"AF",X"AF",X"7F",X"3F",X"0F",X"8F",X"8F",X"4F",X"4F",X"4F",X"8F",X"0F",
		X"0F",X"6F",X"EF",X"4F",X"2F",X"FF",X"FF",X"8F",X"0F",X"0F",X"0F",X"0F",X"4F",X"CF",X"CF",X"4F",
		X"0F",X"1E",X"FF",X"00",X"00",X"00",X"44",X"2A",X"97",X"2F",X"CF",X"33",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
