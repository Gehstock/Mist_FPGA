library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"B0",X"60",X"C0",X"80",X"C0",X"90",X"30",X"70",X"C0",X"80",X"40",X"C0",X"90",X"34",X"74",X"FC",
		X"90",X"30",X"70",X"F0",X"B0",X"B0",X"60",X"30",X"F0",X"F0",X"B0",X"60",X"C0",X"C0",X"90",X"30",
		X"F0",X"70",X"74",X"94",X"94",X"C4",X"44",X"40",X"BC",X"F9",X"F9",X"F9",X"F9",X"79",X"79",X"9C",
		X"80",X"80",X"80",X"C0",X"60",X"60",X"B0",X"B0",X"90",X"C0",X"40",X"40",X"00",X"80",X"80",X"C0",
		X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"9C",X"C4",X"44",X"44",X"00",X"04",X"04",X"04",
		X"30",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"04",X"04",X"0C",X"C9",X"0C",X"09",X"09",X"09",X"07",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"69",X"B9",X"F7",X"F7",X"F7",X"F7",X"F7",X"FF",X"CF",X"6B",X"BB",X"FB",X"FB",X"FB",X"F6",X"F6",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"B0",X"F4",X"F4",X"F4",X"F4",X"F4",X"FC",X"F9",
		X"FF",X"7F",X"9F",X"CB",X"0B",X"0B",X"0B",X"0B",X"F6",X"F6",X"36",X"CC",X"C8",X"08",X"08",X"08",
		X"90",X"C0",X"00",X"04",X"04",X"04",X"04",X"04",X"79",X"99",X"C9",X"09",X"09",X"07",X"07",X"07",
		X"0B",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"08",X"08",X"08",X"00",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"0C",X"0C",X"8C",X"CC",X"CC",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"87",
		X"06",X"06",X"06",X"46",X"46",X"C6",X"96",X"36",X"04",X"44",X"C4",X"94",X"94",X"34",X"74",X"F4",
		X"69",X"B9",X"B9",X"B9",X"B9",X"69",X"C9",X"89",X"8F",X"CF",X"CF",X"CF",X"CF",X"8F",X"4F",X"CF",
		X"76",X"F6",X"F6",X"F6",X"F6",X"B6",X"36",X"66",X"F4",X"F4",X"F4",X"B4",X"34",X"64",X"C4",X"C4",
		X"49",X"C9",X"99",X"39",X"79",X"F9",X"F9",X"FC",X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"B7",
		X"C6",X"C6",X"36",X"F6",X"FB",X"FB",X"FB",X"FB",X"C4",X"C0",X"38",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"6C",X"3C",X"FC",X"F4",X"F4",X"F4",X"F4",X"F4",X"C7",X"67",X"37",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"FB",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"F7",X"F8",X"F8",X"FC",X"F6",X"B6",X"36",X"36",X"36",
		X"F4",X"74",X"74",X"90",X"90",X"40",X"40",X"00",X"F7",X"F9",X"F9",X"F9",X"F9",X"79",X"79",X"9C",
		X"77",X"77",X"97",X"99",X"49",X"49",X"09",X"0C",X"B6",X"BB",X"FB",X"7B",X"3B",X"CF",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"44",X"44",X"04",X"04",X"00",X"00",X"00",
		X"0C",X"04",X"C4",X"34",X"F4",X"F0",X"F0",X"F0",X"07",X"07",X"C7",X"C9",X"39",X"F9",X"FC",X"FC",
		X"80",X"C0",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"C0",X"60",X"B0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"30",X"C0",X"40",X"00",X"F4",X"F4",X"F4",X"F4",X"74",X"94",X"CC",X"0C",
		X"F0",X"F0",X"F0",X"30",X"C0",X"40",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"90",X"C0",X"00",X"00",
		X"34",X"64",X"CC",X"0C",X"09",X"03",X"C7",X"67",X"39",X"99",X"C7",X"07",X"0F",X"0F",X"0F",X"8F",
		X"F0",X"F0",X"30",X"60",X"C0",X"80",X"40",X"C4",X"F0",X"30",X"60",X"C0",X"04",X"04",X"CC",X"39",
		X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"6F",X"3F",X"FF",X"FB",X"FB",X"FF",X"FF",
		X"34",X"74",X"FC",X"FC",X"FC",X"FC",X"3C",X"34",X"F9",X"F3",X"F7",X"F7",X"F7",X"F7",X"77",X"37",
		X"7F",X"3F",X"37",X"B7",X"F3",X"F9",X"FC",X"F4",X"FF",X"FF",X"7F",X"3F",X"BF",X"FF",X"F7",X"F3",
		X"C4",X"C4",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"99",X"C9",X"39",X"FC",X"F4",X"F4",X"F0",X"F0",
		X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F9",X"BC",X"B4",X"B0",X"B0",X"B0",X"B0",X"F0",
		X"F0",X"70",X"30",X"90",X"90",X"C0",X"40",X"40",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"3C",
		X"C0",X"C0",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"34",X"CC",X"C9",X"C7",X"CF",X"3F",X"FB",X"F6",X"69",X"C3",X"9F",X"9F",X"9F",X"33",X"BC",X"B8",
		X"30",X"C0",X"C0",X"04",X"CC",X"C9",X"39",X"F7",X"30",X"C4",X"CC",X"09",X"C3",X"C7",X"3F",X"FF",
		X"F6",X"F6",X"F6",X"F6",X"36",X"93",X"CB",X"0F",X"F0",X"FC",X"F9",X"F9",X"F7",X"7F",X"37",X"93",
		X"F7",X"FF",X"FF",X"FF",X"3F",X"C7",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"3F",X"CF",X"4F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"0C",X"CB",X"4F",X"0F",X"0F",X"0F",X"0F",X"43",X"4C",
		X"07",X"03",X"03",X"89",X"89",X"CC",X"C9",X"67",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"0C",X"8B",
		X"08",X"C0",X"C4",X"34",X"FC",X"F9",X"F9",X"F9",X"49",X"C9",X"93",X"37",X"F7",X"FF",X"FF",X"F3",
		X"67",X"3F",X"3B",X"BB",X"FB",X"FB",X"F6",X"F6",X"86",X"C6",X"CC",X"38",X"F8",X"F8",X"F8",X"F4",
		X"FC",X"FC",X"F3",X"33",X"C3",X"0B",X"CB",X"3F",X"FC",X"FC",X"F8",X"38",X"CC",X"CC",X"9C",X"36",
		X"F6",X"FC",X"FC",X"38",X"C8",X"08",X"08",X"C0",X"F4",X"F4",X"F4",X"3C",X"CC",X"09",X"49",X"C9",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"C3",X"F3",X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"C3",
		X"34",X"74",X"F4",X"F4",X"F4",X"FC",X"F9",X"3C",X"39",X"F7",X"F7",X"F7",X"F7",X"F7",X"37",X"33",
		X"CC",X"00",X"0C",X"CC",X"33",X"3F",X"FF",X"FF",X"0C",X"00",X"08",X"CC",X"C3",X"3F",X"FF",X"FF",
		X"6C",X"6C",X"69",X"39",X"B9",X"F9",X"F9",X"F9",X"CC",X"88",X"CC",X"C3",X"3B",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"33",X"CC",X"0C",X"0C",X"03",X"FF",X"FF",X"FF",X"33",X"9C",X"CC",X"0C",X"03",
		X"F9",X"F9",X"39",X"C9",X"C9",X"0C",X"0C",X"09",X"FF",X"FF",X"7F",X"33",X"CC",X"0C",X"0C",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"06",
		X"C9",X"C9",X"69",X"69",X"39",X"C9",X"C9",X"09",X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",X"8F",X"0F",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"F6",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"79",X"39",X"39",X"99",X"C9",X"49",X"C9",X"9C",X"FF",X"FF",X"FF",X"7F",X"7F",X"77",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F6",X"B6",X"B6",X"36",
		X"9C",X"34",X"74",X"F4",X"F4",X"F4",X"F4",X"F0",X"F7",X"F7",X"F7",X"F3",X"F3",X"F9",X"F9",X"F9",
		X"F7",X"B7",X"37",X"67",X"C3",X"C9",X"C9",X"99",X"66",X"66",X"C3",X"9B",X"9F",X"7F",X"7F",X"FF",
		X"F8",X"F8",X"F8",X"F8",X"7C",X"36",X"66",X"66",X"F9",X"F9",X"FC",X"B4",X"34",X"64",X"C0",X"88",
		X"99",X"74",X"74",X"F4",X"F0",X"F8",X"F8",X"F8",X"F7",X"F7",X"F7",X"F3",X"F9",X"F9",X"F9",X"F4",
		X"66",X"6B",X"8B",X"8B",X"CF",X"CF",X"C7",X"67",X"48",X"48",X"CC",X"9C",X"96",X"96",X"76",X"7B",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",X"30",X"60",
		X"60",X"30",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"BF",X"BF",X"BF",X"B3",X"33",X"3C",X"66",X"6B",X"6B",X"CB",X"CF",X"CF",X"C7",X"83",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",
		X"68",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"8C",X"84",X"80",X"80",X"80",X"80",X"80",X"00",
		X"FF",X"FB",X"F6",X"F6",X"FC",X"FC",X"F6",X"73",X"F6",X"FC",X"F8",X"F0",X"F0",X"F0",X"B8",X"B8",
		X"C0",X"C8",X"0C",X"86",X"C3",X"CB",X"CF",X"CF",X"00",X"00",X"00",X"08",X"0C",X"06",X"0B",X"0F",
		X"3B",X"9F",X"CF",X"4F",X"CF",X"9F",X"9F",X"3F",X"BC",X"36",X"CB",X"CB",X"3F",X"3F",X"BF",X"BF",
		X"CF",X"CF",X"CF",X"CF",X"C7",X"C3",X"CC",X"64",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"89",
		X"77",X"73",X"79",X"FC",X"F4",X"F0",X"F0",X"F0",X"BF",X"BF",X"B7",X"B3",X"B9",X"BC",X"B4",X"F0",
		X"60",X"60",X"60",X"60",X"60",X"60",X"30",X"30",X"8C",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"B0",X"B0",X"B0",X"B0",X"BC",X"FC",X"F3",X"FF",X"C0",X"C0",X"C0",X"60",X"68",X"6C",X"66",X"3B",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"34",X"3C",X"C9",X"F0",X"F0",X"F0",X"F0",X"F4",X"FC",X"73",X"97",
		X"3F",X"CF",X"3F",X"7F",X"77",X"77",X"FF",X"FB",X"6F",X"CF",X"3F",X"BF",X"FF",X"FF",X"F3",X"F6",
		X"07",X"0F",X"0F",X"CF",X"C3",X"33",X"FC",X"FC",X"CF",X"4F",X"4F",X"CF",X"C3",X"33",X"39",X"F7",
		X"FF",X"F0",X"F0",X"F5",X"F5",X"3A",X"C0",X"4F",X"F0",X"FA",X"F5",X"F5",X"F5",X"75",X"3A",X"C0",
		X"F0",X"F5",X"FA",X"FA",X"3A",X"CA",X"05",X"00",X"FF",X"F0",X"F0",X"FA",X"3A",X"C5",X"40",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",
		X"9F",X"4F",X"4F",X"0F",X"0F",X"4F",X"40",X"90",X"70",X"70",X"30",X"90",X"9F",X"9F",X"30",X"70",
		X"0A",X"8A",X"CF",X"6F",X"30",X"F0",X"FF",X"FF",X"0F",X"0F",X"8F",X"CA",X"C0",X"60",X"BF",X"BF",
		X"0F",X"CF",X"CF",X"30",X"F0",X"30",X"95",X"6F",X"05",X"C5",X"C5",X"30",X"F0",X"F0",X"7F",X"3F",
		X"FF",X"70",X"70",X"7F",X"3F",X"3F",X"9A",X"9A",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"B0",X"F0",X"F5",X"FF",X"FF",X"FF",X"FF",X"9F",X"90",X"60",X"6F",X"6F",X"6F",X"65",X"65",
		X"9F",X"90",X"90",X"9F",X"9F",X"90",X"90",X"9F",X"FF",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"30",X"30",X"3F",X"6F",X"60",X"60",X"6F",
		X"70",X"70",X"70",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F0",X"F0",X"FF",
		X"FF",X"BF",X"BF",X"3F",X"65",X"60",X"C0",X"95",X"60",X"C0",X"C0",X"9F",X"9F",X"70",X"70",X"FF",
		X"F0",X"FF",X"FF",X"F0",X"B0",X"B0",X"30",X"60",X"FF",X"BF",X"3A",X"60",X"60",X"CF",X"8F",X"8F",
		X"9F",X"7F",X"75",X"F0",X"F0",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"60",X"C0",X"CF",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"0A",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F5",X"FF",X"FF",X"BF",X"BF",X"BF",X"F0",X"B0",X"BF",X"3F",X"60",X"60",X"C0",X"C0",
		X"0A",X"0F",X"00",X"00",X"05",X"0F",X"0A",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"00",X"00",X"00",
		X"60",X"65",X"6F",X"CA",X"CA",X"C5",X"80",X"80",X"8F",X"8F",X"80",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"00",
		X"80",X"80",X"0F",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"0A",X"0F",X"0F",X"05",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",
		X"05",X"0F",X"0A",X"0A",X"8A",X"8F",X"85",X"80",X"0A",X"0F",X"0F",X"05",X"05",X"00",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"00",
		X"8A",X"CF",X"CF",X"CA",X"6A",X"6A",X"60",X"B0",X"00",X"05",X"0F",X"8F",X"85",X"80",X"C0",X"C0",
		X"0A",X"8F",X"8F",X"CA",X"CA",X"6A",X"6A",X"60",X"00",X"0A",X"0A",X"00",X"00",X"80",X"80",X"C0",
		X"B0",X"FF",X"FF",X"FF",X"F5",X"F0",X"F0",X"70",X"C0",X"6F",X"6F",X"B0",X"BA",X"FF",X"F5",X"F0",
		X"BF",X"BF",X"F0",X"F0",X"F0",X"F5",X"F5",X"F0",X"C0",X"CA",X"6A",X"6A",X"BA",X"BA",X"F0",X"F0",
		X"90",X"9A",X"9A",X"3A",X"3A",X"FF",X"FF",X"F0",X"F5",X"FF",X"7A",X"7A",X"FA",X"FA",X"FA",X"F0",
		X"FF",X"FF",X"F0",X"30",X"90",X"4F",X"0F",X"00",X"F0",X"FA",X"FA",X"FA",X"7A",X"3A",X"90",X"C0",
		X"F0",X"FA",X"FA",X"3A",X"CF",X"C5",X"60",X"30",X"F0",X"F5",X"F5",X"35",X"C5",X"0F",X"8F",X"C0",
		X"80",X"80",X"C0",X"6F",X"6F",X"B0",X"B0",X"B0",X"40",X"00",X"00",X"8A",X"CA",X"C0",X"C0",X"C0",
		X"BF",X"FF",X"FA",X"FA",X"FA",X"FF",X"FF",X"F0",X"C0",X"6A",X"BF",X"F5",X"F0",X"F0",X"F0",X"F0",
		X"BF",X"3F",X"6A",X"6A",X"C0",X"80",X"0F",X"00",X"C0",X"CA",X"8A",X"8A",X"0A",X"0A",X"00",X"00",
		X"F0",X"F5",X"FA",X"FA",X"FA",X"BF",X"35",X"60",X"F0",X"FA",X"F5",X"B5",X"3F",X"6F",X"CA",X"80",
		X"0A",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"00",
		X"C5",X"8F",X"0A",X"0A",X"0A",X"0F",X"05",X"00",X"0F",X"0F",X"05",X"05",X"05",X"0F",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"B0",X"B0",X"F0",X"F0",X"F0",X"F0",X"80",X"85",X"C5",X"C5",X"65",X"65",X"B5",X"B0",
		X"60",X"65",X"6A",X"B0",X"BA",X"B5",X"B0",X"30",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"80",
		X"F0",X"F5",X"F0",X"F0",X"F0",X"F5",X"F0",X"F0",X"F0",X"F0",X"FA",X"F5",X"FA",X"F0",X"F0",X"F0",
		X"65",X"65",X"C5",X"C5",X"85",X"85",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"60",X"FA",X"FA",X"BA",X"BA",X"6A",X"6A",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"60",X"CF",X"8F",X"85",X"00",X"00",X"00",X"00",X"80",X"00",X"0A",X"0F",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"80",X"85",X"CF",X"CA",X"CF",X"65",X"30",X"00",X"00",X"0F",X"05",X"00",X"80",X"8A",X"C0",
		X"80",X"80",X"C0",X"C0",X"60",X"60",X"30",X"B0",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",
		X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"C0",X"60",X"30",X"B0",X"B0",X"F0",X"F0",X"F0",
		X"B3",X"B3",X"6E",X"6E",X"62",X"6F",X"CF",X"C0",X"C2",X"8A",X"88",X"80",X"88",X"0A",X"02",X"00",
		X"30",X"91",X"93",X"92",X"93",X"71",X"70",X"70",X"F3",X"F3",X"FC",X"FC",X"F8",X"BF",X"B7",X"B0",
		X"83",X"8F",X"0C",X"00",X"0C",X"0F",X"03",X"00",X"00",X"02",X"0A",X"0A",X"0A",X"0A",X"02",X"00",
		X"71",X"33",X"C2",X"02",X"0E",X"0F",X"03",X"00",X"32",X"63",X"C5",X"05",X"0D",X"0F",X"03",X"00",
		X"01",X"05",X"00",X"00",X"05",X"0F",X"02",X"00",X"00",X"02",X"0A",X"0A",X"0A",X"00",X"00",X"00",
		X"01",X"03",X"02",X"02",X"03",X"01",X"00",X"00",X"00",X"04",X"0C",X"08",X"0C",X"07",X"03",X"00",
		X"02",X"03",X"0D",X"0C",X"00",X"0F",X"0F",X"00",X"00",X"08",X"0A",X"02",X"0A",X"0A",X"02",X"00",
		X"00",X"01",X"0F",X"0E",X"02",X"03",X"03",X"00",X"03",X"03",X"0C",X"0C",X"04",X"07",X"03",X"00",
		X"00",X"08",X"08",X"08",X"0F",X"0F",X"00",X"00",X"02",X"02",X"0A",X"0A",X"0A",X"02",X"00",X"00",
		X"02",X"02",X"02",X"02",X"03",X"03",X"00",X"00",X"00",X"05",X"09",X"09",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"02",X"00",X"00",
		X"02",X"06",X"0A",X"0E",X"07",X"03",X"00",X"00",X"00",X"01",X"05",X"0D",X"0F",X"07",X"00",X"00",
		X"03",X"07",X"04",X"04",X"0D",X"07",X"02",X"00",X"02",X"0A",X"0E",X"06",X"06",X"08",X"00",X"00",
		X"02",X"06",X"02",X"06",X"07",X"01",X"00",X"00",X"01",X"01",X"0D",X"04",X"0C",X"0F",X"03",X"00",
		X"C3",X"CF",X"CC",X"C0",X"8C",X"0F",X"33",X"30",X"C2",X"CA",X"C8",X"00",X"18",X"3A",X"22",X"30",
		X"03",X"C3",X"C0",X"C0",X"CC",X"CF",X"03",X"30",X"43",X"C3",X"C5",X"C5",X"CD",X"CF",X"03",X"30",
		X"30",X"00",X"C3",X"CF",X"CC",X"C0",X"C0",X"C0",X"32",X"02",X"CA",X"CA",X"CA",X"CA",X"C0",X"C0",
		X"82",X"C2",X"C3",X"C7",X"C6",X"C2",X"C0",X"00",X"00",X"C0",X"C3",X"C7",X"C4",X"C4",X"C0",X"C0",
		X"03",X"3F",X"0C",X"00",X"00",X"01",X"01",X"30",X"00",X"3A",X"3E",X"06",X"06",X"0A",X"00",X"30",
		X"23",X"37",X"04",X"00",X"00",X"00",X"00",X"30",X"03",X"37",X"04",X"00",X"00",X"00",X"00",X"30",
		X"30",X"01",X"C7",X"CB",X"CE",X"CF",X"C3",X"00",X"32",X"0A",X"C2",X"C0",X"C8",X"CA",X"D2",X"D0",
		X"02",X"C3",X"C1",X"C0",X"CC",X"CF",X"C3",X"00",X"10",X"88",X"C6",X"C3",X"CD",X"CF",X"C3",X"00",
		X"20",X"30",X"00",X"3C",X"3F",X"03",X"C0",X"C0",X"02",X"32",X"0A",X"3A",X"3A",X"0A",X"F0",X"F0",
		X"30",X"00",X"00",X"3C",X"0F",X"CB",X"C0",X"C0",X"30",X"30",X"00",X"3C",X"1F",X"83",X"C0",X"C0",
		X"CF",X"CF",X"C0",X"0E",X"30",X"3F",X"3F",X"00",X"FA",X"FA",X"F0",X"08",X"30",X"3A",X"3A",X"00",
		X"C3",X"C3",X"C1",X"00",X"31",X"33",X"33",X"00",X"C7",X"CF",X"CB",X"07",X"3B",X"3F",X"37",X"08",
		X"C3",X"CF",X"CF",X"C2",X"CC",X"CF",X"03",X"30",X"A2",X"FA",X"F8",X"F0",X"F8",X"FA",X"02",X"20",
		X"C3",X"C3",X"C0",X"C0",X"C1",X"C3",X"03",X"30",X"C3",X"C7",X"CD",X"CB",X"CF",X"C7",X"0B",X"30",
		X"33",X"3F",X"3C",X"00",X"CC",X"CF",X"C3",X"C0",X"30",X"32",X"3A",X"0A",X"FA",X"F2",X"F0",X"D0",
		X"31",X"33",X"32",X"02",X"C2",X"C3",X"C1",X"C0",X"33",X"37",X"3C",X"08",X"CC",X"C7",X"C3",X"C0",
		X"C0",X"CA",X"CE",X"06",X"3E",X"0F",X"03",X"00",X"D0",X"D0",X"D0",X"00",X"3C",X"0E",X"02",X"00",
		X"C1",X"C3",X"C2",X"02",X"32",X"03",X"03",X"00",X"C3",X"C7",X"CC",X"08",X"3C",X"07",X"0B",X"00",
		X"02",X"03",X"3F",X"0E",X"C4",X"CF",X"CB",X"C0",X"02",X"30",X"2E",X"0E",X"C2",X"C2",X"C0",X"C0",
		X"21",X"23",X"32",X"02",X"C2",X"C3",X"C1",X"C0",X"03",X"0B",X"34",X"0C",X"C8",X"CF",X"C7",X"C0",
		X"C0",X"81",X"83",X"C3",X"CE",X"CF",X"C3",X"C0",X"C2",X"02",X"02",X"00",X"C8",X"CA",X"C2",X"C0",
		X"C1",X"C3",X"C2",X"C2",X"C2",X"C3",X"43",X"40",X"C3",X"C7",X"C9",X"CC",X"CC",X"C7",X"CB",X"C0",
		X"C3",X"87",X"0C",X"08",X"08",X"81",X"81",X"C0",X"C0",X"02",X"3A",X"3A",X"3A",X"1A",X"10",X"00",
		X"40",X"21",X"23",X"22",X"22",X"13",X"11",X"00",X"C0",X"C1",X"C9",X"C9",X"4D",X"47",X"42",X"20",
		X"30",X"30",X"13",X"2F",X"2C",X"00",X"50",X"50",X"30",X"20",X"0A",X"5A",X"50",X"F0",X"F0",X"A0",
		X"C2",X"82",X"03",X"3F",X"2E",X"02",X"00",X"30",X"00",X"18",X"2B",X"0F",X"1C",X"18",X"30",X"20",
		X"F3",X"F3",X"FC",X"AC",X"A0",X"AF",X"AF",X"A0",X"A0",X"0A",X"0A",X"52",X"FA",X"FA",X"F0",X"F0",
		X"33",X"03",X"C0",X"C0",X"C0",X"C3",X"C3",X"C0",X"23",X"03",X"0C",X"5C",X"50",X"5F",X"5F",X"50",
		X"A0",X"AA",X"AF",X"A7",X"FF",X"FE",X"00",X"10",X"00",X"00",X"50",X"AA",X"A8",X"10",X"10",X"20",
		X"03",X"33",X"30",X"10",X"10",X"03",X"03",X"20",X"53",X"5F",X"51",X"50",X"21",X"2F",X"2F",X"30",
		X"3F",X"1F",X"A3",X"FE",X"F3",X"FF",X"FF",X"F0",X"30",X"3A",X"08",X"F0",X"F8",X"FA",X"F0",X"F0",
		X"33",X"03",X"F0",X"F0",X"F0",X"F3",X"F3",X"F0",X"3F",X"0F",X"F1",X"F3",X"F1",X"FF",X"FF",X"F0",
		X"01",X"33",X"07",X"0E",X"3F",X"0B",X"F1",X"F0",X"02",X"3A",X"08",X"08",X"30",X"0A",X"0A",X"F0",
		X"03",X"33",X"01",X"30",X"31",X"03",X"F3",X"F0",X"00",X"3A",X"07",X"33",X"37",X"0E",X"FC",X"F0",
		X"F0",X"F0",X"FB",X"FF",X"08",X"30",X"00",X"20",X"F0",X"F0",X"F2",X"F2",X"0C",X"34",X"00",X"00",
		X"F3",X"F3",X"F0",X"00",X"03",X"33",X"30",X"30",X"F2",X"FB",X"F5",X"51",X"07",X"3E",X"28",X"30",
		X"10",X"00",X"A0",X"AA",X"FF",X"F7",X"F1",X"F0",X"22",X"3A",X"3A",X"1A",X"1A",X"0A",X"AA",X"A0",
		X"03",X"F3",X"F3",X"F2",X"F2",X"F2",X"F2",X"50",X"00",X"FA",X"FF",X"FF",X"F9",X"F8",X"F8",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"20",X"30",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"50",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F3",X"F0",X"03",X"33",X"00",X"00",X"03",X"F2",X"F2",X"F0",X"00",X"32",X"02",X"02",X"12",
		X"F0",X"F3",X"F0",X"01",X"33",X"02",X"02",X"03",X"F0",X"F3",X"F0",X"02",X"33",X"01",X"01",X"03",
		X"33",X"03",X"50",X"F0",X"F3",X"F0",X"F0",X"F0",X"30",X"02",X"F2",X"F2",X"F0",X"F0",X"F2",X"A2",
		X"01",X"33",X"02",X"F2",X"F1",X"D0",X"D0",X"D0",X"13",X"33",X"00",X"F0",X"F3",X"F0",X"F0",X"F0",
		X"03",X"00",X"A3",X"F3",X"F0",X"F0",X"F3",X"F0",X"A2",X"F0",X"50",X"52",X"F2",X"F2",X"F0",X"F0",
		X"03",X"00",X"31",X"03",X"C2",X"C2",X"C1",X"C0",X"53",X"50",X"03",X"03",X"80",X"D0",X"D3",X"D0",
		X"F0",X"F0",X"00",X"30",X"02",X"03",X"01",X"00",X"F0",X"F0",X"00",X"30",X"10",X"00",X"02",X"02",
		X"C0",X"00",X"30",X"30",X"00",X"21",X"33",X"32",X"C0",X"00",X"20",X"30",X"03",X"03",X"00",X"20",
		X"00",X"0F",X"0F",X"06",X"36",X"36",X"0F",X"0F",X"00",X"0A",X"00",X"32",X"36",X"02",X"00",X"CA",
		X"00",X"00",X"01",X"09",X"0C",X"09",X"01",X"10",X"00",X"05",X"02",X"06",X"0C",X"16",X"32",X"25",
		X"CF",X"CF",X"CF",X"CC",X"CC",X"CF",X"DF",X"DF",X"CF",X"CA",X"D0",X"DC",X"FC",X"F0",X"FA",X"FF",
		X"30",X"20",X"02",X"44",X"C4",X"C2",X"C0",X"C0",X"00",X"45",X"CD",X"CC",X"CC",X"CD",X"C5",X"C0",
		X"03",X"3C",X"3C",X"0C",X"FC",X"FC",X"FC",X"F3",X"02",X"33",X"39",X"09",X"F9",X"F9",X"F3",X"F2",
		X"01",X"33",X"06",X"F6",X"F6",X"F6",X"D3",X"D1",X"03",X"3C",X"3C",X"0C",X"FE",X"FF",X"FC",X"F3",
		X"FC",X"FC",X"56",X"06",X"3B",X"1B",X"0B",X"0F",X"F4",X"F4",X"F0",X"F8",X"08",X"28",X"3C",X"16",
		X"C7",X"C3",X"83",X"03",X"13",X"33",X"27",X"27",X"FB",X"FB",X"0F",X"0F",X"3F",X"0F",X"0F",X"0F",
		X"00",X"10",X"30",X"00",X"C0",X"C0",X"C0",X"CF",X"10",X"30",X"00",X"C0",X"C0",X"C0",X"C0",X"CF",
		X"0A",X"0A",X"3A",X"3A",X"0A",X"CA",X"CA",X"CF",X"00",X"00",X"30",X"20",X"40",X"C0",X"C0",X"CF",
		X"CF",X"C0",X"C0",X"C0",X"C0",X"00",X"30",X"30",X"CF",X"C0",X"C0",X"C0",X"C0",X"00",X"30",X"30",
		X"CF",X"CA",X"CA",X"CA",X"CA",X"0A",X"3A",X"0A",X"CF",X"C0",X"C0",X"C0",X"C0",X"00",X"30",X"30",
		X"00",X"00",X"30",X"30",X"00",X"F0",X"F0",X"FF",X"05",X"35",X"35",X"05",X"F5",X"F5",X"05",X"AF",
		X"00",X"00",X"00",X"30",X"30",X"00",X"C0",X"DF",X"00",X"00",X"00",X"30",X"30",X"00",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",
		X"DF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"30",X"00",X"F0",X"F0",X"F0",X"F0",X"10",X"00",X"30",X"00",X"00",X"F0",X"F0",X"F0",
		X"00",X"20",X"3F",X"0F",X"F0",X"FF",X"FF",X"F0",X"00",X"0A",X"3A",X"00",X"FA",X"FA",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"A0",X"A0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"10",X"00",X"A0",X"F0",
		X"F0",X"FF",X"FF",X"F0",X"FF",X"5F",X"00",X"00",X"F0",X"F0",X"FA",X"FA",X"F0",X"FA",X"FA",X"F0",
		X"F0",X"F0",X"F0",X"D0",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"D0",X"D0",X"80",
		X"20",X"40",X"C0",X"C0",X"CF",X"CF",X"C0",X"C0",X"D0",X"D0",X"C0",X"C0",X"C0",X"CA",X"C0",X"C0",
		X"CF",X"80",X"00",X"10",X"30",X"20",X"00",X"00",X"0A",X"10",X"30",X"20",X"00",X"00",X"00",X"00",
		X"CF",X"C0",X"C0",X"C0",X"8F",X"0F",X"30",X"00",X"CF",X"C0",X"C0",X"80",X"00",X"3A",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"60",X"C0",X"80",X"C0",X"90",X"30",X"70",X"C0",X"80",X"40",X"C0",X"90",X"34",X"74",X"FC",
		X"90",X"30",X"70",X"F0",X"B0",X"B0",X"60",X"30",X"F0",X"F0",X"B0",X"60",X"C0",X"C0",X"90",X"30",
		X"F0",X"70",X"74",X"94",X"94",X"C4",X"44",X"40",X"BC",X"F9",X"F9",X"F9",X"F9",X"79",X"79",X"9C",
		X"80",X"80",X"80",X"C0",X"60",X"60",X"B0",X"B0",X"90",X"C0",X"40",X"40",X"00",X"80",X"80",X"C0",
		X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"9C",X"C4",X"44",X"44",X"00",X"04",X"04",X"04",
		X"30",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"04",X"04",X"0C",X"C9",X"0C",X"09",X"09",X"09",X"07",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"69",X"B9",X"F7",X"F7",X"F7",X"F7",X"F7",X"FF",X"CF",X"6B",X"BB",X"FB",X"FB",X"FB",X"F6",X"F6",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"B0",X"F4",X"F4",X"F4",X"F4",X"F4",X"FC",X"F9",
		X"FF",X"7F",X"9F",X"CB",X"0B",X"0B",X"0B",X"0B",X"F6",X"F6",X"36",X"CC",X"C8",X"08",X"08",X"08",
		X"90",X"C0",X"00",X"04",X"04",X"04",X"04",X"04",X"79",X"99",X"C9",X"09",X"09",X"07",X"07",X"07",
		X"0B",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"08",X"08",X"08",X"00",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"0C",X"0C",X"8C",X"CC",X"CC",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"87",
		X"06",X"06",X"06",X"46",X"46",X"C6",X"96",X"36",X"04",X"44",X"C4",X"94",X"94",X"34",X"74",X"F4",
		X"69",X"B9",X"B9",X"B9",X"B9",X"69",X"C9",X"89",X"8F",X"CF",X"CF",X"CF",X"CF",X"8F",X"4F",X"CF",
		X"76",X"F6",X"F6",X"F6",X"F6",X"B6",X"36",X"66",X"F4",X"F4",X"F4",X"B4",X"34",X"64",X"C4",X"C4",
		X"49",X"C9",X"99",X"39",X"79",X"F9",X"F9",X"FC",X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"B7",
		X"C6",X"C6",X"36",X"F6",X"FB",X"FB",X"FB",X"FB",X"C4",X"C0",X"38",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"6C",X"3C",X"FC",X"F4",X"F4",X"F4",X"F4",X"F4",X"C7",X"67",X"37",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"FB",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"F7",X"F8",X"F8",X"FC",X"F6",X"B6",X"36",X"36",X"36",
		X"F4",X"74",X"74",X"90",X"90",X"40",X"40",X"00",X"F7",X"F9",X"F9",X"F9",X"F9",X"79",X"79",X"9C",
		X"77",X"77",X"97",X"99",X"49",X"49",X"09",X"0C",X"B6",X"BB",X"FB",X"7B",X"3B",X"CF",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"44",X"44",X"04",X"04",X"00",X"00",X"00",
		X"0C",X"04",X"C4",X"34",X"F4",X"F0",X"F0",X"F0",X"07",X"07",X"C7",X"C9",X"39",X"F9",X"FC",X"FC",
		X"80",X"C0",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"C0",X"60",X"B0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"30",X"C0",X"40",X"00",X"F4",X"F4",X"F4",X"F4",X"74",X"94",X"CC",X"0C",
		X"F0",X"F0",X"F0",X"30",X"C0",X"40",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"90",X"C0",X"00",X"00",
		X"34",X"64",X"CC",X"0C",X"09",X"03",X"C7",X"67",X"39",X"99",X"C7",X"07",X"0F",X"0F",X"0F",X"8F",
		X"F0",X"F0",X"30",X"60",X"C0",X"80",X"40",X"C4",X"F0",X"30",X"60",X"C0",X"04",X"04",X"CC",X"39",
		X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"6F",X"3F",X"FF",X"FB",X"FB",X"FF",X"FF",
		X"34",X"74",X"FC",X"FC",X"FC",X"FC",X"3C",X"34",X"F9",X"F3",X"F7",X"F7",X"F7",X"F7",X"77",X"37",
		X"7F",X"3F",X"37",X"B7",X"F3",X"F9",X"FC",X"F4",X"FF",X"FF",X"7F",X"3F",X"BF",X"FF",X"F7",X"F3",
		X"C4",X"C4",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"99",X"C9",X"39",X"FC",X"F4",X"F4",X"F0",X"F0",
		X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F9",X"BC",X"B4",X"B0",X"B0",X"B0",X"B0",X"F0",
		X"F0",X"70",X"30",X"90",X"90",X"C0",X"40",X"40",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"3C",
		X"C0",X"C0",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"34",X"CC",X"C9",X"C7",X"CF",X"3F",X"FB",X"F6",X"69",X"C3",X"9F",X"9F",X"9F",X"33",X"BC",X"B8",
		X"30",X"C0",X"C0",X"04",X"CC",X"C9",X"39",X"F7",X"30",X"C4",X"CC",X"09",X"C3",X"C7",X"3F",X"FF",
		X"F6",X"F6",X"F6",X"F6",X"36",X"93",X"CB",X"0F",X"F0",X"FC",X"F9",X"F9",X"F7",X"7F",X"37",X"93",
		X"F7",X"FF",X"FF",X"FF",X"3F",X"C7",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"3F",X"CF",X"4F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"0C",X"CB",X"4F",X"0F",X"0F",X"0F",X"0F",X"43",X"4C",
		X"07",X"03",X"03",X"89",X"89",X"CC",X"C9",X"67",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"0C",X"8B",
		X"08",X"C0",X"C4",X"34",X"FC",X"F9",X"F9",X"F9",X"49",X"C9",X"93",X"37",X"F7",X"FF",X"FF",X"F3",
		X"67",X"3F",X"3B",X"BB",X"FB",X"FB",X"F6",X"F6",X"86",X"C6",X"CC",X"38",X"F8",X"F8",X"F8",X"F4",
		X"FC",X"FC",X"F3",X"33",X"C3",X"0B",X"CB",X"3F",X"FC",X"FC",X"F8",X"38",X"CC",X"CC",X"9C",X"36",
		X"F6",X"FC",X"FC",X"38",X"C8",X"08",X"08",X"C0",X"F4",X"F4",X"F4",X"3C",X"CC",X"09",X"49",X"C9",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"C3",X"F3",X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"C3",
		X"34",X"74",X"F4",X"F4",X"F4",X"FC",X"F9",X"3C",X"39",X"F7",X"F7",X"F7",X"F7",X"F7",X"37",X"33",
		X"CC",X"00",X"0C",X"CC",X"33",X"3F",X"FF",X"FF",X"0C",X"00",X"08",X"CC",X"C3",X"3F",X"FF",X"FF",
		X"6C",X"6C",X"69",X"39",X"B9",X"F9",X"F9",X"F9",X"CC",X"88",X"CC",X"C3",X"3B",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"33",X"CC",X"0C",X"0C",X"03",X"FF",X"FF",X"FF",X"33",X"9C",X"CC",X"0C",X"03",
		X"F9",X"F9",X"39",X"C9",X"C9",X"0C",X"0C",X"09",X"FF",X"FF",X"7F",X"33",X"CC",X"0C",X"0C",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"06",
		X"C9",X"C9",X"69",X"69",X"39",X"C9",X"C9",X"09",X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",X"8F",X"0F",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"F6",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"79",X"39",X"39",X"99",X"C9",X"49",X"C9",X"9C",X"FF",X"FF",X"FF",X"7F",X"7F",X"77",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F6",X"B6",X"B6",X"36",
		X"9C",X"34",X"74",X"F4",X"F4",X"F4",X"F4",X"F0",X"F7",X"F7",X"F7",X"F3",X"F3",X"F9",X"F9",X"F9",
		X"F7",X"B7",X"37",X"67",X"C3",X"C9",X"C9",X"99",X"66",X"66",X"C3",X"9B",X"9F",X"7F",X"7F",X"FF",
		X"F8",X"F8",X"F8",X"F8",X"7C",X"36",X"66",X"66",X"F9",X"F9",X"FC",X"B4",X"34",X"64",X"C0",X"88",
		X"99",X"74",X"74",X"F4",X"F0",X"F8",X"F8",X"F8",X"F7",X"F7",X"F7",X"F3",X"F9",X"F9",X"F9",X"F4",
		X"66",X"6B",X"8B",X"8B",X"CF",X"CF",X"C7",X"67",X"48",X"48",X"CC",X"9C",X"96",X"96",X"76",X"7B",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",X"30",X"60",
		X"60",X"30",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"BF",X"BF",X"BF",X"B3",X"33",X"3C",X"66",X"6B",X"6B",X"CB",X"CF",X"CF",X"C7",X"83",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",
		X"68",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"8C",X"84",X"80",X"80",X"80",X"80",X"80",X"00",
		X"FF",X"FB",X"F6",X"F6",X"FC",X"FC",X"F6",X"73",X"F6",X"FC",X"F8",X"F0",X"F0",X"F0",X"B8",X"B8",
		X"C0",X"C8",X"0C",X"86",X"C3",X"CB",X"CF",X"CF",X"00",X"00",X"00",X"08",X"0C",X"06",X"0B",X"0F",
		X"3B",X"9F",X"CF",X"4F",X"CF",X"9F",X"9F",X"3F",X"BC",X"36",X"CB",X"CB",X"3F",X"3F",X"BF",X"BF",
		X"CF",X"CF",X"CF",X"CF",X"C7",X"C3",X"CC",X"64",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"89",
		X"77",X"73",X"79",X"FC",X"F4",X"F0",X"F0",X"F0",X"BF",X"BF",X"B7",X"B3",X"B9",X"BC",X"B4",X"F0",
		X"60",X"60",X"60",X"60",X"60",X"60",X"30",X"30",X"8C",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"B0",X"B0",X"B0",X"B0",X"BC",X"FC",X"F3",X"FF",X"C0",X"C0",X"C0",X"60",X"68",X"6C",X"66",X"3B",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"34",X"3C",X"C9",X"F0",X"F0",X"F0",X"F0",X"F4",X"FC",X"73",X"97",
		X"3F",X"CF",X"3F",X"7F",X"77",X"77",X"FF",X"FB",X"6F",X"CF",X"3F",X"BF",X"FF",X"FF",X"F3",X"F6",
		X"07",X"0F",X"0F",X"CF",X"C3",X"33",X"FC",X"FC",X"CF",X"4F",X"4F",X"CF",X"C3",X"33",X"39",X"F7",
		X"FF",X"F0",X"F0",X"F5",X"F5",X"3A",X"C0",X"4F",X"F0",X"FA",X"F5",X"F5",X"F5",X"75",X"3A",X"C0",
		X"F0",X"F5",X"FA",X"FA",X"3A",X"CA",X"05",X"00",X"FF",X"F0",X"F0",X"FA",X"3A",X"C5",X"40",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",
		X"9F",X"4F",X"4F",X"0F",X"0F",X"4F",X"40",X"90",X"70",X"70",X"30",X"90",X"9F",X"9F",X"30",X"70",
		X"0A",X"8A",X"CF",X"6F",X"30",X"F0",X"FF",X"FF",X"0F",X"0F",X"8F",X"CA",X"C0",X"60",X"BF",X"BF",
		X"0F",X"CF",X"CF",X"30",X"F0",X"30",X"95",X"6F",X"05",X"C5",X"C5",X"30",X"F0",X"F0",X"7F",X"3F",
		X"FF",X"70",X"70",X"7F",X"3F",X"3F",X"9A",X"9A",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"B0",X"F0",X"F5",X"FF",X"FF",X"FF",X"FF",X"9F",X"90",X"60",X"6F",X"6F",X"6F",X"65",X"65",
		X"9F",X"90",X"90",X"9F",X"9F",X"90",X"90",X"9F",X"FF",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"30",X"30",X"3F",X"6F",X"60",X"60",X"6F",
		X"70",X"70",X"70",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F0",X"F0",X"FF",
		X"FF",X"BF",X"BF",X"3F",X"65",X"60",X"C0",X"95",X"60",X"C0",X"C0",X"9F",X"9F",X"70",X"70",X"FF",
		X"F0",X"FF",X"FF",X"F0",X"B0",X"B0",X"30",X"60",X"FF",X"BF",X"3A",X"60",X"60",X"CF",X"8F",X"8F",
		X"9F",X"7F",X"75",X"F0",X"F0",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"60",X"C0",X"CF",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"0A",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F5",X"FF",X"FF",X"BF",X"BF",X"BF",X"F0",X"B0",X"BF",X"3F",X"60",X"60",X"C0",X"C0",
		X"0A",X"0F",X"00",X"00",X"05",X"0F",X"0A",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"00",X"00",X"00",
		X"60",X"65",X"6F",X"CA",X"CA",X"C5",X"80",X"80",X"8F",X"8F",X"80",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"00",
		X"80",X"80",X"0F",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"0A",X"0F",X"0F",X"05",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",
		X"05",X"0F",X"0A",X"0A",X"8A",X"8F",X"85",X"80",X"0A",X"0F",X"0F",X"05",X"05",X"00",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"00",
		X"8A",X"CF",X"CF",X"CA",X"6A",X"6A",X"60",X"B0",X"00",X"05",X"0F",X"8F",X"85",X"80",X"C0",X"C0",
		X"0A",X"8F",X"8F",X"CA",X"CA",X"6A",X"6A",X"60",X"00",X"0A",X"0A",X"00",X"00",X"80",X"80",X"C0",
		X"B0",X"FF",X"FF",X"FF",X"F5",X"F0",X"F0",X"70",X"C0",X"6F",X"6F",X"B0",X"BA",X"FF",X"F5",X"F0",
		X"BF",X"BF",X"F0",X"F0",X"F0",X"F5",X"F5",X"F0",X"C0",X"CA",X"6A",X"6A",X"BA",X"BA",X"F0",X"F0",
		X"90",X"9A",X"9A",X"3A",X"3A",X"FF",X"FF",X"F0",X"F5",X"FF",X"7A",X"7A",X"FA",X"FA",X"FA",X"F0",
		X"FF",X"FF",X"F0",X"30",X"90",X"4F",X"0F",X"00",X"F0",X"FA",X"FA",X"FA",X"7A",X"3A",X"90",X"C0",
		X"F0",X"FA",X"FA",X"3A",X"CF",X"C5",X"60",X"30",X"F0",X"F5",X"F5",X"35",X"C5",X"0F",X"8F",X"C0",
		X"80",X"80",X"C0",X"6F",X"6F",X"B0",X"B0",X"B0",X"40",X"00",X"00",X"8A",X"CA",X"C0",X"C0",X"C0",
		X"BF",X"FF",X"FA",X"FA",X"FA",X"FF",X"FF",X"F0",X"C0",X"6A",X"BF",X"F5",X"F0",X"F0",X"F0",X"F0",
		X"BF",X"3F",X"6A",X"6A",X"C0",X"80",X"0F",X"00",X"C0",X"CA",X"8A",X"8A",X"0A",X"0A",X"00",X"00",
		X"F0",X"F5",X"FA",X"FA",X"FA",X"BF",X"35",X"60",X"F0",X"FA",X"F5",X"B5",X"3F",X"6F",X"CA",X"80",
		X"0A",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"00",
		X"C5",X"8F",X"0A",X"0A",X"0A",X"0F",X"05",X"00",X"0F",X"0F",X"05",X"05",X"05",X"0F",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"B0",X"B0",X"F0",X"F0",X"F0",X"F0",X"80",X"85",X"C5",X"C5",X"65",X"65",X"B5",X"B0",
		X"60",X"65",X"6A",X"B0",X"BA",X"B5",X"B0",X"30",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"80",
		X"F0",X"F5",X"F0",X"F0",X"F0",X"F5",X"F0",X"F0",X"F0",X"F0",X"FA",X"F5",X"FA",X"F0",X"F0",X"F0",
		X"65",X"65",X"C5",X"C5",X"85",X"85",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"60",X"FA",X"FA",X"BA",X"BA",X"6A",X"6A",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"60",X"CF",X"8F",X"85",X"00",X"00",X"00",X"00",X"80",X"00",X"0A",X"0F",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"80",X"85",X"CF",X"CA",X"CF",X"65",X"30",X"00",X"00",X"0F",X"05",X"00",X"80",X"8A",X"C0",
		X"80",X"80",X"C0",X"C0",X"60",X"60",X"30",X"B0",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",
		X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"C0",X"60",X"30",X"B0",X"B0",X"F0",X"F0",X"F0",
		X"B3",X"B3",X"6E",X"6E",X"62",X"6F",X"CF",X"C0",X"C2",X"8A",X"88",X"80",X"88",X"0A",X"02",X"00",
		X"30",X"91",X"93",X"92",X"93",X"71",X"70",X"70",X"F3",X"F3",X"FC",X"FC",X"F8",X"BF",X"B7",X"B0",
		X"83",X"8F",X"0C",X"00",X"0C",X"0F",X"03",X"00",X"00",X"02",X"0A",X"0A",X"0A",X"0A",X"02",X"00",
		X"71",X"33",X"C2",X"02",X"0E",X"0F",X"03",X"00",X"32",X"63",X"C5",X"05",X"0D",X"0F",X"03",X"00",
		X"01",X"05",X"00",X"00",X"05",X"0F",X"02",X"00",X"00",X"02",X"0A",X"0A",X"0A",X"00",X"00",X"00",
		X"01",X"03",X"02",X"02",X"03",X"01",X"00",X"00",X"00",X"04",X"0C",X"08",X"0C",X"07",X"03",X"00",
		X"02",X"03",X"0D",X"0C",X"00",X"0F",X"0F",X"00",X"00",X"08",X"0A",X"02",X"0A",X"0A",X"02",X"00",
		X"00",X"01",X"0F",X"0E",X"02",X"03",X"03",X"00",X"03",X"03",X"0C",X"0C",X"04",X"07",X"03",X"00",
		X"00",X"08",X"08",X"08",X"0F",X"0F",X"00",X"00",X"02",X"02",X"0A",X"0A",X"0A",X"02",X"00",X"00",
		X"02",X"02",X"02",X"02",X"03",X"03",X"00",X"00",X"00",X"05",X"09",X"09",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"02",X"00",X"00",
		X"02",X"06",X"0A",X"0E",X"07",X"03",X"00",X"00",X"00",X"01",X"05",X"0D",X"0F",X"07",X"00",X"00",
		X"03",X"07",X"04",X"04",X"0D",X"07",X"02",X"00",X"02",X"0A",X"0E",X"06",X"06",X"08",X"00",X"00",
		X"02",X"06",X"02",X"06",X"07",X"01",X"00",X"00",X"01",X"01",X"0D",X"04",X"0C",X"0F",X"03",X"00",
		X"C3",X"CF",X"CC",X"C0",X"8C",X"0F",X"33",X"30",X"C2",X"CA",X"C8",X"00",X"18",X"3A",X"22",X"30",
		X"03",X"C3",X"C0",X"C0",X"CC",X"CF",X"03",X"30",X"43",X"C3",X"C5",X"C5",X"CD",X"CF",X"03",X"30",
		X"30",X"00",X"C3",X"CF",X"CC",X"C0",X"C0",X"C0",X"32",X"02",X"CA",X"CA",X"CA",X"CA",X"C0",X"C0",
		X"82",X"C2",X"C3",X"C7",X"C6",X"C2",X"C0",X"00",X"00",X"C0",X"C3",X"C7",X"C4",X"C4",X"C0",X"C0",
		X"03",X"3F",X"0C",X"00",X"00",X"01",X"01",X"30",X"00",X"3A",X"3E",X"06",X"06",X"0A",X"00",X"30",
		X"23",X"37",X"04",X"00",X"00",X"00",X"00",X"30",X"03",X"37",X"04",X"00",X"00",X"00",X"00",X"30",
		X"30",X"01",X"C7",X"CB",X"CE",X"CF",X"C3",X"00",X"32",X"0A",X"C2",X"C0",X"C8",X"CA",X"D2",X"D0",
		X"02",X"C3",X"C1",X"C0",X"CC",X"CF",X"C3",X"00",X"10",X"88",X"C6",X"C3",X"CD",X"CF",X"C3",X"00",
		X"20",X"30",X"00",X"3C",X"3F",X"03",X"C0",X"C0",X"02",X"32",X"0A",X"3A",X"3A",X"0A",X"F0",X"F0",
		X"30",X"00",X"00",X"3C",X"0F",X"CB",X"C0",X"C0",X"30",X"30",X"00",X"3C",X"1F",X"83",X"C0",X"C0",
		X"CF",X"CF",X"C0",X"0E",X"30",X"3F",X"3F",X"00",X"FA",X"FA",X"F0",X"08",X"30",X"3A",X"3A",X"00",
		X"C3",X"C3",X"C1",X"00",X"31",X"33",X"33",X"00",X"C7",X"CF",X"CB",X"07",X"3B",X"3F",X"37",X"08",
		X"C3",X"CF",X"CF",X"C2",X"CC",X"CF",X"03",X"30",X"A2",X"FA",X"F8",X"F0",X"F8",X"FA",X"02",X"20",
		X"C3",X"C3",X"C0",X"C0",X"C1",X"C3",X"03",X"30",X"C3",X"C7",X"CD",X"CB",X"CF",X"C7",X"0B",X"30",
		X"33",X"3F",X"3C",X"00",X"CC",X"CF",X"C3",X"C0",X"30",X"32",X"3A",X"0A",X"FA",X"F2",X"F0",X"D0",
		X"31",X"33",X"32",X"02",X"C2",X"C3",X"C1",X"C0",X"33",X"37",X"3C",X"08",X"CC",X"C7",X"C3",X"C0",
		X"C0",X"CA",X"CE",X"06",X"3E",X"0F",X"03",X"00",X"D0",X"D0",X"D0",X"00",X"3C",X"0E",X"02",X"00",
		X"C1",X"C3",X"C2",X"02",X"32",X"03",X"03",X"00",X"C3",X"C7",X"CC",X"08",X"3C",X"07",X"0B",X"00",
		X"02",X"03",X"3F",X"0E",X"C4",X"CF",X"CB",X"C0",X"02",X"30",X"2E",X"0E",X"C2",X"C2",X"C0",X"C0",
		X"21",X"23",X"32",X"02",X"C2",X"C3",X"C1",X"C0",X"03",X"0B",X"34",X"0C",X"C8",X"CF",X"C7",X"C0",
		X"C0",X"81",X"83",X"C3",X"CE",X"CF",X"C3",X"C0",X"C2",X"02",X"02",X"00",X"C8",X"CA",X"C2",X"C0",
		X"C1",X"C3",X"C2",X"C2",X"C2",X"C3",X"43",X"40",X"C3",X"C7",X"C9",X"CC",X"CC",X"C7",X"CB",X"C0",
		X"C3",X"87",X"0C",X"08",X"08",X"81",X"81",X"C0",X"C0",X"02",X"3A",X"3A",X"3A",X"1A",X"10",X"00",
		X"40",X"21",X"23",X"22",X"22",X"13",X"11",X"00",X"C0",X"C1",X"C9",X"C9",X"4D",X"47",X"42",X"20",
		X"30",X"30",X"13",X"2F",X"2C",X"00",X"50",X"50",X"30",X"20",X"0A",X"5A",X"50",X"F0",X"F0",X"A0",
		X"C2",X"82",X"03",X"3F",X"2E",X"02",X"00",X"30",X"00",X"18",X"2B",X"0F",X"1C",X"18",X"30",X"20",
		X"F3",X"F3",X"FC",X"AC",X"A0",X"AF",X"AF",X"A0",X"A0",X"0A",X"0A",X"52",X"FA",X"FA",X"F0",X"F0",
		X"33",X"03",X"C0",X"C0",X"C0",X"C3",X"C3",X"C0",X"23",X"03",X"0C",X"5C",X"50",X"5F",X"5F",X"50",
		X"A0",X"AA",X"AF",X"A7",X"FF",X"FE",X"00",X"10",X"00",X"00",X"50",X"AA",X"A8",X"10",X"10",X"20",
		X"03",X"33",X"30",X"10",X"10",X"03",X"03",X"20",X"53",X"5F",X"51",X"50",X"21",X"2F",X"2F",X"30",
		X"3F",X"1F",X"A3",X"FE",X"F3",X"FF",X"FF",X"F0",X"30",X"3A",X"08",X"F0",X"F8",X"FA",X"F0",X"F0",
		X"33",X"03",X"F0",X"F0",X"F0",X"F3",X"F3",X"F0",X"3F",X"0F",X"F1",X"F3",X"F1",X"FF",X"FF",X"F0",
		X"01",X"33",X"07",X"0E",X"3F",X"0B",X"F1",X"F0",X"02",X"3A",X"08",X"08",X"30",X"0A",X"0A",X"F0",
		X"03",X"33",X"01",X"30",X"31",X"03",X"F3",X"F0",X"00",X"3A",X"07",X"33",X"37",X"0E",X"FC",X"F0",
		X"F0",X"F0",X"FB",X"FF",X"08",X"30",X"00",X"20",X"F0",X"F0",X"F2",X"F2",X"0C",X"34",X"00",X"00",
		X"F3",X"F3",X"F0",X"00",X"03",X"33",X"30",X"30",X"F2",X"FB",X"F5",X"51",X"07",X"3E",X"28",X"30",
		X"10",X"00",X"A0",X"AA",X"FF",X"F7",X"F1",X"F0",X"22",X"3A",X"3A",X"1A",X"1A",X"0A",X"AA",X"A0",
		X"03",X"F3",X"F3",X"F2",X"F2",X"F2",X"F2",X"50",X"00",X"FA",X"FF",X"FF",X"F9",X"F8",X"F8",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"20",X"30",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"50",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F3",X"F0",X"03",X"33",X"00",X"00",X"03",X"F2",X"F2",X"F0",X"00",X"32",X"02",X"02",X"12",
		X"F0",X"F3",X"F0",X"01",X"33",X"02",X"02",X"03",X"F0",X"F3",X"F0",X"02",X"33",X"01",X"01",X"03",
		X"33",X"03",X"50",X"F0",X"F3",X"F0",X"F0",X"F0",X"30",X"02",X"F2",X"F2",X"F0",X"F0",X"F2",X"A2",
		X"01",X"33",X"02",X"F2",X"F1",X"D0",X"D0",X"D0",X"13",X"33",X"00",X"F0",X"F3",X"F0",X"F0",X"F0",
		X"03",X"00",X"A3",X"F3",X"F0",X"F0",X"F3",X"F0",X"A2",X"F0",X"50",X"52",X"F2",X"F2",X"F0",X"F0",
		X"03",X"00",X"31",X"03",X"C2",X"C2",X"C1",X"C0",X"53",X"50",X"03",X"03",X"80",X"D0",X"D3",X"D0",
		X"F0",X"F0",X"00",X"30",X"02",X"03",X"01",X"00",X"F0",X"F0",X"00",X"30",X"10",X"00",X"02",X"02",
		X"C0",X"00",X"30",X"30",X"00",X"21",X"33",X"32",X"C0",X"00",X"20",X"30",X"03",X"03",X"00",X"20",
		X"00",X"0F",X"0F",X"06",X"36",X"36",X"0F",X"0F",X"00",X"0A",X"00",X"32",X"36",X"02",X"00",X"CA",
		X"00",X"00",X"01",X"09",X"0C",X"09",X"01",X"10",X"00",X"05",X"02",X"06",X"0C",X"16",X"32",X"25",
		X"CF",X"CF",X"CF",X"CC",X"CC",X"CF",X"DF",X"DF",X"CF",X"CA",X"D0",X"DC",X"FC",X"F0",X"FA",X"FF",
		X"30",X"20",X"02",X"44",X"C4",X"C2",X"C0",X"C0",X"00",X"45",X"CD",X"CC",X"CC",X"CD",X"C5",X"C0",
		X"03",X"3C",X"3C",X"0C",X"FC",X"FC",X"FC",X"F3",X"02",X"33",X"39",X"09",X"F9",X"F9",X"F3",X"F2",
		X"01",X"33",X"06",X"F6",X"F6",X"F6",X"D3",X"D1",X"03",X"3C",X"3C",X"0C",X"FE",X"FF",X"FC",X"F3",
		X"FC",X"FC",X"56",X"06",X"3B",X"1B",X"0B",X"0F",X"F4",X"F4",X"F0",X"F8",X"08",X"28",X"3C",X"16",
		X"C7",X"C3",X"83",X"03",X"13",X"33",X"27",X"27",X"FB",X"FB",X"0F",X"0F",X"3F",X"0F",X"0F",X"0F",
		X"00",X"10",X"30",X"00",X"C0",X"C0",X"C0",X"CF",X"10",X"30",X"00",X"C0",X"C0",X"C0",X"C0",X"CF",
		X"0A",X"0A",X"3A",X"3A",X"0A",X"CA",X"CA",X"CF",X"00",X"00",X"30",X"20",X"40",X"C0",X"C0",X"CF",
		X"CF",X"C0",X"C0",X"C0",X"C0",X"00",X"30",X"30",X"CF",X"C0",X"C0",X"C0",X"C0",X"00",X"30",X"30",
		X"CF",X"CA",X"CA",X"CA",X"CA",X"0A",X"3A",X"0A",X"CF",X"C0",X"C0",X"C0",X"C0",X"00",X"30",X"30",
		X"00",X"00",X"30",X"30",X"00",X"F0",X"F0",X"FF",X"05",X"35",X"35",X"05",X"F5",X"F5",X"05",X"AF",
		X"00",X"00",X"00",X"30",X"30",X"00",X"C0",X"DF",X"00",X"00",X"00",X"30",X"30",X"00",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",
		X"DF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"30",X"00",X"F0",X"F0",X"F0",X"F0",X"10",X"00",X"30",X"00",X"00",X"F0",X"F0",X"F0",
		X"00",X"20",X"3F",X"0F",X"F0",X"FF",X"FF",X"F0",X"00",X"0A",X"3A",X"00",X"FA",X"FA",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"A0",X"A0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"10",X"00",X"A0",X"F0",
		X"F0",X"FF",X"FF",X"F0",X"FF",X"5F",X"00",X"00",X"F0",X"F0",X"FA",X"FA",X"F0",X"FA",X"FA",X"F0",
		X"F0",X"F0",X"F0",X"D0",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"D0",X"D0",X"80",
		X"20",X"40",X"C0",X"C0",X"CF",X"CF",X"C0",X"C0",X"D0",X"D0",X"C0",X"C0",X"C0",X"CA",X"C0",X"C0",
		X"CF",X"80",X"00",X"10",X"30",X"20",X"00",X"00",X"0A",X"10",X"30",X"20",X"00",X"00",X"00",X"00",
		X"CF",X"C0",X"C0",X"C0",X"8F",X"0F",X"30",X"00",X"CF",X"C0",X"C0",X"80",X"00",X"3A",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
