library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"27",X"76",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"25",X"76",X"75",
		X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"66",X"65",X"52",X"00",X"00",X"FF",X"00",X"02",X"77",
		X"77",X"77",X"72",X"00",X"00",X"FF",X"02",X"66",X"66",X"66",X"66",X"66",X"62",X"00",X"FF",X"00",
		X"E2",X"41",X"23",X"21",X"42",X"E0",X"00",X"FF",X"00",X"02",X"44",X"3A",X"34",X"42",X"00",X"00",
		X"FF",X"00",X"00",X"23",X"37",X"33",X"20",X"00",X"00",X"FF",X"00",X"00",X"24",X"33",X"34",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"02",X"43",X"42",X"00",X"00",X"00",X"FF",X"00",X"02",X"67",X"D7",
		X"D7",X"62",X"00",X"00",X"FF",X"00",X"26",X"67",X"15",X"D7",X"66",X"20",X"00",X"FF",X"00",X"26",
		X"65",X"DD",X"15",X"66",X"20",X"00",X"FF",X"00",X"26",X"65",X"81",X"D5",X"66",X"20",X"00",X"FF",
		X"00",X"23",X"57",X"B9",X"B7",X"53",X"20",X"00",X"FF",X"00",X"23",X"99",X"89",X"89",X"93",X"20",
		X"00",X"FF",X"00",X"02",X"88",X"98",X"98",X"82",X"00",X"00",X"FF",X"00",X"00",X"28",X"82",X"88",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"28",X"92",X"98",X"20",X"00",X"00",X"FF",X"00",X"00",X"22",
		X"22",X"22",X"20",X"00",X"00",X"FF",X"00",X"02",X"19",X"22",X"29",X"12",X"00",X"00",X"FF",X"00",
		X"02",X"22",X"22",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"26",X"66",X"76",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"77",X"20",
		X"00",X"00",X"FF",X"00",X"02",X"77",X"76",X"67",X"62",X"00",X"00",X"FF",X"00",X"02",X"77",X"66",
		X"77",X"72",X"00",X"00",X"FF",X"00",X"02",X"2E",X"E5",X"66",X"66",X"62",X"00",X"FF",X"02",X"2E",
		X"55",X"54",X"12",X"32",X"00",X"00",X"FF",X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",X"FF",
		X"00",X"00",X"23",X"34",X"33",X"32",X"00",X"00",X"FF",X"00",X"00",X"02",X"73",X"33",X"32",X"00",
		X"00",X"FF",X"00",X"02",X"22",X"74",X"47",X"70",X"00",X"00",X"FF",X"00",X"26",X"67",X"5D",X"D5",
		X"20",X"00",X"00",X"FF",X"02",X"66",X"76",X"75",X"11",X"52",X"20",X"00",X"FF",X"23",X"37",X"57",
		X"75",X"DD",X"54",X"42",X"00",X"FF",X"23",X"32",X"77",X"65",X"11",X"24",X"32",X"00",X"FF",X"02",
		X"26",X"66",X"7B",X"BB",X"22",X"20",X"00",X"FF",X"00",X"02",X"77",X"B8",X"8D",X"20",X"00",X"00",
		X"FF",X"02",X"22",X"22",X"88",X"DD",X"D2",X"00",X"00",X"FF",X"28",X"28",X"92",X"98",X"D8",X"DD",
		X"20",X"00",X"FF",X"2B",X"29",X"BB",X"22",X"28",X"D2",X"22",X"20",X"FF",X"22",X"22",X"22",X"B0",
		X"02",X"22",X"B1",X"20",X"FF",X"22",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"02",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",
		X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",
		X"77",X"77",X"72",X"00",X"00",X"FF",X"00",X"02",X"EE",X"66",X"66",X"66",X"62",X"00",X"FF",X"02",
		X"2E",X"55",X"54",X"12",X"32",X"00",X"00",X"FF",X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",
		X"FF",X"00",X"00",X"23",X"34",X"33",X"32",X"00",X"00",X"FF",X"00",X"00",X"02",X"73",X"33",X"32",
		X"00",X"00",X"FF",X"00",X"00",X"02",X"74",X"75",X"20",X"00",X"00",X"FF",X"00",X"00",X"26",X"67",
		X"D5",X"00",X"00",X"00",X"FF",X"00",X"02",X"66",X"75",X"71",X"50",X"00",X"00",X"FF",X"00",X"02",
		X"67",X"25",X"7D",X"50",X"00",X"00",X"FF",X"00",X"23",X"32",X"77",X"71",X"52",X"00",X"00",X"FF",
		X"00",X"24",X"32",X"77",X"99",X"42",X"00",X"00",X"FF",X"00",X"02",X"29",X"99",X"D2",X"20",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"88",X"DD",X"20",X"00",X"00",X"FF",X"00",X"00",X"02",X"2D",X"8D",
		X"82",X"00",X"00",X"FF",X"00",X"00",X"29",X"92",X"82",X"22",X"22",X"00",X"FF",X"00",X"02",X"82",
		X"92",X"22",X"29",X"12",X"00",X"FF",X"00",X"02",X"2B",X"20",X"02",X"22",X"20",X"00",X"FF",X"00",
		X"00",X"22",X"20",X"02",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",
		X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",X"77",X"77",X"72",X"00",X"00",X"FF",X"00",X"02",
		X"EE",X"66",X"66",X"66",X"62",X"00",X"FF",X"02",X"2E",X"55",X"54",X"12",X"32",X"00",X"00",X"FF",
		X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",X"FF",X"00",X"00",X"23",X"34",X"33",X"32",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"73",X"33",X"32",X"00",X"00",X"FF",X"00",X"00",X"02",X"74",X"75",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"57",X"77",X"D5",X"00",X"00",X"00",X"FF",X"00",X"00",X"27",
		X"66",X"71",X"50",X"00",X"00",X"FF",X"00",X"00",X"27",X"6C",X"5D",X"20",X"00",X"00",X"FF",X"00",
		X"00",X"27",X"76",X"51",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"33",X"5B",X"20",X"00",X"00",
		X"FF",X"00",X"00",X"29",X"43",X"82",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"8D",X"82",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"02",X"98",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"8D",
		X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"02",X"2B",X"12",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",
		X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",
		X"77",X"77",X"72",X"00",X"00",X"FF",X"00",X"02",X"EE",X"66",X"66",X"66",X"62",X"00",X"FF",X"02",
		X"2E",X"55",X"54",X"12",X"32",X"00",X"00",X"FF",X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",
		X"FF",X"00",X"00",X"23",X"34",X"33",X"32",X"00",X"00",X"FF",X"00",X"00",X"02",X"73",X"33",X"32",
		X"00",X"00",X"FF",X"00",X"00",X"02",X"74",X"75",X"20",X"00",X"00",X"FF",X"00",X"00",X"57",X"67",
		X"D5",X"00",X"00",X"00",X"FF",X"00",X"00",X"27",X"65",X"51",X"50",X"00",X"00",X"FF",X"00",X"02",
		X"27",X"66",X"62",X"50",X"00",X"00",X"FF",X"00",X"24",X"26",X"56",X"33",X"20",X"00",X"00",X"FF",
		X"00",X"02",X"66",X"65",X"34",X"20",X"00",X"00",X"FF",X"00",X"00",X"29",X"88",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"88",X"D2",X"20",X"00",X"00",X"FF",X"00",X"00",X"02",X"8D",X"D2",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"28",X"98",X"29",X"92",X"00",X"00",X"FF",X"00",X"02",X"22",
		X"82",X"29",X"92",X"20",X"00",X"FF",X"00",X"02",X"12",X"20",X"22",X"B8",X"20",X"00",X"FF",X"00",
		X"00",X"29",X"20",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",X"20",
		X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",X"77",
		X"77",X"72",X"00",X"00",X"FF",X"00",X"02",X"EE",X"66",X"66",X"66",X"62",X"00",X"FF",X"02",X"2E",
		X"55",X"54",X"12",X"32",X"00",X"00",X"FF",X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",X"FF",
		X"00",X"00",X"23",X"34",X"33",X"32",X"00",X"00",X"FF",X"00",X"00",X"02",X"43",X"33",X"32",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"54",X"45",X"20",X"00",X"00",X"FF",X"00",X"02",X"27",X"76",X"62",
		X"00",X"00",X"00",X"FF",X"00",X"27",X"55",X"76",X"6C",X"22",X"00",X"00",X"FF",X"02",X"34",X"26",
		X"75",X"67",X"33",X"20",X"00",X"FF",X"02",X"47",X"26",X"77",X"57",X"34",X"20",X"00",X"FF",X"00",
		X"22",X"66",X"67",X"92",X"22",X"00",X"00",X"FF",X"00",X"00",X"26",X"88",X"89",X"20",X"00",X"00",
		X"FF",X"00",X"22",X"D8",X"8D",X"DB",X"92",X"00",X"00",X"FF",X"02",X"12",X"9D",X"DD",X"B9",X"99",
		X"20",X"00",X"FF",X"02",X"B2",X"88",X"92",X"92",X"99",X"22",X"20",X"FF",X"02",X"22",X"22",X"20",
		X"00",X"2B",X"82",X"20",X"FF",X"02",X"20",X"00",X"00",X"00",X"22",X"22",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"02",X"B0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",
		X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",
		X"77",X"77",X"72",X"20",X"00",X"FF",X"00",X"02",X"EE",X"66",X"66",X"53",X"32",X"00",X"FF",X"02",
		X"2E",X"55",X"54",X"12",X"53",X"42",X"00",X"FF",X"00",X"02",X"53",X"44",X"76",X"65",X"20",X"00",
		X"FF",X"00",X"00",X"23",X"34",X"66",X"52",X"00",X"00",X"FF",X"00",X"00",X"02",X"76",X"66",X"32",
		X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"65",X"B0",X"00",X"00",X"FF",X"00",X"00",X"57",X"77",
		X"55",X"90",X"00",X"00",X"FF",X"00",X"02",X"77",X"77",X"71",X"B0",X"00",X"00",X"FF",X"00",X"26",
		X"67",X"77",X"5D",X"B0",X"00",X"00",X"FF",X"00",X"02",X"66",X"77",X"1B",X"00",X"00",X"00",X"FF",
		X"00",X"22",X"99",X"98",X"29",X"00",X"00",X"00",X"FF",X"22",X"29",X"89",X"82",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"28",X"92",X"20",X"00",X"00",X"00",X"00",X"FF",X"29",X"22",X"20",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"21",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",
		X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",X"77",X"77",X"72",X"20",X"00",X"FF",X"00",X"02",
		X"EE",X"66",X"66",X"53",X"32",X"00",X"FF",X"02",X"2E",X"55",X"54",X"12",X"53",X"42",X"00",X"FF",
		X"00",X"02",X"53",X"44",X"76",X"65",X"20",X"00",X"FF",X"00",X"00",X"23",X"34",X"66",X"52",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"76",X"66",X"32",X"00",X"00",X"FF",X"00",X"00",X"07",X"76",X"65",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"57",X"77",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"27",
		X"77",X"71",X"50",X"00",X"00",X"FF",X"00",X"00",X"27",X"77",X"5D",X"20",X"00",X"00",X"FF",X"00",
		X"02",X"66",X"77",X"5D",X"20",X"00",X"00",X"FF",X"00",X"00",X"26",X"68",X"92",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"29",X"8D",X"92",X"00",X"00",X"00",X"FF",X"00",X"02",X"98",X"99",X"20",X"00",
		X"00",X"00",X"FF",X"00",X"22",X"29",X"82",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"20",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"29",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"12",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",
		X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",
		X"77",X"77",X"72",X"20",X"00",X"FF",X"00",X"02",X"EE",X"66",X"66",X"53",X"32",X"00",X"FF",X"02",
		X"2E",X"55",X"54",X"12",X"53",X"42",X"00",X"FF",X"00",X"02",X"53",X"44",X"76",X"65",X"20",X"00",
		X"FF",X"00",X"00",X"23",X"34",X"66",X"52",X"00",X"00",X"FF",X"00",X"00",X"02",X"76",X"66",X"32",
		X"00",X"00",X"FF",X"00",X"00",X"07",X"76",X"65",X"20",X"00",X"00",X"FF",X"00",X"00",X"57",X"77",
		X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"27",X"77",X"71",X"50",X"00",X"00",X"FF",X"00",X"00",
		X"27",X"77",X"5D",X"20",X"00",X"00",X"FF",X"00",X"02",X"66",X"77",X"51",X"20",X"00",X"00",X"FF",
		X"00",X"00",X"26",X"68",X"9B",X"20",X"00",X"00",X"FF",X"00",X"00",X"02",X"99",X"98",X"22",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"98",X"89",X"82",X"22",X"20",X"FF",X"00",X"00",X"00",X"22",X"98",
		X"22",X"21",X"20",X"FF",X"00",X"00",X"00",X"00",X"22",X"22",X"92",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"02",X"22",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",
		X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",X"77",X"77",X"72",X"20",X"00",X"FF",X"00",X"02",
		X"EE",X"66",X"66",X"53",X"32",X"00",X"FF",X"02",X"2E",X"55",X"54",X"12",X"53",X"42",X"00",X"FF",
		X"00",X"02",X"53",X"44",X"76",X"65",X"20",X"00",X"FF",X"00",X"00",X"23",X"34",X"66",X"52",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"76",X"66",X"32",X"00",X"00",X"FF",X"00",X"00",X"07",X"76",X"65",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"57",X"77",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"27",
		X"77",X"71",X"50",X"00",X"00",X"FF",X"00",X"00",X"27",X"77",X"5D",X"22",X"00",X"22",X"FF",X"00",
		X"02",X"66",X"77",X"79",X"98",X"22",X"12",X"FF",X"00",X"00",X"26",X"68",X"99",X"88",X"22",X"92",
		X"FF",X"00",X"00",X"02",X"B9",X"98",X"99",X"22",X"22",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",
		X"22",X"22",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"26",
		X"66",X"77",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"27",X"76",X"67",X"20",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"02",X"57",X"77",X"77",X"72",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"02",X"EE",X"66",X"66",X"66",X"62",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"2E",
		X"55",X"54",X"12",X"32",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"53",X"44",X"74",
		X"33",X"20",X"00",X"00",X"FF",X"02",X"22",X"00",X"00",X"00",X"23",X"34",X"33",X"32",X"22",X"22",
		X"00",X"FF",X"22",X"2B",X"22",X"02",X"25",X"57",X"43",X"33",X"34",X"47",X"44",X"20",X"FF",X"22",
		X"BB",X"BB",X"B5",X"57",X"77",X"74",X"77",X"77",X"75",X"43",X"20",X"FF",X"22",X"22",X"22",X"97",
		X"77",X"56",X"77",X"75",X"22",X"22",X"22",X"00",X"FF",X"22",X"28",X"88",X"97",X"75",X"66",X"75",
		X"52",X"00",X"00",X"00",X"00",X"FF",X"29",X"29",X"89",X"99",X"76",X"67",X"52",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"21",X"22",X"22",X"23",X"36",X"72",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"00",X"02",X"33",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"27",X"76",X"67",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",
		X"55",X"76",X"66",X"62",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"57",X"77",X"77",
		X"72",X"00",X"00",X"00",X"FF",X"00",X"00",X"20",X"00",X"02",X"EE",X"66",X"66",X"66",X"62",X"00",
		X"00",X"FF",X"00",X"02",X"32",X"02",X"2E",X"55",X"54",X"12",X"32",X"00",X"00",X"00",X"FF",X"00",
		X"02",X"33",X"22",X"22",X"53",X"44",X"74",X"33",X"20",X"00",X"00",X"FF",X"00",X"02",X"33",X"56",
		X"66",X"23",X"34",X"33",X"32",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"56",X"66",X"67",X"43",
		X"33",X"32",X"00",X"00",X"00",X"FF",X"02",X"22",X"BB",X"22",X"76",X"67",X"74",X"47",X"20",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"BB",X"95",X"27",X"75",X"71",X"15",X"20",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"97",X"75",X"57",X"DD",X"27",X"72",X"00",X"00",X"00",X"FF",X"92",X"22",X"99",
		X"99",X"77",X"72",X"22",X"77",X"72",X"00",X"00",X"00",X"FF",X"22",X"28",X"88",X"99",X"22",X"20",
		X"00",X"27",X"77",X"20",X"00",X"00",X"FF",X"22",X"29",X"89",X"82",X"20",X"00",X"00",X"02",X"44",
		X"20",X"00",X"00",X"FF",X"29",X"22",X"22",X"20",X"00",X"00",X"00",X"02",X"44",X"20",X"00",X"00",
		X"FF",X"21",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"FF",X"02",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"22",X"20",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"27",X"72",X"33",X"32",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"02",X"55",X"23",X"44",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"02",X"52",X"27",X"52",X"72",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"E2",X"66",
		X"72",X"66",X"62",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"2E",X"26",X"67",X"22",X"32",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"26",X"72",X"74",X"33",X"20",X"00",X"00",X"FF",
		X"02",X"22",X"20",X"00",X"02",X"77",X"72",X"33",X"32",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",
		X"22",X"26",X"67",X"53",X"33",X"32",X"00",X"00",X"00",X"FF",X"22",X"22",X"99",X"96",X"66",X"77",
		X"75",X"22",X"20",X"00",X"00",X"00",X"FF",X"22",X"29",X"89",X"87",X"66",X"75",X"71",X"20",X"00",
		X"00",X"00",X"00",X"FF",X"22",X"22",X"98",X"97",X"77",X"7D",X"D2",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"22",X"22",X"98",X"89",X"77",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"29",X"22",
		X"22",X"22",X"22",X"25",X"72",X"00",X"00",X"00",X"00",X"00",X"FF",X"21",X"22",X"00",X"00",X"00",
		X"27",X"72",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"20",X"00",X"00",X"02",X"55",X"20",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"44",X"20",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"24",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",
		X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"77",X"20",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"27",X"76",X"67",X"20",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"02",X"57",X"77",X"77",X"72",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"EE",
		X"66",X"66",X"66",X"62",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"2E",X"55",X"54",X"12",X"32",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",X"00",
		X"FF",X"02",X"22",X"00",X"00",X"00",X"23",X"34",X"33",X"32",X"22",X"22",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"25",X"57",X"77",X"66",X"76",X"67",X"33",X"20",X"FF",X"22",X"29",X"82",X"55",X"57",
		X"77",X"76",X"66",X"77",X"75",X"34",X"20",X"FF",X"29",X"28",X"99",X"57",X"67",X"77",X"77",X"75",
		X"22",X"22",X"22",X"00",X"FF",X"21",X"22",X"88",X"97",X"66",X"67",X"77",X"52",X"00",X"00",X"00",
		X"00",X"FF",X"92",X"2B",X"22",X"98",X"77",X"77",X"52",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"2B",X"BB",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"2B",X"00",X"24",
		X"47",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"00",X"00",X"02",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"27",
		X"76",X"67",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"55",X"76",X"66",X"62",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"20",X"02",X"57",X"77",X"77",X"72",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"02",X"42",X"22",X"EE",X"66",X"66",X"66",X"62",X"00",X"00",X"FF",X"00",X"00",
		X"02",X"44",X"2E",X"55",X"54",X"12",X"32",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"44",X"72",
		X"53",X"44",X"74",X"33",X"20",X"00",X"00",X"FF",X"00",X"22",X"20",X"27",X"72",X"23",X"34",X"33",
		X"32",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"02",X"27",X"75",X"43",X"33",X"32",X"00",X"00",
		X"00",X"FF",X"22",X"92",X"22",X"27",X"77",X"77",X"75",X"52",X"20",X"00",X"00",X"00",X"FF",X"21",
		X"22",X"28",X"97",X"77",X"77",X"66",X"20",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"98",X"97",
		X"77",X"55",X"66",X"62",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"29",X"88",X"75",X"52",X"76",
		X"62",X"00",X"00",X"00",X"00",X"FF",X"22",X"2B",X"22",X"99",X"22",X"20",X"26",X"66",X"20",X"00",
		X"00",X"00",X"FF",X"22",X"29",X"B2",X"22",X"00",X"00",X"05",X"57",X"20",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"20",X"00",X"00",X"00",X"02",X"33",X"20",X"00",X"00",X"00",X"FF",X"02",X"20",X"00",
		X"00",X"00",X"00",X"02",X"43",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"77",X"22",X"20",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"27",X"76",X"67",X"24",X"42",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",
		X"55",X"76",X"66",X"62",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"57",X"77",X"77",
		X"72",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"EE",X"66",X"66",X"66",X"62",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"02",X"2E",X"55",X"54",X"12",X"32",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"02",X"53",X"44",X"74",X"33",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"23",X"34",X"33",X"32",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"02",X"27",X"75",X"43",
		X"33",X"32",X"00",X"00",X"00",X"FF",X"22",X"22",X"29",X"96",X"67",X"77",X"75",X"52",X"20",X"00",
		X"00",X"00",X"FF",X"22",X"22",X"89",X"87",X"66",X"77",X"66",X"20",X"00",X"00",X"00",X"00",X"FF",
		X"29",X"22",X"98",X"97",X"77",X"52",X"66",X"20",X"00",X"00",X"00",X"00",X"FF",X"21",X"22",X"28",
		X"89",X"75",X"52",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"00",X"02",X"22",X"22",X"26",
		X"62",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"26",X"62",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"57",X"20",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"23",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"24",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"27",X"76",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"25",X"76",X"75",X"20",
		X"00",X"00",X"FF",X"00",X"02",X"55",X"66",X"65",X"52",X"00",X"00",X"FF",X"00",X"02",X"77",X"77",
		X"77",X"72",X"00",X"00",X"FF",X"02",X"66",X"66",X"66",X"66",X"66",X"62",X"00",X"FF",X"00",X"E2",
		X"41",X"23",X"21",X"42",X"E0",X"00",X"FF",X"00",X"02",X"44",X"37",X"34",X"42",X"00",X"00",X"FF",
		X"00",X"00",X"21",X"D1",X"D1",X"20",X"00",X"00",X"FF",X"02",X"22",X"21",X"D1",X"D1",X"22",X"22",
		X"00",X"FF",X"23",X"77",X"53",X"33",X"33",X"57",X"73",X"20",X"FF",X"24",X"56",X"57",X"D7",X"D7",
		X"56",X"54",X"20",X"FF",X"02",X"22",X"67",X"15",X"D7",X"62",X"22",X"00",X"FF",X"00",X"05",X"65",
		X"DD",X"15",X"65",X"00",X"00",X"FF",X"00",X"05",X"65",X"81",X"D5",X"65",X"00",X"00",X"FF",X"02",
		X"20",X"59",X"B9",X"B9",X"50",X"22",X"00",X"FF",X"02",X"12",X"89",X"98",X"99",X"82",X"12",X"00",
		X"FF",X"02",X"92",X"98",X"99",X"98",X"92",X"92",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",
		X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"52",X"50",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"50",X"23",X"25",X"00",X"00",X"00",X"FF",X"00",X"00",X"52",X"33",X"32",X"50",X"00",X"00",X"FF",
		X"00",X"00",X"24",X"34",X"34",X"20",X"00",X"00",X"FF",X"00",X"22",X"24",X"44",X"44",X"22",X"20",
		X"00",X"FF",X"02",X"67",X"75",X"D1",X"D5",X"77",X"62",X"00",X"FF",X"23",X"61",X"29",X"89",X"89",
		X"21",X"63",X"20",X"FF",X"23",X"29",X"22",X"99",X"92",X"29",X"23",X"20",X"FF",X"22",X"22",X"22",
		X"99",X"92",X"22",X"22",X"20",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",X"20",X"00",X"FF",X"00",
		X"02",X"22",X"00",X"02",X"22",X"00",X"00",X"FF",X"01",X"01",X"10",X"11",X"01",X"10",X"10",X"FF",
		X"16",X"15",X"41",X"23",X"14",X"51",X"71",X"FF",X"11",X"76",X"65",X"55",X"66",X"77",X"11",X"FF",
		X"1C",X"58",X"83",X"D8",X"48",X"86",X"C1",X"FF",X"1C",X"58",X"83",X"88",X"48",X"86",X"C1",X"FF",
		X"16",X"55",X"43",X"23",X"44",X"56",X"71",X"FF",X"11",X"76",X"65",X"55",X"66",X"77",X"11",X"FF",
		X"16",X"65",X"43",X"23",X"44",X"56",X"71",X"FF",X"01",X"65",X"54",X"34",X"45",X"67",X"10",X"FF",
		X"01",X"76",X"55",X"55",X"56",X"71",X"10",X"FF",X"00",X"11",X"66",X"67",X"77",X"11",X"00",X"FF",
		X"00",X"00",X"11",X"61",X"11",X"00",X"00",X"FF",X"00",X"00",X"01",X"67",X"10",X"00",X"00",X"FF",
		X"00",X"01",X"16",X"67",X"71",X"10",X"00",X"FF",X"00",X"16",X"64",X"33",X"47",X"71",X"00",X"FF",
		X"00",X"01",X"11",X"11",X"11",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"B0",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"BB",X"BB",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BB",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"BB",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BB",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0B",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"0B",X"BB",X"B0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"B0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0B",
		X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0B",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"90",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"90",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"90",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"90",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"09",X"99",X"99",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"99",X"99",X"90",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"09",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"25",X"55",X"52",X"22",X"22",X"55",X"52",
		X"22",X"FF",X"55",X"55",X"22",X"22",X"25",X"55",X"52",X"22",X"FF",X"55",X"55",X"22",X"22",X"22",
		X"55",X"55",X"22",X"FF",X"25",X"55",X"52",X"22",X"25",X"55",X"BB",X"22",X"FF",X"22",X"55",X"52",
		X"25",X"55",X"5B",X"BB",X"B2",X"FF",X"22",X"58",X"82",X"22",X"55",X"5B",X"BB",X"BB",X"FF",X"25",
		X"88",X"88",X"82",X"55",X"BB",X"BB",X"BB",X"FF",X"08",X"88",X"88",X"88",X"88",X"BB",X"BB",X"B0",
		X"FF",X"00",X"88",X"88",X"88",X"88",X"BB",X"BB",X"00",X"FF",X"00",X"08",X"88",X"88",X"8B",X"BB",
		X"BB",X"00",X"FF",X"00",X"08",X"88",X"88",X"BB",X"BB",X"BB",X"00",X"FF",X"00",X"00",X"88",X"88",
		X"BB",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"88",X"88",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",
		X"88",X"88",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"08",X"88",X"8B",X"BB",X"B0",X"00",X"FF",
		X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"8B",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"8B",X"BB",
		X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"8B",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"8B",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"25",X"55",X"52",X"22",X"22",X"55",X"52",
		X"22",X"FF",X"55",X"55",X"22",X"22",X"25",X"55",X"52",X"22",X"FF",X"55",X"55",X"22",X"22",X"22",
		X"55",X"55",X"22",X"FF",X"25",X"55",X"52",X"22",X"25",X"55",X"BB",X"22",X"FF",X"22",X"55",X"52",
		X"25",X"55",X"5B",X"BB",X"B2",X"FF",X"22",X"58",X"82",X"22",X"55",X"5B",X"BB",X"BB",X"FF",X"25",
		X"88",X"88",X"82",X"55",X"BB",X"BB",X"EE",X"FF",X"08",X"88",X"88",X"88",X"88",X"BE",X"EE",X"E0",
		X"FF",X"00",X"88",X"88",X"88",X"EE",X"EE",X"BB",X"00",X"FF",X"00",X"08",X"88",X"88",X"8B",X"EB",
		X"BB",X"00",X"FF",X"00",X"08",X"88",X"88",X"BE",X"BB",X"BB",X"00",X"FF",X"00",X"00",X"88",X"88",
		X"BB",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"88",X"88",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",
		X"88",X"88",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"08",X"88",X"8B",X"BB",X"B0",X"00",X"FF",
		X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"8B",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"8B",X"BB",
		X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"8B",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"8B",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"25",X"55",X"52",X"22",X"22",X"55",X"52",
		X"22",X"FF",X"55",X"55",X"22",X"22",X"25",X"55",X"52",X"22",X"FF",X"55",X"55",X"22",X"22",X"22",
		X"55",X"55",X"22",X"FF",X"25",X"55",X"52",X"22",X"25",X"55",X"BB",X"22",X"FF",X"22",X"55",X"52",
		X"25",X"55",X"5B",X"BB",X"B2",X"FF",X"22",X"58",X"82",X"22",X"55",X"5B",X"BB",X"BB",X"FF",X"25",
		X"88",X"88",X"82",X"55",X"BB",X"BB",X"EE",X"FF",X"08",X"88",X"88",X"88",X"BB",X"BE",X"EE",X"00",
		X"FF",X"00",X"88",X"88",X"EE",X"EE",X"E0",X"00",X"00",X"FF",X"00",X"88",X"88",X"8B",X"70",X"00",
		X"00",X"00",X"FF",X"00",X"88",X"88",X"8B",X"BE",X"7B",X"B0",X"00",X"FF",X"00",X"08",X"88",X"88",
		X"E7",X"BB",X"00",X"00",X"FF",X"00",X"08",X"88",X"8E",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"08",
		X"88",X"88",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"08",X"88",X"8B",X"BB",X"B0",X"00",X"00",X"FF",
		X"00",X"08",X"88",X"8B",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"08",X"88",X"BB",X"BB",X"00",X"00",
		X"00",X"FF",X"00",X"08",X"88",X"BB",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"8B",X"BB",X"BB",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"8B",X"BB",X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"88",
		X"BB",X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"88",X"BB",X"B0",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"88",X"8B",X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"8B",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"BB",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"08",X"B0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"B0",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"25",X"55",X"52",X"22",X"22",X"55",X"52",
		X"22",X"FF",X"55",X"55",X"22",X"22",X"25",X"55",X"52",X"22",X"FF",X"55",X"55",X"22",X"22",X"22",
		X"55",X"55",X"22",X"FF",X"25",X"55",X"52",X"22",X"25",X"55",X"BB",X"22",X"FF",X"22",X"55",X"52",
		X"25",X"55",X"5B",X"BB",X"B2",X"FF",X"22",X"58",X"82",X"22",X"55",X"5B",X"BB",X"BB",X"FF",X"25",
		X"88",X"88",X"82",X"55",X"BB",X"BB",X"EE",X"FF",X"08",X"88",X"88",X"88",X"88",X"BE",X"EE",X"E0",
		X"FF",X"00",X"88",X"88",X"88",X"EE",X"E0",X"00",X"00",X"FF",X"00",X"08",X"88",X"80",X"00",X"00",
		X"BB",X"00",X"FF",X"00",X"08",X"88",X"88",X"B0",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"88",X"00",
		X"0B",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"88",X"80",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",
		X"88",X"88",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"08",X"88",X"8B",X"BB",X"B0",X"00",X"FF",
		X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"8B",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"8B",X"BB",
		X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"8B",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"8B",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"25",X"55",X"52",X"22",X"22",X"55",X"52",
		X"22",X"FF",X"55",X"55",X"22",X"22",X"25",X"55",X"52",X"22",X"FF",X"55",X"55",X"22",X"22",X"22",
		X"55",X"55",X"22",X"FF",X"25",X"55",X"52",X"22",X"25",X"55",X"BB",X"22",X"FF",X"22",X"55",X"52",
		X"25",X"55",X"5B",X"BB",X"B2",X"FF",X"22",X"58",X"82",X"22",X"55",X"5B",X"BB",X"BB",X"FF",X"25",
		X"88",X"88",X"82",X"55",X"BB",X"BB",X"EE",X"FF",X"08",X"88",X"88",X"88",X"88",X"BE",X"EE",X"E0",
		X"FF",X"00",X"88",X"88",X"88",X"EE",X"E0",X"00",X"00",X"FF",X"00",X"08",X"88",X"80",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"BB",X"B0",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"0B",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"88",X"00",X"8B",X"BB",X"B0",
		X"00",X"FF",X"00",X"00",X"88",X"88",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"08",X"88",X"8B",
		X"BB",X"B0",X"00",X"FF",X"00",X"00",X"08",X"88",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"08",
		X"88",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"08",X"8B",X"BB",X"B0",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"8B",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"BB",X"B0",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"88",X"8B",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"8B",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",
		X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"08",X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"8B",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"8B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"BB",X"FF",X"00",X"00",X"00",X"BB",X"B0",X"FF",
		X"00",X"00",X"0B",X"BB",X"B0",X"FF",X"88",X"00",X"8B",X"BB",X"B0",X"FF",X"88",X"88",X"8B",X"BB",
		X"B0",X"FF",X"08",X"88",X"8B",X"BB",X"B0",X"FF",X"08",X"88",X"BB",X"BB",X"00",X"FF",X"08",X"88",
		X"BB",X"BB",X"00",X"FF",X"08",X"8B",X"BB",X"B0",X"00",X"FF",X"00",X"8B",X"BB",X"B0",X"00",X"FF",
		X"00",X"88",X"BB",X"B0",X"00",X"FF",X"00",X"88",X"8B",X"B0",X"00",X"FF",X"00",X"88",X"8B",X"00",
		X"00",X"FF",X"00",X"08",X"BB",X"00",X"00",X"FF",X"00",X"08",X"BB",X"00",X"00",X"FF",X"00",X"08",
		X"BB",X"00",X"00",X"FF",X"00",X"08",X"8B",X"00",X"00",X"FF",X"00",X"08",X"8B",X"00",X"00",X"FF",
		X"00",X"00",X"8B",X"00",X"00",X"FF",X"00",X"00",X"80",X"00",X"00",X"FF",X"00",X"00",X"80",X"00",
		X"00",X"FF",X"00",X"00",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"88",X"A8",X"A8",X"00",X"FF",X"00",X"00",X"00",X"88",X"80",X"00",X"08",X"88",X"8A",X"8A",X"AA",
		X"B0",X"FF",X"00",X"00",X"08",X"88",X"8A",X"00",X"88",X"88",X"8A",X"8A",X"AB",X"B0",X"FF",X"00",
		X"00",X"08",X"88",X"AA",X"00",X"88",X"88",X"A8",X"AA",X"AB",X"AA",X"FF",X"00",X"00",X"88",X"8A",
		X"AB",X"08",X"88",X"8A",X"A8",X"AA",X"BA",X"AB",X"FF",X"00",X"00",X"88",X"AB",X"B4",X"0B",X"BA",
		X"AA",X"A8",X"AA",X"BA",X"BB",X"FF",X"00",X"08",X"8A",X"B4",X"40",X"0B",X"BB",X"AA",X"B8",X"AB",
		X"AB",X"BB",X"FF",X"00",X"8A",X"B4",X"40",X"00",X"0B",X"BB",X"BA",X"B8",X"AB",X"AB",X"B4",X"FF",
		X"00",X"8B",X"40",X"08",X"8B",X"00",X"44",X"BB",X"BB",X"8A",X"BB",X"40",X"FF",X"08",X"B4",X"00",
		X"A8",X"AB",X"40",X"00",X"44",X"BB",X"8A",X"B4",X"40",X"FF",X"8B",X"00",X"00",X"0A",X"44",X"00",
		X"8A",X"00",X"44",X"48",X"44",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"FF",X"06",X"56",X"00",X"10",
		X"06",X"56",X"00",X"FF",X"65",X"60",X"00",X"10",X"00",X"65",X"60",X"FF",X"66",X"03",X"11",X"11",
		X"13",X"06",X"60",X"FF",X"70",X"16",X"44",X"45",X"56",X"10",X"70",X"FF",X"01",X"64",X"66",X"66",
		X"65",X"61",X"00",X"FF",X"36",X"56",X"DD",X"DD",X"D6",X"56",X"30",X"FF",X"15",X"6D",X"D2",X"12",
		X"DD",X"65",X"10",X"FF",X"15",X"6D",X"22",X"12",X"2D",X"65",X"10",X"FF",X"15",X"6D",X"22",X"11",
		X"1D",X"65",X"10",X"FF",X"15",X"6D",X"22",X"22",X"2D",X"65",X"10",X"FF",X"15",X"6D",X"D2",X"22",
		X"DD",X"65",X"10",X"FF",X"36",X"56",X"DD",X"DD",X"D6",X"56",X"30",X"FF",X"01",X"65",X"66",X"66",
		X"65",X"61",X"00",X"FF",X"00",X"16",X"55",X"55",X"56",X"10",X"00",X"FF",X"00",X"93",X"11",X"11",
		X"13",X"90",X"00",X"FF",X"09",X"90",X"00",X"00",X"00",X"99",X"00",X"FF",X"00",X"00",X"00",X"99",
		X"22",X"22",X"22",X"22",X"FF",X"02",X"00",X"00",X"09",X"24",X"44",X"44",X"40",X"FF",X"29",X"22",
		X"00",X"02",X"42",X"24",X"44",X"00",X"FF",X"02",X"92",X"21",X"32",X"44",X"42",X"24",X"40",X"FF",
		X"00",X"22",X"22",X"32",X"44",X"44",X"42",X"22",X"FF",X"02",X"72",X"23",X"12",X"24",X"44",X"44",
		X"40",X"FF",X"22",X"22",X"23",X"11",X"24",X"44",X"44",X"00",X"FF",X"08",X"62",X"02",X"21",X"22",
		X"43",X"32",X"10",X"FF",X"00",X"00",X"02",X"22",X"12",X"31",X"11",X"0F",X"FF",X"00",X"00",X"00",
		X"29",X"91",X"12",X"20",X"00",X"FF",X"00",X"00",X"00",X"92",X"29",X"20",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"FF",X"02",X"92",X"20",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"29",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"27",X"22",X"22",X"32",X"20",X"00",X"00",X"FF",X"02",X"22",X"22",X"33",
		X"22",X"22",X"20",X"00",X"FF",X"00",X"86",X"23",X"22",X"44",X"44",X"12",X"00",X"FF",X"00",X"62",
		X"32",X"22",X"24",X"44",X"41",X"22",X"FF",X"09",X"90",X"24",X"44",X"42",X"24",X"41",X"20",X"FF",
		X"00",X"99",X"22",X"44",X"44",X"42",X"44",X"00",X"FF",X"00",X"02",X"44",X"24",X"44",X"44",X"24",
		X"00",X"FF",X"00",X"24",X"44",X"42",X"44",X"00",X"20",X"00",X"FF",X"00",X"24",X"00",X"42",X"40",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"45",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"10",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"FF",X"55",X"5D",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"55",X"55",X"55",
		X"55",X"55",X"00",X"FF",X"55",X"DD",X"EE",X"ED",X"DE",X"EE",X"EE",X"DD",X"EE",X"ED",X"DD",X"EE",
		X"EE",X"DD",X"EE",X"EE",X"ED",X"55",X"55",X"55",X"55",X"50",X"00",X"FF",X"44",X"DE",X"DD",X"DE",
		X"DD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"ED",X"DD",X"ED",X"DD",X"ED",X"DD",X"44",X"44",X"44",
		X"44",X"00",X"00",X"FF",X"55",X"DE",X"DD",X"DD",X"D5",X"DE",X"D5",X"DE",X"DD",X"DE",X"DD",X"ED",
		X"DD",X"ED",X"5D",X"ED",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"FF",X"55",X"DD",X"EE",X"ED",
		X"D5",X"DE",X"D5",X"DE",X"DD",X"DE",X"DD",X"EE",X"EE",X"DD",X"5D",X"ED",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"FF",X"55",X"DD",X"DD",X"DE",X"D5",X"DE",X"D5",X"DE",X"EE",X"EE",X"DD",X"ED",
		X"DE",X"D5",X"5D",X"ED",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"FF",X"44",X"DE",X"DD",X"DE",
		X"D4",X"DE",X"D4",X"DE",X"DD",X"DE",X"DD",X"ED",X"DE",X"DD",X"4D",X"ED",X"44",X"44",X"40",X"00",
		X"00",X"00",X"00",X"FF",X"55",X"DD",X"EE",X"ED",X"D5",X"DE",X"D5",X"DE",X"D5",X"DE",X"DD",X"ED",
		X"DD",X"ED",X"5D",X"ED",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"FF",X"55",X"5D",X"DD",X"DD",
		X"55",X"DD",X"D5",X"DD",X"D5",X"DD",X"DD",X"DD",X"5D",X"DD",X"5D",X"DD",X"55",X"55",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"45",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"00",X"00",X"00",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"00",X"00",X"00",X"FF",X"44",X"33",X"33",X"33",
		X"33",X"33",X"34",X"40",X"00",X"00",X"00",X"FF",X"44",X"33",X"33",X"33",X"33",X"33",X"34",X"40",
		X"00",X"00",X"00",X"FF",X"44",X"00",X"00",X"00",X"43",X"33",X"34",X"40",X"00",X"00",X"00",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"40",X"00",X"00",X"00",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",
		X"00",X"00",X"00",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"00",X"00",X"00",X"FF",
		X"33",X"04",X"43",X"33",X"44",X"33",X"33",X"30",X"00",X"00",X"00",X"FF",X"33",X"44",X"33",X"34",
		X"43",X"33",X"33",X"31",X"00",X"00",X"00",X"FF",X"33",X"43",X"33",X"44",X"33",X"34",X"33",X"35",
		X"00",X"00",X"00",X"FF",X"33",X"33",X"34",X"43",X"33",X"43",X"33",X"35",X"00",X"00",X"44",X"FF",
		X"33",X"33",X"44",X"33",X"34",X"45",X"33",X"35",X"00",X"44",X"44",X"FF",X"33",X"34",X"43",X"33",
		X"54",X"45",X"33",X"35",X"04",X"33",X"34",X"FF",X"33",X"44",X"33",X"34",X"44",X"44",X"33",X"35",
		X"33",X"33",X"34",X"FF",X"33",X"41",X"11",X"11",X"11",X"11",X"11",X"11",X"33",X"30",X"34",X"FF",
		X"33",X"46",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"30",X"00",X"FF",X"33",X"46",X"6E",X"EE",
		X"EE",X"EE",X"EE",X"66",X"33",X"30",X"44",X"FF",X"33",X"46",X"66",X"EE",X"EE",X"EE",X"E6",X"66",
		X"33",X"44",X"44",X"FF",X"33",X"46",X"E6",X"6E",X"EE",X"EE",X"66",X"E6",X"34",X"33",X"34",X"FF",
		X"33",X"46",X"EE",X"66",X"EE",X"E6",X"6E",X"E6",X"43",X"33",X"34",X"FF",X"33",X"46",X"EE",X"E6",
		X"6E",X"66",X"EE",X"E6",X"43",X"30",X"34",X"FF",X"33",X"46",X"EE",X"EE",X"66",X"6E",X"EE",X"E6",
		X"43",X"30",X"00",X"FF",X"33",X"46",X"EE",X"EE",X"66",X"6E",X"EE",X"E6",X"43",X"30",X"00",X"FF",
		X"33",X"46",X"EE",X"E6",X"6E",X"66",X"EE",X"E6",X"43",X"30",X"00",X"FF",X"33",X"46",X"EE",X"66",
		X"EE",X"E6",X"6E",X"E6",X"43",X"30",X"00",X"FF",X"33",X"46",X"E6",X"6E",X"EE",X"EE",X"66",X"E6",
		X"43",X"30",X"00",X"FF",X"33",X"46",X"66",X"EE",X"EE",X"EE",X"E6",X"66",X"43",X"30",X"00",X"FF",
		X"33",X"46",X"6E",X"EE",X"EE",X"EE",X"EE",X"66",X"43",X"30",X"00",X"FF",X"33",X"46",X"66",X"66",
		X"66",X"66",X"66",X"66",X"43",X"30",X"00",X"FF",X"33",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"43",X"30",X"00",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"CC",X"CC",X"9C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"3C",X"CC",X"49",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"CC",X"C4",X"CC",X"C9",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"55",X"55",X"55",X"CC",X"CC",X"C0",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"2A",X"AA",X"A9",X"55",X"CC",X"00",X"54",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"02",X"AA",X"AA",X"99",X"55",X"55",X"54",X"53",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"C2",X"AA",X"AA",X"99",X"AA",X"AA",X"44",X"53",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"54",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"CC",X"24",X"44",X"22",X"22",X"22",X"24",X"44",X"53",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"C2",X"22",X"22",X"88",X"88",X"38",X"82",X"22",X"53",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"C8",X"38",X"38",X"38",X"38",X"83",X"83",X"83",X"9A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"C9",X"C4",X"44",X"44",X"94",X"44",X"44",X"89",X"9A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"C9",X"44",X"11",X"11",X"99",X"41",X"11",X"89",X"A4",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"99",X"41",X"11",X"18",X"94",X"11",X"18",X"99",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"99",X"41",X"11",X"88",X"94",X"11",X"18",X"90",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"99",X"41",X"18",X"99",X"41",X"11",X"88",X"90",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"98",X"88",X"88",X"98",X"88",X"88",X"89",X"94",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"14",X"41",X"00",X"03",X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"B4",X"41",X"00",X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"01",X"10",X"00",X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"CC",X"70",X"00",X"0B",X"90",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"C7",X"0C",X"99",X"A0",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"C5",X"30",X"CC",X"CC",X"77",X"C9",X"9A",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0C",X"C3",X"3C",X"07",X"CC",X"77",X"99",X"AC",X"CC",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"5C",X"CC",X"CC",X"CC",X"77",X"C9",X"9A",X"AC",X"CC",X"CC",X"C0",X"00",X"00",X"FF",
		X"00",X"00",X"55",X"C7",X"CC",X"7C",X"CC",X"C9",X"77",X"79",X"55",X"55",X"70",X"00",X"00",X"FF",
		X"00",X"00",X"09",X"C7",X"CC",X"C5",X"55",X"CC",X"7C",X"79",X"9A",X"A5",X"77",X"00",X"00",X"FF",
		X"00",X"00",X"07",X"CC",X"77",X"58",X"88",X"CC",X"3C",X"CC",X"9A",X"AA",X"50",X"00",X"00",X"FF",
		X"00",X"00",X"77",X"C5",X"55",X"58",X"44",X"CC",X"99",X"CC",X"7A",X"AA",X"55",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"53",X"83",X"44",X"13",X"9C",X"C0",X"C7",X"77",X"7A",X"70",X"00",X"00",X"FF",
		X"00",X"00",X"0C",X"99",X"44",X"11",X"C9",X"CC",X"C9",X"CC",X"77",X"7C",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"CC",X"94",X"41",X"11",X"CC",X"CC",X"CC",X"CC",X"CC",X"70",X"0C",X"00",X"00",X"FF",
		X"00",X"00",X"CC",X"C4",X"11",X"18",X"9C",X"CC",X"44",X"44",X"54",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"55",X"CC",X"C8",X"11",X"8C",X"CC",X"CC",X"54",X"44",X"53",X"9C",X"C0",X"0C",X"00",X"FF",
		X"00",X"54",X"77",X"08",X"18",X"CC",X"C3",X"CC",X"85",X"55",X"53",X"9C",X"C0",X"0C",X"C0",X"FF",
		X"00",X"91",X"10",X"CC",X"C7",X"CC",X"C3",X"93",X"83",X"83",X"9A",X"AC",X"70",X"09",X"B0",X"FF",
		X"00",X"09",X"91",X"CC",X"37",X"C8",X"CC",X"C4",X"44",X"89",X"9A",X"AC",X"70",X"00",X"90",X"FF",
		X"00",X"00",X"0C",X"77",X"CC",X"88",X"CC",X"B1",X"11",X"89",X"A4",X"47",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0C",X"C5",X"1C",X"CC",X"CC",X"B1",X"18",X"C9",X"4C",X"40",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"59",X"41",X"14",X"CC",X"B1",X"18",X"9C",X"4C",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"99",X"48",X"11",X"4C",X"C1",X"88",X"9C",X"47",X"0C",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"11",X"09",X"99",X"11",X"14",X"71",X"19",X"94",X"47",X"0C",X"00",X"00",X"00",X"FF",
		X"00",X"0B",X"44",X"10",X"99",X"11",X"47",X"7C",X"89",X"CC",X"77",X"0C",X"C0",X"00",X"00",X"FF",
		X"00",X"01",X"44",X"10",X"09",X"88",X"77",X"00",X"CC",X"77",X"00",X"01",X"C0",X"00",X"00",X"FF",
		X"00",X"00",X"11",X"00",X"09",X"99",X"70",X"00",X"99",X"00",X"00",X"B4",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"00",X"00",X"14",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"05",X"A5",X"00",X"00",X"55",X"55",X"59",X"4B",X"B5",X"90",X"00",X"FF",
		X"00",X"00",X"00",X"55",X"55",X"A5",X"30",X"00",X"42",X"83",X"99",X"99",X"48",X"90",X"00",X"FF",
		X"00",X"00",X"05",X"AA",X"AA",X"A5",X"30",X"00",X"42",X"88",X"41",X"88",X"98",X"90",X"00",X"FF",
		X"00",X"00",X"04",X"44",X"4A",X"A5",X"80",X"00",X"42",X"83",X"41",X"18",X"99",X"90",X"00",X"FF",
		X"00",X"00",X"00",X"04",X"44",X"A8",X"80",X"00",X"44",X"28",X"41",X"11",X"88",X"90",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"83",X"41",X"11",X"18",X"90",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"88",X"44",X"11",X"18",X"90",X"00",X"FF",
		X"00",X"00",X"B1",X"00",X"00",X"00",X"88",X"90",X"88",X"83",X"94",X"44",X"48",X"90",X"00",X"FF",
		X"00",X"01",X"44",X"10",X"00",X"08",X"99",X"90",X"00",X"88",X"99",X"99",X"98",X"90",X"00",X"FF",
		X"00",X"0B",X"11",X"B0",X"00",X"89",X"94",X"40",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"FF",
		X"00",X"00",X"BB",X"00",X"00",X"99",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",
		X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",
		X"77",X"77",X"72",X"00",X"00",X"FF",X"02",X"77",X"66",X"66",X"66",X"77",X"72",X"00",X"FF",X"00",
		X"27",X"EE",X"55",X"5E",X"E7",X"20",X"00",X"FF",X"00",X"24",X"E5",X"55",X"55",X"E4",X"20",X"00",
		X"FF",X"00",X"02",X"25",X"54",X"55",X"22",X"00",X"00",X"FF",X"00",X"00",X"22",X"43",X"42",X"20",
		X"00",X"00",X"FF",X"00",X"02",X"55",X"66",X"65",X"52",X"00",X"00",X"FF",X"00",X"26",X"56",X"66",
		X"66",X"56",X"20",X"00",X"FF",X"00",X"26",X"76",X"66",X"66",X"76",X"20",X"00",X"FF",X"00",X"26",
		X"56",X"66",X"66",X"56",X"20",X"00",X"FF",X"00",X"26",X"E7",X"6E",X"67",X"E6",X"20",X"00",X"FF",
		X"00",X"23",X"4B",X"6E",X"69",X"43",X"20",X"00",X"FF",X"00",X"02",X"98",X"DA",X"D8",X"92",X"00",
		X"00",X"FF",X"00",X"00",X"28",X"8B",X"88",X"20",X"00",X"00",X"FF",X"00",X"00",X"2A",X"82",X"8A",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"2D",X"82",X"8D",X"20",X"00",X"00",X"FF",X"00",X"00",X"29",
		X"D2",X"D9",X"20",X"00",X"00",X"FF",X"00",X"02",X"19",X"20",X"2B",X"12",X"00",X"00",X"FF",X"00",
		X"02",X"22",X"20",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"77",X"62",X"22",X"00",X"00",X"FF",X"00",X"00",X"02",X"76",X"66",X"75",
		X"20",X"00",X"FF",X"00",X"00",X"26",X"66",X"67",X"55",X"20",X"00",X"FF",X"00",X"00",X"26",X"67",
		X"77",X"75",X"22",X"00",X"FF",X"00",X"02",X"27",X"77",X"66",X"66",X"67",X"20",X"FF",X"00",X"27",
		X"66",X"66",X"55",X"EE",X"72",X"20",X"FF",X"00",X"02",X"4E",X"55",X"55",X"5E",X"42",X"00",X"FF",
		X"00",X"00",X"22",X"55",X"45",X"52",X"22",X"00",X"FF",X"00",X"00",X"22",X"24",X"34",X"22",X"76",
		X"20",X"FF",X"00",X"02",X"65",X"56",X"66",X"55",X"66",X"20",X"FF",X"00",X"26",X"65",X"66",X"66",
		X"65",X"67",X"20",X"FF",X"00",X"26",X"77",X"66",X"66",X"67",X"72",X"00",X"FF",X"00",X"02",X"E6",
		X"66",X"66",X"66",X"20",X"00",X"FF",X"00",X"02",X"56",X"66",X"E6",X"6B",X"20",X"00",X"FF",X"00",
		X"00",X"57",X"99",X"88",X"89",X"20",X"00",X"FF",X"00",X"02",X"92",X"88",X"AA",X"89",X"20",X"00",
		X"FF",X"00",X"02",X"22",X"20",X"B8",X"82",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"28",X"A2",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"28",X"D2",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"2D",X"92",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"22",X"12",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"22",X"20",X"00",X"FF",
		X"00",X"00",X"00",X"22",X"22",X"20",X"00",X"00",X"FF",X"00",X"00",X"02",X"77",X"66",X"62",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"76",X"67",X"72",X"00",X"00",X"FF",X"00",X"00",X"26",X"66",X"67",
		X"55",X"20",X"00",X"FF",X"00",X"00",X"27",X"77",X"77",X"75",X"20",X"00",X"FF",X"00",X"27",X"77",
		X"66",X"66",X"66",X"77",X"20",X"FF",X"00",X"02",X"7E",X"E5",X"55",X"EE",X"72",X"00",X"FF",X"00",
		X"02",X"4E",X"55",X"55",X"5E",X"42",X"00",X"FF",X"00",X"00",X"22",X"55",X"45",X"52",X"EE",X"20",
		X"FF",X"00",X"00",X"02",X"24",X"34",X"22",X"6E",X"20",X"FF",X"00",X"00",X"25",X"56",X"66",X"55",
		X"66",X"20",X"FF",X"00",X"02",X"65",X"66",X"66",X"65",X"67",X"20",X"FF",X"00",X"26",X"77",X"66",
		X"66",X"66",X"72",X"00",X"FF",X"00",X"27",X"E6",X"66",X"66",X"66",X"20",X"00",X"FF",X"00",X"02",
		X"26",X"66",X"E6",X"6E",X"20",X"00",X"FF",X"00",X"00",X"27",X"78",X"88",X"99",X"20",X"00",X"FF",
		X"00",X"02",X"B2",X"88",X"AA",X"89",X"20",X"00",X"FF",X"00",X"02",X"BB",X"29",X"B8",X"82",X"00",
		X"00",X"FF",X"00",X"02",X"89",X"B2",X"28",X"A2",X"00",X"00",X"FF",X"00",X"21",X"92",X"20",X"28",
		X"D2",X"00",X"00",X"FF",X"00",X"22",X"22",X"00",X"2D",X"92",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"91",X"20",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"02",X"22",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"26",X"66",X"77",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",
		X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",X"77",X"77",X"72",X"00",X"00",X"FF",X"02",X"77",
		X"66",X"66",X"66",X"77",X"72",X"00",X"FF",X"00",X"27",X"EE",X"55",X"5E",X"E7",X"20",X"00",X"FF",
		X"00",X"24",X"E5",X"55",X"55",X"E4",X"20",X"00",X"FF",X"02",X"EE",X"25",X"54",X"55",X"2E",X"E2",
		X"00",X"FF",X"02",X"56",X"E2",X"43",X"42",X"E6",X"52",X"00",X"FF",X"02",X"66",X"55",X"66",X"65",
		X"56",X"62",X"00",X"FF",X"00",X"26",X"56",X"66",X"66",X"56",X"20",X"00",X"FF",X"00",X"2E",X"76",
		X"66",X"66",X"7E",X"20",X"00",X"FF",X"00",X"02",X"56",X"66",X"66",X"52",X"00",X"00",X"FF",X"00",
		X"02",X"E6",X"6E",X"66",X"E2",X"00",X"00",X"FF",X"00",X"02",X"B9",X"8A",X"89",X"B2",X"00",X"00",
		X"FF",X"00",X"00",X"28",X"D9",X"D8",X"20",X"00",X"00",X"FF",X"00",X"00",X"28",X"8B",X"88",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"2A",X"82",X"8A",X"20",X"00",X"00",X"FF",X"00",X"00",X"2D",X"82",
		X"8D",X"20",X"00",X"00",X"FF",X"00",X"00",X"29",X"D2",X"D9",X"20",X"00",X"00",X"FF",X"00",X"02",
		X"19",X"20",X"2B",X"12",X"00",X"00",X"FF",X"00",X"02",X"22",X"20",X"22",X"22",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"26",X"77",X"00",X"00",
		X"00",X"FF",X"00",X"02",X"57",X"66",X"67",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",
		X"62",X"00",X"00",X"FF",X"00",X"22",X"57",X"77",X"76",X"62",X"00",X"00",X"FF",X"02",X"76",X"66",
		X"66",X"77",X"72",X"20",X"00",X"FF",X"02",X"27",X"EE",X"55",X"66",X"66",X"72",X"00",X"FF",X"00",
		X"24",X"E5",X"55",X"55",X"E4",X"20",X"00",X"FF",X"00",X"22",X"25",X"54",X"55",X"22",X"00",X"00",
		X"FF",X"02",X"67",X"22",X"43",X"42",X"22",X"00",X"00",X"FF",X"02",X"66",X"55",X"66",X"65",X"56",
		X"20",X"00",X"FF",X"02",X"76",X"56",X"66",X"66",X"56",X"62",X"00",X"FF",X"00",X"27",X"76",X"66",
		X"66",X"77",X"62",X"00",X"FF",X"00",X"02",X"66",X"66",X"66",X"6E",X"20",X"00",X"FF",X"00",X"02",
		X"B6",X"6E",X"66",X"65",X"20",X"00",X"FF",X"00",X"02",X"98",X"88",X"99",X"75",X"00",X"00",X"FF",
		X"00",X"02",X"98",X"AA",X"88",X"29",X"20",X"00",X"FF",X"00",X"00",X"28",X"8B",X"02",X"22",X"20",
		X"00",X"FF",X"00",X"00",X"2A",X"82",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"2D",X"82",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"29",X"D2",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",
		X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"21",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"02",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"26",X"66",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"67",X"20",
		X"00",X"00",X"FF",X"00",X"02",X"55",X"76",X"66",X"62",X"00",X"00",X"FF",X"00",X"02",X"57",X"77",
		X"77",X"72",X"00",X"00",X"FF",X"02",X"77",X"66",X"66",X"66",X"77",X"72",X"00",X"FF",X"00",X"27",
		X"EE",X"55",X"5E",X"E7",X"20",X"00",X"FF",X"00",X"24",X"E5",X"55",X"55",X"E4",X"20",X"00",X"FF",
		X"02",X"EE",X"25",X"54",X"55",X"22",X"00",X"00",X"FF",X"02",X"E6",X"22",X"43",X"42",X"20",X"00",
		X"00",X"FF",X"02",X"66",X"55",X"66",X"65",X"52",X"00",X"00",X"FF",X"02",X"76",X"56",X"66",X"66",
		X"56",X"20",X"00",X"FF",X"00",X"27",X"66",X"66",X"66",X"77",X"62",X"00",X"FF",X"00",X"02",X"66",
		X"66",X"66",X"6E",X"72",X"00",X"FF",X"00",X"02",X"E6",X"6E",X"66",X"62",X"20",X"00",X"FF",X"00",
		X"02",X"99",X"88",X"87",X"72",X"00",X"00",X"FF",X"00",X"02",X"98",X"AA",X"88",X"2B",X"20",X"00",
		X"FF",X"00",X"00",X"28",X"8B",X"92",X"BB",X"20",X"00",X"FF",X"00",X"00",X"2A",X"82",X"2B",X"98",
		X"20",X"00",X"FF",X"00",X"00",X"2D",X"82",X"02",X"29",X"12",X"00",X"FF",X"00",X"00",X"29",X"D2",
		X"00",X"22",X"22",X"00",X"FF",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"19",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",
		X"51",X"16",X"51",X"11",X"11",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",X"11",X"65",
		X"FF",X"51",X"16",X"51",X"11",X"11",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",X"11",
		X"65",X"FF",X"51",X"16",X"51",X"11",X"11",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",
		X"11",X"65",X"FF",X"51",X"16",X"55",X"55",X"55",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",
		X"11",X"11",X"65",X"FF",X"51",X"16",X"56",X"66",X"44",X"51",X"11",X"11",X"11",X"16",X"51",X"11",
		X"11",X"11",X"11",X"65",X"FF",X"51",X"16",X"51",X"11",X"64",X"51",X"11",X"11",X"11",X"16",X"51",
		X"11",X"11",X"11",X"11",X"55",X"FF",X"56",X"16",X"55",X"11",X"13",X"51",X"11",X"11",X"11",X"16",
		X"51",X"11",X"11",X"11",X"55",X"51",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"11",
		X"16",X"51",X"11",X"11",X"15",X"64",X"56",X"FF",X"56",X"66",X"66",X"26",X"32",X"24",X"24",X"45",
		X"51",X"64",X"51",X"11",X"11",X"65",X"11",X"55",X"FF",X"51",X"11",X"11",X"11",X"33",X"21",X"11",
		X"44",X"51",X"65",X"51",X"61",X"64",X"45",X"11",X"15",X"FF",X"51",X"11",X"11",X"11",X"21",X"11",
		X"11",X"14",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"15",X"FF",X"55",X"11",X"11",X"11",X"11",
		X"21",X"11",X"16",X"56",X"32",X"26",X"26",X"64",X"64",X"45",X"65",X"FF",X"15",X"11",X"11",X"11",
		X"11",X"11",X"11",X"16",X"51",X"13",X"21",X"11",X"11",X"11",X"14",X"55",X"FF",X"15",X"11",X"11",
		X"11",X"11",X"21",X"11",X"16",X"51",X"13",X"21",X"11",X"11",X"11",X"11",X"65",X"FF",X"65",X"11",
		X"11",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"31",X"11",X"11",X"11",X"11",X"55",X"FF",X"55",
		X"11",X"11",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",X"11",X"11",X"11",X"51",X"FF",
		X"55",X"11",X"11",X"11",X"11",X"11",X"16",X"55",X"51",X"11",X"11",X"11",X"11",X"11",X"11",X"51",
		X"FF",X"53",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"11",X"11",X"11",X"11",
		X"51",X"FF",X"53",X"22",X"66",X"66",X"46",X"44",X"56",X"66",X"66",X"66",X"44",X"55",X"11",X"11",
		X"11",X"55",X"FF",X"51",X"31",X"11",X"11",X"11",X"64",X"56",X"11",X"11",X"11",X"16",X"65",X"55",
		X"55",X"55",X"55",X"FF",X"52",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",X"11",X"65",
		X"66",X"66",X"64",X"45",X"FF",X"51",X"11",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",X"11",
		X"65",X"61",X"11",X"11",X"45",X"FF",X"55",X"55",X"11",X"11",X"11",X"16",X"51",X"11",X"11",X"11",
		X"11",X"65",X"11",X"11",X"11",X"65",X"FF",X"56",X"64",X"51",X"11",X"11",X"16",X"51",X"11",X"11",
		X"11",X"11",X"55",X"11",X"11",X"11",X"65",X"FF",X"51",X"16",X"51",X"11",X"11",X"16",X"35",X"55",
		X"55",X"55",X"55",X"55",X"61",X"11",X"11",X"65",X"FF",X"51",X"16",X"51",X"11",X"11",X"13",X"32",
		X"25",X"66",X"64",X"55",X"32",X"41",X"11",X"11",X"65",X"FF",X"51",X"16",X"51",X"11",X"11",X"11",
		X"13",X"55",X"61",X"16",X"65",X"32",X"11",X"11",X"11",X"65",X"FF",X"51",X"11",X"55",X"55",X"55",
		X"55",X"55",X"55",X"11",X"11",X"65",X"12",X"11",X"11",X"11",X"65",X"FF",X"51",X"55",X"52",X"16",
		X"66",X"66",X"64",X"45",X"11",X"11",X"65",X"13",X"11",X"11",X"11",X"65",X"FF",X"55",X"33",X"32",
		X"11",X"11",X"11",X"11",X"15",X"11",X"11",X"65",X"11",X"21",X"11",X"11",X"65",X"FF",X"56",X"66",
		X"32",X"11",X"11",X"11",X"11",X"15",X"11",X"11",X"65",X"11",X"11",X"11",X"11",X"65",X"FF",X"51",
		X"11",X"63",X"11",X"11",X"11",X"11",X"14",X"55",X"55",X"55",X"51",X"11",X"11",X"11",X"65",X"FF",
		X"55",X"55",X"55",X"55",X"11",X"11",X"11",X"11",X"46",X"66",X"65",X"55",X"11",X"11",X"11",X"65",
		X"FF",X"56",X"66",X"66",X"45",X"51",X"11",X"11",X"11",X"11",X"65",X"53",X"33",X"35",X"51",X"11",
		X"65",X"FF",X"51",X"11",X"11",X"14",X"65",X"11",X"11",X"11",X"16",X"56",X"33",X"23",X"26",X"65",
		X"55",X"55",X"FF",X"51",X"11",X"11",X"11",X"65",X"11",X"11",X"11",X"16",X"51",X"13",X"32",X"12",
		X"16",X"66",X"65",X"FF",X"52",X"11",X"11",X"11",X"65",X"11",X"11",X"11",X"16",X"51",X"11",X"32",
		X"12",X"11",X"11",X"65",X"FF",X"53",X"21",X"11",X"11",X"65",X"11",X"11",X"11",X"16",X"51",X"12",
		X"13",X"11",X"11",X"16",X"65",X"FF",X"55",X"55",X"13",X"13",X"35",X"51",X"11",X"11",X"66",X"51",
		X"11",X"13",X"11",X"16",X"65",X"55",X"FF",X"11",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"11",X"FF",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"FF",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"10",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",
		X"11",X"16",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"64",X"11",X"10",X"11",X"66",X"66",
		X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"11",X"66",X"66",X"66",X"66",
		X"66",X"41",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"00",X"11",
		X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"FF",X"00",X"01",X"16",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"64",X"11",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"41",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"11",
		X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",
		X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"41",X"FF",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"41",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",
		X"00",X"11",X"16",X"66",X"66",X"66",X"64",X"11",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",
		X"41",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"FF",X"01",
		X"16",X"66",X"66",X"44",X"46",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"64",X"11",X"46",
		X"66",X"66",X"66",X"64",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",
		X"46",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"01",X"16",X"66",X"66",
		X"66",X"64",X"10",X"00",X"00",X"11",X"16",X"66",X"66",X"66",X"64",X"11",X"00",X"00",X"00",X"00",
		X"11",X"16",X"66",X"66",X"66",X"64",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"46",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"64",X"11",X"FF",X"01",X"15",X"55",X"54",X"11",X"14",
		X"55",X"55",X"55",X"44",X"44",X"45",X"55",X"55",X"54",X"11",X"14",X"55",X"55",X"55",X"41",X"11",
		X"55",X"54",X"44",X"45",X"55",X"55",X"54",X"44",X"45",X"55",X"41",X"14",X"55",X"55",X"55",X"44",
		X"44",X"44",X"44",X"45",X"55",X"41",X"00",X"01",X"15",X"55",X"55",X"55",X"54",X"10",X"00",X"00",
		X"01",X"11",X"55",X"55",X"55",X"41",X"10",X"00",X"00",X"00",X"00",X"01",X"11",X"55",X"55",X"55",
		X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"14",X"55",X"55",X"54",X"44",X"45",
		X"55",X"55",X"41",X"10",X"FF",X"11",X"55",X"55",X"41",X"11",X"11",X"55",X"55",X"55",X"41",X"11",
		X"14",X"55",X"55",X"55",X"41",X"11",X"55",X"55",X"55",X"41",X"11",X"55",X"41",X"11",X"15",X"55",
		X"55",X"54",X"11",X"14",X"55",X"41",X"11",X"55",X"55",X"55",X"41",X"11",X"11",X"11",X"14",X"55",
		X"41",X"00",X"01",X"15",X"55",X"55",X"55",X"54",X"10",X"00",X"00",X"00",X"11",X"55",X"55",X"55",
		X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"54",X"11",X"15",X"55",X"55",X"41",X"00",X"FF",
		X"11",X"55",X"55",X"41",X"11",X"11",X"55",X"55",X"55",X"41",X"00",X"11",X"15",X"55",X"55",X"41",
		X"11",X"55",X"55",X"55",X"41",X"01",X"55",X"11",X"01",X"15",X"55",X"55",X"54",X"10",X"11",X"55",
		X"41",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"11",X"55",X"41",X"00",X"11",X"15",X"55",
		X"55",X"55",X"54",X"11",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"55",X"55",X"54",X"10",X"15",X"55",X"55",X"41",X"00",X"FF",X"11",X"33",X"33",X"41",X"11",
		X"11",X"33",X"33",X"33",X"41",X"00",X"01",X"13",X"33",X"33",X"41",X"11",X"33",X"33",X"33",X"41",
		X"01",X"44",X"10",X"01",X"13",X"33",X"33",X"34",X"10",X"01",X"44",X"41",X"11",X"33",X"33",X"33",
		X"41",X"00",X"00",X"00",X"01",X"44",X"41",X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"41",X"00",
		X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"34",X"10",
		X"13",X"33",X"33",X"41",X"00",X"FF",X"11",X"33",X"33",X"41",X"11",X"11",X"33",X"33",X"33",X"41",
		X"00",X"01",X"13",X"33",X"33",X"41",X"11",X"33",X"33",X"33",X"41",X"01",X"11",X"10",X"01",X"13",
		X"33",X"33",X"34",X"10",X"01",X"11",X"11",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"01",
		X"11",X"11",X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"11",X"33",X"33",
		X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"34",X"10",X"13",X"33",X"33",X"41",X"00",
		X"FF",X"11",X"33",X"33",X"34",X"11",X"11",X"33",X"33",X"33",X"41",X"00",X"01",X"13",X"33",X"33",
		X"41",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"01",X"13",X"33",X"33",X"34",X"10",X"00",
		X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"11",X"33",
		X"33",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"33",X"33",X"34",X"10",X"13",X"33",X"33",X"41",X"00",X"FF",X"11",X"33",X"33",X"33",
		X"41",X"11",X"33",X"33",X"33",X"41",X"00",X"01",X"13",X"33",X"33",X"41",X"11",X"33",X"33",X"33",
		X"41",X"00",X"00",X"00",X"01",X"13",X"33",X"33",X"34",X"10",X"00",X"00",X"00",X"11",X"33",X"33",
		X"33",X"41",X"01",X"11",X"11",X"10",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"41",
		X"10",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",
		X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"34",
		X"10",X"13",X"33",X"33",X"41",X"00",X"FF",X"11",X"22",X"22",X"22",X"41",X"11",X"22",X"22",X"22",
		X"41",X"00",X"01",X"12",X"22",X"22",X"41",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"01",
		X"12",X"22",X"22",X"24",X"10",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"11",X"12",X"24",
		X"10",X"00",X"00",X"01",X"12",X"22",X"22",X"44",X"22",X"22",X"24",X"10",X"00",X"00",X"11",X"22",
		X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"24",X"10",X"12",X"22",X"22",X"41",
		X"00",X"FF",X"11",X"22",X"22",X"22",X"41",X"11",X"22",X"22",X"22",X"41",X"00",X"11",X"22",X"22",
		X"22",X"41",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"01",X"12",X"22",X"22",X"24",X"10",
		X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"11",X"22",X"24",X"10",X"00",X"00",X"01",X"12",
		X"22",X"22",X"41",X"22",X"22",X"24",X"10",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"22",X"22",X"24",X"10",X"12",X"22",X"22",X"41",X"00",X"FF",X"11",X"22",X"22",
		X"24",X"11",X"11",X"22",X"22",X"22",X"41",X"11",X"11",X"22",X"22",X"24",X"11",X"11",X"22",X"22",
		X"22",X"41",X"00",X"00",X"00",X"01",X"12",X"22",X"22",X"24",X"10",X"00",X"00",X"00",X"11",X"22",
		X"22",X"22",X"22",X"22",X"22",X"24",X"10",X"00",X"00",X"01",X"12",X"22",X"22",X"41",X"22",X"22",
		X"24",X"10",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",
		X"24",X"10",X"12",X"22",X"22",X"41",X"00",X"FF",X"11",X"42",X"22",X"41",X"10",X"11",X"22",X"22",
		X"22",X"41",X"11",X"12",X"22",X"22",X"24",X"10",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",
		X"01",X"12",X"22",X"22",X"24",X"10",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"22",X"22",X"22",
		X"24",X"10",X"00",X"00",X"01",X"12",X"22",X"22",X"41",X"22",X"22",X"24",X"11",X"00",X"00",X"11",
		X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"24",X"10",X"12",X"22",X"22",
		X"41",X"00",X"FF",X"01",X"14",X"44",X"11",X"00",X"11",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"41",X"10",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"01",X"12",X"22",X"22",X"24",
		X"10",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"22",X"22",X"22",X"24",X"10",X"00",X"00",X"11",
		X"22",X"22",X"24",X"11",X"12",X"22",X"22",X"41",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"22",X"22",X"24",X"10",X"12",X"22",X"22",X"41",X"00",X"FF",X"00",X"11",
		X"11",X"00",X"00",X"11",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"24",X"11",X"00",X"11",X"22",
		X"22",X"22",X"41",X"00",X"00",X"00",X"01",X"12",X"22",X"22",X"24",X"10",X"00",X"00",X"00",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"24",X"10",X"00",X"00",X"11",X"22",X"22",X"24",X"11",X"12",
		X"22",X"22",X"41",X"00",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",
		X"22",X"24",X"10",X"12",X"22",X"22",X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"41",X"10",X"00",X"11",X"22",X"22",X"22",X"41",X"00",X"00",
		X"00",X"01",X"12",X"22",X"22",X"24",X"10",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"44",X"44",
		X"22",X"24",X"10",X"00",X"00",X"11",X"22",X"22",X"24",X"11",X"12",X"22",X"22",X"41",X"00",X"00",
		X"11",X"22",X"22",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"24",X"10",X"12",X"22",
		X"22",X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"11",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"01",X"13",X"33",X"33",
		X"34",X"10",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"11",X"43",X"34",X"10",X"00",X"00",
		X"11",X"33",X"33",X"34",X"11",X"13",X"33",X"33",X"41",X"10",X"00",X"11",X"33",X"33",X"33",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"34",X"10",X"13",X"33",X"33",X"41",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"44",X"44",X"44",X"11",X"10",X"00",X"00",X"11",
		X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"01",X"13",X"33",X"33",X"34",X"10",X"00",X"00",X"00",
		X"11",X"33",X"33",X"33",X"41",X"01",X"14",X"44",X"10",X"00",X"01",X"13",X"33",X"33",X"41",X"11",
		X"11",X"33",X"33",X"34",X"10",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"33",X"33",X"34",X"10",X"13",X"33",X"33",X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",
		X"33",X"33",X"33",X"41",X"11",X"11",X"10",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",
		X"00",X"00",X"01",X"13",X"33",X"33",X"34",X"10",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",
		X"00",X"11",X"11",X"10",X"00",X"01",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"34",X"10",
		X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",
		X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"34",X"10",X"13",
		X"33",X"33",X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"01",X"13",X"33",
		X"33",X"34",X"10",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"00",X"00",
		X"01",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"34",X"10",X"00",X"11",X"33",X"33",X"33",
		X"41",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"33",X"33",X"33",X"41",X"00",X"00",X"00",X"01",
		X"11",X"11",X"00",X"00",X"00",X"11",X"33",X"33",X"34",X"10",X"13",X"33",X"33",X"41",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"01",X"15",X"55",X"55",X"54",X"10",X"00",X"00",
		X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",X"00",X"01",X"15",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"54",X"11",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"01",
		X"11",X"11",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",
		X"11",X"55",X"55",X"54",X"10",X"15",X"55",X"55",X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",
		X"00",X"00",X"00",X"01",X"15",X"55",X"55",X"54",X"10",X"00",X"00",X"00",X"11",X"55",X"55",X"55",
		X"41",X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"41",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"11",X"55",X"41",X"11",X"55",X"55",
		X"55",X"41",X"00",X"00",X"00",X"11",X"55",X"41",X"00",X"00",X"00",X"11",X"55",X"55",X"54",X"10",
		X"15",X"55",X"55",X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"01",X"15",
		X"55",X"55",X"54",X"10",X"00",X"00",X"00",X"11",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",
		X"00",X"11",X"55",X"55",X"54",X"44",X"44",X"44",X"45",X"55",X"55",X"41",X"01",X"11",X"55",X"55",
		X"55",X"41",X"11",X"11",X"11",X"11",X"55",X"41",X"11",X"55",X"55",X"55",X"41",X"11",X"11",X"11",
		X"11",X"55",X"41",X"00",X"00",X"00",X"11",X"55",X"55",X"54",X"11",X"15",X"55",X"55",X"41",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"41",X"10",X"00",X"00",X"00",X"00",
		X"00",X"11",X"66",X"66",X"66",X"41",X"10",X"00",X"00",X"01",X"16",X"66",X"66",X"64",X"11",X"00",
		X"00",X"00",X"11",X"66",X"66",X"66",X"41",X"10",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"64",
		X"11",X"11",X"11",X"16",X"66",X"66",X"41",X"11",X"16",X"66",X"66",X"66",X"41",X"11",X"11",X"11",
		X"16",X"66",X"41",X"16",X"66",X"66",X"66",X"41",X"11",X"11",X"11",X"16",X"66",X"41",X"00",X"00",
		X"01",X"11",X"66",X"66",X"64",X"11",X"16",X"66",X"66",X"41",X"10",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"16",X"66",X"66",X"66",X"64",X"11",X"00",X"00",X"00",X"00",X"01",X"16",X"66",X"66",X"66",
		X"64",X"11",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"41",X"10",X"00",X"01",X"16",X"66",X"66",
		X"66",X"64",X"11",X"00",X"00",X"00",X"01",X"16",X"66",X"66",X"64",X"11",X"00",X"01",X"16",X"66",
		X"66",X"64",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"11",X"16",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"64",X"11",X"FF",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",
		X"66",X"41",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"01",X"16",
		X"66",X"66",X"66",X"66",X"64",X"10",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",
		X"00",X"11",X"66",X"66",X"66",X"66",X"41",X"00",X"01",X"66",X"66",X"66",X"66",X"41",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"41",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"41",X"FF",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",
		X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"01",X"16",X"66",X"66",X"66",X"66",X"64",
		X"10",X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"11",X"66",X"66",X"66",
		X"66",X"41",X"00",X"01",X"66",X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"00",
		X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"FF",X"00",X"00",X"00",
		X"00",X"11",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"00",X"11",X"66",X"66",X"66",
		X"66",X"66",X"41",X"00",X"01",X"16",X"66",X"66",X"66",X"66",X"64",X"10",X"00",X"11",X"66",X"66",
		X"66",X"66",X"66",X"41",X"00",X"00",X"00",X"11",X"66",X"66",X"66",X"66",X"41",X"00",X"01",X"66",
		X"66",X"66",X"66",X"41",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"00",X"00",X"11",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"41",X"FF",X"00",X"00",X"00",X"00",X"11",X"44",X"44",X"44",
		X"44",X"44",X"41",X"00",X"00",X"00",X"00",X"11",X"44",X"44",X"44",X"44",X"44",X"41",X"00",X"01",
		X"14",X"44",X"44",X"44",X"44",X"44",X"10",X"00",X"11",X"44",X"44",X"44",X"44",X"44",X"41",X"00",
		X"00",X"00",X"11",X"44",X"44",X"44",X"44",X"41",X"00",X"01",X"44",X"44",X"44",X"44",X"41",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"41",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"41",X"00",X"00",X"11",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"41",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"11",X"11",X"11",X"11",X"11",
		X"11",X"10",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"11",X"11",X"11",
		X"11",X"11",X"11",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",
		X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"01",X"11",X"01",X"10",X"11",X"00",X"00",X"FF",
		X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"FF",X"00",X"01",X"11",X"11",X"11",X"11",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"77",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"25",X"76",X"75",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",
		X"66",X"65",X"52",X"00",X"00",X"FF",X"00",X"02",X"77",X"77",X"77",X"72",X"00",X"00",X"FF",X"02",
		X"66",X"66",X"66",X"66",X"66",X"62",X"00",X"FF",X"02",X"E2",X"41",X"23",X"21",X"42",X"E2",X"00",
		X"FF",X"21",X"12",X"44",X"37",X"34",X"42",X"11",X"20",X"FF",X"21",X"11",X"21",X"D1",X"D1",X"21",
		X"1A",X"20",X"FF",X"02",X"11",X"21",X"D1",X"D1",X"2A",X"A2",X"00",X"FF",X"23",X"77",X"53",X"33",
		X"33",X"57",X"73",X"20",X"FF",X"24",X"56",X"57",X"D7",X"D7",X"56",X"54",X"20",X"FF",X"02",X"22",
		X"67",X"15",X"D7",X"62",X"22",X"00",X"FF",X"00",X"05",X"65",X"DD",X"15",X"65",X"00",X"00",X"FF",
		X"00",X"05",X"65",X"81",X"D5",X"65",X"00",X"00",X"FF",X"02",X"20",X"59",X"B9",X"B9",X"50",X"22",
		X"00",X"FF",X"02",X"12",X"89",X"98",X"99",X"82",X"12",X"00",X"FF",X"02",X"92",X"98",X"99",X"98",
		X"92",X"92",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",X"20",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"01",X"11",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"FF",X"00",X"01",X"11",X"10",X"11",X"01",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"11",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"27",X"76",X"77",X"20",X"00",X"00",X"FF",X"00",X"00",X"25",X"76",
		X"75",X"20",X"00",X"00",X"FF",X"00",X"02",X"55",X"66",X"65",X"52",X"00",X"00",X"FF",X"00",X"02",
		X"77",X"77",X"77",X"72",X"00",X"00",X"FF",X"02",X"66",X"66",X"66",X"66",X"66",X"62",X"00",X"FF",
		X"02",X"E2",X"42",X"13",X"12",X"42",X"E2",X"00",X"FF",X"00",X"02",X"44",X"37",X"34",X"42",X"00",
		X"00",X"FF",X"02",X"21",X"21",X"D1",X"D1",X"21",X"22",X"00",X"FF",X"21",X"11",X"21",X"D1",X"D1",
		X"2A",X"11",X"20",X"FF",X"23",X"77",X"53",X"33",X"33",X"57",X"73",X"20",X"FF",X"24",X"56",X"57",
		X"D7",X"D7",X"56",X"54",X"20",X"FF",X"02",X"22",X"67",X"15",X"D7",X"62",X"22",X"00",X"FF",X"00",
		X"05",X"65",X"DD",X"15",X"65",X"00",X"00",X"FF",X"00",X"05",X"65",X"81",X"D5",X"65",X"00",X"00",
		X"FF",X"02",X"20",X"59",X"B9",X"B9",X"50",X"22",X"00",X"FF",X"02",X"12",X"89",X"98",X"99",X"82",
		X"12",X"00",X"FF",X"02",X"92",X"98",X"99",X"98",X"92",X"92",X"00",X"FF",X"00",X"22",X"22",X"22",
		X"22",X"22",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"10",X"00",X"FF",X"01",X"13",X"41",X"10",X"FF",X"13",X"37",X"84",X"41",X"FF",X"13",
		X"48",X"84",X"61",X"FF",X"12",X"44",X"44",X"61",X"FF",X"12",X"44",X"84",X"61",X"FF",X"13",X"47",
		X"44",X"61",X"FF",X"01",X"44",X"46",X"10",X"FF",X"00",X"13",X"51",X"00",X"FF",X"00",X"13",X"51",
		X"00",X"FF",X"00",X"12",X"51",X"10",X"FF",X"00",X"14",X"55",X"61",X"FF",X"00",X"14",X"56",X"10",
		X"FF",X"00",X"15",X"61",X"00",X"FF",X"00",X"15",X"61",X"00",X"FF",X"00",X"01",X"10",X"00",X"FF",
		X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"01",X"2A",X"22",X"2A",X"10",X"00",X"FF",
		X"00",X"01",X"22",X"2A",X"AA",X"10",X"00",X"FF",X"00",X"00",X"19",X"B9",X"91",X"00",X"00",X"FF",
		X"00",X"01",X"19",X"BB",X"91",X"10",X"00",X"FF",X"00",X"12",X"AA",X"2A",X"2A",X"A1",X"00",X"FF",
		X"01",X"2A",X"22",X"2A",X"22",X"2A",X"10",X"FF",X"01",X"22",X"22",X"12",X"12",X"22",X"10",X"FF",
		X"1A",X"22",X"11",X"11",X"11",X"1A",X"21",X"FF",X"1A",X"22",X"12",X"12",X"12",X"2A",X"21",X"FF",
		X"12",X"A2",X"11",X"11",X"11",X"12",X"21",X"FF",X"12",X"22",X"22",X"12",X"12",X"12",X"A1",X"FF",
		X"12",X"A2",X"11",X"11",X"11",X"12",X"A1",X"FF",X"01",X"22",X"22",X"12",X"12",X"2A",X"10",X"FF",
		X"00",X"11",X"A2",X"22",X"2A",X"11",X"00",X"FF",X"00",X"01",X"11",X"11",X"11",X"10",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",
		X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"01",X"44",X"10",X"01",X"44",X"10",X"00",X"FF",X"00",
		X"15",X"44",X"51",X"15",X"44",X"51",X"00",X"FF",X"00",X"15",X"44",X"51",X"15",X"44",X"51",X"00",
		X"FF",X"00",X"15",X"44",X"51",X"15",X"45",X"51",X"00",X"FF",X"01",X"45",X"66",X"55",X"45",X"66",
		X"54",X"10",X"FF",X"15",X"46",X"66",X"65",X"46",X"66",X"64",X"51",X"FF",X"15",X"46",X"66",X"65",
		X"46",X"66",X"64",X"51",X"FF",X"15",X"47",X"77",X"75",X"47",X"77",X"74",X"51",X"FF",X"15",X"66",
		X"57",X"56",X"65",X"75",X"66",X"51",X"FF",X"16",X"66",X"67",X"66",X"66",X"76",X"66",X"61",X"FF",
		X"16",X"66",X"67",X"66",X"66",X"76",X"66",X"61",X"FF",X"17",X"77",X"77",X"77",X"77",X"77",X"77",
		X"71",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"FF",X"00",X"00",X"22",
		X"00",X"20",X"02",X"20",X"00",X"FF",X"00",X"00",X"02",X"00",X"00",X"02",X"00",X"00",X"FF",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"FF",X"02",X"20",X"11",X"00",X"00",X"11",X"02",X"20",
		X"FF",X"00",X"01",X"22",X"10",X"01",X"22",X"10",X"00",X"FF",X"00",X"14",X"22",X"41",X"14",X"22",
		X"41",X"00",X"FF",X"00",X"14",X"22",X"41",X"14",X"22",X"41",X"00",X"FF",X"00",X"14",X"22",X"41",
		X"14",X"22",X"41",X"00",X"FF",X"01",X"24",X"66",X"44",X"24",X"66",X"42",X"10",X"FF",X"14",X"26",
		X"66",X"64",X"26",X"66",X"62",X"41",X"FF",X"14",X"26",X"66",X"64",X"26",X"66",X"62",X"41",X"FF",
		X"14",X"27",X"77",X"74",X"27",X"77",X"72",X"41",X"FF",X"14",X"66",X"47",X"46",X"64",X"74",X"66",
		X"41",X"FF",X"16",X"66",X"67",X"66",X"66",X"76",X"66",X"61",X"FF",X"16",X"66",X"67",X"66",X"66",
		X"76",X"66",X"61",X"FF",X"17",X"77",X"77",X"77",X"77",X"77",X"77",X"71",X"FF",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"09",X"2A",X"90",X"00",X"00",X"FF",X"09",X"90",X"92",X"ED",X"A9",X"09",X"90",X"FF",X"9A",X"B9",
		X"92",X"ED",X"A9",X"92",X"29",X"FF",X"92",X"AB",X"AE",X"DD",X"AB",X"BE",X"A9",X"FF",X"92",X"AB",
		X"AD",X"DA",X"BB",X"ED",X"A9",X"FF",X"9D",X"2A",X"BD",X"AA",X"9E",X"DA",X"90",X"FF",X"09",X"DA",
		X"BA",X"BA",X"BA",X"D9",X"00",X"FF",X"09",X"BD",X"AB",X"2B",X"BD",X"A9",X"99",X"FF",X"09",X"AB",
		X"B2",X"EA",X"BA",X"B2",X"29",X"FF",X"9B",X"BA",X"9E",X"AB",X"AB",X"2D",X"A9",X"FF",X"92",X"EB",
		X"AE",X"AB",X"9D",X"DA",X"B9",X"FF",X"9A",X"DE",X"BA",X"AB",X"DD",X"A9",X"90",X"FF",X"09",X"AA",
		X"DA",X"BA",X"DA",X"B9",X"00",X"FF",X"00",X"9B",X"AB",X"9B",X"BB",X"90",X"00",X"FF",X"00",X"09",
		X"99",X"09",X"99",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"66",X"99",X"96",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"66",X"99",X"A8",X"96",X"00",X"00",X"FF",X"00",X"00",X"00",X"66",X"99",X"A1",X"88",X"A6",X"00",
		X"00",X"FF",X"00",X"00",X"66",X"99",X"A1",X"11",X"88",X"A6",X"00",X"00",X"FF",X"00",X"66",X"99",
		X"A1",X"11",X"15",X"88",X"A6",X"00",X"00",X"FF",X"06",X"A9",X"91",X"11",X"15",X"55",X"88",X"A6",
		X"00",X"00",X"FF",X"6A",X"A3",X"91",X"15",X"55",X"55",X"58",X"A6",X"00",X"00",X"FF",X"6A",X"34",
		X"A5",X"55",X"55",X"55",X"5A",X"A6",X"60",X"00",X"FF",X"6A",X"44",X"A5",X"55",X"55",X"52",X"D2",
		X"89",X"96",X"60",X"FF",X"6A",X"44",X"A5",X"55",X"52",X"E2",X"EC",X"22",X"C9",X"96",X"FF",X"6B",
		X"A4",X"A5",X"5A",X"2D",X"2C",X"2D",X"E2",X"99",X"A6",X"FF",X"06",X"BA",X"AA",X"A2",X"2E",X"2E",
		X"2C",X"99",X"3A",X"A6",X"FF",X"00",X"6B",X"A9",X"DE",X"22",X"CD",X"99",X"AA",X"33",X"A6",X"FF",
		X"00",X"06",X"AA",X"99",X"C2",X"99",X"3A",X"6A",X"34",X"A6",X"FF",X"00",X"06",X"A3",X"3A",X"99",
		X"AA",X"3A",X"6A",X"44",X"A6",X"FF",X"00",X"06",X"A3",X"43",X"A9",X"A4",X"3A",X"A4",X"44",X"A6",
		X"FF",X"00",X"06",X"A3",X"44",X"49",X"A4",X"44",X"A4",X"44",X"A6",X"FF",X"00",X"06",X"A3",X"44",
		X"49",X"A4",X"44",X"A4",X"AA",X"A6",X"FF",X"00",X"06",X"AA",X"44",X"49",X"A4",X"44",X"AA",X"A6",
		X"60",X"FF",X"00",X"06",X"6A",X"AA",X"49",X"A4",X"AA",X"A6",X"60",X"00",X"FF",X"00",X"00",X"06",
		X"6A",X"A9",X"AA",X"A6",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"69",X"A6",X"60",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",
		X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"12",X"22",X"22",X"2D",X"10",X"00",X"FF",X"01",X"EA",
		X"2E",X"EE",X"DA",X"B1",X"00",X"FF",X"1A",X"DD",X"A2",X"ED",X"AA",X"AB",X"10",X"FF",X"12",X"EE",
		X"EA",X"AA",X"BB",X"BB",X"10",X"FF",X"01",X"AD",X"DE",X"EA",X"BA",X"B1",X"00",X"FF",X"00",X"1A",
		X"DA",X"2B",X"AB",X"10",X"00",X"FF",X"00",X"01",X"BA",X"EA",X"91",X"00",X"00",X"FF",X"01",X"88",
		X"1B",X"E9",X"18",X"81",X"00",X"FF",X"01",X"8C",X"C1",X"B1",X"CC",X"81",X"00",X"FF",X"18",X"88",
		X"1C",X"CC",X"1C",X"C8",X"10",X"FF",X"18",X"81",X"CC",X"CC",X"C1",X"88",X"10",X"FF",X"18",X"8C",
		X"88",X"88",X"8C",X"88",X"10",X"FF",X"1C",X"CC",X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",
		X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"01",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"12",
		X"22",X"22",X"2E",X"10",X"00",X"FF",X"01",X"EA",X"2E",X"EE",X"EA",X"B1",X"00",X"FF",X"1A",X"EE",
		X"A2",X"EE",X"AA",X"AB",X"10",X"FF",X"12",X"EE",X"EA",X"AA",X"BB",X"BB",X"10",X"FF",X"01",X"AE",
		X"EE",X"EA",X"BA",X"B1",X"00",X"FF",X"00",X"1A",X"EA",X"2B",X"AB",X"10",X"00",X"FF",X"00",X"01",
		X"BA",X"EA",X"91",X"00",X"00",X"FF",X"01",X"88",X"1B",X"E9",X"18",X"81",X"00",X"FF",X"01",X"8C",
		X"C1",X"B1",X"CC",X"81",X"00",X"FF",X"18",X"88",X"1C",X"CC",X"1C",X"C8",X"10",X"FF",X"18",X"81",
		X"CC",X"CC",X"C1",X"88",X"10",X"FF",X"18",X"8C",X"88",X"88",X"8C",X"88",X"10",X"FF",X"1C",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"01",
		X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"12",X"22",X"22",X"22",X"10",X"00",X"FF",X"01",X"EE",
		X"2E",X"EE",X"2E",X"B1",X"00",X"FF",X"1E",X"22",X"E2",X"E2",X"EE",X"EB",X"10",X"FF",X"12",X"EE",
		X"EE",X"EE",X"BB",X"BB",X"10",X"FF",X"01",X"E2",X"2E",X"EE",X"BE",X"B1",X"00",X"FF",X"00",X"1E",
		X"2E",X"2B",X"EB",X"10",X"00",X"FF",X"00",X"01",X"BE",X"EE",X"91",X"00",X"00",X"FF",X"01",X"88",
		X"1B",X"E9",X"18",X"81",X"00",X"FF",X"01",X"8C",X"C1",X"B1",X"CC",X"81",X"00",X"FF",X"18",X"88",
		X"1C",X"CC",X"1C",X"C8",X"10",X"FF",X"18",X"81",X"CC",X"CC",X"C1",X"88",X"10",X"FF",X"18",X"8C",
		X"88",X"88",X"8C",X"88",X"10",X"FF",X"1C",X"CC",X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",
		X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"01",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"12",
		X"22",X"22",X"24",X"10",X"00",X"FF",X"01",X"EA",X"2E",X"EE",X"4A",X"B1",X"00",X"FF",X"1A",X"44",
		X"A2",X"E4",X"AA",X"AB",X"10",X"FF",X"12",X"EE",X"EA",X"AA",X"BB",X"BB",X"10",X"FF",X"01",X"A4",
		X"4E",X"EA",X"BA",X"B1",X"00",X"FF",X"00",X"1A",X"4A",X"2B",X"AB",X"10",X"00",X"FF",X"00",X"01",
		X"BA",X"EA",X"91",X"00",X"00",X"FF",X"01",X"88",X"1B",X"E9",X"18",X"81",X"00",X"FF",X"01",X"8C",
		X"C1",X"B1",X"CC",X"81",X"00",X"FF",X"18",X"88",X"1C",X"CC",X"1C",X"C8",X"10",X"FF",X"18",X"81",
		X"CC",X"CC",X"C1",X"88",X"10",X"FF",X"18",X"8C",X"88",X"88",X"8C",X"88",X"10",X"FF",X"1C",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"00",
		X"01",X"11",X"00",X"00",X"00",X"FF",X"00",X"01",X"1A",X"AB",X"11",X"00",X"00",X"FF",X"00",X"1A",
		X"AA",X"AA",X"BB",X"10",X"00",X"FF",X"01",X"AA",X"EE",X"DA",X"AB",X"B1",X"00",X"FF",X"01",X"AE",
		X"2E",X"ED",X"AA",X"91",X"00",X"FF",X"1A",X"AE",X"E2",X"ED",X"AA",X"B9",X"10",X"FF",X"1B",X"AA",
		X"EE",X"DD",X"AA",X"B9",X"10",X"FF",X"01",X"BA",X"DD",X"DA",X"AB",X"91",X"00",X"FF",X"01",X"BB",
		X"AA",X"AA",X"BB",X"91",X"00",X"FF",X"00",X"19",X"BB",X"BB",X"99",X"10",X"00",X"FF",X"01",X"CC",
		X"19",X"99",X"11",X"C1",X"00",X"FF",X"01",X"88",X"C1",X"11",X"CC",X"81",X"00",X"FF",X"18",X"81",
		X"1C",X"CC",X"88",X"88",X"10",X"FF",X"18",X"88",X"88",X"88",X"88",X"88",X"10",X"FF",X"1C",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"00",
		X"01",X"11",X"00",X"00",X"00",X"FF",X"00",X"01",X"1D",X"DA",X"11",X"00",X"00",X"FF",X"00",X"1D",
		X"DD",X"DD",X"AA",X"10",X"00",X"FF",X"01",X"DD",X"22",X"ED",X"DA",X"A1",X"00",X"FF",X"01",X"D2",
		X"22",X"2E",X"DD",X"B1",X"00",X"FF",X"1D",X"D2",X"22",X"2E",X"DD",X"AB",X"10",X"FF",X"1A",X"DD",
		X"22",X"EE",X"DD",X"AB",X"10",X"FF",X"01",X"AD",X"EE",X"ED",X"DA",X"B1",X"00",X"FF",X"01",X"AA",
		X"DD",X"DD",X"AA",X"B1",X"00",X"FF",X"00",X"1B",X"AA",X"AA",X"BB",X"10",X"00",X"FF",X"01",X"CC",
		X"1B",X"BB",X"11",X"C1",X"00",X"FF",X"01",X"88",X"C1",X"11",X"CC",X"81",X"00",X"FF",X"18",X"81",
		X"1C",X"CC",X"88",X"88",X"10",X"FF",X"18",X"88",X"88",X"88",X"88",X"88",X"10",X"FF",X"1C",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"00",
		X"01",X"11",X"00",X"00",X"00",X"FF",X"00",X"01",X"1E",X"ED",X"11",X"00",X"00",X"FF",X"00",X"1E",
		X"EE",X"EE",X"DD",X"10",X"00",X"FF",X"01",X"EE",X"22",X"2E",X"ED",X"D1",X"00",X"FF",X"01",X"E2",
		X"22",X"22",X"EE",X"A1",X"00",X"FF",X"1E",X"E2",X"22",X"22",X"EE",X"DA",X"10",X"FF",X"1D",X"EE",
		X"22",X"22",X"EE",X"DA",X"10",X"FF",X"01",X"DE",X"22",X"2E",X"ED",X"A1",X"00",X"FF",X"01",X"DD",
		X"EE",X"EE",X"DD",X"A1",X"00",X"FF",X"00",X"1A",X"DD",X"DD",X"AA",X"10",X"00",X"FF",X"01",X"CC",
		X"1A",X"AA",X"11",X"C1",X"00",X"FF",X"01",X"88",X"C1",X"11",X"CC",X"81",X"00",X"FF",X"18",X"81",
		X"1C",X"CC",X"88",X"88",X"10",X"FF",X"18",X"88",X"88",X"88",X"88",X"88",X"10",X"FF",X"1C",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"00",
		X"01",X"11",X"00",X"00",X"00",X"FF",X"00",X"01",X"12",X"2E",X"11",X"00",X"00",X"FF",X"00",X"12",
		X"22",X"22",X"EE",X"10",X"00",X"FF",X"01",X"22",X"22",X"22",X"2E",X"E1",X"00",X"FF",X"01",X"22",
		X"22",X"22",X"22",X"D1",X"00",X"FF",X"12",X"22",X"22",X"22",X"22",X"ED",X"10",X"FF",X"1E",X"22",
		X"22",X"22",X"22",X"ED",X"10",X"FF",X"01",X"E2",X"22",X"22",X"2E",X"D1",X"00",X"FF",X"01",X"EE",
		X"22",X"22",X"EE",X"D1",X"00",X"FF",X"00",X"1D",X"EE",X"EE",X"DD",X"10",X"00",X"FF",X"01",X"CC",
		X"1D",X"DD",X"11",X"C1",X"00",X"FF",X"01",X"88",X"C1",X"11",X"CC",X"81",X"00",X"FF",X"18",X"81",
		X"1C",X"CC",X"88",X"88",X"10",X"FF",X"18",X"88",X"88",X"88",X"88",X"88",X"10",X"FF",X"1C",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"10",X"FF",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"02",X"00",X"FF",X"00",X"00",X"00",X"00",X"15",X"A5",
		X"10",X"00",X"00",X"02",X"00",X"FF",X"02",X"00",X"00",X"11",X"5B",X"89",X"51",X"10",X"00",X"02",
		X"00",X"FF",X"00",X"00",X"01",X"23",X"35",X"95",X"34",X"41",X"00",X"02",X"00",X"FF",X"00",X"00",
		X"12",X"46",X"C2",X"34",X"C6",X"44",X"12",X"22",X"22",X"FF",X"00",X"01",X"36",X"C8",X"43",X"6C",
		X"8C",X"64",X"10",X"02",X"00",X"FF",X"00",X"01",X"4C",X"88",X"82",X"3C",X"88",X"C4",X"10",X"02",
		X"00",X"FF",X"00",X"01",X"6C",X"88",X"88",X"34",X"C8",X"C6",X"10",X"02",X"00",X"FF",X"00",X"01",
		X"6C",X"88",X"86",X"4C",X"88",X"C6",X"10",X"02",X"00",X"FF",X"00",X"01",X"6C",X"88",X"84",X"4C",
		X"88",X"C6",X"10",X"02",X"00",X"FF",X"00",X"00",X"16",X"C8",X"85",X"58",X"8C",X"61",X"00",X"02",
		X"00",X"FF",X"00",X"00",X"16",X"CC",X"C6",X"6C",X"CC",X"61",X"00",X"00",X"00",X"FF",X"00",X"01",
		X"65",X"54",X"43",X"24",X"45",X"56",X"10",X"00",X"00",X"FF",X"00",X"11",X"69",X"5B",X"4A",X"3B",
		X"49",X"56",X"11",X"00",X"00",X"FF",X"01",X"81",X"65",X"54",X"23",X"34",X"45",X"56",X"1C",X"10",
		X"00",X"FF",X"18",X"88",X"11",X"11",X"11",X"11",X"11",X"11",X"C8",X"C1",X"00",X"FF",X"18",X"88",
		X"C1",X"1C",X"CC",X"CC",X"C1",X"1C",X"88",X"C1",X"00",X"FF",X"18",X"8C",X"1C",X"88",X"88",X"88",
		X"2C",X"C1",X"C8",X"C1",X"00",X"FF",X"1C",X"88",X"88",X"88",X"88",X"82",X"22",X"CC",X"C8",X"C1",
		X"00",X"FF",X"1C",X"C8",X"88",X"8C",X"CC",X"CC",X"28",X"88",X"8C",X"C1",X"00",X"FF",X"01",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"2C",X"CC",X"CC",X"10",X"00",X"FF",X"00",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"00",X"00",X"00",X"15",X"A5",X"10",X"00",X"00",X"00",X"00",X"FF",X"22",X"20",
		X"00",X"11",X"5B",X"89",X"51",X"10",X"00",X"02",X"00",X"FF",X"02",X"00",X"01",X"23",X"35",X"95",
		X"34",X"41",X"00",X"02",X"00",X"FF",X"00",X"00",X"12",X"46",X"C2",X"34",X"C6",X"44",X"10",X"22",
		X"20",X"FF",X"00",X"01",X"36",X"C8",X"43",X"6C",X"8C",X"64",X"10",X"02",X"00",X"FF",X"00",X"01",
		X"4C",X"88",X"82",X"3C",X"88",X"C4",X"10",X"02",X"00",X"FF",X"00",X"01",X"6C",X"88",X"88",X"34",
		X"C8",X"C6",X"10",X"02",X"00",X"FF",X"00",X"01",X"6C",X"88",X"86",X"4C",X"88",X"C6",X"10",X"00",
		X"00",X"FF",X"00",X"01",X"6C",X"88",X"84",X"4C",X"88",X"C6",X"10",X"00",X"00",X"FF",X"00",X"00",
		X"16",X"C8",X"85",X"58",X"8C",X"61",X"00",X"00",X"00",X"FF",X"00",X"00",X"16",X"CC",X"C6",X"6C",
		X"CC",X"61",X"00",X"00",X"00",X"FF",X"00",X"01",X"65",X"54",X"43",X"24",X"45",X"56",X"10",X"00",
		X"00",X"FF",X"00",X"11",X"69",X"5B",X"4A",X"3B",X"49",X"56",X"11",X"00",X"00",X"FF",X"01",X"81",
		X"65",X"54",X"23",X"34",X"45",X"56",X"1C",X"10",X"00",X"FF",X"18",X"88",X"11",X"11",X"11",X"11",
		X"11",X"11",X"C8",X"C1",X"00",X"FF",X"18",X"88",X"C1",X"1C",X"CC",X"CC",X"21",X"1C",X"88",X"C1",
		X"00",X"FF",X"18",X"8C",X"1C",X"88",X"88",X"88",X"2C",X"C1",X"C8",X"C1",X"00",X"FF",X"1C",X"88",
		X"88",X"88",X"88",X"22",X"22",X"2C",X"C8",X"C1",X"00",X"FF",X"1C",X"C8",X"88",X"8C",X"CC",X"CC",
		X"28",X"88",X"8C",X"C1",X"00",X"FF",X"01",X"CC",X"CC",X"CC",X"CC",X"CC",X"2C",X"CC",X"CC",X"10",
		X"00",X"FF",X"00",X"11",X"11",X"11",X"11",X"11",X"21",X"11",X"11",X"00",X"00",X"FF",X"02",X"00",
		X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"00",X"00",X"00",X"15",X"A5",
		X"10",X"00",X"00",X"00",X"00",X"FF",X"22",X"20",X"00",X"11",X"5B",X"89",X"51",X"10",X"00",X"00",
		X"00",X"FF",X"02",X"00",X"01",X"23",X"35",X"95",X"34",X"41",X"00",X"00",X"00",X"FF",X"02",X"00",
		X"12",X"46",X"C2",X"34",X"C6",X"44",X"10",X"02",X"00",X"FF",X"02",X"01",X"36",X"C8",X"43",X"6C",
		X"8C",X"64",X"10",X"00",X"00",X"FF",X"00",X"01",X"4C",X"88",X"82",X"3C",X"88",X"C4",X"10",X"00",
		X"00",X"FF",X"00",X"01",X"6C",X"88",X"88",X"34",X"C8",X"C6",X"10",X"00",X"00",X"FF",X"00",X"01",
		X"6C",X"88",X"86",X"4C",X"88",X"C6",X"10",X"00",X"00",X"FF",X"00",X"01",X"6C",X"88",X"84",X"4C",
		X"88",X"C6",X"10",X"00",X"00",X"FF",X"00",X"00",X"16",X"C8",X"85",X"58",X"8C",X"61",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"16",X"CC",X"C6",X"6C",X"CC",X"61",X"00",X"00",X"00",X"FF",X"00",X"01",
		X"65",X"54",X"43",X"24",X"45",X"56",X"10",X"00",X"00",X"FF",X"00",X"11",X"69",X"5B",X"4A",X"3B",
		X"49",X"56",X"11",X"00",X"00",X"FF",X"01",X"81",X"65",X"54",X"23",X"34",X"45",X"56",X"1C",X"10",
		X"00",X"FF",X"18",X"88",X"11",X"11",X"11",X"11",X"11",X"11",X"C8",X"C1",X"00",X"FF",X"18",X"88",
		X"C1",X"1C",X"CC",X"CC",X"C1",X"1C",X"88",X"C1",X"00",X"FF",X"18",X"8C",X"1C",X"88",X"88",X"88",
		X"2C",X"C1",X"C8",X"C1",X"00",X"FF",X"1C",X"88",X"88",X"88",X"88",X"82",X"22",X"CC",X"C8",X"C1",
		X"00",X"FF",X"1C",X"C8",X"88",X"8C",X"CC",X"CC",X"28",X"88",X"8C",X"C1",X"00",X"FF",X"01",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"2C",X"CC",X"CC",X"10",X"00",X"FF",X"00",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"00",X"00",X"00",X"15",X"A5",X"10",X"00",X"00",X"00",X"00",X"FF",X"22",X"20",
		X"00",X"11",X"5B",X"89",X"51",X"10",X"00",X"02",X"00",X"FF",X"02",X"00",X"01",X"23",X"35",X"95",
		X"34",X"41",X"00",X"02",X"00",X"FF",X"00",X"00",X"12",X"46",X"C2",X"34",X"C6",X"44",X"10",X"22",
		X"20",X"FF",X"00",X"01",X"36",X"C8",X"43",X"6C",X"8C",X"64",X"10",X"02",X"00",X"FF",X"00",X"01",
		X"4C",X"88",X"82",X"3C",X"88",X"C4",X"10",X"02",X"00",X"FF",X"00",X"01",X"6C",X"88",X"88",X"34",
		X"C8",X"C6",X"10",X"02",X"00",X"FF",X"00",X"01",X"6C",X"88",X"86",X"4C",X"88",X"C6",X"10",X"00",
		X"00",X"FF",X"00",X"01",X"6C",X"88",X"84",X"4C",X"88",X"C6",X"10",X"00",X"00",X"FF",X"00",X"00",
		X"16",X"C8",X"85",X"58",X"8C",X"61",X"00",X"00",X"00",X"FF",X"00",X"00",X"16",X"CC",X"C6",X"6C",
		X"CC",X"61",X"00",X"00",X"00",X"FF",X"00",X"01",X"65",X"54",X"43",X"24",X"45",X"56",X"10",X"00",
		X"00",X"FF",X"00",X"11",X"69",X"5B",X"4A",X"3B",X"49",X"56",X"11",X"00",X"00",X"FF",X"01",X"81",
		X"65",X"54",X"23",X"34",X"45",X"56",X"1C",X"10",X"00",X"FF",X"18",X"88",X"11",X"11",X"11",X"11",
		X"11",X"11",X"C8",X"C1",X"00",X"FF",X"18",X"88",X"C1",X"1C",X"CC",X"CC",X"C1",X"1C",X"88",X"C1",
		X"00",X"FF",X"18",X"8C",X"1C",X"88",X"88",X"88",X"CC",X"C1",X"C8",X"C1",X"00",X"FF",X"1C",X"88",
		X"88",X"88",X"88",X"88",X"28",X"CC",X"C8",X"C1",X"00",X"FF",X"1C",X"C8",X"88",X"8C",X"CC",X"CC",
		X"88",X"88",X"8C",X"C1",X"00",X"FF",X"01",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"10",
		X"00",X"FF",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"FF",
		X"00",X"44",X"44",X"00",X"00",X"44",X"42",X"E4",X"30",X"00",X"FF",X"04",X"41",X"54",X"44",X"44",
		X"44",X"28",X"2E",X"44",X"00",X"FF",X"44",X"45",X"54",X"45",X"54",X"44",X"42",X"D4",X"44",X"00",
		X"FF",X"31",X"11",X"44",X"41",X"11",X"11",X"44",X"44",X"55",X"30",X"FF",X"16",X"65",X"11",X"16",
		X"66",X"66",X"11",X"14",X"45",X"40",X"FF",X"55",X"55",X"66",X"65",X"55",X"55",X"66",X"64",X"44",
		X"3A",X"FF",X"0A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"4A",X"A0",X"FF",X"90",X"A0",X"A0",
		X"29",X"0A",X"A0",X"A0",X"90",X"A0",X"02",X"FF",X"00",X"02",X"00",X"A0",X"A0",X"A9",X"0A",X"02",
		X"09",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"04",X"55",X"13",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"04",X"34",X"44",X"44",X"43",X"04",X"44",X"44",X"00",X"00",X"FF",
		X"00",X"73",X"33",X"54",X"44",X"44",X"42",X"E4",X"30",X"00",X"FF",X"00",X"00",X"78",X"33",X"34",
		X"44",X"21",X"2E",X"44",X"00",X"FF",X"00",X"00",X"00",X"08",X"84",X"44",X"42",X"D4",X"44",X"00",
		X"FF",X"00",X"82",X"88",X"82",X"87",X"11",X"44",X"44",X"55",X"30",X"FF",X"46",X"65",X"82",X"86",
		X"66",X"66",X"11",X"14",X"45",X"40",X"FF",X"55",X"55",X"66",X"65",X"55",X"55",X"66",X"64",X"44",
		X"30",X"FF",X"0A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"4A",X"B9",X"FF",X"0B",X"A2",X"A9",
		X"0B",X"00",X"A0",X"A0",X"B0",X"C2",X"90",X"FF",X"09",X"00",X"90",X"A0",X"20",X"B0",X"0A",X"29",
		X"00",X"00",X"FF",X"00",X"0B",X"00",X"09",X"0C",X"00",X"20",X"00",X"C0",X"00",X"FF",X"00",X"44",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"04",X"55",X"14",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"04",X"33",X"34",X"54",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"70",X"84",X"45",X"44",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"78",X"43",X"44",X"44",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"78",X"44",X"44",X"44",X"44",X"40",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"84",X"44",X"44",X"2E",X"34",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",
		X"44",X"42",X"12",X"E4",X"00",X"FF",X"00",X"00",X"00",X"08",X"88",X"34",X"44",X"2D",X"E4",X"30",
		X"FF",X"00",X"82",X"88",X"82",X"82",X"88",X"84",X"44",X"55",X"30",X"FF",X"46",X"65",X"82",X"86",
		X"66",X"66",X"11",X"14",X"45",X"40",X"FF",X"45",X"55",X"66",X"65",X"55",X"55",X"66",X"64",X"44",
		X"30",X"FF",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"4B",X"0A",X"FF",X"09",X"C0",X"BC",
		X"AA",X"C0",X"00",X"B9",X"A0",X"BA",X"90",X"FF",X"00",X"A0",X"90",X"B0",X"B9",X"2A",X"00",X"0A",
		X"90",X"20",X"FF",X"00",X"00",X"20",X"09",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",
		X"00",X"24",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"45",X"00",X"FF",X"00",X"24",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"45",X"39",X"FF",X"89",X"24",X"4A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A4",X"45",X"39",X"FF",X"28",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"45",X"44",X"FF",X"28",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"45",X"39",
		X"FF",X"B9",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"25",X"39",X"FF",X"8A",X"99",
		X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"39",X"AA",X"FF",X"00",X"99",X"44",X"44",X"44",
		X"49",X"94",X"44",X"44",X"48",X"99",X"AA",X"FF",X"00",X"09",X"41",X"11",X"11",X"18",X"94",X"11",
		X"11",X"18",X"9A",X"44",X"FF",X"00",X"09",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"94",
		X"04",X"FF",X"00",X"AA",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",
		X"A0",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"AA",X"98",X"88",
		X"88",X"88",X"98",X"88",X"88",X"89",X"44",X"00",X"FF",X"00",X"00",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"B4",X"41",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"14",X"4B",X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"01",X"10",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",X"00",X"24",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"45",X"00",X"FF",X"00",X"24",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"45",X"39",X"FF",X"89",X"24",X"4A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A4",
		X"45",X"39",X"FF",X"28",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"45",X"44",X"FF",
		X"28",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"45",X"39",X"FF",X"B9",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"25",X"39",X"FF",X"8A",X"99",X"38",X"38",X"38",X"38",
		X"38",X"38",X"38",X"38",X"39",X"AA",X"FF",X"00",X"99",X"44",X"44",X"44",X"49",X"94",X"44",X"44",
		X"48",X"99",X"AA",X"FF",X"00",X"09",X"41",X"11",X"11",X"18",X"94",X"11",X"11",X"18",X"9A",X"44",
		X"FF",X"00",X"09",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"94",X"04",X"FF",X"00",X"AA",
		X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"A0",X"94",X"11",X"11",
		X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"AA",X"98",X"88",X"88",X"88",X"98",X"88",
		X"88",X"89",X"44",X"00",X"FF",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"14",X"41",X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",
		X"41",X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"00",X"00",
		X"0B",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"25",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",X"00",X"24",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"45",X"00",X"FF",X"00",X"24",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"45",
		X"39",X"FF",X"89",X"24",X"4A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A4",X"45",X"39",X"FF",X"28",
		X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"45",X"44",X"FF",X"28",X"24",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"45",X"39",X"FF",X"B9",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"25",X"39",X"FF",X"8A",X"99",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"39",X"AA",X"FF",X"00",X"99",X"44",X"44",X"44",X"49",X"94",X"44",X"44",X"48",X"99",X"AA",X"FF",
		X"00",X"09",X"41",X"11",X"11",X"18",X"94",X"11",X"11",X"18",X"9A",X"44",X"FF",X"00",X"09",X"94",
		X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"94",X"04",X"FF",X"00",X"AA",X"94",X"11",X"11",X"18",
		X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"A0",X"94",X"11",X"11",X"18",X"94",X"11",X"11",
		X"89",X"04",X"04",X"FF",X"00",X"AA",X"98",X"88",X"88",X"88",X"98",X"88",X"88",X"89",X"44",X"00",
		X"FF",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"B4",X"41",
		X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"14",
		X"4B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"01",X"10",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"FF",X"00",X"24",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"45",X"00",
		X"FF",X"00",X"24",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"45",X"39",X"FF",X"89",X"24",
		X"4A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A4",X"45",X"39",X"FF",X"28",X"24",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"44",X"FF",X"28",X"24",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"45",X"39",X"FF",X"B9",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"25",
		X"39",X"FF",X"8A",X"99",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"39",X"AA",X"FF",X"00",
		X"99",X"44",X"44",X"44",X"49",X"94",X"44",X"44",X"48",X"99",X"AA",X"FF",X"00",X"09",X"41",X"11",
		X"11",X"18",X"94",X"11",X"11",X"18",X"9A",X"44",X"FF",X"00",X"09",X"94",X"11",X"11",X"18",X"94",
		X"11",X"11",X"89",X"94",X"04",X"FF",X"00",X"AA",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",
		X"04",X"04",X"FF",X"00",X"A0",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",
		X"00",X"AA",X"98",X"88",X"88",X"88",X"98",X"88",X"88",X"89",X"44",X"00",X"FF",X"00",X"00",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"14",X"41",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"14",X"41",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"0B",X"10",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",
		X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"47",X"66",X"66",X"40",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"46",X"66",X"77",X"40",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"04",X"66",X"66",X"7D",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"04",X"77",X"77",X"77",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"04",X"66",
		X"66",X"66",X"77",X"44",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0D",X"C4",X"2E",X"ED",
		X"D4",X"44",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"EE",X"EC",X"D4",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"55",X"55",X"5D",X"CC",X"CC",X"CC",X"45",X"55",X"55",X"55",X"00",X"FF",
		X"00",X"CC",X"AA",X"AD",X"CC",X"CC",X"74",X"AA",X"AA",X"AA",X"45",X"00",X"FF",X"00",X"EC",X"EA",
		X"AA",X"44",X"EE",X"74",X"AA",X"AA",X"AA",X"45",X"39",X"FF",X"89",X"4E",X"E7",X"AA",X"7D",X"D7",
		X"77",X"DA",X"AA",X"A4",X"45",X"39",X"FF",X"28",X"CC",X"47",X"77",X"37",X"66",X"77",X"D4",X"44",
		X"44",X"45",X"44",X"FF",X"28",X"EC",X"E4",X"47",X"76",X"67",X"7D",X"D4",X"44",X"44",X"45",X"39",
		X"FF",X"B9",X"44",X"35",X"52",X"22",X"22",X"22",X"22",X"22",X"22",X"25",X"39",X"FF",X"8A",X"99",
		X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"39",X"AA",X"FF",X"00",X"99",X"44",X"44",X"44",
		X"49",X"94",X"44",X"44",X"48",X"99",X"AA",X"FF",X"00",X"09",X"41",X"11",X"11",X"18",X"94",X"11",
		X"11",X"18",X"9A",X"44",X"FF",X"00",X"09",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"94",
		X"04",X"FF",X"00",X"AA",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",
		X"A0",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"AA",X"98",X"88",
		X"88",X"88",X"98",X"88",X"88",X"89",X"44",X"00",X"FF",X"00",X"00",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"B4",X"41",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"14",X"4B",X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"01",X"10",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"47",X"66",X"66",X"40",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"46",X"66",X"77",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"04",X"66",X"66",X"7D",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"77",
		X"77",X"77",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"04",X"66",X"66",X"66",X"77",X"44",
		X"40",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0D",X"C4",X"2E",X"ED",X"D4",X"44",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"EE",X"EC",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"55",X"55",X"5D",X"CC",X"CC",X"CC",X"45",X"55",X"55",X"55",X"00",X"FF",X"00",X"CC",X"AA",X"AD",
		X"CC",X"CC",X"74",X"AA",X"AA",X"AA",X"45",X"00",X"FF",X"00",X"EC",X"EA",X"AA",X"44",X"EE",X"74",
		X"AA",X"AA",X"AA",X"45",X"39",X"FF",X"89",X"4E",X"E7",X"AA",X"7D",X"D7",X"77",X"DA",X"AA",X"A4",
		X"45",X"39",X"FF",X"28",X"CC",X"47",X"77",X"37",X"66",X"77",X"D4",X"44",X"44",X"45",X"44",X"FF",
		X"28",X"EC",X"E4",X"47",X"76",X"67",X"7D",X"D4",X"44",X"44",X"45",X"39",X"FF",X"B9",X"44",X"35",
		X"52",X"22",X"22",X"22",X"22",X"22",X"22",X"25",X"39",X"FF",X"8A",X"99",X"38",X"38",X"38",X"38",
		X"38",X"38",X"38",X"38",X"39",X"AA",X"FF",X"00",X"99",X"44",X"44",X"44",X"49",X"94",X"44",X"44",
		X"48",X"99",X"AA",X"FF",X"00",X"09",X"41",X"11",X"11",X"18",X"94",X"11",X"11",X"18",X"9A",X"44",
		X"FF",X"00",X"09",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"94",X"04",X"FF",X"00",X"AA",
		X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"A0",X"94",X"11",X"11",
		X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"AA",X"98",X"88",X"88",X"88",X"98",X"88",
		X"88",X"89",X"44",X"00",X"FF",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"14",X"41",X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",
		X"41",X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"00",X"00",
		X"0B",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"47",X"66",X"66",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"46",X"66",X"77",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"66",X"66",
		X"7D",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"77",X"77",X"77",X"D4",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"04",X"66",X"66",X"66",X"77",X"44",X"40",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"0D",X"C4",X"2E",X"ED",X"D4",X"44",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"DC",X"CC",X"EE",X"EC",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",X"55",X"55",X"5D",X"CC",
		X"CC",X"CC",X"45",X"55",X"55",X"55",X"00",X"FF",X"00",X"CC",X"AA",X"AD",X"CC",X"CC",X"74",X"AA",
		X"AA",X"AA",X"45",X"00",X"FF",X"00",X"EC",X"EA",X"AA",X"44",X"EE",X"74",X"AA",X"AA",X"AA",X"45",
		X"39",X"FF",X"89",X"4E",X"E7",X"AA",X"7D",X"D7",X"77",X"DA",X"AA",X"A4",X"45",X"39",X"FF",X"28",
		X"CC",X"47",X"77",X"37",X"66",X"77",X"D4",X"44",X"44",X"45",X"44",X"FF",X"28",X"EC",X"E4",X"47",
		X"76",X"67",X"7D",X"D4",X"44",X"44",X"45",X"39",X"FF",X"B9",X"44",X"35",X"52",X"22",X"22",X"22",
		X"22",X"22",X"22",X"25",X"39",X"FF",X"8A",X"99",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"39",X"AA",X"FF",X"00",X"99",X"44",X"44",X"44",X"49",X"94",X"44",X"44",X"48",X"99",X"AA",X"FF",
		X"00",X"09",X"41",X"11",X"11",X"18",X"94",X"11",X"11",X"18",X"9A",X"44",X"FF",X"00",X"09",X"94",
		X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"94",X"04",X"FF",X"00",X"AA",X"94",X"11",X"11",X"18",
		X"94",X"11",X"11",X"89",X"04",X"04",X"FF",X"00",X"A0",X"94",X"11",X"11",X"18",X"94",X"11",X"11",
		X"89",X"04",X"04",X"FF",X"00",X"AA",X"98",X"88",X"88",X"88",X"98",X"88",X"88",X"89",X"44",X"00",
		X"FF",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"B4",X"41",
		X"00",X"00",X"14",X"41",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"14",
		X"4B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"01",X"10",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"47",X"66",X"66",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"46",X"66",X"77",
		X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"66",X"66",X"7D",X"D4",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"77",X"77",X"77",X"D4",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"04",X"66",X"66",X"66",X"77",X"44",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"0D",X"C4",X"2E",X"ED",X"D4",X"44",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"EE",
		X"EC",X"D4",X"00",X"00",X"00",X"00",X"FF",X"00",X"55",X"55",X"5D",X"CC",X"CC",X"CC",X"45",X"55",
		X"55",X"55",X"00",X"FF",X"00",X"CC",X"AA",X"AD",X"CC",X"CC",X"74",X"AA",X"AA",X"AA",X"45",X"00",
		X"FF",X"00",X"EC",X"EA",X"AA",X"44",X"EE",X"74",X"AA",X"AA",X"AA",X"45",X"39",X"FF",X"89",X"4E",
		X"E7",X"AA",X"7D",X"D7",X"77",X"DA",X"AA",X"A4",X"45",X"39",X"FF",X"28",X"CC",X"47",X"77",X"37",
		X"66",X"77",X"D4",X"44",X"44",X"45",X"44",X"FF",X"28",X"EC",X"E4",X"47",X"76",X"67",X"7D",X"D4",
		X"44",X"44",X"45",X"39",X"FF",X"B9",X"44",X"35",X"52",X"22",X"22",X"22",X"22",X"22",X"22",X"25",
		X"39",X"FF",X"8A",X"99",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"39",X"AA",X"FF",X"00",
		X"99",X"44",X"44",X"44",X"49",X"94",X"44",X"44",X"48",X"99",X"AA",X"FF",X"00",X"09",X"41",X"11",
		X"11",X"18",X"94",X"11",X"11",X"18",X"9A",X"44",X"FF",X"00",X"09",X"94",X"11",X"11",X"18",X"94",
		X"11",X"11",X"89",X"94",X"04",X"FF",X"00",X"AA",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",
		X"04",X"04",X"FF",X"00",X"A0",X"94",X"11",X"11",X"18",X"94",X"11",X"11",X"89",X"04",X"04",X"FF",
		X"00",X"AA",X"98",X"88",X"88",X"88",X"98",X"88",X"88",X"89",X"44",X"00",X"FF",X"00",X"00",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"14",X"41",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"14",X"41",X"00",X"00",X"14",X"41",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"0B",X"10",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"45",X"09",X"90",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"AA",X"45",X"59",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"AA",X"AA",X"44",X"54",X"49",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"44",
		X"55",X"99",X"FF",X"00",X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"45",X"9A",X"FF",
		X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"29",X"AA",X"FF",X"00",X"00",X"55",
		X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"39",X"44",X"FF",X"00",X"55",X"AA",X"AA",X"AA",X"A4",
		X"44",X"42",X"28",X"38",X"99",X"04",X"FF",X"22",X"4A",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"34",
		X"48",X"94",X"04",X"FF",X"02",X"44",X"4A",X"A4",X"44",X"42",X"28",X"34",X"41",X"18",X"94",X"40",
		X"FF",X"02",X"24",X"44",X"44",X"42",X"28",X"39",X"41",X"11",X"18",X"90",X"40",X"FF",X"00",X"24",
		X"44",X"42",X"28",X"34",X"89",X"41",X"11",X"11",X"99",X"44",X"FF",X"09",X"22",X"42",X"28",X"34",
		X"44",X"89",X"44",X"11",X"88",X"99",X"40",X"FF",X"88",X"92",X"28",X"34",X"41",X"11",X"18",X"94",
		X"88",X"89",X"99",X"00",X"FF",X"B2",X"82",X"88",X"44",X"11",X"11",X"18",X"94",X"89",X"99",X"00",
		X"00",X"FF",X"0B",X"89",X"99",X"94",X"11",X"11",X"88",X"99",X"99",X"33",X"10",X"00",X"FF",X"00",
		X"8A",X"09",X"94",X"41",X"88",X"89",X"99",X"03",X"44",X"10",X"00",X"FF",X"00",X"00",X"00",X"99",
		X"48",X"89",X"99",X"00",X"0B",X"44",X"10",X"00",X"FF",X"00",X"00",X"0A",X"A9",X"99",X"99",X"00",
		X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"AA",X"09",X"99",X"33",X"10",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",X"03",X"44",X"B0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"45",X"09",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"AA",X"45",X"59",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"AA",X"AA",X"44",X"54",
		X"49",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"44",X"55",X"99",X"FF",X"00",
		X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"45",X"9A",X"FF",X"00",X"00",X"00",X"55",
		X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"29",X"AA",X"FF",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",
		X"44",X"42",X"28",X"39",X"44",X"FF",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"38",
		X"99",X"04",X"FF",X"22",X"4A",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"34",X"48",X"94",X"04",X"FF",
		X"02",X"44",X"4A",X"A4",X"44",X"42",X"28",X"34",X"41",X"18",X"94",X"40",X"FF",X"02",X"24",X"44",
		X"44",X"42",X"28",X"39",X"41",X"11",X"18",X"90",X"40",X"FF",X"00",X"24",X"44",X"42",X"28",X"34",
		X"89",X"41",X"11",X"11",X"99",X"44",X"FF",X"09",X"22",X"42",X"28",X"34",X"44",X"89",X"44",X"11",
		X"88",X"99",X"40",X"FF",X"88",X"92",X"28",X"34",X"41",X"11",X"18",X"94",X"88",X"89",X"99",X"00",
		X"FF",X"B2",X"82",X"88",X"44",X"11",X"11",X"18",X"94",X"89",X"99",X"00",X"00",X"FF",X"0B",X"89",
		X"99",X"94",X"11",X"11",X"88",X"99",X"99",X"33",X"10",X"00",X"FF",X"00",X"8A",X"09",X"94",X"41",
		X"88",X"89",X"99",X"03",X"44",X"10",X"00",X"FF",X"00",X"00",X"00",X"99",X"48",X"89",X"99",X"00",
		X"01",X"44",X"10",X"00",X"FF",X"00",X"00",X"0A",X"A9",X"99",X"99",X"00",X"00",X"00",X"1B",X"00",
		X"00",X"FF",X"00",X"00",X"AA",X"09",X"99",X"33",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0A",X"AA",X"03",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"45",X"09",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"AA",X"45",X"59",X"40",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"AA",X"AA",X"44",X"54",X"49",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"44",X"55",X"99",X"FF",X"00",X"00",X"00",X"00",X"55",
		X"AA",X"AA",X"AA",X"A4",X"44",X"45",X"9A",X"FF",X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",
		X"44",X"42",X"29",X"AA",X"FF",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"39",
		X"44",X"FF",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"38",X"99",X"04",X"FF",X"22",
		X"4A",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"34",X"48",X"94",X"04",X"FF",X"02",X"44",X"4A",X"A4",
		X"44",X"42",X"28",X"34",X"41",X"18",X"94",X"40",X"FF",X"02",X"24",X"44",X"44",X"42",X"28",X"39",
		X"41",X"11",X"18",X"90",X"40",X"FF",X"00",X"24",X"44",X"42",X"28",X"34",X"89",X"41",X"11",X"11",
		X"99",X"44",X"FF",X"09",X"22",X"42",X"28",X"34",X"44",X"89",X"44",X"11",X"88",X"99",X"40",X"FF",
		X"88",X"92",X"28",X"34",X"41",X"11",X"18",X"94",X"88",X"89",X"99",X"00",X"FF",X"B2",X"82",X"88",
		X"44",X"11",X"11",X"18",X"94",X"89",X"99",X"00",X"00",X"FF",X"0B",X"89",X"99",X"94",X"11",X"11",
		X"88",X"99",X"99",X"33",X"10",X"00",X"FF",X"00",X"8A",X"09",X"94",X"41",X"88",X"89",X"99",X"03",
		X"44",X"B0",X"00",X"FF",X"00",X"00",X"00",X"99",X"48",X"89",X"99",X"00",X"01",X"44",X"10",X"00",
		X"FF",X"00",X"00",X"0A",X"A9",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",
		X"AA",X"09",X"99",X"33",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",X"03",
		X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",X"44",X"10",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"45",X"09",X"90",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"AA",X"45",X"59",X"40",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"AA",X"AA",X"44",X"54",X"49",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",
		X"AA",X"AA",X"AA",X"44",X"55",X"99",X"FF",X"00",X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",
		X"44",X"45",X"9A",X"FF",X"00",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"29",X"AA",
		X"FF",X"00",X"00",X"55",X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"39",X"44",X"FF",X"00",X"55",
		X"AA",X"AA",X"AA",X"A4",X"44",X"42",X"28",X"38",X"99",X"04",X"FF",X"22",X"4A",X"AA",X"AA",X"A4",
		X"44",X"42",X"28",X"34",X"48",X"94",X"04",X"FF",X"02",X"44",X"4A",X"A4",X"44",X"42",X"28",X"34",
		X"41",X"18",X"94",X"40",X"FF",X"02",X"24",X"44",X"44",X"42",X"28",X"39",X"41",X"11",X"18",X"90",
		X"40",X"FF",X"00",X"24",X"44",X"42",X"28",X"34",X"89",X"41",X"11",X"11",X"99",X"44",X"FF",X"09",
		X"22",X"42",X"28",X"34",X"44",X"89",X"44",X"11",X"88",X"99",X"40",X"FF",X"88",X"92",X"28",X"34",
		X"41",X"11",X"18",X"94",X"88",X"89",X"99",X"00",X"FF",X"B2",X"82",X"88",X"44",X"11",X"11",X"18",
		X"94",X"89",X"99",X"00",X"00",X"FF",X"0B",X"89",X"99",X"94",X"11",X"11",X"88",X"99",X"99",X"33",
		X"10",X"00",X"FF",X"00",X"8A",X"09",X"94",X"41",X"88",X"89",X"99",X"03",X"44",X"10",X"00",X"FF",
		X"00",X"00",X"00",X"99",X"48",X"89",X"99",X"00",X"01",X"44",X"10",X"00",X"FF",X"00",X"00",X"0A",
		X"A9",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"AA",X"09",X"99",X"33",
		X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",X"03",X"44",X"10",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"76",
		X"66",X"64",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"66",X"67",X"74",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"46",X"66",X"67",X"DD",X"40",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"47",X"77",X"77",X"7D",X"40",X"00",X"55",X"00",X"00",X"FF",X"00",
		X"00",X"46",X"66",X"66",X"67",X"74",X"44",X"55",X"45",X"09",X"90",X"FF",X"00",X"00",X"00",X"DC",
		X"42",X"EE",X"DD",X"44",X"4A",X"45",X"59",X"40",X"FF",X"00",X"00",X"0D",X"CC",X"CE",X"EE",X"CD",
		X"4A",X"AA",X"44",X"54",X"49",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"CC",X"C4",X"AA",X"AA",X"44",
		X"55",X"99",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"C7",X"4A",X"AA",X"A4",X"44",X"45",X"9A",X"FF",
		X"00",X"00",X"00",X"54",X"4E",X"E7",X"4A",X"A4",X"44",X"42",X"29",X"AA",X"FF",X"00",X"00",X"55",
		X"AA",X"AD",X"77",X"7D",X"44",X"42",X"28",X"39",X"44",X"FF",X"00",X"55",X"AA",X"AA",X"A7",X"66",
		X"74",X"42",X"28",X"38",X"99",X"04",X"FF",X"22",X"4A",X"AA",X"AA",X"77",X"66",X"42",X"28",X"34",
		X"48",X"94",X"04",X"FF",X"0C",X"CC",X"4A",X"67",X"46",X"62",X"28",X"34",X"41",X"18",X"94",X"40",
		X"FF",X"0C",X"EE",X"E4",X"74",X"62",X"28",X"39",X"41",X"11",X"18",X"90",X"40",X"FF",X"00",X"4C",
		X"C4",X"65",X"58",X"34",X"89",X"41",X"11",X"11",X"99",X"44",X"FF",X"09",X"EE",X"E3",X"58",X"34",
		X"44",X"89",X"44",X"11",X"88",X"99",X"40",X"FF",X"88",X"94",X"48",X"34",X"41",X"11",X"18",X"94",
		X"88",X"89",X"99",X"00",X"FF",X"B2",X"84",X"88",X"44",X"11",X"11",X"18",X"94",X"89",X"99",X"00",
		X"00",X"FF",X"0B",X"89",X"99",X"94",X"11",X"11",X"88",X"99",X"99",X"33",X"10",X"00",X"FF",X"00",
		X"8A",X"09",X"94",X"41",X"88",X"89",X"99",X"03",X"44",X"10",X"00",X"FF",X"00",X"00",X"00",X"99",
		X"48",X"89",X"99",X"00",X"0B",X"44",X"10",X"00",X"FF",X"00",X"00",X"0A",X"A9",X"99",X"99",X"00",
		X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"AA",X"09",X"99",X"33",X"10",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",X"03",X"44",X"B0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"44",X"44",
		X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"76",X"66",X"64",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"66",X"67",X"74",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"46",X"66",X"67",X"DD",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"47",X"77",X"77",X"7D",X"40",X"00",X"55",X"00",X"00",X"FF",X"00",X"00",X"46",X"66",X"66",
		X"67",X"74",X"44",X"55",X"45",X"09",X"90",X"FF",X"00",X"00",X"00",X"DC",X"42",X"EE",X"DD",X"44",
		X"4A",X"45",X"59",X"40",X"FF",X"00",X"00",X"0D",X"CC",X"CE",X"EE",X"CD",X"4A",X"AA",X"44",X"54",
		X"49",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"CC",X"C4",X"AA",X"AA",X"44",X"55",X"99",X"FF",X"00",
		X"00",X"00",X"DC",X"CC",X"C7",X"4A",X"AA",X"A4",X"44",X"45",X"9A",X"FF",X"00",X"00",X"00",X"54",
		X"4E",X"E7",X"4A",X"A4",X"44",X"42",X"29",X"AA",X"FF",X"00",X"00",X"55",X"AA",X"AD",X"77",X"7D",
		X"44",X"42",X"28",X"39",X"44",X"FF",X"00",X"55",X"AA",X"AA",X"A7",X"66",X"74",X"42",X"28",X"38",
		X"99",X"04",X"FF",X"22",X"4A",X"AA",X"AA",X"77",X"66",X"42",X"28",X"34",X"48",X"94",X"04",X"FF",
		X"0C",X"CC",X"4A",X"67",X"46",X"62",X"28",X"34",X"41",X"18",X"94",X"40",X"FF",X"0C",X"EE",X"E4",
		X"74",X"62",X"28",X"39",X"41",X"11",X"18",X"90",X"40",X"FF",X"00",X"4C",X"C4",X"65",X"58",X"34",
		X"89",X"41",X"11",X"11",X"99",X"44",X"FF",X"09",X"EE",X"E3",X"58",X"34",X"44",X"89",X"44",X"11",
		X"88",X"99",X"40",X"FF",X"88",X"94",X"48",X"34",X"41",X"11",X"18",X"94",X"88",X"89",X"99",X"00",
		X"FF",X"B2",X"84",X"88",X"44",X"11",X"11",X"18",X"94",X"89",X"99",X"00",X"00",X"FF",X"0B",X"89",
		X"99",X"94",X"11",X"11",X"88",X"99",X"99",X"33",X"10",X"00",X"FF",X"00",X"8A",X"09",X"94",X"41",
		X"88",X"89",X"99",X"03",X"44",X"10",X"00",X"FF",X"00",X"00",X"00",X"99",X"48",X"89",X"99",X"00",
		X"01",X"44",X"10",X"00",X"FF",X"00",X"00",X"0A",X"A9",X"99",X"99",X"00",X"00",X"00",X"1B",X"00",
		X"00",X"FF",X"00",X"00",X"AA",X"09",X"99",X"33",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0A",X"AA",X"03",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"76",X"66",X"64",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"04",X"66",X"67",X"74",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"46",X"66",X"67",X"DD",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"47",X"77",X"77",
		X"7D",X"40",X"00",X"55",X"00",X"00",X"FF",X"00",X"00",X"46",X"66",X"66",X"67",X"74",X"44",X"55",
		X"45",X"09",X"90",X"FF",X"00",X"00",X"00",X"DC",X"42",X"EE",X"DD",X"44",X"4A",X"45",X"59",X"40",
		X"FF",X"00",X"00",X"0D",X"CC",X"CE",X"EE",X"CD",X"4A",X"AA",X"44",X"54",X"49",X"FF",X"00",X"00",
		X"00",X"DC",X"CC",X"CC",X"C4",X"AA",X"AA",X"44",X"55",X"99",X"FF",X"00",X"00",X"00",X"DC",X"CC",
		X"C7",X"4A",X"AA",X"A4",X"44",X"45",X"9A",X"FF",X"00",X"00",X"00",X"54",X"4E",X"E7",X"4A",X"A4",
		X"44",X"42",X"29",X"AA",X"FF",X"00",X"00",X"55",X"AA",X"AD",X"77",X"7D",X"44",X"42",X"28",X"39",
		X"44",X"FF",X"00",X"55",X"AA",X"AA",X"A7",X"66",X"74",X"42",X"28",X"38",X"99",X"04",X"FF",X"22",
		X"4A",X"AA",X"AA",X"77",X"66",X"42",X"28",X"34",X"48",X"94",X"04",X"FF",X"0C",X"CC",X"4A",X"67",
		X"46",X"62",X"28",X"34",X"41",X"18",X"94",X"40",X"FF",X"0C",X"EE",X"E4",X"74",X"62",X"28",X"39",
		X"41",X"11",X"18",X"90",X"40",X"FF",X"00",X"4C",X"C4",X"65",X"58",X"34",X"89",X"41",X"11",X"11",
		X"99",X"44",X"FF",X"09",X"EE",X"E3",X"58",X"34",X"44",X"89",X"44",X"11",X"88",X"99",X"40",X"FF",
		X"88",X"94",X"48",X"34",X"41",X"11",X"18",X"94",X"88",X"89",X"99",X"00",X"FF",X"B2",X"84",X"88",
		X"44",X"11",X"11",X"18",X"94",X"89",X"99",X"00",X"00",X"FF",X"0B",X"89",X"99",X"94",X"11",X"11",
		X"88",X"99",X"99",X"33",X"10",X"00",X"FF",X"00",X"8A",X"09",X"94",X"41",X"88",X"89",X"99",X"03",
		X"44",X"B0",X"00",X"FF",X"00",X"00",X"00",X"99",X"48",X"89",X"99",X"00",X"01",X"44",X"10",X"00",
		X"FF",X"00",X"00",X"0A",X"A9",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",
		X"AA",X"09",X"99",X"33",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",X"03",
		X"44",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",X"44",X"10",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"04",X"76",X"66",X"64",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",
		X"66",X"67",X"74",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"46",X"66",X"67",X"DD",
		X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"47",X"77",X"77",X"7D",X"40",X"00",X"55",
		X"00",X"00",X"FF",X"00",X"00",X"46",X"66",X"66",X"67",X"74",X"44",X"55",X"45",X"09",X"90",X"FF",
		X"00",X"00",X"00",X"DC",X"42",X"EE",X"DD",X"44",X"4A",X"45",X"59",X"40",X"FF",X"00",X"00",X"0D",
		X"CC",X"CE",X"EE",X"CD",X"4A",X"AA",X"44",X"54",X"49",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"CC",
		X"C4",X"AA",X"AA",X"44",X"55",X"99",X"FF",X"00",X"00",X"00",X"DC",X"CC",X"C7",X"4A",X"AA",X"A4",
		X"44",X"45",X"9A",X"FF",X"00",X"00",X"00",X"54",X"4E",X"E7",X"4A",X"A4",X"44",X"42",X"29",X"AA",
		X"FF",X"00",X"00",X"55",X"AA",X"AD",X"77",X"7D",X"44",X"42",X"28",X"39",X"44",X"FF",X"00",X"55",
		X"AA",X"AA",X"A7",X"66",X"74",X"42",X"28",X"38",X"99",X"04",X"FF",X"22",X"4A",X"AA",X"AA",X"77",
		X"66",X"42",X"28",X"34",X"48",X"94",X"04",X"FF",X"0C",X"CC",X"4A",X"67",X"46",X"62",X"28",X"34",
		X"41",X"18",X"94",X"40",X"FF",X"0C",X"EE",X"E4",X"74",X"62",X"28",X"39",X"41",X"11",X"18",X"90",
		X"40",X"FF",X"00",X"4C",X"C4",X"65",X"58",X"34",X"89",X"41",X"11",X"11",X"99",X"44",X"FF",X"09",
		X"EE",X"E3",X"58",X"34",X"44",X"89",X"44",X"11",X"88",X"99",X"40",X"FF",X"88",X"94",X"48",X"34",
		X"41",X"11",X"18",X"94",X"88",X"89",X"99",X"00",X"FF",X"B2",X"84",X"88",X"44",X"11",X"11",X"18",
		X"94",X"89",X"99",X"00",X"00",X"FF",X"0B",X"89",X"99",X"94",X"11",X"11",X"88",X"99",X"99",X"33",
		X"10",X"00",X"FF",X"00",X"8A",X"09",X"94",X"41",X"88",X"89",X"99",X"03",X"44",X"10",X"00",X"FF",
		X"00",X"00",X"00",X"99",X"48",X"89",X"99",X"00",X"01",X"44",X"10",X"00",X"FF",X"00",X"00",X"0A",
		X"A9",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"AA",X"09",X"99",X"33",
		X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",X"03",X"44",X"10",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"44",X"10",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"21",X"FF",
		X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",
		X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",
		X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",X"21",X"FF",
		X"21",X"FF",X"21",X"FF",X"00",X"FF",X"00",X"21",X"FF",X"00",X"21",X"FF",X"00",X"21",X"FF",X"00",
		X"21",X"FF",X"00",X"21",X"FF",X"00",X"21",X"FF",X"00",X"21",X"FF",X"00",X"21",X"FF",X"00",X"21",
		X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",
		X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",X"10",X"FF",X"02",
		X"10",X"FF",X"21",X"00",X"FF",X"21",X"00",X"FF",X"21",X"00",X"FF",X"21",X"00",X"FF",X"21",X"00",
		X"FF",X"21",X"00",X"FF",X"21",X"00",X"FF",X"21",X"00",X"FF",X"00",X"00",X"21",X"FF",X"00",X"02",
		X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",
		X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"21",
		X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",
		X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",
		X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",
		X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",
		X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",
		X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",
		X"00",X"21",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",
		X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"21",X"00",
		X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",
		X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",
		X"21",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"FF",X"02",X"10",
		X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"FF",X"21",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"21",X"FF",X"00",X"00",X"21",X"FF",X"00",X"00",X"21",X"FF",X"00",X"00",
		X"21",X"FF",X"00",X"00",X"21",X"FF",X"00",X"00",X"21",X"FF",X"00",X"00",X"21",X"FF",X"00",X"02",
		X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",
		X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"02",X"10",X"FF",X"00",X"21",
		X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",
		X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"21",X"00",X"FF",X"00",X"10",X"00",X"FF",X"02",X"10",
		X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",X"00",X"FF",X"02",X"10",
		X"00",X"FF",X"02",X"10",X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",
		X"00",X"FF",X"21",X"00",X"00",X"FF",X"21",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",
		X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",
		X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"21",
		X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"02",X"10",X"00",
		X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",
		X"00",X"21",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"FF",X"02",
		X"10",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"FF",X"21",X"00",
		X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"10",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"02",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",
		X"21",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"21",
		X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",
		X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"02",X"10",X"FF",X"00",
		X"00",X"21",X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",
		X"21",X"00",X"FF",X"00",X"00",X"21",X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",
		X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",X"00",X"FF",X"00",X"02",X"10",X"00",
		X"FF",X"00",X"21",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"21",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"FF",X"02",
		X"10",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"FF",X"21",X"00",
		X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"10",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"02",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"10",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"02",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"02",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",
		X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"02",X"10",
		X"00",X"FF",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",
		X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"21",X"FF",
		X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"02",
		X"10",X"FF",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",
		X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"02",X"20",X"FF",X"00",X"00",X"00",X"21",X"00",X"FF",
		X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"21",
		X"00",X"FF",X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",
		X"02",X"10",X"00",X"FF",X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"02",X"10",X"00",
		X"00",X"FF",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"21",
		X"00",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"00",X"FF",
		X"02",X"10",X"00",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"00",X"FF",X"21",X"00",X"00",X"00",
		X"00",X"FF",X"21",X"00",X"00",X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"02",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"21",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"02",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"21",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"02",X"21",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"21",X"10",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"02",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"21",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"10",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"02",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"20",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"60",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"80",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"FF",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"55",X"23",X"43",X"55",X"00",X"00",X"FF",X"00",X"05",X"22",X"22",X"23",X"44",X"50",X"00",X"FF",
		X"00",X"52",X"21",X"11",X"22",X"34",X"45",X"00",X"FF",X"05",X"22",X"11",X"11",X"12",X"23",X"44",
		X"50",X"FF",X"05",X"32",X"11",X"11",X"12",X"23",X"34",X"50",X"FF",X"53",X"32",X"11",X"11",X"12",
		X"33",X"34",X"45",X"FF",X"53",X"32",X"21",X"11",X"22",X"33",X"34",X"45",X"FF",X"53",X"32",X"22",
		X"22",X"22",X"33",X"34",X"45",X"FF",X"53",X"33",X"22",X"22",X"23",X"33",X"44",X"45",X"FF",X"53",
		X"33",X"32",X"33",X"33",X"33",X"44",X"45",X"FF",X"05",X"33",X"33",X"33",X"33",X"34",X"44",X"50",
		X"FF",X"05",X"44",X"33",X"33",X"33",X"44",X"44",X"50",X"FF",X"00",X"54",X"44",X"43",X"44",X"44",
		X"45",X"00",X"FF",X"00",X"05",X"44",X"44",X"44",X"44",X"50",X"00",X"FF",X"00",X"00",X"55",X"44",
		X"44",X"55",X"00",X"00",X"FF",X"00",X"00",X"05",X"66",X"65",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"05",X"24",X"45",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"56",X"50",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"FF",X"00",X"00",X"07",X"00",X"07",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"77",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"04",X"00",X"00",
		X"40",X"00",X"00",X"FF",X"22",X"20",X"00",X"42",X"24",X"00",X"02",X"22",X"FF",X"04",X"42",X"00",
		X"72",X"27",X"00",X"24",X"40",X"FF",X"02",X"44",X"21",X"64",X"26",X"12",X"44",X"20",X"FF",X"22",
		X"22",X"42",X"15",X"51",X"24",X"22",X"22",X"FF",X"00",X"22",X"22",X"21",X"12",X"22",X"22",X"00",
		X"FF",X"02",X"24",X"42",X"12",X"21",X"24",X"42",X"20",X"FF",X"00",X"02",X"24",X"22",X"22",X"42",
		X"20",X"00",X"FF",X"00",X"00",X"24",X"12",X"21",X"42",X"00",X"00",X"FF",X"00",X"02",X"00",X"21",
		X"12",X"00",X"20",X"00",X"FF",X"00",X"00",X"00",X"20",X"02",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"04",X"00",X"00",X"40",X"00",X"00",X"FF",X"00",X"00",X"00",X"42",X"24",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"72",X"27",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"68",X"C6",X"20",X"00",
		X"00",X"FF",X"00",X"02",X"22",X"15",X"51",X"22",X"20",X"00",X"FF",X"00",X"22",X"44",X"21",X"12",
		X"44",X"22",X"00",X"FF",X"00",X"24",X"22",X"12",X"21",X"22",X"42",X"00",X"FF",X"02",X"42",X"02",
		X"12",X"21",X"20",X"24",X"20",X"FF",X"02",X"20",X"20",X"21",X"12",X"02",X"02",X"20",X"FF",X"00",
		X"20",X"00",X"20",X"02",X"00",X"02",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"48",
		X"88",X"80",X"00",X"00",X"FF",X"00",X"00",X"48",X"44",X"44",X"48",X"80",X"10",X"FF",X"00",X"08",
		X"84",X"44",X"88",X"84",X"48",X"01",X"FF",X"00",X"04",X"44",X"88",X"88",X"18",X"D8",X"00",X"FF",
		X"00",X"04",X"47",X"87",X"44",X"82",X"24",X"80",X"FF",X"00",X"84",X"74",X"77",X"44",X"81",X"2D",
		X"80",X"FF",X"00",X"84",X"47",X"77",X"74",X"48",X"24",X"10",X"FF",X"00",X"84",X"47",X"77",X"74",
		X"48",X"22",X"80",X"FF",X"00",X"08",X"44",X"77",X"44",X"88",X"21",X"01",X"FF",X"00",X"0D",X"84",
		X"44",X"48",X"80",X"21",X"00",X"FF",X"00",X"00",X"0D",X"D8",X"80",X"00",X"10",X"10",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"20",X"20",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",
		X"81",X"80",X"00",X"00",X"FF",X"00",X"00",X"08",X"84",X"D4",X"31",X"10",X"00",X"FF",X"00",X"00",
		X"84",X"D2",X"22",X"30",X"00",X"00",X"FF",X"00",X"00",X"88",X"82",X"18",X"88",X"00",X"30",X"FF",
		X"00",X"08",X"84",X"18",X"84",X"48",X"80",X"00",X"FF",X"00",X"08",X"44",X"D4",X"44",X"44",X"80",
		X"10",X"FF",X"00",X"08",X"4D",X"D4",X"47",X"74",X"48",X"01",X"FF",X"00",X"0D",X"44",X"84",X"77",
		X"74",X"48",X"01",X"FF",X"00",X"0D",X"44",X"74",X"77",X"77",X"4D",X"00",X"FF",X"00",X"00",X"84",
		X"47",X"77",X"74",X"8D",X"00",X"FF",X"00",X"00",X"48",X"44",X"74",X"48",X"D0",X"00",X"FF",X"00",
		X"00",X"08",X"DD",X"48",X"8D",X"D0",X"00",X"FF",X"00",X"00",X"00",X"0D",X"8D",X"80",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"88",X"DD",X"00",X"00",X"FF",X"00",X"03",X"00",X"88",X"44",X"48",X"DD",X"00",X"FF",X"00",X"01",
		X"08",X"84",X"44",X"74",X"8D",X"00",X"FF",X"00",X"00",X"08",X"44",X"77",X"77",X"48",X"80",X"FF",
		X"00",X"10",X"08",X"44",X"77",X"77",X"44",X"D0",X"FF",X"00",X"01",X"D0",X"84",X"47",X"77",X"74",
		X"80",X"FF",X"00",X"01",X"1D",X"84",X"44",X"77",X"4D",X"D0",X"FF",X"00",X"01",X"18",X"11",X"48",
		X"44",X"4D",X"80",X"FF",X"00",X"00",X"18",X"44",X"D4",X"44",X"88",X"00",X"FF",X"00",X"00",X"18",
		X"84",X"44",X"88",X"48",X"00",X"FF",X"00",X"00",X"08",X"11",X"88",X"8D",X"D0",X"00",X"FF",X"00",
		X"00",X"00",X"0D",X"DD",X"D0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"33",X"00",X"FF",X"00",X"00",X"00",X"03",X"33",X"30",X"3A",X"AB",X"A0",X"FF",X"00",X"00",
		X"00",X"33",X"30",X"0B",X"A9",X"30",X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"CA",X"9A",X"BA",
		X"00",X"FF",X"00",X"00",X"00",X"33",X"30",X"A3",X"99",X"00",X"00",X"FF",X"00",X"00",X"03",X"33",
		X"3B",X"99",X"AB",X"A0",X"00",X"FF",X"00",X"03",X"37",X"D3",X"3A",X"9A",X"90",X"00",X"00",X"FF",
		X"00",X"38",X"E3",X"33",X"39",X"99",X"B3",X"33",X"00",X"FF",X"03",X"11",X"1E",X"33",X"33",X"33",
		X"33",X"30",X"30",X"FF",X"00",X"32",X"23",X"33",X"33",X"33",X"33",X"33",X"00",X"FF",X"00",X"00",
		X"00",X"03",X"33",X"34",X"E3",X"03",X"30",X"FF",X"00",X"00",X"00",X"00",X"0E",X"4E",X"30",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"00",X"30",X"FF",X"00",X"03",X"33",X"33",X"33",X"33",X"00",X"33",X"00",X"FF",X"00",X"3E",
		X"37",X"D3",X"33",X"33",X"33",X"30",X"30",X"FF",X"03",X"8E",X"13",X"33",X"A3",X"AA",X"33",X"33",
		X"00",X"FF",X"00",X"06",X"62",X"3B",X"CA",X"3A",X"A3",X"30",X"00",X"FF",X"00",X"03",X"23",X"33",
		X"3C",X"CB",X"BB",X"33",X"00",X"FF",X"00",X"00",X"00",X"33",X"33",X"E4",X"E3",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"32",X"23",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"33",X"03",X"33",X"30",X"00",X"00",X"03",X"30",X"FF",X"03",X"8E",X"37",X"D3",
		X"33",X"33",X"03",X"33",X"00",X"FF",X"38",X"1E",X"13",X"33",X"33",X"33",X"33",X"33",X"30",X"FF",
		X"31",X"05",X"61",X"39",X"A3",X"33",X"33",X"30",X"00",X"FF",X"00",X"56",X"42",X"3B",X"A3",X"AA",
		X"33",X"03",X"30",X"FF",X"00",X"04",X"20",X"BA",X"93",X"3A",X"B0",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"BA",X"93",X"A3",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CA",X"A9",X"9A",X"B0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0C",X"AA",X"99",X"90",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"CC",X"CB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"66",X"16",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"61",X"B1",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"66",X"66",X"16",X"66",X"00",X"FF",X"00",X"00",X"00",X"66",X"66",X"26",
		X"66",X"63",X"00",X"FF",X"00",X"00",X"66",X"66",X"22",X"26",X"22",X"30",X"00",X"FF",X"00",X"00",
		X"66",X"22",X"22",X"26",X"23",X"00",X"00",X"FF",X"00",X"06",X"26",X"66",X"67",X"76",X"60",X"00",
		X"00",X"FF",X"00",X"06",X"77",X"77",X"66",X"27",X"60",X"00",X"00",X"FF",X"00",X"07",X"66",X"66",
		X"76",X"60",X"60",X"00",X"00",X"FF",X"00",X"06",X"22",X"66",X"62",X"60",X"60",X"00",X"00",X"FF",
		X"00",X"00",X"77",X"22",X"22",X"00",X"06",X"00",X"00",X"FF",X"00",X"00",X"00",X"77",X"72",X"26",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"66",X"1B",X"16",
		X"60",X"FF",X"00",X"00",X"00",X"06",X"66",X"66",X"61",X"66",X"66",X"FF",X"00",X"00",X"00",X"66",
		X"66",X"22",X"66",X"62",X"30",X"FF",X"00",X"00",X"06",X"62",X"22",X"22",X"66",X"23",X"00",X"FF",
		X"00",X"00",X"06",X"67",X"22",X"22",X"36",X"30",X"00",X"FF",X"00",X"00",X"06",X"62",X"72",X"32",
		X"36",X"00",X"00",X"FF",X"00",X"00",X"06",X"62",X"33",X"33",X"36",X"70",X"00",X"FF",X"00",X"00",
		X"06",X"27",X"73",X"30",X"06",X"07",X"00",X"FF",X"00",X"00",X"66",X"27",X"00",X"00",X"00",X"60",
		X"00",X"FF",X"00",X"00",X"62",X"77",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"20",X"70",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"27",X"70",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"06",X"20",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"60",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"06",X"66",X"60",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"00",X"00",X"26",X"00",X"00",X"22",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"66",X"00",X"07",X"70",X"00",X"00",X"00",X"FF",X"00",X"06",
		X"60",X"00",X"00",X"77",X"00",X"00",X"00",X"FF",X"00",X"66",X"00",X"06",X"66",X"66",X"60",X"00",
		X"00",X"FF",X"00",X"66",X"66",X"66",X"62",X"66",X"66",X"00",X"00",X"FF",X"00",X"02",X"72",X"72",
		X"72",X"26",X"66",X"66",X"60",X"FF",X"00",X"00",X"00",X"03",X"32",X"22",X"26",X"62",X"16",X"FF",
		X"00",X"00",X"00",X"03",X"33",X"22",X"76",X"21",X"B1",X"FF",X"00",X"00",X"00",X"00",X"33",X"37",
		X"62",X"66",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"37",X"22",X"26",X"60",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"76",X"03",X"32",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"70",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"07",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"0C",X"00",X"00",X"FF",X"00",X"CB",X"00",X"BC",X"05",X"00",
		X"FF",X"00",X"0C",X"B0",X"9D",X"5B",X"B0",X"FF",X"0B",X"0D",X"BD",X"5D",X"BC",X"0B",X"FF",X"0C",
		X"55",X"DB",X"9D",X"CB",X"BC",X"FF",X"00",X"DC",X"BC",X"5C",X"9D",X"D0",X"FF",X"0B",X"59",X"55",
		X"CD",X"55",X"9B",X"FF",X"CC",X"CC",X"BC",X"9C",X"BC",X"D0",X"FF",X"00",X"BB",X"DB",X"5B",X"DB",
		X"B0",X"FF",X"0B",X"0C",X"9D",X"5C",X"9C",X"CB",X"FF",X"00",X"0C",X"BD",X"BC",X"B0",X"C0",X"FF",
		X"00",X"CB",X"0C",X"B0",X"CB",X"0C",X"FF",X"00",X"00",X"0C",X"00",X"0C",X"00",X"FF",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"FF",X"00",X"00",X"DD",X"E4",X"45",X"C0",X"FF",X"00",X"DD",X"3D",X"EC",
		X"46",X"5C",X"FF",X"0D",X"38",X"3D",X"BC",X"DD",X"45",X"FF",X"0D",X"87",X"83",X"33",X"22",X"D5",
		X"FF",X"D3",X"87",X"78",X"81",X"32",X"DC",X"FF",X"D1",X"7C",X"88",X"1C",X"12",X"3C",X"FF",X"D1",
		X"78",X"C1",X"C1",X"12",X"DC",X"FF",X"D3",X"78",X"11",X"11",X"13",X"DC",X"FF",X"D3",X"18",X"CC",
		X"C1",X"23",X"C0",X"FF",X"0D",X"3C",X"A1",X"AC",X"3D",X"C0",X"FF",X"0D",X"32",X"12",X"22",X"DC",
		X"00",X"FF",X"00",X"D3",X"DC",X"DD",X"C0",X"00",X"FF",X"00",X"0C",X"C0",X"CC",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"05",X"45",X"35",X"55",X"00",X"55",X"33",X"55",X"00",X"55",X"00",
		X"FF",X"00",X"55",X"33",X"33",X"35",X"55",X"53",X"00",X"03",X"35",X"00",X"00",X"FF",X"05",X"53",
		X"30",X"00",X"03",X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"55",X"53",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"54",X"55",X"33",X"35",X"50",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"55",X"33",
		X"00",X"33",X"50",X"00",X"00",X"05",X"55",X"50",X"FF",X"00",X"05",X"53",X"00",X"00",X"03",X"35",
		X"50",X"00",X"53",X"00",X"05",X"FF",X"00",X"55",X"03",X"00",X"00",X"00",X"33",X"55",X"55",X"30",
		X"00",X"00",X"FF",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"33",X"30",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",X"53",X"33",X"33",X"55",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"55",X"33",X"00",X"00",X"33",X"50",X"00",X"00",X"00",X"FF",X"00",X"54",
		X"53",X"53",X"30",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"FF",X"55",X"55",X"33",X"33",X"00",
		X"00",X"00",X"00",X"35",X"00",X"00",X"00",X"FF",X"03",X"33",X"30",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"50",X"00",X"FF",X"00",
		X"00",X"08",X"00",X"00",X"00",X"FF",X"00",X"88",X"83",X"88",X"80",X"00",X"FF",X"08",X"43",X"33",
		X"72",X"28",X"00",X"FF",X"84",X"44",X"73",X"33",X"22",X"80",X"FF",X"84",X"74",X"44",X"73",X"72",
		X"80",X"FF",X"84",X"44",X"74",X"43",X"33",X"80",X"FF",X"08",X"65",X"55",X"54",X"48",X"00",X"FF",
		X"08",X"68",X"55",X"48",X"48",X"00",X"FF",X"08",X"68",X"85",X"88",X"48",X"00",X"FF",X"08",X"65",
		X"55",X"44",X"48",X"00",X"FF",X"08",X"65",X"55",X"54",X"48",X"00",X"FF",X"08",X"61",X"81",X"81",
		X"48",X"00",X"FF",X"08",X"61",X"81",X"81",X"48",X"00",X"FF",X"08",X"66",X"64",X"44",X"48",X"00",
		X"FF",X"00",X"86",X"65",X"44",X"80",X"00",X"FF",X"00",X"08",X"85",X"88",X"00",X"00",X"FF",X"00",
		X"00",X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"62",X"66",X"00",X"FF",
		X"06",X"33",X"26",X"60",X"FF",X"66",X"43",X"26",X"27",X"FF",X"62",X"42",X"22",X"27",X"FF",X"66",
		X"42",X"32",X"66",X"FF",X"62",X"32",X"32",X"26",X"FF",X"62",X"32",X"22",X"66",X"FF",X"61",X"44",
		X"44",X"27",X"FF",X"61",X"42",X"24",X"47",X"FF",X"44",X"14",X"42",X"44",X"FF",X"42",X"44",X"24",
		X"24",X"FF",X"42",X"42",X"24",X"11",X"FF",X"44",X"24",X"42",X"44",X"FF",X"04",X"42",X"24",X"40",
		X"FF",X"00",X"44",X"44",X"00",X"FF",X"00",X"62",X"66",X"00",X"FF",X"06",X"32",X"26",X"60",X"FF",
		X"73",X"42",X"36",X"26",X"FF",X"64",X"22",X"22",X"26",X"FF",X"24",X"23",X"26",X"66",X"FF",X"24",
		X"23",X"26",X"26",X"FF",X"23",X"22",X"22",X"66",X"FF",X"62",X"44",X"44",X"16",X"FF",X"64",X"42",
		X"24",X"16",X"FF",X"44",X"24",X"41",X"44",X"FF",X"42",X"42",X"14",X"24",X"FF",X"42",X"42",X"24",
		X"24",X"FF",X"11",X"24",X"42",X"44",X"FF",X"04",X"42",X"24",X"40",X"FF",X"00",X"44",X"44",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"62",X"66",X"00",X"FF",
		X"06",X"26",X"23",X"60",X"FF",X"76",X"26",X"34",X"26",X"FF",X"66",X"22",X"43",X"26",X"FF",X"62",
		X"63",X"43",X"62",X"FF",X"66",X"12",X"32",X"26",X"FF",X"76",X"12",X"32",X"26",X"FF",X"76",X"14",
		X"44",X"62",X"FF",X"74",X"12",X"24",X"46",X"FF",X"44",X"21",X"42",X"44",X"FF",X"42",X"42",X"24",
		X"24",X"FF",X"42",X"42",X"24",X"24",X"FF",X"44",X"24",X"42",X"44",X"FF",X"04",X"41",X"24",X"40",
		X"FF",X"00",X"41",X"44",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"07",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"07",X"46",X"47",
		X"44",X"00",X"00",X"FF",X"00",X"00",X"00",X"46",X"70",X"06",X"47",X"60",X"00",X"FF",X"00",X"00",
		X"00",X"46",X"00",X"00",X"04",X"44",X"00",X"FF",X"00",X"00",X"01",X"60",X"00",X"00",X"06",X"70",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"46",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"66",X"00",X"FF",X"00",X"00",X"00",X"03",X"55",X"56",X"67",X"70",X"00",X"FF",
		X"00",X"00",X"53",X"22",X"34",X"47",X"44",X"00",X"00",X"FF",X"00",X"95",X"22",X"23",X"54",X"67",
		X"00",X"66",X"00",X"FF",X"07",X"55",X"93",X"35",X"46",X"44",X"00",X"00",X"00",X"FF",X"00",X"77",
		X"55",X"56",X"67",X"04",X"00",X"00",X"00",X"FF",X"44",X"60",X"77",X"76",X"74",X"06",X"60",X"00",
		X"00",X"FF",X"00",X"46",X"70",X"46",X"04",X"00",X"00",X"00",X"00",X"FF",X"06",X"64",X"74",X"60",
		X"06",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"07",X"44",X"70",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"04",X"46",X"67",X"46",X"00",X"FF",X"00",X"00",X"00",X"00",X"16",X"60",
		X"00",X"46",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"46",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"74",X"46",X"70",X"00",X"FF",X"00",X"00",X"00",X"05",
		X"55",X"67",X"66",X"00",X"00",X"FF",X"00",X"00",X"03",X"54",X"44",X"74",X"70",X"00",X"00",X"FF",
		X"00",X"03",X"22",X"35",X"46",X"60",X"40",X"00",X"00",X"FF",X"04",X"92",X"23",X"54",X"67",X"40",
		X"66",X"00",X"00",X"FF",X"07",X"54",X"95",X"66",X"60",X"04",X"00",X"00",X"00",X"FF",X"00",X"77",
		X"67",X"67",X"74",X"06",X"60",X"00",X"00",X"FF",X"04",X"46",X"04",X"40",X"04",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"04",X"74",X"60",X"06",X"60",X"00",X"00",X"00",X"FF",X"00",X"66",X"67",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"62",X"33",X"22",X"00",X"00",X"FF",X"00",X"66",
		X"23",X"32",X"36",X"26",X"00",X"FF",X"06",X"22",X"63",X"22",X"36",X"66",X"60",X"FF",X"06",X"62",
		X"44",X"44",X"44",X"26",X"10",X"FF",X"66",X"44",X"33",X"22",X"22",X"44",X"17",X"FF",X"64",X"43",
		X"44",X"44",X"44",X"21",X"47",X"FF",X"64",X"34",X"43",X"32",X"24",X"12",X"47",X"FF",X"44",X"04",
		X"30",X"44",X"00",X"42",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"63",X"32",X"66",X"00",X"00",X"FF",X"00",X"62",
		X"63",X"62",X"32",X"66",X"00",X"FF",X"06",X"66",X"23",X"21",X"36",X"26",X"70",X"FF",X"06",X"62",
		X"44",X"41",X"44",X"26",X"70",X"FF",X"76",X"44",X"22",X"21",X"22",X"44",X"67",X"FF",X"74",X"40",
		X"44",X"04",X"04",X"24",X"47",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"66",X"32",X"66",X"00",X"00",X"FF",X"00",X"76",
		X"13",X"32",X"26",X"67",X"00",X"FF",X"07",X"62",X"14",X"44",X"42",X"67",X"70",X"FF",X"07",X"70",
		X"41",X"22",X"00",X"47",X"70",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"FF",X"00",X"00",X"0E",X"11",X"10",X"00",X"00",X"FF",X"00",X"00",
		X"22",X"21",X"22",X"EE",X"01",X"FF",X"00",X"12",X"22",X"12",X"22",X"2E",X"00",X"FF",X"0E",X"22",
		X"55",X"5E",X"2E",X"22",X"10",X"FF",X"0E",X"25",X"58",X"E8",X"E2",X"22",X"30",X"FF",X"E2",X"2E",
		X"8E",X"78",X"E8",X"23",X"31",X"FF",X"E2",X"25",X"67",X"E6",X"72",X"22",X"31",X"FF",X"12",X"28",
		X"87",X"88",X"68",X"23",X"21",X"FF",X"13",X"21",X"E8",X"78",X"68",X"23",X"30",X"FF",X"03",X"22",
		X"28",X"62",X"83",X"23",X"10",X"FF",X"01",X"32",X"32",X"22",X"23",X"33",X"10",X"FF",X"01",X"33",
		X"22",X"32",X"33",X"33",X"00",X"FF",X"00",X"13",X"33",X"33",X"32",X"30",X"00",X"FF",X"00",X"00",
		X"11",X"33",X"30",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"0D",X"12",X"20",X"FF",X"D5",X"D1",
		X"22",X"FF",X"1D",X"21",X"33",X"FF",X"12",X"12",X"13",X"FF",X"32",X"32",X"39",X"FF",X"03",X"23",
		X"30",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0D",X"D1",X"00",X"00",X"10",X"FF",X"00",X"01",
		X"33",X"32",X"31",X"10",X"00",X"FF",X"00",X"E2",X"23",X"23",X"33",X"32",X"0E",X"FF",X"00",X"22",
		X"22",X"52",X"22",X"33",X"30",X"FF",X"00",X"2E",X"58",X"28",X"83",X"33",X"20",X"FF",X"01",X"25",
		X"5E",X"76",X"68",X"23",X"22",X"FF",X"01",X"2E",X"88",X"68",X"82",X"12",X"32",X"FF",X"02",X"15",
		X"E7",X"E8",X"76",X"23",X"33",X"FF",X"02",X"22",X"5E",X"77",X"88",X"22",X"31",X"FF",X"02",X"21",
		X"18",X"68",X"E2",X"32",X"30",X"FF",X"00",X"22",X"1E",X"58",X"32",X"23",X"10",X"FF",X"00",X"12",
		X"22",X"22",X"22",X"33",X"00",X"FF",X"00",X"0E",X"E3",X"32",X"33",X"21",X"00",X"FF",X"00",X"00",
		X"0E",X"E1",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"02",X"23",X"10",X"01",X"0D",X"FF",X"00",X"03",X"22",X"33",X"33",X"10",X"00",X"FF",X"00",X"23",
		X"33",X"23",X"22",X"33",X"10",X"FF",X"01",X"23",X"32",X"12",X"23",X"23",X"20",X"FF",X"01",X"32",
		X"38",X"26",X"82",X"3E",X"30",X"FF",X"03",X"32",X"86",X"87",X"8E",X"33",X"3E",X"FF",X"12",X"32",
		X"86",X"88",X"78",X"82",X"21",X"FF",X"D2",X"25",X"27",X"6E",X"76",X"23",X"3E",X"FF",X"12",X"32",
		X"8E",X"87",X"E8",X"E3",X"30",X"FF",X"01",X"22",X"55",X"8E",X"21",X"23",X"E0",X"FF",X"00",X"22",
		X"E5",X"E2",X"21",X"32",X"00",X"FF",X"00",X"E2",X"22",X"21",X"22",X"21",X"00",X"FF",X"00",X"00",
		X"21",X"12",X"11",X"00",X"00",X"FF",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"09",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",X"CC",
		X"CC",X"CC",X"CC",X"9C",X"C9",X"9C",X"99",X"9C",X"C9",X"FF",X"09",X"99",X"9E",X"EE",X"EE",X"AE",
		X"EA",X"AE",X"AA",X"AE",X"00",X"FF",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"07",X"00",X"70",X"00",X"00",X"FF",X"00",X"00",X"7C",X"D7",X"CD",X"00",
		X"00",X"FF",X"00",X"00",X"0D",X"99",X"D9",X"07",X"00",X"FF",X"00",X"00",X"04",X"49",X"99",X"90",
		X"00",X"FF",X"00",X"00",X"0E",X"CE",X"CE",X"90",X"00",X"FF",X"00",X"00",X"09",X"99",X"9C",X"47",
		X"00",X"FF",X"00",X"00",X"00",X"44",X"44",X"90",X"00",X"FF",X"00",X"00",X"00",X"07",X"76",X"97",
		X"00",X"FF",X"00",X"00",X"00",X"44",X"49",X"C0",X"00",X"FF",X"00",X"00",X"00",X"76",X"49",X"C0",
		X"00",X"FF",X"00",X"00",X"04",X"44",X"9C",X"07",X"00",X"FF",X"00",X"00",X"07",X"69",X"9C",X"00",
		X"00",X"FF",X"00",X"00",X"44",X"99",X"C0",X"70",X"00",X"FF",X"00",X"00",X"76",X"9C",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"44",X"9C",X"70",X"00",X"00",X"FF",X"00",X"00",X"09",X"C0",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"FF",X"00",X"00",X"70",X"07",X"00",X"00",
		X"00",X"FF",X"00",X"07",X"6D",X"76",X"D0",X"70",X"00",X"FF",X"00",X"00",X"D4",X"9D",X"99",X"00",
		X"00",X"FF",X"00",X"00",X"04",X"49",X"99",X"90",X"00",X"FF",X"00",X"00",X"EC",X"EC",X"EC",X"90",
		X"70",X"FF",X"00",X"00",X"00",X"99",X"99",X"49",X"00",X"FF",X"00",X"00",X"00",X"04",X"44",X"99",
		X"00",X"FF",X"00",X"00",X"00",X"07",X"74",X"9C",X"70",X"FF",X"00",X"00",X"00",X"04",X"46",X"9C",
		X"00",X"FF",X"00",X"00",X"00",X"47",X"49",X"C0",X"70",X"FF",X"00",X"00",X"74",X"74",X"69",X"C0",
		X"00",X"FF",X"00",X"09",X"64",X"64",X"9C",X"07",X"00",X"FF",X"00",X"09",X"99",X"99",X"C0",X"00",
		X"00",X"FF",X"00",X"00",X"CC",X"CC",X"07",X"00",X"00",X"FF",X"00",X"00",X"07",X"07",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0E",X"E3",X"31",X"1E",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"E4",X"48",X"31",X"13",X"1E",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"4A",X"86",X"33",
		X"A6",X"83",X"E0",X"00",X"00",X"FF",X"00",X"0E",X"E8",X"A8",X"65",X"63",X"65",X"6A",X"8E",X"E0",
		X"00",X"FF",X"0E",X"EA",X"8A",X"AA",X"86",X"3A",X"A6",X"83",X"A8",X"3E",X"E0",X"FF",X"E5",X"AA",
		X"A5",X"55",X"8A",X"AA",X"AA",X"55",X"5A",X"83",X"5E",X"FF",X"0E",X"55",X"5E",X"EE",X"55",X"55",
		X"55",X"EE",X"E5",X"55",X"E0",X"FF",X"00",X"EE",X"E0",X"00",X"EE",X"EE",X"EE",X"00",X"0E",X"EE",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"EE",X"33",X"EE",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"33",X"11",
		X"13",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"E8",X"3A",X"31",X"11",X"3E",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0E",X"E3",X"A6",X"83",X"A6",X"3E",X"E0",X"00",X"00",X"FF",X"00",X"00",
		X"EE",X"33",X"67",X"63",X"67",X"68",X"EE",X"00",X"00",X"FF",X"00",X"0E",X"88",X"38",X"A6",X"A8",
		X"86",X"AA",X"83",X"E0",X"00",X"FF",X"00",X"EA",X"55",X"38",X"AA",X"55",X"58",X"8A",X"A5",X"5E",
		X"00",X"FF",X"0E",X"85",X"EE",X"5A",X"A5",X"EE",X"E5",X"8A",X"5E",X"E5",X"E0",X"FF",X"0E",X"5E",
		X"00",X"E5",X"5E",X"00",X"0E",X"55",X"E0",X"0E",X"5E",X"FF",X"00",X"E0",X"00",X"0E",X"E0",X"00",
		X"00",X"EE",X"00",X"00",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"EE",
		X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"E3",X"31",X"3E",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0E",X"33",X"11",X"13",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"E8",X"88",X"83",X"13",X"3E",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"E8",X"A6",X"88",
		X"36",X"3E",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"8A",X"65",X"6A",X"65",X"63",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"0E",X"4A",X"86",X"8A",X"A6",X"33",X"E0",X"00",X"00",X"FF",X"00",X"00",
		X"E8",X"A8",X"38",X"88",X"A8",X"83",X"3E",X"00",X"00",X"FF",X"00",X"EE",X"88",X"A5",X"58",X"88",
		X"AA",X"A5",X"58",X"EE",X"00",X"FF",X"0E",X"58",X"8A",X"5E",X"E5",X"88",X"8A",X"5E",X"E5",X"A5",
		X"E0",X"FF",X"00",X"E5",X"55",X"E0",X"0E",X"55",X"55",X"E0",X"0E",X"5E",X"00",X"FF",X"00",X"0E",
		X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
