library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kroozr_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kroozr_sp_bits is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"AA",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"07",X"77",X"00",X"0A",X"00",X"77",
		X"00",X"0A",X"77",X"70",X"00",X"00",X"07",X"77",X"00",X"AA",X"00",X"07",X"00",X"00",X"00",X"77",
		X"00",X"06",X"00",X"77",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"67",X"00",X"00",X"F0",X"07",
		X"FF",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"76",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A6",X"66",X"00",X"00",X"00",X"70",X"00",
		X"00",X"FA",X"77",X"0A",X"00",X"AA",X"70",X"0A",X"00",X"AA",X"76",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"A0",X"66",X"00",X"00",X"00",X"AA",X"00",X"00",X"06",X"6A",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"66",
		X"00",X"00",X"00",X"00",X"00",X"F6",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"06",X"7A",X"00",
		X"00",X"00",X"A0",X"0A",X"00",X"00",X"A7",X"A6",X"00",X"00",X"F0",X"00",X"00",X"06",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"70",X"00",X"FF",X"66",X"00",X"00",X"FF",X"00",X"00",X"60",X"00",X"00",
		X"00",X"A0",X"F0",X"00",X"00",X"00",X"A7",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"66",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"0A",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A7",X"00",X"00",X"00",X"A0",X"60",
		X"00",X"00",X"FA",X"00",X"00",X"0A",X"7A",X"00",X"00",X"00",X"77",X"00",X"00",X"07",X"F7",X"00",
		X"60",X"76",X"FF",X"00",X"00",X"07",X"F7",X"00",X"00",X"66",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"06",X"7A",X"00",X"00",X"00",X"7A",X"60",X"00",X"00",X"FA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"A7",X"00",
		X"00",X"00",X"FA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"67",X"00",
		X"00",X"00",X"70",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"07",X"00",X"6C",X"00",X"7A",
		X"00",X"66",X"06",X"77",X"00",X"06",X"66",X"17",X"00",X"00",X"55",X"00",X"00",X"00",X"35",X"55",
		X"00",X"72",X"35",X"A5",X"00",X"27",X"35",X"A5",X"00",X"77",X"35",X"A5",X"00",X"70",X"35",X"A5",
		X"06",X"70",X"35",X"AA",X"06",X"00",X"35",X"AA",X"0A",X"C5",X"33",X"AA",X"0A",X"C5",X"33",X"AA",
		X"06",X"C1",X"31",X"A1",X"06",X"C1",X"33",X"A1",X"06",X"C1",X"30",X"AA",X"01",X"C1",X"30",X"AA",
		X"00",X"C1",X"30",X"AA",X"00",X"C1",X"3C",X"AA",X"00",X"1C",X"30",X"1A",X"00",X"0C",X"30",X"0A",
		X"00",X"0C",X"31",X"0A",X"00",X"0C",X"00",X"0A",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"00",X"06",X"60",X"D6",X"00",X"66",X"60",X"00",X"00",X"A3",X"66",X"00",X"00",
		X"A3",X"06",X"02",X"00",X"AA",X"0A",X"07",X"00",X"5A",X"AD",X"07",X"00",X"5A",X"5D",X"07",X"00",
		X"5A",X"5D",X"07",X"60",X"5A",X"D5",X"00",X"60",X"5A",X"DD",X"53",X"66",X"5C",X"5D",X"53",X"66",
		X"5C",X"5D",X"53",X"56",X"55",X"5D",X"33",X"5A",X"25",X"5D",X"33",X"AA",X"26",X"55",X"33",X"A5",
		X"61",X"25",X"33",X"A5",X"61",X"22",X"33",X"A5",X"61",X"22",X"53",X"A1",X"E1",X"12",X"53",X"A1",
		X"E1",X"12",X"53",X"11",X"E1",X"11",X"53",X"10",X"E1",X"11",X"53",X"10",X"E0",X"11",X"53",X"00",
		X"E0",X"11",X"53",X"00",X"E0",X"11",X"60",X"00",X"E0",X"11",X"60",X"00",X"E0",X"00",X"60",X"00",
		X"E0",X"00",X"60",X"00",X"E0",X"00",X"63",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"E3",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"EE",X"00",X"00",X"0D",X"AA",X"00",
		X"00",X"0D",X"FF",X"00",X"00",X"0D",X"FF",X"00",X"00",X"DD",X"9F",X"00",X"00",X"DE",X"09",X"EC",
		X"00",X"DE",X"09",X"DC",X"00",X"EC",X"9F",X"DE",X"0C",X"EC",X"FF",X"00",X"0C",X"6C",X"55",X"00",
		X"CC",X"6C",X"55",X"00",X"C0",X"CC",X"00",X"00",X"C0",X"CE",X"AA",X"C0",X"EC",X"CE",X"EE",X"C0",
		X"0C",X"E0",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"E6",
		X"00",X"00",X"EE",X"60",X"00",X"0E",X"EE",X"00",X"00",X"EE",X"06",X"00",X"00",X"0E",X"66",X"00",
		X"00",X"00",X"6E",X"00",X"00",X"07",X"EE",X"00",X"00",X"0A",X"EE",X"00",X"00",X"00",X"6E",X"00",
		X"00",X"66",X"6E",X"00",X"00",X"66",X"66",X"00",X"00",X"11",X"61",X"00",X"00",X"01",X"10",X"00",
		X"00",X"00",X"10",X"19",X"00",X"00",X"11",X"49",X"00",X"00",X"14",X"99",X"00",X"00",X"07",X"94",
		X"00",X"00",X"E0",X"44",X"00",X"0E",X"E0",X"44",X"00",X"EE",X"0E",X"44",X"00",X"E7",X"0E",X"45",
		X"00",X"E4",X"77",X"45",X"00",X"14",X"44",X"54",X"00",X"44",X"44",X"44",X"01",X"44",X"45",X"44",
		X"01",X"44",X"44",X"11",X"11",X"44",X"44",X"10",X"7A",X"44",X"11",X"00",X"01",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",
		X"00",X"00",X"EE",X"E6",X"00",X"00",X"EE",X"60",X"00",X"0E",X"60",X"00",X"00",X"60",X"06",X"00",
		X"00",X"E0",X"6E",X"00",X"00",X"E0",X"6E",X"00",X"00",X"E0",X"6E",X"00",X"00",X"60",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"16",X"66",X"00",X"00",X"01",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"61",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"E6",X"00",X"00",X"11",X"EE",X"10",
		X"00",X"14",X"EE",X"11",X"00",X"44",X"00",X"44",X"00",X"47",X"E6",X"44",X"00",X"41",X"66",X"44",
		X"00",X"44",X"77",X"44",X"00",X"44",X"11",X"44",X"00",X"44",X"44",X"41",X"00",X"14",X"44",X"11",
		X"00",X"11",X"A4",X"10",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"7A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0A",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"E6",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"7E",X"99",
		X"00",X"00",X"7E",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"E1",X"99",X"00",X"00",X"11",X"09",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6E",X"50",X"00",X"00",X"66",X"50",X"00",X"AA",X"66",X"50",
		X"00",X"AA",X"66",X"50",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"66",
		X"00",X"00",X"55",X"AA",X"00",X"00",X"55",X"AA",X"00",X"00",X"55",X"AA",X"00",X"05",X"55",X"AA",
		X"00",X"AA",X"55",X"AA",X"00",X"AA",X"50",X"A9",X"00",X"10",X"06",X"90",X"00",X"11",X"6A",X"00",
		X"00",X"A1",X"99",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"0E",X"AA",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"77",X"EC",X"00",X"00",X"00",X"00",X"00",X"EE",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"DC",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"DD",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"2B",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"22",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0A",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"E6",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"7E",X"99",
		X"00",X"00",X"7E",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"E1",X"99",X"00",X"00",X"11",X"09",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6E",X"50",X"00",X"00",X"66",X"50",X"00",X"AA",X"66",X"50",
		X"00",X"AA",X"66",X"50",X"00",X"AA",X"66",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"66",
		X"00",X"55",X"55",X"AA",X"00",X"AA",X"35",X"AA",X"00",X"A1",X"55",X"AA",X"00",X"11",X"55",X"AA",
		X"00",X"10",X"55",X"AA",X"00",X"00",X"55",X"A9",X"00",X"00",X"50",X"90",X"00",X"00",X"50",X"00",
		X"00",X"40",X"09",X"00",X"00",X"44",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"66",
		X"00",X"00",X"DD",X"66",X"00",X"00",X"DD",X"66",X"00",X"00",X"00",X"06",X"00",X"D9",X"ED",X"C0",
		X"00",X"ED",X"00",X"CC",X"00",X"9E",X"ED",X"DC",X"00",X"99",X"00",X"DD",X"00",X"9D",X"DD",X"DD",
		X"00",X"DE",X"DD",X"DD",X"00",X"00",X"CC",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"88",X"88",X"88",X"77",X"77",X"77",X"88",X"88",X"88",X"77",X"88",X"87",X"8F",X"77",
		X"88",X"77",X"87",X"77",X"88",X"88",X"88",X"77",X"88",X"77",X"8F",X"77",X"88",X"77",X"87",X"77",
		X"88",X"7F",X"88",X"87",X"88",X"77",X"77",X"77",X"88",X"77",X"77",X"77",X"88",X"00",X"88",X"88",
		X"88",X"00",X"88",X"88",X"88",X"88",X"BB",X"88",X"88",X"8B",X"33",X"88",X"88",X"B8",X"33",X"88",
		X"88",X"8B",X"33",X"88",X"88",X"88",X"BB",X"88",X"88",X"8D",X"88",X"88",X"88",X"83",X"33",X"88",
		X"88",X"8D",X"33",X"88",X"88",X"8D",X"33",X"88",X"88",X"8B",X"33",X"88",X"88",X"88",X"BB",X"88",
		X"88",X"8D",X"88",X"88",X"88",X"8D",X"33",X"88",X"88",X"8D",X"33",X"88",X"88",X"8D",X"33",X"88",
		X"88",X"8D",X"33",X"88",X"88",X"8D",X"33",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"38",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"73",X"5E",X"00",X"00",X"EE",X"55",
		X"00",X"00",X"5E",X"55",X"00",X"00",X"5E",X"55",X"00",X"55",X"55",X"EE",X"00",X"15",X"55",X"55",
		X"00",X"15",X"55",X"55",X"00",X"11",X"55",X"55",X"00",X"10",X"55",X"55",X"00",X"00",X"55",X"55",
		X"00",X"00",X"55",X"55",X"00",X"10",X"55",X"55",X"00",X"11",X"55",X"55",X"00",X"15",X"55",X"55",
		X"00",X"45",X"55",X"55",X"00",X"55",X"55",X"66",X"00",X"00",X"56",X"55",X"00",X"00",X"46",X"55",
		X"00",X"00",X"66",X"44",X"00",X"00",X"64",X"46",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"55",X"EE",X"0E",
		X"00",X"55",X"5E",X"33",X"00",X"11",X"5E",X"55",X"00",X"11",X"55",X"55",X"00",X"66",X"55",X"55",
		X"00",X"66",X"55",X"55",X"00",X"66",X"55",X"EE",X"00",X"E6",X"55",X"55",X"F5",X"56",X"55",X"55",
		X"54",X"41",X"55",X"55",X"00",X"16",X"55",X"55",X"00",X"66",X"55",X"66",X"00",X"66",X"55",X"55",
		X"00",X"66",X"55",X"55",X"00",X"11",X"55",X"55",X"00",X"11",X"56",X"44",X"00",X"55",X"56",X"44",
		X"00",X"44",X"66",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"4E",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E6",X"00",X"00",X"F5",X"56",X"00",
		X"00",X"54",X"41",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"46",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"70",X"00",X"00",X"60",X"07",X"00",
		X"00",X"60",X"07",X"00",X"00",X"06",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"06",X"60",X"00",X"00",X"60",X"60",X"60",X"00",X"60",X"00",X"60",
		X"00",X"66",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"06",X"70",X"00",X"00",X"00",X"07",X"00",
		X"00",X"06",X"07",X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"60",X"00",X"00",X"60",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"0C",X"AA",X"9C",X"AA",X"00",X"00",X"00",X"00",X"00",X"AA",X"99",X"AC",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"99",X"00",X"D9",X"09",X"90",X"00",X"DD",X"09",X"90",
		X"00",X"9D",X"99",X"99",X"00",X"09",X"9C",X"90",X"00",X"09",X"9F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"BF",X"00",X"09",X"99",X"9F",X"99",X"B9",X"FF",X"F9",X"FB",X"09",X"99",X"B9",X"99",
		X"00",X"DB",X"9F",X"CB",X"00",X"99",X"9B",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"D0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"09",
		X"00",X"09",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9B",X"00",
		X"00",X"00",X"9B",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9B",X"99",X"00",X"00",X"9B",X"9D",
		X"00",X"00",X"9F",X"DD",X"00",X"90",X"9F",X"D9",X"00",X"C9",X"9F",X"90",X"00",X"9B",X"F9",X"9B",
		X"00",X"99",X"9F",X"B0",X"00",X"99",X"F9",X"00",X"00",X"09",X"9B",X"00",X"00",X"00",X"F9",X"90",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"FF",X"9C",X"00",X"00",X"9F",X"FF",
		X"00",X"00",X"9F",X"99",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9B",X"9B",X"00",X"0C",X"9B",X"BB",
		X"00",X"09",X"9F",X"99",X"00",X"90",X"9B",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9F",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"66",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"07",
		X"00",X"00",X"00",X"07",X"00",X"70",X"00",X"70",X"00",X"77",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"10",X"00",X"60",X"00",X"10",
		X"00",X"00",X"00",X"01",X"00",X"00",X"07",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"70",X"0F",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"F0",X"00",
		X"20",X"00",X"F0",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"22",
		X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"21",X"00",X"00",X"09",X"11",X"00",X"00",X"A9",X"21",X"00",X"00",X"A9",X"41",
		X"00",X"AA",X"E9",X"11",X"00",X"AA",X"A9",X"22",X"00",X"AA",X"E9",X"42",X"00",X"AA",X"AA",X"42",
		X"00",X"EE",X"AA",X"44",X"00",X"DE",X"AA",X"14",X"00",X"0D",X"AA",X"91",X"00",X"00",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"86",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"42",
		X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"84",
		X"00",X"00",X"00",X"01",X"00",X"00",X"09",X"11",X"00",X"00",X"A9",X"11",X"00",X"00",X"A9",X"11",
		X"00",X"AA",X"E9",X"11",X"00",X"AA",X"A9",X"11",X"00",X"AA",X"E9",X"44",X"00",X"AA",X"AA",X"42",
		X"00",X"EE",X"AA",X"44",X"00",X"DE",X"AA",X"11",X"00",X"0D",X"AA",X"91",X"00",X"00",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"00",X"09",X"18",X"00",X"00",X"A9",X"18",X"00",X"00",X"A9",X"18",
		X"00",X"AA",X"E9",X"22",X"00",X"AA",X"A9",X"22",X"00",X"AA",X"E9",X"22",X"00",X"AA",X"AA",X"24",
		X"00",X"EE",X"AA",X"28",X"00",X"DE",X"AA",X"81",X"00",X"0D",X"AA",X"91",X"00",X"00",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"DD",
		X"06",X"00",X"00",X"00",X"60",X"88",X"00",X"00",X"60",X"88",X"00",X"00",X"66",X"68",X"00",X"00",
		X"62",X"08",X"00",X"00",X"26",X"02",X"00",X"00",X"FF",X"62",X"00",X"00",X"0F",X"22",X"00",X"00",
		X"00",X"12",X"00",X"00",X"00",X"42",X"00",X"00",X"22",X"12",X"00",X"00",X"22",X"42",X"00",X"00",
		X"22",X"42",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"00",X"00",X"00",X"24",X"00",X"00",X"00",
		X"41",X"EE",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"AE",X"00",X"00",X"88",X"EE",X"00",
		X"00",X"88",X"AA",X"00",X"82",X"88",X"AA",X"A0",X"82",X"88",X"EA",X"AA",X"22",X"88",X"EE",X"AD",
		X"24",X"88",X"AA",X"D0",X"44",X"99",X"AA",X"00",X"46",X"9A",X"AA",X"00",X"66",X"AA",X"AA",X"00",
		X"99",X"AA",X"AD",X"00",X"AA",X"AA",X"DD",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"0D",X"CC",X"00",X"00",X"D0",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"C0",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"00",X"00",X"CC",X"0C",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"D0",X"90",X"0C",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"C0",X"00",
		X"00",X"D0",X"0D",X"00",X"0D",X"DD",X"00",X"00",X"CD",X"C0",X"0C",X"00",X"0C",X"CC",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"D0",X"00",X"00",X"90",X"CD",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"0D",X"CD",X"00",X"00",X"C0",X"C0",
		X"00",X"00",X"0C",X"0C",X"00",X"C0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"CD",X"00",
		X"00",X"00",X"00",X"DD",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"0C",X"C0",
		X"DC",X"00",X"00",X"C0",X"CD",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0D",X"00",X"00",X"00",X"0C",
		X"DC",X"00",X"00",X"00",X"C0",X"00",X"00",X"CD",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"DD",X"00",X"C0",X"CC",X"CC",X"00",X"D0",X"0C",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"D0",X"00",X"00",X"00",X"0C",X"CD",X"0C",X"90",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"66",X"80",X"00",X"00",X"66",X"82",X"00",X"00",X"26",X"82",X"00",
		X"00",X"61",X"82",X"00",X"88",X"FF",X"22",X"00",X"08",X"0F",X"22",X"00",X"88",X"00",X"24",X"00",
		X"00",X"00",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"22",X"00",X"20",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"88",X"12",X"00",X"40",
		X"08",X"01",X"22",X"00",X"08",X"00",X"00",X"00",X"08",X"02",X"22",X"00",X"00",X"22",X"22",X"00",
		X"04",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"22",
		X"08",X"00",X"42",X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"66",X"80",X"00",X"00",X"66",X"82",X"00",X"00",X"26",X"82",X"00",
		X"00",X"61",X"82",X"00",X"88",X"FF",X"22",X"00",X"08",X"0F",X"22",X"00",X"88",X"00",X"24",X"00",
		X"00",X"00",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"02",X"00",X"88",X"12",X"22",X"00",
		X"08",X"01",X"24",X"00",X"08",X"00",X"41",X"00",X"08",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"42",X"22",X"22",
		X"08",X"22",X"22",X"20",X"00",X"24",X"42",X"00",X"00",X"22",X"04",X"00",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"66",X"80",X"00",X"00",X"66",X"82",X"00",X"00",X"26",X"82",X"00",
		X"00",X"61",X"82",X"00",X"88",X"FF",X"22",X"00",X"08",X"0F",X"22",X"00",X"88",X"00",X"24",X"00",
		X"00",X"00",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"22",X"11",X"00",X"00",X"22",X"22",X"00",X"00",X"21",X"21",X"00",X"88",X"12",X"22",X"24",
		X"08",X"01",X"42",X"22",X"08",X"00",X"14",X"22",X"08",X"00",X"11",X"22",X"00",X"00",X"01",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"41",
		X"08",X"00",X"01",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"A9",X"11",X"00",X"00",X"A9",X"11",
		X"00",X"AA",X"E9",X"11",X"00",X"AA",X"A9",X"11",X"00",X"AA",X"E9",X"11",X"00",X"AA",X"AA",X"11",
		X"00",X"EE",X"AA",X"11",X"00",X"DE",X"AA",X"11",X"00",X"0D",X"AA",X"91",X"00",X"00",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"08",X"AF",X"00",X"00",X"08",X"AF",X"00",X"00",X"80",X"AA",X"00",
		X"00",X"80",X"AA",X"00",X"00",X"0A",X"AA",X"00",X"EE",X"AA",X"AA",X"00",X"11",X"01",X"AA",X"00",
		X"11",X"EE",X"AA",X"00",X"11",X"11",X"AA",X"00",X"11",X"11",X"1A",X"00",X"11",X"D1",X"11",X"D0",
		X"11",X"D1",X"A1",X"DD",X"11",X"D1",X"AA",X"AD",X"11",X"D1",X"EA",X"AA",X"11",X"D1",X"EE",X"AD",
		X"11",X"D1",X"AA",X"D0",X"11",X"99",X"AA",X"00",X"66",X"9A",X"AA",X"00",X"66",X"AA",X"AA",X"00",
		X"99",X"AA",X"AD",X"00",X"AA",X"AA",X"DD",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"50",X"00",X"00",X"0D",X"55",X"00",X"00",X"D9",X"00",X"10",X"00",X"99",X"00",X"99",
		X"00",X"91",X"00",X"11",X"00",X"D9",X"55",X"71",X"00",X"99",X"11",X"D1",X"00",X"FF",X"99",X"D1",
		X"00",X"AA",X"D9",X"D9",X"00",X"AA",X"9D",X"D9",X"00",X"AA",X"99",X"99",X"00",X"AA",X"19",X"9B",
		X"00",X"1A",X"19",X"BD",X"00",X"1A",X"19",X"D9",X"00",X"1A",X"19",X"99",X"00",X"AA",X"19",X"99",
		X"00",X"AA",X"99",X"9D",X"00",X"AF",X"99",X"D1",X"00",X"AA",X"DD",X"10",X"00",X"AF",X"1D",X"10",
		X"00",X"11",X"D1",X"00",X"00",X"0D",X"10",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"00",X"00",X"A7",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"A7",X"EE",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"A8",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"0A",X"88",X"88",X"88",X"1A",X"88",X"88",X"88",X"1A",X"88",X"88",X"88",X"1A",X"58",X"88",
		X"88",X"15",X"55",X"88",X"88",X"15",X"55",X"88",X"88",X"55",X"11",X"88",X"88",X"15",X"11",X"88",
		X"88",X"15",X"55",X"18",X"88",X"15",X"B5",X"18",X"81",X"15",X"5B",X"A8",X"8A",X"15",X"5A",X"A8",
		X"8A",X"15",X"1A",X"88",X"81",X"15",X"5A",X"88",X"88",X"15",X"5A",X"88",X"88",X"15",X"11",X"88",
		X"88",X"15",X"81",X"88",X"88",X"A5",X"88",X"88",X"88",X"A5",X"18",X"88",X"88",X"A5",X"A1",X"88",
		X"88",X"A5",X"AA",X"88",X"88",X"A5",X"AA",X"88",X"88",X"15",X"11",X"88",X"88",X"81",X"88",X"88",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"06",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",
		X"00",X"00",X"00",X"6E",X"00",X"00",X"05",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"11",X"6E",
		X"00",X"00",X"11",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"10",X"6E",X"00",X"00",X"11",X"6E",
		X"00",X"00",X"01",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"40",X"6E",X"00",X"00",X"46",X"6E",
		X"00",X"00",X"46",X"6E",X"00",X"00",X"06",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"11",X"6E",X"00",X"00",X"01",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",
		X"00",X"11",X"00",X"6E",X"00",X"13",X"00",X"6E",X"00",X"10",X"06",X"6E",X"00",X"1F",X"66",X"6E",
		X"00",X"41",X"00",X"6E",X"00",X"41",X"00",X"6E",X"00",X"44",X"00",X"6E",X"00",X"44",X"10",X"6E",
		X"00",X"44",X"40",X"6E",X"00",X"07",X"40",X"6E",X"00",X"07",X"40",X"6E",X"00",X"01",X"41",X"6E",
		X"00",X"11",X"44",X"6E",X"00",X"AA",X"44",X"6E",X"00",X"4D",X"44",X"6E",X"00",X"44",X"44",X"6E",
		X"00",X"44",X"14",X"6E",X"00",X"14",X"01",X"6E",X"00",X"01",X"41",X"6E",X"00",X"00",X"46",X"6E",
		X"00",X"00",X"46",X"6E",X"00",X"00",X"06",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"11",X"6E",X"00",X"00",X"01",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",
		X"00",X"11",X"00",X"6E",X"00",X"13",X"00",X"6E",X"00",X"43",X"06",X"6E",X"00",X"10",X"66",X"6E",
		X"00",X"4F",X"00",X"6E",X"00",X"41",X"00",X"6E",X"04",X"44",X"00",X"6E",X"04",X"44",X"10",X"6E",
		X"01",X"71",X"40",X"6E",X"00",X"70",X"40",X"6E",X"00",X"00",X"40",X"6E",X"00",X"01",X"41",X"6E",
		X"00",X"1A",X"44",X"6E",X"00",X"AD",X"44",X"6E",X"00",X"AD",X"44",X"6E",X"00",X"41",X"44",X"6E",
		X"00",X"44",X"14",X"6E",X"00",X"44",X"01",X"6E",X"00",X"14",X"41",X"6E",X"00",X"11",X"46",X"6E",
		X"00",X"00",X"46",X"6E",X"00",X"00",X"06",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"6E",
		X"00",X"00",X"11",X"6E",X"00",X"00",X"01",X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E6",X"00",X"00",X"66",X"60",X"00",
		X"00",X"66",X"60",X"0D",X"00",X"6A",X"66",X"E0",X"00",X"60",X"EE",X"E0",X"00",X"AA",X"66",X"EE",
		X"00",X"60",X"66",X"EE",X"00",X"6A",X"E6",X"EE",X"00",X"6A",X"66",X"EE",X"00",X"6A",X"0E",X"EE",
		X"00",X"A0",X"D0",X"EE",X"00",X"00",X"00",X"6E",X"00",X"A0",X"0A",X"6E",X"00",X"A0",X"AA",X"EE",
		X"00",X"66",X"A0",X"EE",X"00",X"66",X"AA",X"60",X"00",X"66",X"AA",X"60",X"00",X"AA",X"AA",X"60",
		X"00",X"66",X"0A",X"60",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"0F",X"FB",X"00",
		X"00",X"0F",X"FB",X"00",X"00",X"0F",X"BA",X"00",X"00",X"0F",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"06",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"7A",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0F",X"99",X"00",X"00",X"0F",X"09",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"09",X"00",X"00",X"0F",X"99",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"06",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"FB",X"00",
		X"00",X"0F",X"BB",X"00",X"00",X"0F",X"B5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"06",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"FB",X"00",X"00",X"0F",X"FB",X"00",
		X"00",X"0F",X"BB",X"00",X"00",X"0F",X"B5",X"00",X"00",X"0F",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"06",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",
		X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",
		X"00",X"00",X"30",X"09",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"39",X"00",X"00",X"33",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"30",X"00",X"99",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"99",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",
		X"33",X"90",X"00",X"00",X"99",X"00",X"03",X"00",X"00",X"00",X"39",X"00",X"33",X"33",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",
		X"00",X"30",X"00",X"33",X"00",X"30",X"00",X"99",X"00",X"33",X"00",X"09",X"00",X"99",X"00",X"09",
		X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"33",X"00",X"00",X"03",X"99",X"00",X"00",X"03",X"90",X"00",
		X"03",X"33",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"99",X"00",X"39",X"33",X"00",X"00",X"99",X"99",X"00",X"03",X"90",
		X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"00",
		X"00",X"33",X"00",X"00",X"33",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"0A",X"00",X"00",X"09",X"AA",
		X"00",X"00",X"09",X"0E",X"00",X"00",X"9B",X"00",X"00",X"90",X"99",X"90",X"00",X"09",X"09",X"99",
		X"00",X"99",X"99",X"99",X"00",X"9B",X"B9",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"09",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"90",X"99",X"00",X"90",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"99",X"9B",X"B9",X"00",X"00",X"09",X"99",X"00",X"00",X"90",X"99",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AF",X"A0",X"00",X"60",X"AA",X"A0",X"00",X"0A",X"00",X"A0",
		X"06",X"6A",X"00",X"00",X"00",X"AA",X"00",X"0A",X"00",X"00",X"70",X"6A",X"00",X"00",X"00",X"0A",
		X"F0",X"60",X"60",X"0A",X"00",X"00",X"70",X"70",X"66",X"67",X"00",X"00",X"00",X"77",X"00",X"00",
		X"0A",X"00",X"00",X"06",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"77",X"00",X"07",X"00",X"07",
		X"66",X"00",X"0F",X"77",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"66",X"60",X"66",X"0A",X"00",X"00",X"77",X"00",
		X"00",X"A0",X"77",X"AA",X"00",X"00",X"07",X"A0",X"00",X"A0",X"67",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"6A",X"6A",X"06",X"00",X"0A",X"AA",X"00",X"00",X"60",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"06",X"06",X"A0",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"F0",X"00",X"00",X"7A",X"77",X"00",
		X"00",X"00",X"FA",X"00",X"00",X"00",X"FA",X"00",X"00",X"A0",X"FA",X"00",X"00",X"77",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"00",X"00",X"0F",X"00",X"00",X"E0",X"F6",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"06",X"76",X"00",X"00",X"00",X"07",X"00",X"00",X"A7",X"FA",X"60",X"00",X"0A",X"7F",X"00",
		X"00",X"6F",X"77",X"00",X"00",X"00",X"70",X"06",X"00",X"7F",X"AA",X"00",X"00",X"67",X"0F",X"00",
		X"00",X"06",X"F6",X"00",X"00",X"0A",X"00",X"00",X"60",X"A0",X"60",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"00",X"C0",X"00",X"77",
		X"00",X"CC",X"66",X"77",X"00",X"66",X"55",X"7A",X"00",X"66",X"55",X"1A",X"00",X"06",X"55",X"5A",
		X"00",X"06",X"55",X"AA",X"00",X"0C",X"55",X"AA",X"00",X"0C",X"55",X"AA",X"66",X"0C",X"35",X"AA",
		X"5C",X"0C",X"33",X"AA",X"55",X"CD",X"33",X"AA",X"55",X"CD",X"33",X"AA",X"55",X"CD",X"30",X"AA",
		X"AA",X"CD",X"30",X"AA",X"AA",X"CD",X"30",X"AA",X"1A",X"CD",X"30",X"A1",X"1A",X"CD",X"11",X"A1",
		X"1A",X"CD",X"11",X"A1",X"0A",X"C1",X"11",X"A1",X"0A",X"C1",X"01",X"A1",X"0A",X"00",X"01",X"A1",
		X"0A",X"00",X"01",X"A1",X"0A",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A1",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"60",X"00",X"A0",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"07",X"00",X"00",X"00",
		X"07",X"A0",X"70",X"00",X"00",X"6D",X"27",X"00",X"3A",X"3D",X"AA",X"00",X"3A",X"3D",X"7A",X"00",
		X"3A",X"3D",X"77",X"00",X"AA",X"DD",X"07",X"00",X"AA",X"DD",X"00",X"60",X"AA",X"DD",X"AA",X"60",
		X"AC",X"DD",X"3A",X"66",X"AC",X"D3",X"5A",X"66",X"A5",X"D3",X"5A",X"56",X"A6",X"D3",X"5A",X"55",
		X"A1",X"DD",X"5A",X"55",X"A1",X"DD",X"6A",X"55",X"A1",X"DD",X"6A",X"50",X"A1",X"1D",X"6A",X"00",
		X"A1",X"1D",X"66",X"00",X"A1",X"1D",X"66",X"00",X"A1",X"1D",X"60",X"00",X"A1",X"1D",X"60",X"00",
		X"A0",X"1D",X"00",X"00",X"A0",X"1D",X"00",X"00",X"A0",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"00",X"00",X"0D",X"44",X"00",X"00",X"DC",X"AA",X"00",
		X"00",X"DA",X"0A",X"00",X"00",X"EA",X"F0",X"00",X"00",X"E0",X"FF",X"00",X"00",X"E0",X"FF",X"CC",
		X"0C",X"C0",X"FF",X"CC",X"CC",X"C0",X"FF",X"EE",X"CC",X"C0",X"55",X"00",X"E0",X"E0",X"50",X"00",
		X"00",X"EA",X"00",X"00",X"00",X"EE",X"0A",X"00",X"00",X"06",X"AE",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"06",X"0E",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"6E",X"00",
		X"00",X"0E",X"61",X"00",X"00",X"00",X"16",X"00",X"00",X"0E",X"1E",X"00",X"00",X"0E",X"1E",X"00",
		X"00",X"66",X"6E",X"00",X"00",X"66",X"00",X"09",X"00",X"66",X"00",X"09",X"00",X"11",X"00",X"99",
		X"00",X"00",X"01",X"9A",X"00",X"00",X"11",X"AA",X"00",X"00",X"77",X"AA",X"00",X"0E",X"91",X"4A",
		X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"54",X"00",X"0E",X"09",X"54",X"00",X"1E",X"07",X"44",
		X"00",X"71",X"74",X"44",X"01",X"44",X"44",X"44",X"11",X"44",X"44",X"41",X"14",X"44",X"45",X"11",
		X"4A",X"44",X"44",X"10",X"AA",X"44",X"44",X"00",X"AA",X"44",X"00",X"00",X"11",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"E0",X"60",
		X"00",X"00",X"E0",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"6E",X"00",X"00",X"EE",X"E6",X"00",
		X"00",X"00",X"E6",X"00",X"00",X"0A",X"E1",X"00",X"00",X"07",X"E1",X"00",X"00",X"00",X"E1",X"00",
		X"00",X"66",X"E6",X"00",X"00",X"66",X"60",X"00",X"00",X"16",X"10",X"00",X"00",X"01",X"90",X"00",
		X"00",X"00",X"A9",X"00",X"00",X"00",X"A9",X"00",X"00",X"11",X"A9",X"00",X"00",X"14",X"67",X"00",
		X"00",X"47",X"E6",X"10",X"00",X"79",X"0E",X"10",X"00",X"19",X"0E",X"11",X"00",X"77",X"60",X"41",
		X"00",X"41",X"77",X"41",X"00",X"44",X"11",X"11",X"00",X"44",X"44",X"10",X"00",X"44",X"44",X"00",
		X"00",X"14",X"44",X"00",X"00",X"11",X"44",X"00",X"00",X"01",X"A4",X"00",X"00",X"00",X"11",X"00",
		X"00",X"E1",X"00",X"00",X"00",X"6E",X"10",X"00",X"00",X"1E",X"11",X"00",X"00",X"16",X"E6",X"00",
		X"00",X"11",X"66",X"00",X"00",X"1E",X"6E",X"00",X"00",X"1E",X"EE",X"00",X"00",X"1E",X"E6",X"00",
		X"00",X"01",X"E1",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"E1",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"6E",X"00",
		X"00",X"AA",X"1E",X"90",X"00",X"A0",X"16",X"90",X"00",X"A0",X"06",X"09",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"AA",X"00",X"55",X"55",X"AA",X"00",X"55",X"55",X"AA",X"00",X"55",X"50",X"AA",
		X"00",X"A5",X"06",X"AA",X"00",X"AA",X"66",X"99",X"00",X"AA",X"AA",X"00",X"00",X"0A",X"A9",X"00",
		X"00",X"1A",X"90",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"06",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"AE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"7E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"7E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E7",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"00",X"DD",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"B2",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"22",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E1",X"00",X"00",X"00",X"6E",X"10",X"00",X"00",X"1E",X"11",X"00",X"00",X"16",X"E6",X"00",
		X"00",X"11",X"66",X"00",X"00",X"1E",X"6E",X"00",X"00",X"1E",X"EE",X"00",X"00",X"1E",X"E6",X"00",
		X"00",X"01",X"E1",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"E1",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"6E",X"00",
		X"00",X"AA",X"1E",X"90",X"00",X"A0",X"16",X"90",X"00",X"00",X"06",X"09",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"AA",X"00",X"AA",X"55",X"AA",X"00",X"AA",X"55",X"AA",X"00",X"1A",X"50",X"AA",
		X"00",X"01",X"06",X"AA",X"00",X"00",X"06",X"99",X"00",X"00",X"6A",X"00",X"00",X"00",X"A9",X"00",
		X"00",X"01",X"90",X"00",X"00",X"11",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"65",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"6E",X"10",X"00",X"00",X"1E",X"11",
		X"00",X"00",X"16",X"E6",X"00",X"00",X"11",X"66",X"00",X"00",X"1E",X"6E",X"00",X"00",X"1E",X"EE",
		X"00",X"00",X"1E",X"E6",X"00",X"00",X"01",X"E1",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"00",X"00",X"DC",X"EE",
		X"00",X"00",X"DC",X"6E",X"00",X"00",X"DD",X"6E",X"00",X"09",X"0D",X"60",X"00",X"99",X"DD",X"0C",
		X"00",X"09",X"00",X"CC",X"00",X"D9",X"DD",X"CD",X"99",X"D0",X"0D",X"DD",X"99",X"E9",X"DD",X"DC",
		X"00",X"99",X"DD",X"D9",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"88",X"88",X"80",X"77",X"77",X"88",X"80",X"78",X"88",X"88",X"80",X"F8",X"FF",X"88",
		X"80",X"F8",X"77",X"88",X"80",X"F8",X"88",X"88",X"80",X"F8",X"FF",X"88",X"80",X"F8",X"77",X"88",
		X"80",X"F8",X"88",X"88",X"80",X"77",X"77",X"88",X"88",X"77",X"77",X"88",X"88",X"80",X"88",X"88",
		X"88",X"00",X"88",X"88",X"88",X"0B",X"88",X"88",X"88",X"BB",X"38",X"88",X"88",X"8B",X"33",X"88",
		X"88",X"B8",X"38",X"88",X"88",X"BB",X"88",X"88",X"88",X"88",X"33",X"88",X"88",X"DD",X"33",X"88",
		X"88",X"D3",X"33",X"88",X"88",X"DD",X"33",X"88",X"88",X"D3",X"38",X"88",X"88",X"BD",X"88",X"88",
		X"88",X"88",X"33",X"88",X"88",X"DD",X"33",X"88",X"88",X"DD",X"33",X"88",X"88",X"DD",X"33",X"88",
		X"88",X"DD",X"33",X"88",X"88",X"DD",X"33",X"88",X"88",X"DD",X"38",X"88",X"88",X"83",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"55",X"30",X"00",X"00",X"55",X"EE",
		X"00",X"00",X"55",X"5E",X"00",X"00",X"E5",X"5E",X"00",X"05",X"E5",X"E5",X"00",X"51",X"EE",X"5E",
		X"00",X"55",X"EE",X"55",X"00",X"55",X"E5",X"55",X"00",X"55",X"E5",X"55",X"00",X"05",X"E5",X"55",
		X"00",X"05",X"E5",X"55",X"00",X"55",X"65",X"55",X"00",X"55",X"65",X"55",X"00",X"55",X"65",X"55",
		X"00",X"51",X"66",X"56",X"00",X"04",X"65",X"64",X"00",X"00",X"65",X"56",X"00",X"00",X"55",X"56",
		X"00",X"00",X"45",X"66",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",
		X"00",X"50",X"53",X"E3",X"00",X"55",X"E5",X"5E",X"00",X"15",X"E5",X"5E",X"00",X"15",X"E5",X"55",
		X"00",X"11",X"EE",X"EE",X"0E",X"61",X"E5",X"55",X"0E",X"61",X"E5",X"55",X"55",X"61",X"E5",X"55",
		X"44",X"61",X"E5",X"55",X"06",X"61",X"65",X"55",X"0E",X"61",X"65",X"55",X"00",X"11",X"66",X"66",
		X"00",X"15",X"65",X"55",X"00",X"15",X"65",X"56",X"00",X"55",X"64",X"46",X"00",X"50",X"44",X"64",
		X"00",X"00",X"40",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"0E",X"66",X"00",X"00",X"0E",X"66",X"00",X"00",X"55",X"66",X"00",
		X"00",X"44",X"66",X"00",X"00",X"06",X"61",X"00",X"00",X"0E",X"16",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"06",X"60",X"00",X"00",X"60",X"60",X"00",
		X"00",X"60",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"66",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A6",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",X"00",X"06",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7E",X"06",X"EE",X"00",X"00",X"00",X"00",X"00",X"E1",X"0E",X"E6",X"00",X"00",X"00",X"00",
		X"00",X"6E",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"0E",X"0A",X"00",X"00",X"00",X"00",X"AA",X"EA",X"AE",X"AA",X"00",X"00",X"00",X"00",
		X"CA",X"CA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"A9",X"9C",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"B0",X"9B",X"00",X"00",X"0B",X"CF",X"00",X"00",X"99",X"9F",X"00",
		X"00",X"D0",X"F9",X"00",X"00",X"DD",X"F9",X"00",X"00",X"9B",X"99",X"00",X"00",X"09",X"9B",X"00",
		X"00",X"00",X"9F",X"00",X"99",X"99",X"9C",X"99",X"FB",X"F9",X"FF",X"BF",X"99",X"9F",X"F9",X"99",
		X"09",X"D9",X"9D",X"DB",X"00",X"99",X"DD",X"99",X"00",X"00",X"9D",X"00",X"00",X"99",X"09",X"00",
		X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"C9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"9D",X"00",X"00",X"90",X"D9",X"09",X"00",X"90",X"90",
		X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"00",X"00",X"99",X"90",X"B0",X"00",X"9F",X"90",X"00",
		X"00",X"B0",X"99",X"00",X"00",X"9B",X"9B",X"00",X"00",X"9B",X"CC",X"00",X"00",X"99",X"F9",X"90",
		X"00",X"09",X"9B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"CF",X"B9",
		X"00",X"09",X"BC",X"99",X"00",X"0C",X"99",X"F9",X"00",X"99",X"99",X"9F",X"00",X"D9",X"90",X"B9",
		X"00",X"9D",X"90",X"99",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"00",X"10",X"00",X"07",X"00",X"01",X"00",X"07",
		X"00",X"00",X"06",X"07",X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"10",X"F0",X"00",X"00",X"10",X"00",X"00",X"70",X"01",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"02",X"BB",X"00",
		X"00",X"B2",X"00",X"B0",X"BB",X"02",X"00",X"0B",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"22",X"02",X"00",X"02",X"00",X"22",X"0B",X"20",
		X"00",X"00",X"22",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"F0",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"E6",X"00",X"00",X"08",X"16",X"00",X"00",X"08",X"21",
		X"00",X"00",X"08",X"44",X"00",X"00",X"08",X"44",X"00",X"00",X"08",X"42",X"00",X"00",X"08",X"14",
		X"00",X"00",X"08",X"02",X"00",X"00",X"88",X"04",X"00",X"00",X"80",X"01",X"00",X"00",X"80",X"08",
		X"00",X"00",X"80",X"10",X"00",X"00",X"EE",X"10",X"00",X"00",X"11",X"11",X"00",X"0A",X"11",X"11",
		X"00",X"AA",X"11",X"11",X"00",X"AA",X"11",X"21",X"00",X"AA",X"91",X"22",X"00",X"AE",X"99",X"42",
		X"00",X"EE",X"A9",X"44",X"00",X"EE",X"AA",X"44",X"00",X"EA",X"AA",X"46",X"00",X"DD",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"8E",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"22",X"00",X"00",X"08",X"21",X"00",X"00",X"08",X"24",
		X"00",X"00",X"08",X"24",X"00",X"00",X"08",X"24",X"00",X"00",X"08",X"22",X"00",X"00",X"08",X"24",
		X"00",X"00",X"08",X"28",X"00",X"00",X"88",X"81",X"00",X"00",X"80",X"24",X"00",X"00",X"80",X"48",
		X"00",X"00",X"80",X"40",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",X"11",X"00",X"0A",X"11",X"11",
		X"00",X"AA",X"11",X"11",X"00",X"AA",X"11",X"44",X"00",X"AA",X"91",X"22",X"00",X"AE",X"99",X"42",
		X"00",X"EE",X"A9",X"44",X"00",X"EE",X"AA",X"11",X"00",X"EA",X"AA",X"46",X"00",X"DD",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"82",
		X"00",X"00",X"00",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"84",X"00",X"00",X"0E",X"80",X"00",X"00",X"11",X"80",X"00",X"0A",X"11",X"80",
		X"00",X"AA",X"11",X"80",X"00",X"AA",X"11",X"28",X"00",X"AA",X"91",X"22",X"00",X"AE",X"99",X"42",
		X"00",X"EE",X"A9",X"44",X"00",X"EE",X"AA",X"84",X"00",X"EA",X"AA",X"86",X"00",X"DD",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"66",X"02",X"00",X"00",X"61",X"22",X"00",X"00",
		X"22",X"24",X"00",X"00",X"12",X"21",X"00",X"00",X"F1",X"20",X"00",X"00",X"FF",X"20",X"00",X"00",
		X"FF",X"40",X"00",X"00",X"FF",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"24",X"10",X"00",X"00",
		X"24",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"44",X"E0",X"00",X"00",X"14",X"1E",X"00",X"00",X"14",X"11",X"E0",X"00",X"42",X"11",X"AA",X"00",
		X"42",X"11",X"AA",X"00",X"22",X"81",X"AA",X"00",X"24",X"81",X"AA",X"00",X"44",X"81",X"EE",X"00",
		X"44",X"99",X"EE",X"00",X"46",X"9A",X"AA",X"00",X"66",X"AA",X"AA",X"00",X"99",X"AA",X"AD",X"00",
		X"9A",X"AA",X"DD",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"DD",X"00",X"00",X"DD",X"D0",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"C0",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"D0",X"00",X"0C",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CD",
		X"00",X"00",X"00",X"D0",X"00",X"C0",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"D0",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"D0",X"00",X"00",X"00",X"0C",X"0D",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"D0",X"0C",X"00",X"00",X"DD",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"0C",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"0C",X"00",X"0D",X"DD",X"00",X"00",
		X"CC",X"D0",X"09",X"00",X"0C",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"0D",X"00",X"CD",X"00",X"00",X"00",X"0D",X"90",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",
		X"00",X"00",X"DC",X"00",X"00",X"00",X"00",X"CD",X"00",X"00",X"0C",X"0C",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"CD",X"00",X"D0",X"09",X"00",X"00",X"CD",X"00",X"90",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"CD",X"00",X"00",X"C0",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"0C",
		X"CC",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"DC",X"00",X"C0",X"0D",X"00",X"0D",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"02",X"66",X"00",X"00",
		X"02",X"22",X"00",X"00",X"02",X"66",X"00",X"00",X"02",X"F6",X"00",X"00",X"08",X"F2",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"02",X"41",X"00",X"00",
		X"02",X"21",X"00",X"00",X"02",X"12",X"00",X"00",X"04",X"22",X"00",X"00",X"04",X"24",X"22",X"00",
		X"08",X"11",X"20",X"00",X"08",X"00",X"00",X"00",X"08",X"22",X"40",X"00",X"42",X"44",X"22",X"00",
		X"22",X"00",X"22",X"00",X"48",X"00",X"22",X"01",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"20",
		X"00",X"00",X"22",X"40",X"00",X"00",X"22",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"02",X"66",X"00",X"00",
		X"02",X"22",X"00",X"00",X"02",X"66",X"00",X"00",X"02",X"F6",X"00",X"00",X"08",X"F2",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"02",X"41",X"00",X"00",
		X"02",X"21",X"00",X"00",X"02",X"12",X"00",X"00",X"04",X"22",X"22",X"00",X"04",X"24",X"41",X"00",
		X"08",X"11",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"40",X"00",X"00",X"00",X"22",X"00",
		X"08",X"00",X"22",X"00",X"08",X"02",X"22",X"01",X"00",X"02",X"22",X"24",X"00",X"02",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"11",X"22",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"02",X"66",X"00",X"00",
		X"02",X"22",X"00",X"00",X"02",X"66",X"00",X"00",X"02",X"F6",X"00",X"00",X"08",X"F2",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"22",X"00",X"00",X"04",X"12",X"00",X"00",X"02",X"41",X"00",X"00",
		X"02",X"21",X"00",X"00",X"02",X"12",X"24",X"00",X"04",X"22",X"22",X"00",X"04",X"24",X"12",X"40",
		X"08",X"11",X"21",X"40",X"08",X"00",X"21",X"21",X"08",X"00",X"21",X"21",X"00",X"00",X"21",X"22",
		X"00",X"00",X"21",X"24",X"00",X"00",X"24",X"41",X"00",X"00",X"24",X"11",X"00",X"02",X"22",X"40",
		X"00",X"02",X"22",X"40",X"00",X"22",X"21",X"24",X"00",X"42",X"21",X"22",X"00",X"42",X"24",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"EE",
		X"00",X"00",X"80",X"11",X"00",X"00",X"EE",X"11",X"00",X"00",X"11",X"11",X"00",X"0A",X"11",X"11",
		X"00",X"AA",X"11",X"11",X"00",X"AA",X"11",X"11",X"00",X"AA",X"91",X"11",X"00",X"AE",X"99",X"11",
		X"00",X"EE",X"A9",X"11",X"00",X"EE",X"AA",X"11",X"00",X"EA",X"AA",X"16",X"00",X"DD",X"AA",X"99",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"DA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"00",X"DD",
		X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"88",X"AA",X"00",X"00",X"08",X"FA",X"00",X"00",X"0A",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"EE",X"AA",X"AA",X"00",X"11",X"1A",X"AA",X"00",
		X"11",X"E1",X"AA",X"00",X"11",X"1E",X"A1",X"00",X"11",X"11",X"A1",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"A1",X"D0",X"11",X"11",X"AA",X"D0",X"11",X"11",X"EE",X"00",
		X"11",X"99",X"EE",X"00",X"16",X"9A",X"AA",X"00",X"66",X"AA",X"AA",X"00",X"99",X"AA",X"AD",X"00",
		X"9A",X"AA",X"DD",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"DD",X"00",X"00",X"DD",X"D0",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"53",X"00",X"00",X"05",X"55",X"00",X"00",X"05",X"55",X"00",
		X"00",X"05",X"05",X"00",X"00",X"D5",X"59",X"00",X"00",X"95",X"50",X"00",X"00",X"55",X"50",X"70",
		X"00",X"11",X"51",X"D0",X"00",X"99",X"11",X"D0",X"0D",X"99",X"19",X"DD",X"0D",X"F9",X"11",X"99",
		X"0D",X"F9",X"91",X"99",X"0D",X"F1",X"DD",X"9B",X"01",X"A1",X"DD",X"BD",X"01",X"A1",X"D9",X"D9",
		X"00",X"AA",X"1D",X"99",X"00",X"1A",X"91",X"99",X"00",X"A1",X"99",X"9D",X"00",X"A1",X"99",X"D1",
		X"00",X"11",X"99",X"10",X"00",X"11",X"91",X"00",X"00",X"19",X"DD",X"00",X"00",X"19",X"11",X"00",
		X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"88",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"77",X"09",X"99",X"09",
		X"00",X"00",X"00",X"00",X"77",X"66",X"99",X"00",X"00",X"00",X"00",X"00",X"A7",X"00",X"09",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8A",X"88",X"88",X"88",X"8A",X"88",X"88",X"88",X"AA",X"88",X"88",X"88",X"AA",X"88",X"88",
		X"88",X"A9",X"88",X"88",X"8A",X"AA",X"88",X"88",X"8A",X"9A",X"88",X"88",X"8A",X"9A",X"88",X"88",
		X"81",X"9A",X"51",X"88",X"81",X"95",X"B5",X"88",X"81",X"95",X"55",X"88",X"85",X"95",X"15",X"88",
		X"85",X"95",X"11",X"88",X"15",X"95",X"51",X"88",X"AA",X"95",X"AA",X"88",X"AA",X"95",X"BB",X"88",
		X"11",X"95",X"AA",X"88",X"88",X"95",X"AA",X"88",X"88",X"95",X"AA",X"88",X"88",X"95",X"AA",X"88",
		X"88",X"95",X"11",X"88",X"88",X"95",X"88",X"88",X"88",X"95",X"88",X"88",X"88",X"95",X"88",X"88",
		X"88",X"95",X"18",X"88",X"88",X"9A",X"A8",X"88",X"88",X"55",X"18",X"88",X"88",X"55",X"88",X"88",
		X"88",X"11",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"EE",X"00",X"00",X"66",X"1E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"50",X"EE",X"00",X"00",X"51",X"EE",X"00",X"00",X"01",X"1E",X"00",X"00",X"11",X"EE",
		X"00",X"00",X"11",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"11",X"EE",
		X"00",X"00",X"11",X"EE",X"00",X"00",X"10",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"1E",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"EE",X"00",X"01",X"66",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"11",X"1E",X"00",X"00",X"01",X"EE",X"00",X"00",X"00",X"E1",
		X"00",X"33",X"00",X"00",X"00",X"33",X"06",X"EE",X"00",X"00",X"66",X"1E",X"00",X"0F",X"00",X"EE",
		X"00",X"FF",X"00",X"EE",X"04",X"11",X"00",X"EE",X"44",X"14",X"00",X"EE",X"44",X"44",X"00",X"EE",
		X"17",X"44",X"00",X"EE",X"07",X"11",X"00",X"EE",X"00",X"11",X"00",X"1E",X"00",X"AA",X"00",X"EE",
		X"00",X"A1",X"00",X"EE",X"00",X"A1",X"00",X"EE",X"00",X"D1",X"00",X"EE",X"00",X"44",X"40",X"EE",
		X"00",X"44",X"44",X"EE",X"00",X"41",X"44",X"EE",X"00",X"11",X"41",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"1E",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"EE",X"00",X"01",X"66",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"11",X"1E",X"00",X"00",X"01",X"EE",X"00",X"00",X"00",X"E1",
		X"00",X"33",X"00",X"00",X"00",X"33",X"06",X"EE",X"00",X"FF",X"66",X"1E",X"00",X"0F",X"00",X"EE",
		X"04",X"0F",X"00",X"EE",X"44",X"FF",X"00",X"EE",X"44",X"14",X"00",X"EE",X"44",X"44",X"00",X"EE",
		X"71",X"44",X"00",X"EE",X"70",X"14",X"00",X"EE",X"00",X"11",X"00",X"1E",X"00",X"A1",X"00",X"EE",
		X"00",X"DD",X"00",X"EE",X"00",X"1D",X"00",X"EE",X"00",X"71",X"00",X"EE",X"00",X"74",X"40",X"EE",
		X"00",X"44",X"44",X"EE",X"00",X"44",X"44",X"EE",X"00",X"44",X"41",X"EE",X"00",X"11",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"1E",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"EE",X"00",X"01",X"66",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"11",X"1E",X"00",X"00",X"01",X"EE",X"00",X"00",X"00",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"66",X"00",X"00",X"66",X"06",X"00",
		X"00",X"E6",X"00",X"0D",X"00",X"00",X"0D",X"00",X"00",X"E6",X"66",X"0D",X"00",X"A6",X"6E",X"00",
		X"00",X"AA",X"6E",X"00",X"C0",X"66",X"6E",X"00",X"00",X"CA",X"6E",X"00",X"00",X"AA",X"66",X"00",
		X"00",X"AA",X"66",X"0D",X"00",X"0A",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"06",X"00",X"00",X"A0",X"AA",X"00",X"00",X"AA",X"AA",X"0D",X"00",X"AA",X"00",X"00",
		X"00",X"6A",X"00",X"00",X"00",X"6A",X"0A",X"00",X"00",X"66",X"AA",X"D0",X"00",X"06",X"66",X"00",
		X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0B",X"FB",X"00",X"00",X"B0",X"FB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"B5",X"00",X"00",X"99",X"B5",X"00",X"00",X"FF",X"B5",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"A5",X"00",X"00",X"FB",X"A5",X"00",
		X"00",X"BB",X"55",X"00",X"00",X"05",X"A5",X"00",X"00",X"60",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0A",X"FB",X"00",X"00",X"AF",X"FB",X"00",
		X"00",X"FF",X"BB",X"00",X"00",X"FF",X"B5",X"00",X"00",X"FF",X"95",X"00",X"00",X"FF",X"95",X"00",
		X"00",X"FF",X"95",X"00",X"00",X"FF",X"95",X"00",X"00",X"FF",X"55",X"00",X"00",X"FB",X"55",X"00",
		X"00",X"BB",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"60",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"FB",X"00",X"00",X"FF",X"FB",X"00",
		X"00",X"FF",X"BB",X"00",X"00",X"FF",X"B5",X"00",X"00",X"FF",X"B5",X"00",X"00",X"FF",X"B5",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"59",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"90",X"00",
		X"00",X"0B",X"90",X"00",X"00",X"05",X"99",X"00",X"00",X"60",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"FB",X"00",X"00",X"FF",X"FB",X"00",
		X"00",X"FF",X"BB",X"00",X"00",X"FF",X"B5",X"00",X"00",X"FF",X"B5",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FB",X"55",X"00",
		X"00",X"BB",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"60",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"90",X"03",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"99",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"99",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"03",X"00",X"99",X"00",X"39",X"00",X"00",X"00",X"90",X"00",X"33",X"33",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"33",X"00",X"33",X"00",X"99",X"00",X"93",
		X"00",X"00",X"30",X"99",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"93",X"30",X"00",X"00",X"99",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"03",X"00",
		X"99",X"00",X"33",X"00",X"00",X"00",X"39",X"00",X"00",X"33",X"99",X"00",X"00",X"99",X"00",X"00",
		X"33",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"30",X"33",X"99",X"00",X"90",X"39",X"00",X"00",X"00",X"99",X"00",X"33",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"99",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"9B",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"A5",X"00",X"00",X"B9",X"E5",X"00",X"00",X"99",X"05",
		X"00",X"90",X"90",X"AA",X"00",X"09",X"99",X"EE",X"00",X"90",X"99",X"00",X"00",X"0B",X"99",X"90",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"90",X"09",X"99",X"09",X"B9",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"9B",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"90",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"60",X"00",X"AA",X"00",X"00",
		X"66",X"FA",X"77",X"00",X"00",X"0A",X"07",X"0A",X"06",X"66",X"67",X"0A",X"00",X"07",X"77",X"A0",
		X"00",X"07",X"00",X"00",X"0A",X"07",X"00",X"00",X"60",X"00",X"00",X"0A",X"00",X"70",X"00",X"AA",
		X"A0",X"00",X"00",X"AA",X"0A",X"00",X"00",X"A0",X"0A",X"70",X"00",X"AA",X"0A",X"70",X"00",X"00",
		X"AA",X"00",X"00",X"6A",X"00",X"70",X"00",X"0A",X"0F",X"77",X"00",X"FA",X"00",X"70",X"00",X"AA",
		X"00",X"70",X"00",X"0A",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"AA",X"00",X"00",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",X"06",X"A0",X"77",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"07",
		X"00",X"00",X"F0",X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",X"00",X"0A",X"77",X"77",X"00",
		X"00",X"AF",X"0A",X"00",X"00",X"00",X"A7",X"00",X"00",X"AF",X"0A",X"00",X"0A",X"77",X"76",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F7",X"70",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"07",X"00",X"00",X"0A",X"00",X"E0",X"60",X"60",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"7A",X"6A",X"00",X"60",X"7A",X"A0",X"00",X"00",X"6F",X"67",X"00",X"00",X"FA",X"A0",X"00",
		X"00",X"77",X"FA",X"00",X"00",X"A7",X"00",X"00",X"00",X"67",X"F6",X"00",X"00",X"FA",X"A0",X"00",
		X"00",X"AF",X"A7",X"00",X"00",X"70",X"7A",X"00",X"00",X"07",X"76",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"7A",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"03",X"A0",X"00",X"00",X"AA",X"A0",
		X"00",X"C0",X"63",X"A5",X"00",X"C6",X"53",X"A5",X"06",X"C5",X"53",X"A5",X"00",X"C5",X"53",X"A5",
		X"00",X"CC",X"F3",X"A5",X"07",X"C3",X"33",X"A5",X"02",X"D3",X"33",X"A5",X"07",X"D3",X"33",X"55",
		X"02",X"DD",X"33",X"52",X"00",X"5D",X"03",X"52",X"AC",X"5D",X"33",X"52",X"AC",X"5D",X"33",X"62",
		X"AA",X"1D",X"33",X"12",X"AA",X"11",X"13",X"12",X"1A",X"11",X"13",X"12",X"1A",X"11",X"13",X"12",
		X"1A",X"11",X"11",X"12",X"0A",X"11",X"11",X"12",X"0A",X"11",X"11",X"12",X"00",X"01",X"11",X"12",
		X"00",X"00",X"11",X"02",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"77",X"0D",X"66",X"00",X"77",X"DD",X"06",X"00",
		X"A7",X"D0",X"00",X"00",X"A0",X"66",X"20",X"00",X"AC",X"56",X"72",X"00",X"AA",X"56",X"A7",X"00",
		X"AA",X"53",X"27",X"00",X"AA",X"3D",X"70",X"00",X"CA",X"3D",X"00",X"00",X"CA",X"3D",X"A5",X"00",
		X"5A",X"DD",X"AA",X"00",X"5A",X"DD",X"5A",X"00",X"5A",X"DD",X"5A",X"60",X"2A",X"D5",X"5A",X"60",
		X"2A",X"D5",X"5A",X"60",X"2A",X"D5",X"6A",X"00",X"2A",X"55",X"6A",X"00",X"21",X"55",X"6A",X"00",
		X"21",X"15",X"6A",X"00",X"21",X"15",X"1A",X"00",X"11",X"00",X"1A",X"00",X"11",X"00",X"1A",X"00",
		X"11",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"01",X"00",X"0A",X"00",X"11",X"00",X"0A",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D3",X"00",X"00",X"00",X"44",X"D0",X"00",X"00",X"AA",X"DD",X"00",
		X"00",X"A0",X"AD",X"00",X"00",X"0F",X"AE",X"00",X"00",X"FF",X"0E",X"00",X"0C",X"FF",X"0E",X"00",
		X"CC",X"FF",X"0C",X"CC",X"CC",X"FF",X"0C",X"EC",X"E0",X"55",X"0C",X"0E",X"00",X"05",X"0E",X"00",
		X"00",X"00",X"AE",X"00",X"00",X"A0",X"EE",X"00",X"00",X"EA",X"60",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",
		X"CE",X"00",X"00",X"00",X"CE",X"00",X"0E",X"00",X"CC",X"00",X"CC",X"00",X"0C",X"00",X"C0",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"E0",X"EE",X"00",X"00",X"6E",X"EE",X"EE",X"00",X"06",X"EE",X"E6",X"00",X"00",X"EE",X"16",X"00",
		X"00",X"00",X"6E",X"00",X"00",X"07",X"EE",X"09",X"00",X"0A",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"66",X"00",X"9A",X"00",X"66",X"00",X"9A",X"00",X"66",X"00",X"AA",X"00",X"16",X"00",X"AA",
		X"00",X"11",X"11",X"AA",X"00",X"01",X"44",X"AA",X"00",X"06",X"74",X"AA",X"00",X"E6",X"77",X"A9",
		X"00",X"00",X"99",X"44",X"00",X"E0",X"99",X"41",X"00",X"EE",X"97",X"41",X"00",X"1E",X"74",X"41",
		X"01",X"7E",X"44",X"11",X"14",X"41",X"44",X"10",X"44",X"44",X"45",X"10",X"44",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"11",X"00",X"A4",X"44",X"00",X"00",X"11",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"E6",X"EE",X"00",X"00",X"06",X"EE",X"0E",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"E1",X"00",
		X"00",X"E0",X"16",X"00",X"00",X"00",X"6E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"E0",X"00",
		X"00",X"66",X"E0",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"19",X"10",X"00",X"00",X"19",X"11",X"00",X"00",X"47",X"44",X"00",
		X"00",X"96",X"97",X"00",X"00",X"9E",X"99",X"00",X"01",X"EE",X"E9",X"00",X"01",X"90",X"97",X"00",
		X"01",X"77",X"71",X"00",X"01",X"11",X"14",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"41",X"00",X"00",X"14",X"11",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"E1",X"00",X"00",X"0E",X"E1",X"00",
		X"00",X"EE",X"E1",X"00",X"00",X"0E",X"61",X"00",X"00",X"00",X"10",X"00",X"00",X"07",X"10",X"00",
		X"00",X"E7",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"55",X"90",X"00",X"00",X"05",X"99",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"06",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"05",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"AA",X"00",X"55",X"06",X"AA",X"00",X"55",X"66",X"AA",
		X"00",X"53",X"6A",X"99",X"00",X"55",X"AA",X"00",X"00",X"55",X"AA",X"00",X"00",X"55",X"99",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"06",X"EE",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"06",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"DE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"42",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"44",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"09",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"E1",X"00",X"00",X"0E",X"E1",X"00",
		X"00",X"EE",X"E1",X"00",X"00",X"0E",X"61",X"00",X"00",X"00",X"10",X"00",X"00",X"07",X"10",X"00",
		X"00",X"E7",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"55",X"90",X"00",X"00",X"05",X"99",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"06",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"05",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"AA",X"00",X"A5",X"06",X"AA",X"00",X"AA",X"66",X"AA",
		X"00",X"AA",X"6A",X"99",X"00",X"1A",X"AA",X"00",X"00",X"1A",X"AA",X"00",X"00",X"1A",X"99",X"00",
		X"00",X"1A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"E1",
		X"00",X"00",X"0E",X"E1",X"00",X"00",X"EE",X"E1",X"00",X"00",X"0E",X"61",X"00",X"00",X"00",X"10",
		X"00",X"00",X"71",X"10",X"00",X"00",X"EE",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"CC",X"AC",X"00",X"00",X"6A",X"1A",
		X"00",X"00",X"A1",X"1A",X"00",X"E5",X"CC",X"1A",X"00",X"90",X"0C",X"1A",X"00",X"99",X"DD",X"CC",
		X"00",X"00",X"D0",X"DD",X"99",X"99",X"DD",X"C9",X"99",X"00",X"0D",X"90",X"99",X"99",X"DD",X"90",
		X"00",X"EE",X"DD",X"00",X"00",X"00",X"CC",X"0A",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"88",X"08",X"88",X"88",X"07",X"77",X"77",X"88",X"07",X"77",X"FA",X"88",X"07",X"77",X"F8",X"88",
		X"07",X"77",X"F8",X"88",X"07",X"77",X"F8",X"88",X"07",X"77",X"F8",X"88",X"07",X"77",X"F8",X"88",
		X"07",X"88",X"F8",X"88",X"07",X"77",X"77",X"88",X"07",X"77",X"77",X"88",X"80",X"08",X"88",X"88",
		X"80",X"08",X"88",X"88",X"80",X"08",X"88",X"88",X"80",X"88",X"88",X"88",X"88",X"B8",X"88",X"88",
		X"88",X"B3",X"88",X"88",X"88",X"BB",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"33",X"88",X"88",
		X"88",X"D3",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"D3",X"88",X"88",X"88",X"DB",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"D3",X"88",X"88",X"88",X"DD",X"88",X"88",X"88",X"D3",X"88",X"88",
		X"88",X"DD",X"88",X"88",X"88",X"D3",X"88",X"88",X"88",X"DD",X"88",X"88",X"88",X"33",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"55",X"00",X"00",X"03",X"55",X"30",
		X"00",X"35",X"55",X"30",X"00",X"55",X"55",X"53",X"00",X"55",X"5E",X"E5",X"00",X"55",X"E5",X"E5",
		X"00",X"15",X"55",X"E5",X"05",X"55",X"55",X"5E",X"05",X"55",X"55",X"5E",X"05",X"55",X"55",X"5E",
		X"05",X"55",X"55",X"5E",X"05",X"54",X"55",X"56",X"00",X"14",X"55",X"56",X"00",X"14",X"55",X"65",
		X"00",X"44",X"65",X"64",X"00",X"44",X"56",X"64",X"00",X"44",X"55",X"44",X"00",X"44",X"55",X"40",
		X"00",X"04",X"55",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"35",X"30",X"30",X"00",X"15",X"53",X"53",X"00",X"51",X"55",X"E5",X"0E",X"55",X"55",X"E5",
		X"EE",X"55",X"55",X"E5",X"E7",X"55",X"E5",X"5E",X"7E",X"45",X"5E",X"5E",X"EE",X"45",X"55",X"5E",
		X"EE",X"45",X"55",X"5E",X"E6",X"45",X"56",X"56",X"66",X"55",X"65",X"56",X"66",X"55",X"55",X"65",
		X"06",X"55",X"55",X"65",X"00",X"51",X"54",X"64",X"00",X"11",X"44",X"44",X"00",X"44",X"40",X"40",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"E7",X"60",X"00",X"00",X"7E",X"60",X"00",X"00",X"EE",X"55",X"00",
		X"00",X"EE",X"44",X"00",X"00",X"E6",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"06",X"60",X"00",
		X"00",X"60",X"06",X"00",X"00",X"6A",X"60",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"60",X"60",X"00",X"00",X"06",X"6A",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"EE",X"00",X"E6",X"00",X"00",X"00",X"00",
		X"01",X"E1",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"6E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"4E",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"4E",X"0E",X"0E",X"00",X"00",X"00",X"00",
		X"A0",X"EE",X"0E",X"6E",X"00",X"00",X"00",X"00",X"AA",X"EA",X"A0",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AC",X"AC",X"00",X"00",X"00",X"00",X"0C",X"C9",X"9A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"55",
		X"00",X"00",X"50",X"55",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"D0",X"00",X"00",X"00",X"09",X"00",X"99",X"00",
		X"9D",X"00",X"99",X"00",X"99",X"00",X"9F",X"00",X"00",X"00",X"9F",X"00",X"00",X"B0",X"9F",X"00",
		X"00",X"9B",X"9B",X"00",X"00",X"D9",X"FB",X"00",X"00",X"DC",X"FC",X"00",X"00",X"DC",X"BB",X"00",
		X"00",X"9B",X"C9",X"00",X"99",X"99",X"B9",X"90",X"BF",X"F9",X"FF",X"99",X"99",X"9F",X"99",X"99",
		X"DD",X"9B",X"DD",X"DD",X"99",X"9B",X"D9",X"99",X"00",X"99",X"DD",X"00",X"00",X"FB",X"DD",X"00",
		X"00",X"0B",X"9C",X"00",X"00",X"B9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"09",X"90",X"09",X"00",X"00",X"90",X"9B",X"00",
		X"00",X"F9",X"DD",X"00",X"00",X"B9",X"CC",X"00",X"00",X"BB",X"C9",X"00",X"00",X"9B",X"90",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"99",X"FF",X"00",X"00",X"09",X"99",X"99",X"00",X"9D",X"B9",X"00",
		X"00",X"DD",X"BF",X"90",X"00",X"DD",X"BC",X"90",X"00",X"9D",X"99",X"90",X"00",X"D0",X"09",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"10",X"66",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"10",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"07",X"00",X"00",X"70",X"70",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"60",X"07",X"00",X"10",X"60",X"70",X"70",X"10",X"60",X"00",X"07",X"10",X"60",X"00",X"00",X"70",
		X"67",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"BB",X"B0",X"00",
		X"0B",X"00",X"BB",X"00",X"B0",X"00",X"B0",X"BB",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"20",X"00",X"B0",X"22",X"02",X"20",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"8E",X"00",X"00",X"08",X"66",X"00",X"00",X"08",X"EE",X"00",X"00",X"08",X"6E",
		X"00",X"00",X"08",X"6E",X"00",X"00",X"08",X"66",X"00",X"00",X"88",X"66",X"00",X"00",X"88",X"61",
		X"00",X"00",X"88",X"62",X"00",X"00",X"88",X"12",X"00",X"00",X"80",X"22",X"00",X"00",X"80",X"22",
		X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"44",
		X"00",X"00",X"0E",X"01",X"00",X"00",X"E1",X"80",X"00",X"0E",X"11",X"88",X"00",X"AA",X"11",X"18",
		X"00",X"AA",X"12",X"12",X"00",X"AA",X"22",X"22",X"00",X"AA",X"22",X"22",X"00",X"EE",X"44",X"22",
		X"00",X"EE",X"99",X"C2",X"00",X"AA",X"A9",X"62",X"00",X"AA",X"AA",X"66",X"00",X"DA",X"AA",X"99",
		X"00",X"DD",X"AA",X"A9",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"08",X"8E",X"00",X"00",X"08",X"6E",X"00",X"00",X"08",X"66",X"00",X"00",X"08",X"26",
		X"00",X"00",X"08",X"41",X"00",X"00",X"08",X"1F",X"00",X"00",X"88",X"FF",X"00",X"00",X"88",X"F8",
		X"00",X"00",X"88",X"F0",X"00",X"00",X"88",X"F0",X"00",X"00",X"80",X"24",X"00",X"00",X"80",X"22",
		X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"0E",X"42",X"00",X"00",X"E1",X"84",X"00",X"0E",X"11",X"88",X"00",X"AA",X"11",X"18",
		X"00",X"AA",X"17",X"44",X"00",X"AA",X"12",X"22",X"00",X"AA",X"12",X"22",X"00",X"EE",X"12",X"14",
		X"00",X"EE",X"99",X"14",X"00",X"AA",X"A9",X"64",X"00",X"AA",X"AA",X"66",X"00",X"DA",X"AA",X"99",
		X"00",X"DD",X"AA",X"A9",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"08",X"80",X"00",X"00",X"08",X"06",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"4F",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"08",X"42",X"00",X"00",X"E1",X"11",X"00",X"0E",X"11",X"88",X"00",X"AA",X"11",X"88",
		X"00",X"AA",X"11",X"88",X"00",X"AA",X"11",X"88",X"00",X"AA",X"88",X"88",X"00",X"EE",X"12",X"28",
		X"00",X"EE",X"99",X"22",X"00",X"AA",X"A9",X"62",X"00",X"AA",X"AA",X"64",X"00",X"DA",X"AA",X"99",
		X"00",X"DD",X"AA",X"A9",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"42",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"48",X"E0",X"00",X"00",X"22",X"11",X"00",X"00",X"22",X"11",X"A0",X"00",
		X"22",X"11",X"AA",X"00",X"24",X"11",X"AA",X"00",X"44",X"19",X"AA",X"00",X"4C",X"99",X"EA",X"00",
		X"22",X"9A",X"EE",X"00",X"22",X"AA",X"EE",X"00",X"62",X"AA",X"AE",X"00",X"99",X"AA",X"DD",X"00",
		X"AA",X"AA",X"00",X"00",X"AA",X"AD",X"00",X"00",X"AA",X"DD",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"D0",X"DD",
		X"0C",X"00",X"CC",X"C0",X"00",X"C0",X"C0",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"C0",X"00",X"DD",X"00",X"00",X"00",X"CC",X"00",X"0C",X"0D",X"00",X"00",X"9C",X"0C",X"00",
		X"00",X"C0",X"DC",X"00",X"00",X"CC",X"CC",X"DD",X"00",X"C0",X"C0",X"CC",X"00",X"0C",X"CD",X"00",
		X"C0",X"0C",X"0D",X"0C",X"00",X"0C",X"CC",X"CD",X"00",X"00",X"0C",X"C0",X"00",X"00",X"0C",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0C",X"09",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"90",X"00",X"00",X"0C",X"00",X"00",X"D0",X"00",X"00",X"C0",X"D0",X"C0",X"0C",X"00",
		X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"0D",X"00",
		X"0D",X"00",X"0D",X"09",X"CD",X"0D",X"0C",X"00",X"C0",X"CD",X"00",X"00",X"0C",X"C0",X"0C",X"00",
		X"C0",X"00",X"00",X"0C",X"D0",X"00",X"00",X"00",X"00",X"D0",X"90",X"D0",X"00",X"00",X"00",X"CD",
		X"00",X"00",X"00",X"0C",X"C0",X"00",X"D0",X"00",X"00",X"00",X"0D",X"0D",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"CD",
		X"00",X"D0",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"CC",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",
		X"C0",X"0D",X"00",X"00",X"00",X"DC",X"00",X"00",X"90",X"0D",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"CC",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"CD",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",
		X"06",X"26",X"00",X"00",X"02",X"26",X"00",X"00",X"2F",X"22",X"00",X"00",X"20",X"22",X"00",X"00",
		X"40",X"42",X"00",X"00",X"12",X"22",X"00",X"00",X"22",X"24",X"00",X"00",X"22",X"11",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"04",X"00",X"22",X"28",X"42",X"00",X"42",X"42",X"22",X"00",
		X"11",X"42",X"00",X"00",X"88",X"42",X"00",X"00",X"80",X"42",X"00",X"00",X"22",X"44",X"24",X"00",
		X"22",X"04",X"22",X"00",X"82",X"01",X"22",X"22",X"24",X"00",X"22",X"22",X"40",X"00",X"22",X"04",
		X"00",X"00",X"22",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"26",X"00",X"00",
		X"06",X"26",X"00",X"00",X"02",X"26",X"00",X"00",X"2F",X"22",X"00",X"00",X"20",X"22",X"00",X"00",
		X"40",X"42",X"00",X"00",X"12",X"22",X"00",X"00",X"22",X"24",X"00",X"00",X"22",X"11",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"22",X"00",X"22",X"28",X"22",X"00",X"42",X"48",X"24",X"00",
		X"81",X"28",X"22",X"00",X"88",X"22",X"11",X"00",X"80",X"42",X"00",X"00",X"00",X"42",X"40",X"00",
		X"88",X"44",X"24",X"00",X"88",X"21",X"22",X"22",X"88",X"00",X"22",X"22",X"00",X"00",X"22",X"02",
		X"00",X"00",X"24",X"22",X"00",X"00",X"20",X"22",X"00",X"00",X"40",X"11",X"00",X"00",X"22",X"00",
		X"00",X"00",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",
		X"06",X"26",X"00",X"00",X"02",X"26",X"00",X"00",X"2F",X"22",X"00",X"00",X"20",X"22",X"00",X"00",
		X"40",X"42",X"00",X"00",X"12",X"22",X"00",X"00",X"22",X"24",X"00",X"00",X"22",X"11",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"44",X"00",X"22",X"28",X"22",X"00",X"42",X"40",X"22",X"22",
		X"11",X"00",X"22",X"42",X"88",X"00",X"22",X"02",X"80",X"00",X"42",X"42",X"00",X"00",X"42",X"22",
		X"00",X"00",X"14",X"00",X"00",X"02",X"14",X"00",X"00",X"22",X"01",X"02",X"00",X"22",X"20",X"02",
		X"00",X"22",X"20",X"02",X"00",X"12",X"22",X"20",X"00",X"02",X"22",X"20",X"00",X"02",X"24",X"40",
		X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",
		X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",
		X"00",X"00",X"0E",X"11",X"00",X"00",X"E1",X"11",X"00",X"0E",X"11",X"11",X"00",X"AA",X"11",X"11",
		X"00",X"AA",X"11",X"11",X"00",X"AA",X"11",X"11",X"00",X"AA",X"11",X"11",X"00",X"EE",X"11",X"11",
		X"00",X"EE",X"99",X"11",X"00",X"AA",X"A9",X"61",X"00",X"AA",X"AA",X"66",X"00",X"DA",X"AA",X"99",
		X"00",X"DD",X"AA",X"A9",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"AA",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"8A",X"00",X"00",X"00",X"8A",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"A0",X"00",X"EE",X"AA",X"00",X"00",
		X"11",X"1A",X"00",X"00",X"11",X"EE",X"1D",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"19",X"AA",X"00",X"11",X"99",X"EA",X"00",
		X"11",X"9A",X"EE",X"00",X"11",X"AA",X"EE",X"00",X"61",X"AA",X"AE",X"00",X"99",X"AA",X"DD",X"00",
		X"AA",X"AA",X"00",X"00",X"AA",X"AD",X"00",X"00",X"AA",X"DD",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"50",X"55",X"00",X"00",X"55",X"59",X"00",
		X"00",X"05",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"35",X"00",X"00",X"50",X"51",X"00",
		X"0D",X"15",X"11",X"00",X"DD",X"11",X"19",X"00",X"99",X"99",X"11",X"00",X"99",X"DD",X"99",X"D0",
		X"99",X"99",X"11",X"BD",X"99",X"99",X"71",X"DD",X"DD",X"11",X"91",X"9D",X"11",X"AA",X"91",X"9D",
		X"01",X"AA",X"91",X"D0",X"00",X"AA",X"D9",X"D0",X"00",X"AA",X"1D",X"10",X"00",X"11",X"11",X"00",
		X"00",X"19",X"1D",X"00",X"00",X"99",X"1D",X"00",X"00",X"99",X"DD",X"00",X"00",X"99",X"11",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",
		X"00",X"D1",X"00",X"00",X"88",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"92",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"42",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"7E",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"77",X"66",X"99",X"96",X"00",X"00",X"00",X"00",X"77",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"A8",X"88",X"88",X"88",X"A8",X"88",X"88",X"88",X"AA",X"88",X"88",X"88",X"BA",X"88",X"88",
		X"88",X"AB",X"88",X"88",X"88",X"AA",X"88",X"88",X"A8",X"AB",X"88",X"88",X"AA",X"AA",X"88",X"88",
		X"AA",X"A5",X"88",X"88",X"AB",X"AB",X"18",X"88",X"55",X"55",X"55",X"88",X"55",X"5B",X"5A",X"88",
		X"55",X"55",X"AA",X"88",X"51",X"5B",X"11",X"88",X"A5",X"55",X"A1",X"88",X"11",X"5B",X"A8",X"88",
		X"88",X"55",X"BA",X"88",X"88",X"5B",X"AB",X"88",X"88",X"5B",X"AA",X"88",X"88",X"5B",X"AA",X"88",
		X"88",X"5B",X"88",X"88",X"88",X"5B",X"88",X"88",X"88",X"5B",X"88",X"88",X"88",X"5B",X"88",X"88",
		X"81",X"5B",X"88",X"88",X"8A",X"5B",X"88",X"88",X"81",X"5B",X"88",X"88",X"88",X"51",X"88",X"88",
		X"88",X"18",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",
		X"00",X"06",X"00",X"EE",X"00",X"66",X"00",X"EE",X"00",X"60",X"00",X"EE",X"00",X"60",X"01",X"EE",
		X"00",X"60",X"15",X"EE",X"00",X"60",X"55",X"EE",X"00",X"60",X"00",X"EE",X"00",X"60",X"11",X"EE",
		X"00",X"60",X"11",X"EE",X"00",X"60",X"01",X"EE",X"00",X"60",X"00",X"EE",X"00",X"60",X"11",X"EE",
		X"00",X"60",X"00",X"EE",X"00",X"60",X"40",X"EE",X"00",X"60",X"44",X"EE",X"00",X"64",X"44",X"EE",
		X"00",X"60",X"40",X"EE",X"00",X"66",X"46",X"EE",X"00",X"66",X"06",X"EE",X"00",X"66",X"66",X"EE",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"EE",X"00",X"11",X"66",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"E1",X"00",X"00",X"11",X"11",X"00",X"00",X"01",X"10",
		X"00",X"11",X"06",X"00",X"03",X"31",X"66",X"00",X"10",X"31",X"00",X"E0",X"1F",X"F1",X"00",X"EE",
		X"14",X"14",X"00",X"EE",X"44",X"14",X"00",X"EE",X"44",X"44",X"00",X"EE",X"44",X"44",X"00",X"EE",
		X"11",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"00",X"11",X"00",X"EE",X"00",X"A1",X"00",X"EE",
		X"00",X"71",X"00",X"EE",X"04",X"74",X"00",X"EE",X"01",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",
		X"00",X"41",X"00",X"EE",X"00",X"10",X"40",X"EE",X"00",X"60",X"44",X"EE",X"00",X"64",X"44",X"EE",
		X"00",X"60",X"40",X"EE",X"00",X"66",X"46",X"EE",X"00",X"66",X"06",X"EE",X"00",X"66",X"66",X"EE",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"EE",X"00",X"11",X"66",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"E1",X"00",X"00",X"11",X"11",X"00",X"00",X"01",X"10",
		X"00",X"11",X"06",X"00",X"0F",X"31",X"66",X"00",X"1F",X"F1",X"00",X"E0",X"1F",X"F1",X"00",X"EE",
		X"14",X"F4",X"00",X"EE",X"44",X"14",X"00",X"EE",X"44",X"44",X"00",X"EE",X"44",X"44",X"00",X"EE",
		X"01",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",
		X"00",X"14",X"00",X"EE",X"00",X"14",X"00",X"EE",X"07",X"44",X"00",X"EE",X"47",X"44",X"00",X"EE",
		X"14",X"41",X"00",X"EE",X"01",X"40",X"40",X"EE",X"00",X"10",X"44",X"EE",X"00",X"14",X"44",X"EE",
		X"00",X"60",X"40",X"EE",X"00",X"66",X"46",X"EE",X"00",X"66",X"06",X"EE",X"00",X"66",X"66",X"EE",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"EE",X"00",X"11",X"66",X"EE",X"00",X"00",X"66",X"EE",
		X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"E1",X"00",X"00",X"11",X"11",X"00",X"00",X"01",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"DE",X"00",X"00",X"60",X"6E",X"00",
		X"00",X"0E",X"6E",X"00",X"00",X"66",X"6E",X"00",X"00",X"E6",X"6E",X"00",X"00",X"60",X"EE",X"00",
		X"00",X"A0",X"EE",X"00",X"00",X"AA",X"E0",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"A0",X"66",X"00",X"0C",X"AA",X"66",X"00",X"00",X"AA",X"A0",X"00",
		X"00",X"0D",X"6E",X"00",X"00",X"0A",X"AE",X"00",X"C0",X"AA",X"AE",X"00",X"00",X"00",X"AE",X"00",
		X"00",X"00",X"A6",X"00",X"00",X"A0",X"A6",X"00",X"00",X"A0",X"06",X"00",X"00",X"AA",X"66",X"00",
		X"00",X"66",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"00",X"99",X"B0",X"00",X"00",X"09",X"50",X"00",
		X"00",X"09",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"9F",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"BB",X"55",X"00",X"00",X"B5",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"00",X"FF",X"B0",X"00",X"00",X"FF",X"50",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"F9",X"55",X"00",X"00",X"F9",X"55",X"00",
		X"00",X"F9",X"55",X"00",X"00",X"F9",X"55",X"00",X"00",X"BB",X"55",X"00",X"00",X"B5",X"55",X"00",
		X"00",X"55",X"5A",X"00",X"00",X"55",X"A0",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"00",X"FA",X"B0",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FA",X"55",X"00",X"00",X"FA",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"99",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"B5",X"09",X"00",X"00",X"55",X"90",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"00",X"FF",X"B0",X"00",X"00",X"FF",X"50",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"BB",X"55",X"00",X"00",X"B5",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"93",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"09",X"00",X"00",X"93",X"00",X"33",
		X"00",X"93",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"33",X"00",X"39",X"00",X"99",X"00",X"90",X"00",X"00",X"33",X"00",X"00",X"33",X"99",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"30",
		X"00",X"33",X"00",X"93",X"00",X"93",X"00",X"09",X"00",X"99",X"33",X"00",X"03",X"00",X"99",X"00",
		X"09",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"33",X"00",X"00",X"00",X"93",X"00",X"33",
		X"00",X"93",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"00",X"33",X"90",X"00",X"00",X"99",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",
		X"33",X"90",X"00",X"00",X"39",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"B9",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"07",X"00",X"00",X"99",X"07",X"00",X"00",X"99",X"07",X"00",X"00",X"09",X"75",
		X"00",X"00",X"99",X"7A",X"00",X"00",X"9B",X"7E",X"00",X"00",X"99",X"70",X"00",X"00",X"99",X"70",
		X"00",X"09",X"99",X"A0",X"00",X"00",X"99",X"AA",X"00",X"99",X"99",X"EE",X"09",X"90",X"B9",X"07",
		X"00",X"99",X"99",X"07",X"09",X"90",X"99",X"07",X"90",X"99",X"99",X"05",X"09",X"99",X"99",X"00",
		X"99",X"9B",X"99",X"90",X"00",X"99",X"99",X"90",X"09",X"90",X"B9",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"09",X"99",
		X"F0",X"0A",X"0A",X"06",X"00",X"0A",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"AA",X"AF",X"0A",
		X"00",X"A6",X"AA",X"A0",X"00",X"A0",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"07",X"77",X"00",
		X"0A",X"77",X"66",X"A0",X"00",X"70",X"00",X"00",X"0A",X"00",X"00",X"A0",X"0A",X"F0",X"07",X"A0",
		X"00",X"00",X"67",X"A0",X"A0",X"00",X"00",X"AA",X"A0",X"00",X"60",X"AA",X"A0",X"00",X"00",X"A0",
		X"A0",X"00",X"00",X"A6",X"00",X"00",X"00",X"00",X"A6",X"00",X"76",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"70",X"00",X"0A",X"00",X"70",X"00",X"AA",X"66",X"00",X"00",X"A0",X"77",X"00",X"00",
		X"00",X"77",X"00",X"00",X"AA",X"07",X"00",X"60",X"A6",X"67",X"A0",X"00",X"A0",X"AA",X"AF",X"00",
		X"AA",X"6A",X"AA",X"00",X"00",X"0A",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"6F",X"00",X"00",X"00",X"F0",X"00",X"0A",X"6A",X"60",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"7A",X"00",X"0E",X"00",X"0F",X"0A",X"00",X"00",X"FF",X"A6",X"00",
		X"00",X"FF",X"00",X"00",X"06",X"0F",X"77",X"07",X"00",X"FF",X"00",X"00",X"00",X"F0",X"A0",X"00",
		X"00",X"7F",X"00",X"00",X"00",X"7A",X"00",X"00",X"A0",X"00",X"00",X"0E",X"00",X"07",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"70",X"00",X"00",X"0A",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"6A",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"7F",X"70",X"00",
		X"00",X"FF",X"AA",X"00",X"00",X"7F",X"07",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"00",
		X"60",X"A7",X"60",X"00",X"00",X"AF",X"00",X"00",X"60",X"66",X"A0",X"00",X"00",X"77",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"7A",X"00",X"00",X"00",X"AF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"7A",X"00",X"00",X"00",X"67",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"36",X"66",X"00",X"00",X"60",X"06",X"00",X"00",X"00",X"3A",
		X"06",X"00",X"A0",X"35",X"66",X"66",X"A0",X"33",X"00",X"55",X"AA",X"53",X"00",X"3D",X"AA",X"53",
		X"72",X"CD",X"AA",X"53",X"27",X"CD",X"AA",X"53",X"AA",X"CC",X"AA",X"53",X"27",X"3C",X"AA",X"55",
		X"77",X"3C",X"AA",X"35",X"00",X"3C",X"AA",X"52",X"CA",X"3C",X"AA",X"52",X"DA",X"3C",X"AA",X"22",
		X"DA",X"3C",X"AA",X"22",X"AA",X"31",X"AA",X"22",X"DA",X"31",X"AA",X"26",X"DA",X"33",X"A1",X"26",
		X"DA",X"30",X"A1",X"26",X"DA",X"30",X"A1",X"26",X"D1",X"30",X"A1",X"1E",X"D0",X"30",X"A0",X"0E",
		X"D0",X"30",X"10",X"0E",X"D0",X"30",X"10",X"0E",X"D0",X"00",X"00",X"0E",X"D0",X"00",X"00",X"0E",
		X"D0",X"00",X"00",X"0E",X"0D",X"00",X"00",X"0E",X"D0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",
		X"60",X"06",X"00",X"00",X"06",X"0D",X"00",X"00",X"00",X"DD",X"60",X"00",X"70",X"0D",X"66",X"00",
		X"60",X"0D",X"66",X"00",X"0C",X"DD",X"06",X"00",X"0C",X"D0",X"06",X"00",X"AA",X"D0",X"06",X"00",
		X"AC",X"D0",X"06",X"00",X"AD",X"D3",X"06",X"00",X"C5",X"D3",X"66",X"00",X"C5",X"D3",X"66",X"00",
		X"C5",X"D3",X"A5",X"00",X"C5",X"D3",X"A5",X"00",X"C5",X"D5",X"AA",X"00",X"C5",X"D5",X"5A",X"00",
		X"C1",X"D5",X"5A",X"00",X"C1",X"D5",X"5A",X"00",X"C1",X"D5",X"6A",X"00",X"C1",X"55",X"1A",X"00",
		X"C1",X"55",X"1A",X"00",X"C1",X"55",X"1A",X"00",X"1C",X"55",X"1A",X"00",X"C1",X"55",X"0A",X"00",
		X"C1",X"05",X"0A",X"00",X"01",X"05",X"0A",X"00",X"11",X"05",X"0A",X"00",X"10",X"05",X"0A",X"00",
		X"00",X"05",X"0A",X"00",X"00",X"05",X"0A",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"0A",X"00",
		X"00",X"3E",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"AA",X"D0",X"00",
		X"00",X"FF",X"D0",X"00",X"00",X"FF",X"D0",X"00",X"00",X"F9",X"DD",X"00",X"CC",X"90",X"ED",X"00",
		X"CD",X"90",X"ED",X"00",X"ED",X"F9",X"CE",X"C0",X"00",X"FF",X"CE",X"C0",X"00",X"55",X"C6",X"C0",
		X"00",X"55",X"C6",X"C0",X"00",X"00",X"CC",X"EC",X"0C",X"AA",X"EC",X"0C",X"CC",X"EE",X"EC",X"0C",
		X"CC",X"00",X"0C",X"0C",X"CE",X"00",X"0C",X"0C",X"E0",X"00",X"0C",X"0E",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"E0",X"EE",X"E6",X"00",X"00",X"E6",X"60",X"00",X"06",X"00",X"00",X"09",
		X"0E",X"06",X"00",X"99",X"0E",X"06",X"00",X"99",X"0E",X"06",X"00",X"A9",X"06",X"06",X"00",X"A9",
		X"06",X"66",X"00",X"A9",X"01",X"66",X"00",X"A9",X"00",X"66",X"00",X"A9",X"00",X"66",X"00",X"A9",
		X"00",X"11",X"11",X"A9",X"00",X"61",X"44",X"A9",X"00",X"66",X"44",X"A9",X"00",X"6E",X"44",X"99",
		X"00",X"0E",X"74",X"10",X"00",X"00",X"74",X"10",X"00",X"E0",X"44",X"00",X"0E",X"1E",X"44",X"00",
		X"E1",X"71",X"44",X"00",X"44",X"44",X"45",X"00",X"44",X"44",X"54",X"00",X"44",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"11",X"00",X"44",X"11",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"6E",X"00",X"EE",X"EE",X"E6",X"00",X"60",X"EE",X"66",X"00",X"00",X"E0",X"60",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0A",X"E0",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"10",X"00",X"00",X"6E",X"11",X"00",
		X"11",X"EE",X"44",X"00",X"14",X"00",X"74",X"00",X"14",X"06",X"17",X"00",X"44",X"66",X"74",X"00",
		X"44",X"77",X"44",X"00",X"14",X"11",X"44",X"00",X"11",X"44",X"44",X"00",X"01",X"44",X"44",X"00",
		X"00",X"44",X"11",X"00",X"00",X"4A",X"10",X"00",X"00",X"AA",X"00",X"00",X"00",X"1A",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"0E",X"10",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"09",X"00",
		X"00",X"E0",X"09",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",X"50",X"00",
		X"00",X"00",X"55",X"00",X"00",X"11",X"55",X"A0",X"0A",X"16",X"53",X"00",X"0A",X"66",X"55",X"00",
		X"09",X"60",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"50",X"55",X"00",X"00",X"55",X"50",X"00",
		X"00",X"55",X"06",X"00",X"00",X"55",X"6A",X"A0",X"00",X"53",X"6A",X"AA",X"00",X"35",X"AA",X"99",
		X"00",X"55",X"AA",X"00",X"0A",X"55",X"AA",X"00",X"0A",X"55",X"99",X"00",X"0A",X"50",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"EE",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"66",X"A7",X"EE",X"00",X"00",X"00",X"00",X"00",X"60",X"77",X"6C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"DD",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"E0",X"42",X"44",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"0E",X"10",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"09",X"00",
		X"00",X"E0",X"09",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",X"50",X"00",
		X"00",X"00",X"55",X"00",X"00",X"11",X"55",X"A0",X"0A",X"16",X"53",X"00",X"0A",X"66",X"55",X"00",
		X"09",X"60",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"50",X"55",X"00",X"00",X"55",X"50",X"00",
		X"00",X"35",X"06",X"00",X"05",X"53",X"6A",X"A0",X"5A",X"55",X"6A",X"AA",X"AA",X"55",X"AA",X"99",
		X"A1",X"55",X"AA",X"00",X"14",X"55",X"AA",X"00",X"14",X"55",X"99",X"00",X"14",X"55",X"00",X"00",
		X"14",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"0E",X"10",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E7",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"C0",X"00",X"00",X"16",X"CC",
		X"00",X"00",X"16",X"AC",X"00",X"ED",X"00",X"CC",X"00",X"50",X"C0",X"C9",X"00",X"EE",X"CC",X"C9",
		X"99",X"05",X"DC",X"90",X"99",X"EE",X"DD",X"9A",X"99",X"50",X"0D",X"00",X"99",X"EE",X"DD",X"A0",
		X"09",X"DD",X"DD",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"77",X"77",X"77",X"88",X"78",X"8F",X"77",X"88",X"78",X"8F",X"77",X"88",
		X"78",X"8F",X"77",X"88",X"78",X"8F",X"77",X"88",X"78",X"8F",X"77",X"88",X"78",X"8F",X"77",X"88",
		X"78",X"8F",X"88",X"88",X"77",X"77",X"77",X"88",X"77",X"77",X"77",X"88",X"00",X"88",X"88",X"88",
		X"00",X"78",X"88",X"88",X"00",X"70",X"88",X"88",X"88",X"78",X"88",X"88",X"88",X"F8",X"88",X"88",
		X"88",X"33",X"88",X"88",X"88",X"BB",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"33",X"88",X"88",
		X"88",X"33",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"BB",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"D3",X"88",X"88",
		X"88",X"3D",X"88",X"88",X"88",X"D3",X"88",X"88",X"88",X"33",X"88",X"88",X"88",X"33",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"EE",X"55",X"00",X"00",X"33",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"05",X"55",X"EE",X"00",X"05",X"55",X"55",X"30",
		X"55",X"55",X"55",X"50",X"51",X"55",X"55",X"50",X"51",X"55",X"55",X"5A",X"11",X"55",X"55",X"5F",
		X"41",X"55",X"55",X"5F",X"51",X"55",X"55",X"5A",X"54",X"55",X"55",X"50",X"55",X"55",X"55",X"40",
		X"05",X"55",X"55",X"40",X"05",X"55",X"66",X"00",X"00",X"45",X"55",X"00",X"00",X"44",X"55",X"00",
		X"00",X"44",X"55",X"00",X"00",X"66",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"00",X"00",
		X"05",X"55",X"03",X"00",X"05",X"55",X"35",X"00",X"51",X"55",X"55",X"00",X"E5",X"15",X"55",X"30",
		X"7E",X"15",X"55",X"50",X"EE",X"55",X"55",X"50",X"EE",X"55",X"EE",X"5A",X"EF",X"55",X"55",X"5F",
		X"65",X"55",X"55",X"5F",X"66",X"54",X"66",X"5A",X"66",X"45",X"55",X"50",X"66",X"15",X"55",X"50",
		X"66",X"15",X"55",X"40",X"51",X"45",X"45",X"00",X"05",X"55",X"44",X"00",X"05",X"55",X"04",X"00",
		X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"7E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EF",X"55",X"00",
		X"00",X"65",X"44",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"65",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"06",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"07",X"60",X"00",X"00",X"70",X"60",X"00",
		X"00",X"70",X"00",X"00",X"60",X"07",X"60",X"00",X"06",X"00",X"60",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"60",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"77",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"E7",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"E6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"06",X"00",X"00",X"00",X"00",X"00",X"0E",X"66",X"E6",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"46",X"66",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"C9",X"AA",X"C0",X"00",X"00",X"00",X"00",X"CA",X"99",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"05",X"50",
		X"00",X"00",X"05",X"55",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"99",X"00",
		X"90",X"00",X"F9",X"00",X"D9",X"09",X"9B",X"00",X"9D",X"00",X"BB",X"00",X"99",X"09",X"9B",X"00",
		X"00",X"00",X"B9",X"00",X"00",X"09",X"B9",X"00",X"00",X"90",X"99",X"00",X"00",X"C9",X"90",X"00",
		X"00",X"C9",X"90",X"00",X"99",X"CF",X"99",X"00",X"BB",X"B9",X"BB",X"00",X"99",X"9F",X"99",X"99",
		X"DD",X"BB",X"DD",X"C9",X"99",X"0C",X"99",X"99",X"00",X"BB",X"D0",X"00",X"00",X"B9",X"9D",X"00",
		X"00",X"B9",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"90",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",
		X"90",X"9D",X"09",X"00",X"F9",X"9B",X"9D",X"00",X"99",X"9D",X"DD",X"00",X"99",X"99",X"D0",X"00",
		X"09",X"99",X"D9",X"00",X"00",X"BB",X"9B",X"00",X"00",X"0B",X"00",X"00",X"00",X"CB",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"BF",X"C9",X"00",X"00",X"D9",X"FF",X"00",X"00",X"DD",X"99",X"00",
		X"00",X"DD",X"F9",X"90",X"00",X"9D",X"BB",X"00",X"00",X"9D",X"BB",X"00",X"00",X"9D",X"99",X"90",
		X"00",X"9C",X"99",X"00",X"00",X"9B",X"09",X"90",X"00",X"9D",X"00",X"00",X"00",X"9B",X"00",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"11",X"00",X"00",X"70",X"00",X"00",X"00",X"07",X"06",X"00",X"00",
		X"07",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"70",X"00",X"00",X"60",X"07",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"0F",X"07",X"00",
		X"77",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"F0",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"BB",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"0F",X"00",X"0B",
		X"00",X"0F",X"00",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E8",X"00",X"00",X"02",X"E0",X"00",X"00",X"02",X"EE",X"00",X"00",X"04",X"66",
		X"00",X"00",X"04",X"66",X"00",X"00",X"04",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"80",X"16",
		X"00",X"00",X"80",X"61",X"00",X"00",X"80",X"62",X"00",X"00",X"80",X"12",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"0C",X"42",X"00",X"00",X"22",X"24",
		X"00",X"00",X"2C",X"44",X"00",X"00",X"2C",X"01",X"00",X"EA",X"2C",X"04",X"00",X"EE",X"2C",X"82",
		X"00",X"AA",X"24",X"22",X"0A",X"AA",X"41",X"22",X"AA",X"AE",X"22",X"22",X"DA",X"EE",X"44",X"24",
		X"0D",X"AA",X"11",X"44",X"00",X"AA",X"99",X"41",X"00",X"AA",X"A9",X"66",X"00",X"AA",X"AA",X"66",
		X"00",X"DA",X"AA",X"99",X"00",X"DD",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"20",X"E8",X"00",X"00",X"22",X"EE",X"00",X"00",X"22",X"44",X"00",X"00",X"42",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"42",X"00",X"00",X"84",X"F2",X"00",X"00",X"84",X"82",
		X"00",X"00",X"84",X"02",X"00",X"00",X"82",X"52",X"00",X"00",X"84",X"22",X"00",X"00",X"08",X"22",
		X"00",X"00",X"08",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"EE",X"22",X"00",X"00",X"11",X"22",X"00",X"EA",X"C1",X"42",X"00",X"EE",X"C1",X"11",
		X"00",X"AA",X"77",X"24",X"0A",X"AA",X"22",X"24",X"AA",X"AE",X"1C",X"22",X"DA",X"EE",X"22",X"22",
		X"0D",X"AA",X"0C",X"22",X"00",X"AA",X"99",X"44",X"00",X"AA",X"A9",X"66",X"00",X"AA",X"AA",X"66",
		X"00",X"DA",X"AA",X"99",X"00",X"DD",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"60",X"00",X"00",X"88",X"06",X"00",X"00",X"88",X"64",
		X"00",X"00",X"08",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"08",X"F2",X"00",X"00",X"00",X"02",
		X"00",X"00",X"88",X"02",X"00",X"00",X"88",X"22",X"00",X"00",X"88",X"22",X"00",X"00",X"80",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"08",X"24",X"00",X"00",X"11",X"11",X"00",X"EA",X"81",X"88",X"00",X"EE",X"88",X"08",
		X"00",X"AA",X"42",X"80",X"0A",X"AA",X"42",X"88",X"AA",X"AE",X"42",X"88",X"DA",X"EE",X"42",X"82",
		X"0D",X"AA",X"44",X"22",X"00",X"AA",X"99",X"28",X"00",X"AA",X"A9",X"44",X"00",X"AA",X"AA",X"66",
		X"00",X"DA",X"AA",X"99",X"00",X"DD",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"DD",
		X"06",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"26",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"24",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"81",X"90",X"00",X"00",X"81",X"9A",X"00",X"00",X"20",X"9A",X"00",X"00",
		X"28",X"9E",X"AA",X"00",X"28",X"9A",X"AA",X"00",X"28",X"9E",X"AA",X"00",X"28",X"AA",X"AA",X"00",
		X"28",X"AA",X"EE",X"00",X"88",X"AA",X"ED",X"00",X"19",X"AA",X"D0",X"00",X"99",X"AA",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"AA",X"DD",X"00",X"00",X"AA",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"DD",X"0D",
		X"00",X"00",X"C0",X"CD",X"00",X"00",X"00",X"C0",X"00",X"D0",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"0C",X"0D",X"0D",X"00",X"C0",X"DC",X"CD",X"C0",X"C0",X"0C",X"C0",X"00",X"00",X"C0",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"D0",X"00",X"CC",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"D0",X"CD",X"00",X"CD",X"00",X"0C",X"00",X"C0",X"D0",X"00",X"00",X"0C",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"C0",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"C0",X"00",X"0D",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"0C",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"0C",X"C0",X"C0",X"C0",X"00",X"0C",X"0C",X"00",X"C0",X"00",X"00",
		X"C0",X"00",X"90",X"CD",X"00",X"DC",X"00",X"0C",X"90",X"00",X"D0",X"00",X"00",X"00",X"0D",X"0D",
		X"00",X"00",X"C0",X"CC",X"C0",X"00",X"0C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CD",X"00",X"C0",X"00",X"C0",X"00",X"D0",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"90",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"D0",X"0D",X"00",X"0D",X"DD",X"0C",X"00",X"CD",X"CD",X"0C",X"00",X"C0",X"CD",X"00",X"00",
		X"CD",X"C0",X"00",X"00",X"90",X"CD",X"90",X"00",X"D0",X"C0",X"00",X"00",X"0C",X"CD",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DC",X"00",X"0C",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"08",X"00",X"00",X"66",X"00",X"00",X"00",X"62",X"60",X"00",X"00",
		X"22",X"60",X"00",X"00",X"62",X"66",X"00",X"00",X"F2",X"64",X"00",X"00",X"02",X"62",X"00",X"00",
		X"02",X"24",X"00",X"00",X"22",X"24",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"24",X"00",X"00",
		X"22",X"20",X"42",X"00",X"22",X"40",X"22",X"00",X"22",X"80",X"20",X"00",X"21",X"80",X"22",X"00",
		X"11",X"02",X"00",X"00",X"80",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"24",X"22",X"40",X"00",X"40",X"42",X"24",X"00",X"00",X"44",X"22",X"22",X"00",X"84",X"22",X"22",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"66",X"00",X"00",X"00",X"62",X"60",X"00",X"00",
		X"22",X"60",X"00",X"00",X"62",X"66",X"00",X"00",X"F2",X"64",X"00",X"00",X"02",X"62",X"00",X"00",
		X"02",X"24",X"00",X"00",X"22",X"24",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"24",X"00",X"00",
		X"22",X"20",X"00",X"00",X"22",X"40",X"20",X"00",X"22",X"80",X"22",X"00",X"21",X"80",X"22",X"00",
		X"11",X"02",X"11",X"00",X"80",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"88",X"22",X"00",X"00",X"80",X"22",X"40",X"00",X"02",X"42",X"40",X"00",X"22",X"82",X"22",X"00",
		X"22",X"04",X"42",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"08",X"00",X"00",X"66",X"00",X"00",X"00",X"62",X"60",X"00",X"00",
		X"22",X"60",X"00",X"00",X"62",X"66",X"00",X"00",X"F2",X"64",X"00",X"00",X"02",X"62",X"00",X"00",
		X"02",X"24",X"00",X"00",X"22",X"24",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"24",X"00",X"00",
		X"22",X"21",X"00",X"00",X"22",X"12",X"00",X"00",X"22",X"42",X"44",X"00",X"24",X"44",X"22",X"22",
		X"11",X"41",X"22",X"42",X"80",X"21",X"22",X"04",X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",
		X"00",X"20",X"22",X"00",X"00",X"20",X"42",X"00",X"00",X"40",X"14",X"00",X"00",X"00",X"11",X"20",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",
		X"00",X"00",X"EE",X"11",X"00",X"00",X"11",X"11",X"00",X"EA",X"11",X"11",X"00",X"EE",X"1D",X"11",
		X"00",X"AA",X"1D",X"11",X"0A",X"AA",X"1D",X"11",X"AA",X"AE",X"1D",X"11",X"DA",X"EE",X"0D",X"11",
		X"0D",X"AA",X"1D",X"11",X"00",X"AA",X"99",X"11",X"00",X"AA",X"A9",X"66",X"00",X"AA",X"AA",X"66",
		X"00",X"DA",X"AA",X"99",X"00",X"DD",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"08",X"AA",X"A0",X"00",X"08",X"AA",X"A0",X"00",X"08",X"AA",X"00",X"00",X"EE",X"AA",X"00",X"00",
		X"11",X"AA",X"00",X"00",X"11",X"1A",X"D0",X"00",X"11",X"91",X"1D",X"00",X"11",X"9A",X"11",X"00",
		X"11",X"9E",X"11",X"00",X"11",X"9A",X"1A",X"00",X"11",X"9E",X"AA",X"00",X"11",X"AA",X"AA",X"00",
		X"11",X"AA",X"EE",X"00",X"11",X"AA",X"ED",X"00",X"19",X"AA",X"D0",X"00",X"99",X"AA",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"AA",X"DD",X"00",X"00",X"AA",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"90",X"00",
		X"00",X"55",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"11",X"00",X"DD",X"00",X"99",X"00",
		X"99",X"55",X"11",X"00",X"DD",X"11",X"99",X"00",X"99",X"91",X"11",X"00",X"99",X"99",X"71",X"00",
		X"9A",X"DD",X"D1",X"00",X"9A",X"99",X"D1",X"00",X"91",X"11",X"D9",X"00",X"D1",X"FF",X"D9",X"00",
		X"D1",X"AA",X"99",X"00",X"19",X"AF",X"9B",X"00",X"01",X"AA",X"BD",X"00",X"11",X"11",X"D9",X"00",
		X"1A",X"99",X"99",X"00",X"1A",X"99",X"99",X"00",X"1A",X"9D",X"DD",X"00",X"1A",X"D1",X"11",X"00",
		X"11",X"11",X"00",X"00",X"00",X"1D",X"00",X"00",X"00",X"D1",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"22",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"24",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"EE",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"7E",X"60",X"99",X"66",X"00",X"00",X"00",X"00",X"EE",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"A8",X"88",X"88",X"88",X"AA",X"88",X"88",X"88",X"AA",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"55",X"A8",X"88",X"88",X"85",X"A8",X"88",X"88",X"85",X"A8",X"88",X"88",X"88",X"A8",X"88",X"88",
		X"A1",X"51",X"88",X"88",X"51",X"51",X"88",X"88",X"B5",X"51",X"18",X"88",X"5B",X"51",X"A1",X"88",
		X"55",X"51",X"AA",X"88",X"55",X"51",X"AA",X"88",X"15",X"51",X"1A",X"88",X"55",X"51",X"81",X"88",
		X"11",X"51",X"88",X"88",X"88",X"51",X"88",X"88",X"88",X"51",X"A8",X"88",X"88",X"51",X"A8",X"88",
		X"88",X"51",X"88",X"88",X"81",X"5A",X"88",X"88",X"81",X"5A",X"88",X"88",X"1A",X"5A",X"88",X"88",
		X"AA",X"5A",X"88",X"88",X"AA",X"5A",X"88",X"88",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"E0",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"EE",X"00",X"00",X"11",X"EE",
		X"00",X"00",X"51",X"EE",X"00",X"00",X"51",X"EE",X"00",X"00",X"51",X"EE",X"00",X"00",X"11",X"EE",
		X"00",X"01",X"11",X"1E",X"00",X"00",X"11",X"EE",X"00",X"00",X"01",X"EE",X"00",X"00",X"10",X"EE",
		X"00",X"00",X"01",X"EE",X"00",X"00",X"40",X"EE",X"00",X"44",X"40",X"EE",X"00",X"44",X"46",X"1E",
		X"00",X"40",X"46",X"EE",X"00",X"06",X"46",X"EE",X"00",X"66",X"06",X"EE",X"00",X"66",X"66",X"EE",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"1E",X"00",X"11",X"66",X"E1",
		X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"10",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",
		X"31",X"00",X"66",X"00",X"33",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F4",X"06",X"00",X"00",
		X"44",X"46",X"00",X"E0",X"44",X"41",X"00",X"1E",X"44",X"44",X"00",X"EE",X"44",X"44",X"00",X"EE",
		X"11",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"70",X"44",X"00",X"EE",
		X"70",X"44",X"00",X"1E",X"41",X"44",X"00",X"EE",X"44",X"41",X"00",X"EE",X"14",X"11",X"00",X"EE",
		X"01",X"00",X"00",X"EE",X"00",X"00",X"40",X"EE",X"00",X"44",X"40",X"EE",X"00",X"44",X"46",X"1E",
		X"00",X"40",X"46",X"EE",X"00",X"06",X"46",X"EE",X"00",X"66",X"06",X"EE",X"00",X"66",X"66",X"EE",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"1E",X"00",X"11",X"66",X"E1",
		X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"10",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",
		X"31",X"00",X"66",X"00",X"F3",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"04",X"06",X"00",X"00",
		X"44",X"46",X"00",X"E0",X"44",X"41",X"00",X"1E",X"44",X"44",X"00",X"EE",X"44",X"44",X"00",X"EE",
		X"11",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",X"00",X"44",X"00",X"EE",
		X"00",X"44",X"00",X"1E",X"01",X"44",X"00",X"EE",X"1A",X"41",X"00",X"EE",X"44",X"11",X"00",X"EE",
		X"44",X"00",X"00",X"EE",X"11",X"00",X"40",X"EE",X"01",X"44",X"40",X"EE",X"00",X"44",X"46",X"1E",
		X"00",X"40",X"46",X"EE",X"00",X"06",X"46",X"EE",X"00",X"66",X"06",X"EE",X"00",X"66",X"66",X"EE",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"1E",X"00",X"11",X"66",X"E1",
		X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"10",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"C0",X"EE",X"00",X"00",X"00",X"66",X"EE",X"00",
		X"00",X"06",X"0E",X"00",X"06",X"66",X"EE",X"00",X"06",X"60",X"E0",X"00",X"66",X"66",X"EE",X"00",
		X"6A",X"E6",X"EE",X"00",X"66",X"AA",X"0E",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"D0",
		X"6C",X"00",X"00",X"00",X"6A",X"00",X"0E",X"00",X"6A",X"00",X"66",X"00",X"6A",X"A0",X"66",X"00",
		X"66",X"AA",X"EA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"A0",X"00",X"00",X"AA",X"66",X"00",
		X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",X"FF",X"50",X"00",
		X"00",X"FF",X"50",X"00",X"00",X"FB",X"50",X"00",X"00",X"BB",X"50",X"00",X"00",X"5A",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"50",X"00",X"00",X"B0",X"50",X"00",
		X"00",X"00",X"50",X"00",X"00",X"90",X"50",X"00",X"00",X"99",X"50",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",X"AF",X"50",X"00",X"00",X"FF",X"50",X"00",
		X"00",X"FF",X"50",X"00",X"00",X"FB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"55",X"90",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",X"FF",X"50",X"00",
		X"00",X"FF",X"50",X"00",X"00",X"FB",X"50",X"00",X"00",X"BB",X"50",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"09",X"33",
		X"00",X"33",X"00",X"93",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"39",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"39",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"39",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"99",X"00",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"99",X"00",X"99",X"30",X"00",X"00",X"09",X"30",X"00",
		X"33",X"00",X"33",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"33",
		X"00",X"33",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"39",X"00",X"33",X"00",X"99",X"00",X"33",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"B9",X"00",X"00",X"00",X"99",X"07",X"00",X"00",X"09",X"75",X"00",X"00",X"99",X"70",
		X"00",X"00",X"99",X"50",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"0B",X"99",X"AA",X"00",X"00",X"99",X"EE",X"00",X"00",X"90",X"00",X"00",X"B0",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"90",X"99",X"AA",X"00",X"99",X"99",X"EE",X"09",X"99",X"99",X"00",
		X"90",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"70",X"B9",X"90",X"99",X"70",
		X"99",X"99",X"99",X"57",X"90",X"99",X"99",X"05",X"09",X"99",X"99",X"00",X"09",X"9B",X"99",X"99",
		X"90",X"99",X"99",X"99",X"00",X"99",X"09",X"99",X"00",X"09",X"99",X"99",X"00",X"90",X"99",X"99");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
