library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kbe2_IC5 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kbe2_IC5 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"97",X"01",X"05",X"8F",X"FF",X"DB",X"30",X"00",X"68",X"FF",X"FB",X"C2",X"30",X"36",X"AF",
		X"FE",X"C8",X"42",X"03",X"5D",X"DF",X"CF",X"55",X"02",X"37",X"ED",X"FC",X"E3",X"30",X"14",X"BF",
		X"FF",X"E8",X"50",X"00",X"5D",X"EF",X"CF",X"45",X"01",X"27",X"EE",X"FC",X"C4",X"40",X"14",X"AF",
		X"FF",X"F6",X"60",X"11",X"6C",X"EF",X"EC",X"63",X"11",X"39",X"DF",X"FF",X"67",X"02",X"07",X"CF",
		X"FF",X"C5",X"30",X"13",X"9C",X"FE",X"F5",X"60",X"11",X"7D",X"FF",X"FB",X"61",X"00",X"4A",X"EF",
		X"FF",X"44",X"01",X"38",X"DF",X"FF",X"85",X"00",X"06",X"CF",X"FF",X"E4",X"20",X"02",X"9F",X"FF",
		X"F7",X"60",X"00",X"6C",X"FF",X"FE",X"52",X"00",X"27",X"FF",X"FF",X"77",X"00",X"05",X"CF",X"FF",
		X"E6",X"10",X"03",X"8F",X"FF",X"F6",X"50",X"00",X"5C",X"FF",X"FB",X"60",X"00",X"5A",X"FF",X"FF",
		X"45",X"01",X"27",X"DF",X"FF",X"85",X"00",X"05",X"BF",X"FF",X"F5",X"20",X"02",X"8E",X"FF",X"F9",
		X"50",X"00",X"5B",X"FF",X"FF",X"62",X"00",X"37",X"EF",X"FF",X"85",X"00",X"05",X"BF",X"FF",X"E6",
		X"20",X"02",X"7D",X"FF",X"FA",X"50",X"00",X"5B",X"FF",X"FD",X"71",X"00",X"37",X"EF",X"FF",X"95",
		X"00",X"14",X"BE",X"FF",X"E7",X"10",X"03",X"7D",X"FF",X"FB",X"60",X"00",X"49",X"DF",X"FE",X"73",
		X"01",X"36",X"CF",X"FF",X"B6",X"10",X"14",X"9D",X"FF",X"F9",X"41",X"03",X"5B",X"EF",X"FD",X"72",
		X"00",X"48",X"CF",X"FF",X"A5",X"10",X"25",X"AD",X"FF",X"D8",X"31",X"24",X"8C",X"FF",X"EA",X"41",
		X"02",X"6B",X"FF",X"FB",X"62",X"01",X"59",X"EF",X"FD",X"73",X"01",X"38",X"DF",X"FF",X"93",X"00",
		X"26",X"CF",X"FF",X"A4",X"10",X"26",X"AF",X"FF",X"C6",X"10",X"15",X"9E",X"FF",X"D7",X"20",X"14",
		X"8D",X"FF",X"E9",X"30",X"13",X"7C",X"FF",X"FA",X"41",X"02",X"6B",X"FF",X"FB",X"51",X"02",X"5A",
		X"FF",X"FC",X"72",X"01",X"5A",X"EF",X"FC",X"73",X"12",X"59",X"DF",X"FC",X"83",X"11",X"48",X"DF",
		X"FD",X"84",X"11",X"38",X"CF",X"FD",X"94",X"21",X"37",X"BF",X"FE",X"95",X"21",X"37",X"BE",X"FE",
		X"A5",X"21",X"36",X"BE",X"FE",X"B6",X"31",X"36",X"AE",X"FF",X"B6",X"31",X"25",X"9D",X"FF",X"C8",
		X"42",X"25",X"9D",X"FF",X"C8",X"42",X"24",X"8C",X"FF",X"D9",X"52",X"24",X"7B",X"EF",X"DA",X"52",
		X"13",X"7B",X"EF",X"EA",X"62",X"13",X"6A",X"DF",X"EB",X"73",X"23",X"59",X"CF",X"FD",X"84",X"22",
		X"48",X"CF",X"FE",X"A5",X"21",X"36",X"AE",X"FE",X"B7",X"31",X"25",X"9D",X"FF",X"D9",X"42",X"24",
		X"7B",X"EF",X"EB",X"63",X"23",X"69",X"DF",X"FC",X"84",X"22",X"47",X"BE",X"FE",X"B7",X"32",X"35",
		X"9C",X"EE",X"D9",X"53",X"24",X"7A",X"CE",X"EB",X"85",X"33",X"57",X"AC",X"DD",X"A8",X"54",X"46",
		X"8A",X"CC",X"CA",X"75",X"55",X"78",X"AB",X"BB",X"A8",X"76",X"67",X"88",X"99",X"AA",X"98",X"87",
		X"77",X"78",X"8A",X"AB",X"A8",X"76",X"66",X"78",X"9B",X"CB",X"A8",X"76",X"55",X"78",X"AC",X"CB",
		X"97",X"65",X"56",X"7A",X"BC",X"CA",X"86",X"55",X"67",X"9A",X"BC",X"B9",X"75",X"56",X"78",X"AB",
		X"BA",X"98",X"76",X"78",X"99",X"99",X"88",X"88",X"89",X"99",X"98",X"77",X"78",X"9A",X"AA",X"A8",
		X"76",X"66",X"89",X"AB",X"BA",X"87",X"66",X"67",X"9A",X"BB",X"A9",X"87",X"66",X"78",X"9A",X"AA",
		X"98",X"77",X"78",X"89",X"99",X"98",X"88",X"88",X"98",X"88",X"88",X"88",X"89",X"99",X"98",X"77",
		X"77",X"89",X"9A",X"A9",X"87",X"77",X"88",X"9A",X"A9",X"98",X"77",X"78",X"9A",X"AA",X"98",X"77",
		X"77",X"89",X"AA",X"A9",X"87",X"77",X"88",X"9A",X"A9",X"88",X"77",X"88",X"99",X"99",X"98",X"88",
		X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",
		X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",
		X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"87",X"88",X"89",X"99",
		X"99",X"88",X"77",X"88",X"99",X"99",X"98",X"77",X"78",X"89",X"99",X"98",X"87",X"77",X"88",X"99",
		X"99",X"88",X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",
		X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"88",
		X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"99",X"99",
		X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"88",X"89",
		X"98",X"88",X"88",X"88",X"88",X"89",X"98",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"98",X"88",
		X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",
		X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"99",X"99",X"88",
		X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"89",X"98",X"89",X"88",
		X"88",X"89",X"89",X"89",X"99",X"87",X"88",X"89",X"88",X"88",X"89",X"89",X"88",X"88",X"89",X"99",
		X"88",X"88",X"88",X"88",X"98",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",
		X"98",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"99",X"99",X"98",X"88",X"98",X"98",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"98",
		X"88",X"77",X"77",X"78",X"89",X"9A",X"AA",X"AA",X"99",X"87",X"77",X"66",X"77",X"88",X"9A",X"AA",
		X"AA",X"A9",X"88",X"77",X"66",X"67",X"78",X"89",X"AA",X"BB",X"AA",X"99",X"87",X"66",X"66",X"67",
		X"78",X"9A",X"AB",X"BB",X"A9",X"87",X"76",X"66",X"66",X"78",X"89",X"AB",X"BB",X"BB",X"A9",X"87",
		X"66",X"66",X"67",X"78",X"9A",X"AB",X"BB",X"BA",X"98",X"77",X"66",X"66",X"67",X"77",X"99",X"AA",
		X"BB",X"BA",X"A9",X"87",X"76",X"66",X"67",X"78",X"89",X"AB",X"BB",X"BA",X"A8",X"97",X"87",X"87",
		X"88",X"88",X"77",X"77",X"78",X"89",X"AA",X"AA",X"A9",X"99",X"98",X"88",X"87",X"66",X"66",X"68",
		X"8A",X"BB",X"CB",X"B9",X"A8",X"97",X"87",X"87",X"77",X"66",X"67",X"79",X"9B",X"AC",X"BB",X"A9",
		X"88",X"87",X"87",X"87",X"76",X"76",X"77",X"99",X"BB",X"CB",X"BA",X"99",X"78",X"78",X"78",X"78",
		X"77",X"77",X"78",X"99",X"BA",X"CA",X"B9",X"98",X"87",X"88",X"78",X"78",X"77",X"67",X"78",X"9A",
		X"BB",X"CA",X"B9",X"A7",X"87",X"87",X"88",X"88",X"77",X"67",X"78",X"99",X"BA",X"CA",X"B8",X"97",
		X"87",X"87",X"88",X"78",X"77",X"66",X"77",X"99",X"CB",X"DA",X"C9",X"97",X"87",X"78",X"78",X"78",
		X"67",X"66",X"77",X"A8",X"CA",X"DA",X"B9",X"88",X"77",X"68",X"79",X"79",X"77",X"66",X"76",X"99",
		X"BC",X"CD",X"AB",X"79",X"68",X"68",X"88",X"88",X"87",X"75",X"57",X"6A",X"9D",X"BD",X"BB",X"97",
		X"86",X"86",X"87",X"98",X"88",X"66",X"56",X"77",X"B9",X"EA",X"E9",X"B8",X"77",X"68",X"69",X"79",
		X"89",X"86",X"65",X"67",X"7A",X"9D",X"AD",X"AA",X"97",X"86",X"86",X"87",X"98",X"88",X"66",X"56",
		X"77",X"9A",X"BD",X"BD",X"9B",X"69",X"67",X"77",X"88",X"98",X"97",X"76",X"56",X"87",X"BA",X"EB",
		X"DB",X"A9",X"68",X"57",X"68",X"88",X"A8",X"96",X"85",X"65",X"87",X"B9",X"EB",X"DB",X"A9",X"68",
		X"47",X"68",X"89",X"A9",X"A7",X"75",X"54",X"86",X"BA",X"EC",X"CD",X"8A",X"47",X"47",X"77",X"A8",
		X"B9",X"A7",X"75",X"44",X"57",X"8D",X"AF",X"AF",X"9A",X"65",X"65",X"77",X"8A",X"9C",X"9A",X"77",
		X"54",X"46",X"78",X"DA",X"FB",X"F9",X"A6",X"56",X"47",X"88",X"B9",X"C9",X"A7",X"65",X"33",X"37",
		X"6D",X"BF",X"ED",X"D7",X"A2",X"63",X"67",X"8B",X"BC",X"C9",X"95",X"63",X"33",X"48",X"8F",X"CF",
		X"DE",X"A7",X"72",X"43",X"68",X"AC",X"CC",X"C9",X"84",X"52",X"22",X"59",X"9F",X"DF",X"FD",X"C4",
		X"70",X"42",X"78",X"CB",X"FC",X"D8",X"85",X"33",X"12",X"47",X"AC",X"FD",X"FA",X"E5",X"52",X"14",
		X"59",X"BE",X"EF",X"BB",X"66",X"23",X"22",X"35",X"9B",X"EF",X"DF",X"8D",X"36",X"23",X"56",X"AC",
		X"DE",X"DB",X"96",X"53",X"34",X"34",X"58",X"BA",X"FB",X"FA",X"C8",X"55",X"24",X"68",X"CC",X"EE",
		X"CB",X"76",X"44",X"44",X"35",X"4B",X"8F",X"FD",X"F9",X"D5",X"54",X"24",X"68",X"DC",X"FD",X"BB",
		X"67",X"34",X"44",X"34",X"3A",X"7E",X"FD",X"F9",X"D7",X"44",X"24",X"67",X"CE",X"DF",X"BC",X"76",
		X"43",X"44",X"44",X"46",X"B9",X"FE",X"EF",X"9C",X"54",X"43",X"59",X"8E",X"DD",X"F8",X"B4",X"54",
		X"35",X"65",X"64",X"7A",X"8E",X"ED",X"F9",X"C6",X"55",X"45",X"88",X"CE",X"BE",X"8A",X"65",X"54",
		X"57",X"56",X"44",X"98",X"AF",X"BF",X"E9",X"C3",X"64",X"56",X"98",X"EB",X"CB",X"79",X"57",X"56",
		X"67",X"45",X"25",X"88",X"EF",X"FF",X"CB",X"85",X"44",X"37",X"7A",X"CB",X"DB",X"A8",X"76",X"66",
		X"55",X"33",X"25",X"99",X"FF",X"FF",X"DB",X"75",X"34",X"36",X"8A",X"DD",X"DC",X"A9",X"76",X"55",
		X"45",X"44",X"34",X"9A",X"EF",X"FF",X"DB",X"75",X"23",X"35",X"9A",X"DD",X"DD",X"A9",X"76",X"45",
		X"55",X"54",X"54",X"8B",X"CF",X"FF",X"FB",X"87",X"33",X"44",X"79",X"AE",X"CC",X"C8",X"86",X"54",
		X"55",X"65",X"55",X"59",X"AC",X"FF",X"EF",X"A9",X"64",X"34",X"47",X"AA",X"ED",X"DC",X"97",X"64",
		X"46",X"57",X"66",X"55",X"7A",X"AE",X"FE",X"FB",X"97",X"43",X"44",X"69",X"AD",X"ED",X"CA",X"76",
		X"54",X"56",X"67",X"66",X"55",X"8A",X"BF",X"FE",X"FA",X"85",X"32",X"44",X"8A",X"BE",X"EC",X"B8",
		X"65",X"55",X"68",X"78",X"75",X"44",X"8A",X"BF",X"FF",X"FB",X"85",X"31",X"43",X"8A",X"CE",X"FC",
		X"B9",X"56",X"45",X"68",X"79",X"76",X"54",X"5A",X"9D",X"FD",X"FC",X"A5",X"50",X"35",X"6B",X"CD",
		X"DE",X"9A",X"65",X"56",X"78",X"98",X"96",X"53",X"24",X"99",X"EF",X"EF",X"D9",X"56",X"13",X"56",
		X"AC",X"EC",X"EA",X"97",X"65",X"77",X"79",X"78",X"75",X"33",X"26",X"AB",X"FF",X"FF",X"D7",X"64",
		X"14",X"58",X"AD",X"CD",X"CA",X"88",X"66",X"77",X"88",X"77",X"64",X"32",X"26",X"BD",X"FF",X"FF",
		X"C7",X"32",X"01",X"57",X"BE",X"FE",X"EB",X"86",X"54",X"56",X"78",X"88",X"76",X"53",X"24",X"9D",
		X"FF",X"FF",X"E9",X"41",X"10",X"36",X"BD",X"FF",X"DB",X"85",X"34",X"46",X"8A",X"AA",X"96",X"54",
		X"22",X"49",X"EF",X"FF",X"FC",X"73",X"01",X"05",X"9E",X"FF",X"FB",X"95",X"52",X"56",X"8A",X"BA",
		X"88",X"55",X"44",X"35",X"7C",X"FF",X"FF",X"D8",X"62",X"13",X"48",X"AF",X"EF",X"C9",X"65",X"54",
		X"68",X"AA",X"BA",X"87",X"54",X"45",X"45",X"69",X"DE",X"FF",X"EC",X"87",X"43",X"56",X"8A",X"CB",
		X"B9",X"85",X"56",X"78",X"AB",X"AA",X"97",X"55",X"55",X"56",X"66",X"8B",X"EE",X"FF",X"DA",X"76",
		X"23",X"35",X"7A",X"CC",X"DB",X"A7",X"76",X"76",X"89",X"99",X"98",X"77",X"76",X"67",X"65",X"79",
		X"DE",X"FF",X"C9",X"65",X"23",X"47",X"AC",X"FE",X"C9",X"84",X"34",X"57",X"9C",X"CC",X"A9",X"76",
		X"65",X"55",X"66",X"56",X"8C",X"DE",X"FE",X"C9",X"74",X"33",X"67",X"9B",X"CC",X"BA",X"86",X"56",
		X"78",X"AA",X"BA",X"97",X"66",X"66",X"67",X"77",X"67",X"9E",X"EE",X"FD",X"95",X"53",X"34",X"8B",
		X"CE",X"EC",X"87",X"54",X"35",X"79",X"CC",X"CA",X"97",X"66",X"66",X"67",X"77",X"66",X"7A",X"DC",
		X"ED",X"D8",X"76",X"55",X"6A",X"AB",X"BC",X"97",X"65",X"54",X"79",X"BD",X"DD",X"A9",X"65",X"44",
		X"45",X"68",X"98",X"88",X"AD",X"CC",X"CD",X"97",X"66",X"55",X"89",X"AA",X"CB",X"98",X"77",X"67",
		X"89",X"AA",X"BA",X"98",X"87",X"77",X"76",X"66",X"66",X"66",X"AD",X"DD",X"DD",X"97",X"65",X"55",
		X"89",X"AA",X"BA",X"87",X"67",X"67",X"8A",X"BB",X"CB",X"96",X"65",X"55",X"67",X"78",X"88",X"76",
		X"9C",X"CD",X"DE",X"A7",X"55",X"44",X"79",X"BB",X"CB",X"97",X"55",X"56",X"69",X"BC",X"CC",X"B8",
		X"75",X"55",X"56",X"78",X"88",X"87",X"9C",X"DD",X"CD",X"B8",X"55",X"55",X"68",X"AB",X"BB",X"A8",
		X"66",X"67",X"78",X"AB",X"BA",X"A8",X"76",X"66",X"66",X"78",X"87",X"77",X"79",X"CD",X"DC",X"DA",
		X"85",X"56",X"67",X"8B",X"BB",X"A9",X"76",X"55",X"77",X"9B",X"DC",X"BA",X"87",X"55",X"56",X"67",
		X"89",X"98",X"87",X"8B",X"CC",X"BC",X"B8",X"65",X"66",X"78",X"BC",X"BA",X"98",X"66",X"57",X"89",
		X"9B",X"CB",X"A8",X"87",X"66",X"67",X"77",X"78",X"78",X"77",X"AC",X"DC",X"CC",X"A8",X"56",X"67",
		X"78",X"BB",X"A8",X"87",X"76",X"78",X"99",X"9B",X"BA",X"87",X"77",X"66",X"78",X"88",X"78",X"87",
		X"66",X"8C",X"DC",X"BC",X"B9",X"65",X"67",X"88",X"AB",X"A9",X"87",X"77",X"67",X"89",X"AA",X"AA",
		X"A8",X"88",X"87",X"67",X"77",X"66",X"78",X"88",X"79",X"CD",X"CA",X"BA",X"96",X"56",X"78",X"79",
		X"AA",X"98",X"88",X"87",X"77",X"88",X"89",X"9A",X"AA",X"99",X"87",X"66",X"66",X"66",X"78",X"99",
		X"89",X"AB",X"BB",X"AA",X"98",X"66",X"77",X"88",X"9A",X"A9",X"88",X"88",X"77",X"89",X"99",X"99");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
