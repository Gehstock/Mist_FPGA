library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prg_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prg_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FB",X"E5",X"76",X"39",X"88",X"58",X"3F",X"3A",X"C6",X"48",X"6B",X"B3",X"88",X"2F",X"20",X"42",
		X"55",X"53",X"54",X"59",X"20",X"2F",X"2F",X"20",X"46",X"4C",X"49",X"50",X"50",X"59",X"20",X"2F",
		X"DC",X"23",X"CC",X"7A",X"20",X"53",X"45",X"47",X"41",X"20",X"31",X"39",X"38",X"34",X"2F",X"30",
		X"35",X"2F",X"32",X"34",X"35",X"50",X"B7",X"69",X"4B",X"2D",X"3E",X"CD",X"60",X"AA",X"6D",X"F1",
		X"AC",X"C5",X"0F",X"22",X"3F",X"D3",X"AC",X"AF",X"67",X"66",X"AF",X"F6",X"AF",X"28",X"89",X"17",
		X"92",X"DA",X"E8",X"50",X"46",X"50",X"AF",X"0F",X"AF",X"0F",X"76",X"AF",X"80",X"89",X"1F",X"32",
		X"DD",X"48",X"3F",X"D3",X"98",X"C3",X"D7",X"A8",X"8A",X"D3",X"AD",X"AF",X"B2",X"2C",X"48",X"C5",
		X"64",X"D4",X"6D",X"56",X"0B",X"CD",X"FF",X"AB",X"6D",X"1D",X"0A",X"CD",X"9A",X"AA",X"6D",X"43",
		X"AB",X"BE",X"8B",X"3A",X"88",X"48",X"3F",X"3A",X"89",X"48",X"4D",X"A3",X"AC",X"BA",X"D8",X"48",
		X"07",X"CA",X"96",X"88",X"1F",X"DB",X"08",X"CB",X"DF",X"CA",X"7B",X"8D",X"6B",X"67",X"A0",X"CB",
		X"4B",X"EF",X"6A",X"84",X"88",X"BA",X"D8",X"48",X"DE",X"2A",X"B0",X"A8",X"92",X"2E",X"48",X"C3",
		X"C7",X"20",X"30",X"CB",X"E7",X"00",X"2F",X"12",X"78",X"48",X"76",X"8A",X"90",X"AE",X"B2",X"E7",
		X"48",X"BC",X"DE",X"2B",X"90",X"29",X"3F",X"3A",X"E7",X"48",X"10",X"BC",X"4D",X"12",X"AB",X"17",
		X"92",X"88",X"E8",X"CD",X"AB",X"AB",X"92",X"8B",X"E8",X"16",X"29",X"32",X"2D",X"48",X"B6",X"8A",
		X"6B",X"C5",X"88",X"17",X"B2",X"52",X"48",X"3A",X"88",X"48",X"B2",X"2D",X"48",X"3A",X"89",X"48",
		X"1F",X"32",X"47",X"48",X"92",X"8E",X"E8",X"CD",X"9A",X"AA",X"6D",X"3A",X"0B",X"EB",X"2D",X"89",
		X"96",X"29",X"B2",X"28",X"40",X"C5",X"03",X"23",X"B2",X"2A",X"40",X"BA",X"08",X"48",X"EE",X"29",
		X"20",X"25",X"21",X"47",X"E8",X"39",X"F8",X"48",X"36",X"28",X"29",X"2D",X"28",X"C5",X"B0",X"12",
		X"0C",X"48",X"EE",X"29",X"80",X"20",X"92",X"29",X"40",X"76",X"00",X"3A",X"09",X"48",X"96",X"29",
		X"32",X"50",X"E8",X"76",X"21",X"20",X"E8",X"36",X"28",X"39",X"09",X"48",X"29",X"68",X"28",X"C5",
		X"B8",X"BA",X"0A",X"48",X"B2",X"21",X"40",X"29",X"00",X"48",X"31",X"09",X"40",X"3E",X"08",X"09",
		X"68",X"28",X"C5",X"B0",X"12",X"2B",X"E8",X"32",X"A9",X"48",X"21",X"28",X"CC",X"39",X"29",X"44",
		X"B6",X"28",X"21",X"A8",X"08",X"E5",X"B8",X"C5",X"8D",X"23",X"92",X"E7",X"40",X"27",X"96",X"28",
		X"20",X"3E",X"12",X"28",X"E8",X"E6",X"29",X"00",X"3D",X"12",X"46",X"48",X"14",X"32",X"46",X"48",
		X"EE",X"29",X"96",X"2D",X"A0",X"2A",X"96",X"A9",X"B2",X"3C",X"40",X"43",X"17",X"29",X"4D",X"0D",
		X"27",X"12",X"3C",X"48",X"32",X"04",X"E8",X"CD",X"01",X"25",X"12",X"3B",X"E8",X"32",X"8B",X"48",
		X"A1",X"28",X"43",X"19",X"08",X"46",X"21",X"28",X"09",X"E5",X"B8",X"C5",X"F9",X"24",X"96",X"29",
		X"32",X"50",X"E8",X"76",X"CD",X"A9",X"6D",X"CD",X"03",X"24",X"CD",X"9C",X"0C",X"21",X"20",X"48",
		X"B6",X"28",X"31",X"A9",X"40",X"09",X"AF",X"28",X"CD",X"30",X"4D",X"12",X"8A",X"C5",X"15",X"22",
		X"21",X"28",X"28",X"22",X"0A",X"48",X"BF",X"32",X"04",X"48",X"32",X"4C",X"E8",X"12",X"18",X"48",
		X"94",X"4F",X"EE",X"2B",X"DE",X"2B",X"A0",X"AB",X"96",X"29",X"B2",X"A4",X"40",X"F8",X"EE",X"B4",
		X"0F",X"D6",X"18",X"10",X"08",X"FE",X"3E",X"D6",X"18",X"10",X"2A",X"FE",X"3E",X"4F",X"2E",X"28",
		X"A1",X"16",X"9D",X"89",X"46",X"2B",X"E6",X"E9",X"A2",X"6A",X"48",X"BE",X"77",X"3A",X"97",X"48",
		X"6D",X"91",X"24",X"2E",X"28",X"21",X"FE",X"9A",X"B2",X"B8",X"E8",X"D6",X"3F",X"10",X"0D",X"D6",
		X"A7",X"B8",X"8C",X"F6",X"CF",X"B8",X"8D",X"0E",X"89",X"29",X"86",X"3B",X"D0",X"3A",X"BD",X"48",
		X"99",X"C0",X"DC",X"29",X"38",X"88",X"65",X"B0",X"99",X"00",X"DC",X"29",X"38",X"88",X"65",X"B0",
		X"31",X"C8",X"7C",X"09",X"98",X"28",X"CD",X"30",X"31",X"A8",X"7D",X"09",X"98",X"28",X"CD",X"30",
		X"99",X"C0",X"DD",X"29",X"38",X"88",X"65",X"B0",X"B2",X"B2",X"E8",X"15",X"EF",X"2E",X"28",X"21",
		X"F5",X"3E",X"92",X"35",X"48",X"27",X"80",X"2B",X"A1",X"0B",X"9E",X"89",X"D6",X"3A",X"A7",X"54",
		X"92",X"77",X"DD",X"12",X"12",X"48",X"B5",X"2F",X"8F",X"2F",X"EF",X"2E",X"28",X"21",X"F6",X"9B",
		X"92",X"35",X"48",X"27",X"80",X"2B",X"A1",X"AE",X"9C",X"89",X"31",X"30",X"7C",X"09",X"A8",X"28",
		X"65",X"B0",X"A2",X"BA",X"E8",X"29",X"08",X"88",X"A9",X"22",X"43",X"48",X"81",X"70",X"29",X"22",
		X"BA",X"48",X"4D",X"17",X"BE",X"C5",X"73",X"21",X"4D",X"75",X"AB",X"BA",X"E7",X"48",X"DE",X"2A",
		X"80",X"AB",X"8E",X"80",X"81",X"7A",X"31",X"39",X"28",X"4B",X"4B",X"5B",X"2A",X"2E",X"18",X"39",
		X"88",X"4C",X"A1",X"E2",X"91",X"BA",X"A4",X"48",X"AF",X"A8",X"A8",X"29",X"3A",X"B9",X"31",X"28",
		X"EB",X"2E",X"20",X"50",X"8E",X"88",X"6D",X"9F",X"0B",X"16",X"30",X"32",X"C3",X"4E",X"B6",X"8A",
		X"B2",X"C4",X"4E",X"BA",X"40",X"4E",X"4B",X"97",X"B2",X"C8",X"4E",X"17",X"B2",X"DA",X"4E",X"3A",
		X"F3",X"4E",X"92",X"A0",X"E8",X"16",X"D7",X"32",X"11",X"48",X"B2",X"A4",X"E8",X"A7",X"A0",X"8D",
		X"96",X"17",X"6B",X"38",X"0B",X"BA",X"1C",X"48",X"47",X"0E",X"08",X"29",X"52",X"3B",X"01",X"FE",
		X"32",X"21",X"EC",X"16",X"29",X"32",X"08",X"4C",X"32",X"A9",X"E8",X"16",X"A9",X"32",X"1A",X"4C",
		X"96",X"EF",X"B2",X"AD",X"40",X"BE",X"C7",X"3A",X"2E",X"48",X"3F",X"3A",X"0F",X"4C",X"B2",X"3D",
		X"E8",X"12",X"47",X"48",X"D6",X"2A",X"20",X"22",X"BF",X"32",X"6C",X"48",X"CD",X"A3",X"08",X"EB",
		X"81",X"2C",X"92",X"A4",X"40",X"27",X"80",X"B2",X"96",X"40",X"B2",X"21",X"43",X"3A",X"A9",X"4B",
		X"21",X"10",X"28",X"22",X"2F",X"4B",X"21",X"00",X"29",X"22",X"27",X"4B",X"16",X"99",X"32",X"A8",
		X"43",X"D5",X"A1",X"28",X"43",X"C5",X"93",X"32",X"5D",X"29",X"28",X"4B",X"4D",X"13",X"9A",X"C5",
		X"92",X"6C",X"DD",X"21",X"68",X"4B",X"CD",X"12",X"7A",X"DD",X"21",X"E8",X"EB",X"CD",X"9A",X"7A",
		X"96",X"21",X"FD",X"C5",X"CD",X"23",X"5D",X"FE",X"0D",X"F6",X"88",X"38",X"5E",X"AA",X"EB",X"48",
		X"5D",X"7C",X"DD",X"46",X"2F",X"DD",X"66",X"20",X"B7",X"C5",X"7A",X"54",X"E6",X"29",X"DD",X"77",
		X"88",X"D5",X"F5",X"2F",X"5D",X"FE",X"0D",X"0F",X"27",X"0F",X"5D",X"7F",X"18",X"29",X"79",X"B3",
		X"DD",X"75",X"2B",X"DD",X"74",X"2C",X"DD",X"36",X"0D",X"28",X"12",X"30",X"E8",X"E6",X"D4",X"0F",
		X"DE",X"2C",X"90",X"2A",X"96",X"2C",X"CD",X"4C",X"6E",X"2F",X"5D",X"4E",X"0D",X"B0",X"B0",X"2C",
		X"DD",X"36",X"0D",X"29",X"21",X"9C",X"33",X"DD",X"75",X"29",X"DD",X"74",X"2A",X"CD",X"9B",X"32",
		X"6B",X"70",X"0C",X"F6",X"88",X"A8",X"EE",X"BA",X"AC",X"48",X"AF",X"A8",X"E8",X"D5",X"D6",X"2D",
		X"D6",X"36",X"30",X"E9",X"12",X"30",X"E8",X"14",X"D6",X"38",X"10",X"29",X"BF",X"E6",X"0C",X"0F",
		X"47",X"0E",X"88",X"29",X"DE",X"3C",X"01",X"CE",X"A3",X"6E",X"C1",X"D5",X"D6",X"2D",X"7E",X"21",
		X"8F",X"2F",X"EF",X"09",X"F6",X"DD",X"D7",X"8F",X"83",X"56",X"7D",X"77",X"08",X"23",X"F6",X"DD",
		X"F7",X"3A",X"4B",X"FF",X"A0",X"2C",X"94",X"43",X"A3",X"2C",X"95",X"D5",X"F7",X"23",X"5D",X"3E",
		X"1C",X"88",X"6B",X"57",X"A0",X"A8",X"7D",X"CB",X"28",X"4E",X"7D",X"CB",X"1C",X"4E",X"83",X"56",
		X"5D",X"7F",X"9C",X"D5",X"B6",X"21",X"69",X"D5",X"B6",X"32",X"88",X"D5",X"B6",X"24",X"88",X"C5",
		X"9B",X"BA",X"4B",X"F8",X"2C",X"CD",X"9A",X"C3",X"6D",X"F5",X"6C",X"F1",X"B4",X"D6",X"20",X"DA",
		X"0A",X"2B",X"5D",X"65",X"96",X"28",X"FD",X"C5",X"ED",X"23",X"5D",X"C3",X"88",X"F6",X"80",X"23",
		X"81",X"F3",X"2C",X"E5",X"7D",X"46",X"2B",X"DD",X"C6",X"8C",X"61",X"F1",X"B4",X"D6",X"08",X"20",
		X"8A",X"BE",X"A9",X"F6",X"BE",X"28",X"7F",X"D5",X"E9",X"17",X"B2",X"50",X"48",X"BA",X"88",X"48",
		X"46",X"89",X"4A",X"8C",X"2D",X"12",X"04",X"48",X"8E",X"09",X"07",X"20",X"2A",X"2E",X"AA",X"50",
		X"4D",X"BD",X"CD",X"BA",X"A4",X"48",X"AF",X"A8",X"9A",X"29",X"6A",X"38",X"31",X"5C",X"60",X"C5",
		X"FE",X"AA",X"6D",X"88",X"0B",X"CD",X"28",X"AB",X"4B",X"8C",X"2D",X"16",X"29",X"32",X"36",X"48",
		X"26",X"2C",X"92",X"28",X"48",X"66",X"08",X"28",X"BF",X"45",X"A1",X"8F",X"98",X"19",X"5A",X"C2",
		X"B2",X"89",X"E8",X"E6",X"29",X"00",X"2B",X"21",X"B6",X"98",X"6B",X"68",X"80",X"8E",X"6D",X"5E",
		X"AA",X"43",X"47",X"2C",X"4D",X"C5",X"AA",X"41",X"6D",X"F8",X"DE",X"2B",X"90",X"2E",X"4D",X"28",
		X"0B",X"EB",X"D5",X"8C",X"6D",X"14",X"0D",X"CD",X"28",X"AB",X"6D",X"14",X"0D",X"CD",X"28",X"AB",
		X"69",X"0D",X"A0",X"96",X"92",X"28",X"40",X"76",X"00",X"3A",X"08",X"48",X"B1",X"28",X"50",X"F3",
		X"BF",X"32",X"EB",X"48",X"21",X"28",X"EB",X"39",X"20",X"28",X"CB",X"56",X"20",X"21",X"14",X"D6",
		X"28",X"A8",X"A9",X"99",X"6B",X"32",X"0D",X"65",X"5D",X"61",X"B2",X"4B",X"40",X"19",X"B9",X"2D",
		X"FD",X"04",X"04",X"04",X"5E",X"04",X"7E",X"C3",X"C1",X"12",X"EB",X"48",X"14",X"D6",X"20",X"00",
		X"8B",X"19",X"28",X"28",X"5D",X"99",X"5D",X"65",X"E9",X"43",X"9A",X"2D",X"92",X"51",X"40",X"27",
		X"CA",X"E4",X"2D",X"CD",X"F6",X"23",X"CD",X"5F",X"0B",X"CD",X"1D",X"6D",X"CD",X"28",X"0B",X"CD",
		X"B4",X"66",X"3F",X"3A",X"D1",X"48",X"4D",X"F1",X"8C",X"43",X"7A",X"28",X"92",X"A4",X"40",X"27",
		X"CA",X"DF",X"2D",X"12",X"13",X"48",X"D6",X"3C",X"DA",X"E9",X"2F",X"12",X"14",X"48",X"A7",X"CA",
		X"86",X"2E",X"DE",X"A8",X"A0",X"32",X"A1",X"35",X"1E",X"19",X"1A",X"C3",X"4D",X"5E",X"8A",X"8E",
		X"09",X"21",X"03",X"3E",X"39",X"12",X"C3",X"CD",X"D8",X"22",X"29",X"28",X"38",X"CD",X"A2",X"3F",
		X"A1",X"2F",X"1E",X"19",X"5A",X"C2",X"4D",X"5E",X"8A",X"BA",X"BC",X"48",X"A1",X"64",X"E2",X"C5",
		X"EF",X"25",X"12",X"B5",X"E8",X"E6",X"2B",X"4F",X"2E",X"28",X"21",X"01",X"3E",X"09",X"5E",X"12",
		X"BD",X"48",X"EE",X"34",X"07",X"8F",X"AF",X"5F",X"80",X"20",X"6E",X"B8",X"C7",X"2E",X"89",X"2A",
		X"42",X"C2",X"53",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"EE",X"30",X"47",X"26",X"21",X"22",X"E4",
		X"E2",X"FB",X"EE",X"27",X"6E",X"B8",X"C7",X"2A",X"EE",X"C2",X"96",X"21",X"B2",X"F9",X"E2",X"CB",
		X"6A",X"CD",X"A2",X"3F",X"EB",X"06",X"2E",X"12",X"47",X"48",X"D6",X"2A",X"20",X"ED",X"12",X"6C",
		X"48",X"27",X"4A",X"E9",X"8F",X"BA",X"AA",X"48",X"DE",X"2F",X"5A",X"E9",X"8F",X"28",X"EC",X"BA",
		X"6C",X"48",X"76",X"8A",X"6A",X"C1",X"2F",X"16",X"2A",X"32",X"6C",X"48",X"6D",X"3A",X"0A",X"DD",
		X"ED",X"D5",X"A1",X"28",X"4C",X"C5",X"A2",X"6C",X"5D",X"C3",X"88",X"96",X"5D",X"29",X"C8",X"4B",
		X"6D",X"A2",X"6C",X"DD",X"6B",X"88",X"96",X"DD",X"81",X"88",X"ED",X"CD",X"02",X"CC",X"7D",X"CB",
		X"88",X"96",X"5D",X"29",X"80",X"4D",X"4D",X"A2",X"CC",X"D5",X"4B",X"28",X"36",X"D5",X"E9",X"C5",
		X"D3",X"A9",X"81",X"1C",X"C2",X"CD",X"EC",X"F0",X"4B",X"C1",X"2F",X"D6",X"0E",X"DA",X"61",X"8F",
		X"6B",X"FA",X"88",X"BA",X"9B",X"48",X"DE",X"D7",X"6A",X"E9",X"8F",X"BA",X"40",X"4D",X"EE",X"08",
		X"4A",X"C1",X"2F",X"21",X"28",X"4B",X"89",X"80",X"28",X"1E",X"08",X"CB",X"F6",X"EA",X"61",X"8F",
		X"15",X"A8",X"8C",X"89",X"6B",X"F3",X"8E",X"BA",X"96",X"48",X"AF",X"42",X"C1",X"2F",X"96",X"D7",
		X"92",X"97",X"E8",X"12",X"47",X"48",X"46",X"89",X"A0",X"AA",X"8E",X"8C",X"6D",X"88",X"0B",X"38",
		X"73",X"43",X"D2",X"28",X"92",X"A3",X"48",X"C5",X"CD",X"E9",X"96",X"06",X"4D",X"BD",X"CD",X"BA",
		X"04",X"48",X"07",X"EA",X"05",X"8F",X"B6",X"8F",X"92",X"E5",X"E8",X"21",X"64",X"61",X"B2",X"99",
		X"48",X"C5",X"4F",X"25",X"A1",X"F8",X"61",X"BA",X"98",X"48",X"4D",X"4F",X"AD",X"29",X"D6",X"3B",
		X"99",X"EC",X"C1",X"CD",X"FE",X"AA",X"81",X"08",X"3B",X"39",X"40",X"61",X"6D",X"5E",X"0A",X"21",
		X"0D",X"3B",X"31",X"FC",X"61",X"C5",X"5E",X"22",X"A1",X"10",X"98",X"19",X"EC",X"C2",X"4D",X"5E",
		X"0A",X"0E",X"2D",X"12",X"39",X"48",X"07",X"20",X"3A",X"12",X"38",X"48",X"46",X"D0",X"AF",X"0F",
		X"07",X"8F",X"AF",X"8E",X"08",X"F6",X"0A",X"B8",X"0A",X"CF",X"05",X"0E",X"08",X"C3",X"21",X"29",
		X"71",X"3E",X"09",X"ED",X"4E",X"23",X"6E",X"CD",X"A2",X"3F",X"E9",X"21",X"EE",X"3B",X"09",X"56",
		X"A3",X"6E",X"C7",X"0E",X"8A",X"8E",X"89",X"19",X"EA",X"C2",X"4D",X"52",X"8A",X"29",X"08",X"28",
		X"22",X"38",X"E8",X"12",X"E8",X"48",X"E6",X"24",X"0F",X"0F",X"4F",X"2E",X"28",X"21",X"2E",X"B8",
		X"01",X"FE",X"B2",X"E5",X"40",X"7E",X"92",X"38",X"40",X"F6",X"0C",X"B8",X"66",X"C5",X"76",X"23",
		X"CD",X"5F",X"0B",X"CD",X"9A",X"22",X"16",X"D7",X"32",X"E5",X"E8",X"CD",X"F3",X"24",X"EB",X"86",
		X"09",X"BA",X"E8",X"48",X"AF",X"28",X"09",X"7E",X"3F",X"3A",X"E8",X"48",X"92",X"28",X"40",X"66",
		X"29",X"CA",X"0C",X"2D",X"CD",X"99",X"0B",X"21",X"ED",X"48",X"CB",X"6E",X"23",X"EA",X"EF",X"2F",
		X"B5",X"FE",X"DE",X"C8",X"7A",X"2F",X"88",X"BA",X"58",X"48",X"AF",X"A8",X"89",X"C5",X"47",X"23",
		X"CD",X"5E",X"0A",X"EB",X"D3",X"2F",X"12",X"E7",X"E8",X"D6",X"29",X"20",X"3D",X"21",X"AA",X"38",
		X"31",X"3E",X"E2",X"C5",X"56",X"22",X"A1",X"04",X"18",X"19",X"14",X"C1",X"4D",X"5E",X"8A",X"43",
		X"D3",X"2F",X"21",X"0A",X"38",X"39",X"FE",X"C4",X"CD",X"5E",X"0A",X"21",X"8C",X"38",X"39",X"7C",
		X"E4",X"C5",X"56",X"22",X"6B",X"D3",X"0F",X"3D",X"D6",X"F6",X"60",X"52",X"0F",X"20",X"31",X"3E",
		X"C2",X"21",X"AA",X"38",X"CD",X"C5",X"0A",X"21",X"AA",X"38",X"39",X"5E",X"C4",X"CD",X"C5",X"22",
		X"31",X"1C",X"E1",X"29",X"84",X"38",X"4D",X"C5",X"8A",X"29",X"84",X"38",X"31",X"7C",X"E4",X"C5",
		X"C5",X"22",X"21",X"72",X"38",X"39",X"0C",X"C2",X"CD",X"C5",X"0A",X"BF",X"32",X"4E",X"E8",X"12",
		X"4D",X"48",X"CE",X"29",X"B2",X"4D",X"48",X"BA",X"D8",X"48",X"AF",X"C2",X"AC",X"2D",X"3F",X"D3",
		X"08",X"07",X"92",X"8E",X"E8",X"CB",X"C7",X"6F",X"4A",X"D2",X"28",X"12",X"78",X"48",X"76",X"89",
		X"4A",X"24",X"8D",X"C3",X"C0",X"42",X"D2",X"28",X"6B",X"24",X"8D",X"D5",X"ED",X"29",X"88",X"4B",
		X"1F",X"F5",X"45",X"DD",X"41",X"E5",X"7D",X"4E",X"2D",X"2E",X"28",X"CB",X"89",X"21",X"40",X"A8",
		X"92",X"6C",X"48",X"27",X"80",X"2B",X"A1",X"1C",X"A8",X"89",X"46",X"2B",X"E6",X"E9",X"21",X"7B",
		X"08",X"ED",X"61",X"12",X"6C",X"48",X"07",X"CC",X"9B",X"BA",X"41",X"29",X"20",X"88",X"A9",X"F1",
		X"94",X"F6",X"9B",X"28",X"6C",X"D5",X"E9",X"C1",X"E5",X"72",X"2E",X"20",X"A3",X"21",X"A3",X"21",
		X"03",X"A9",X"03",X"A9",X"03",X"A9",X"03",X"A9",X"09",X"A9",X"52",X"FA",X"8B",X"FA",X"A2",X"FA",
		X"31",X"72",X"58",X"72",X"47",X"72",X"76",X"72",X"A6",X"73",X"BD",X"73",X"B7",X"73",X"96",X"46",
		X"7D",X"77",X"09",X"C9",X"E9",X"A8",X"E9",X"A8",X"C0",X"A8",X"E9",X"A8",X"E9",X"A8",X"E9",X"A8",
		X"49",X"20",X"49",X"20",X"69",X"20",X"49",X"20",X"32",X"20",X"07",X"BC",X"07",X"BC",X"07",X"BC",
		X"A7",X"94",X"A7",X"94",X"6F",X"C0",X"33",X"C0",X"E9",X"A8",X"1F",X"32",X"0A",X"48",X"4B",X"19",
		X"C0",X"C5",X"A2",X"6C",X"5D",X"C3",X"88",X"96",X"49",X"C5",X"1D",X"22",X"A1",X"E8",X"88",X"2A",
		X"2F",X"4C",X"B6",X"C4",X"92",X"A9",X"EC",X"BF",X"7D",X"77",X"0D",X"21",X"1C",X"95",X"82",X"8B",
		X"4C",X"29",X"94",X"BC",X"A2",X"29",X"4C",X"C1",X"A1",X"A8",X"89",X"D5",X"F5",X"2F",X"5D",X"7C",
		X"08",X"16",X"64",X"DD",X"D7",X"A9",X"81",X"C1",X"15",X"DD",X"D5",X"89",X"7D",X"74",X"2A",X"21",
		X"5C",X"B3",X"5D",X"7D",X"0B",X"D5",X"F4",X"2C",X"49",X"BE",X"47",X"3A",X"89",X"4C",X"A1",X"A8",
		X"2A",X"22",X"2F",X"4C",X"16",X"C6",X"32",X"3A",X"EC",X"BF",X"32",X"24",X"EC",X"32",X"3F",X"4C",
		X"96",X"99",X"B2",X"28",X"44",X"BE",X"09",X"3A",X"4D",X"48",X"49",X"43",X"FD",X"6C",X"92",X"28",
		X"E8",X"E6",X"57",X"32",X"28",X"48",X"12",X"A4",X"E8",X"A7",X"00",X"2E",X"CD",X"DB",X"0C",X"EB",
		X"A5",X"21",X"92",X"2C",X"40",X"66",X"8C",X"F6",X"8C",X"C2",X"A5",X"21",X"A1",X"2A",X"40",X"BA",
		X"29",X"48",X"E6",X"29",X"00",X"2B",X"21",X"2B",X"E8",X"35",X"EA",X"85",X"09",X"12",X"28",X"48",
		X"EE",X"29",X"A0",X"3D",X"96",X"0F",X"4D",X"BD",X"4D",X"29",X"02",X"38",X"31",X"5E",X"E4",X"C5",
		X"FE",X"22",X"2E",X"21",X"CD",X"28",X"0B",X"38",X"D3",X"CD",X"CC",X"24",X"CD",X"DE",X"0B",X"CD",
		X"57",X"23",X"4D",X"1D",X"8A",X"C5",X"92",X"22",X"A1",X"47",X"40",X"BA",X"09",X"48",X"EE",X"29",
		X"00",X"2B",X"21",X"5A",X"E8",X"CD",X"84",X"FC",X"CD",X"35",X"6D",X"12",X"29",X"48",X"E6",X"2A",
		X"4A",X"FA",X"08",X"C5",X"E4",X"21",X"4A",X"FA",X"08",X"0E",X"09",X"98",X"0A",X"0E",X"0C",X"C5",
		X"28",X"23",X"38",X"D3",X"CD",X"35",X"6D",X"16",X"29",X"32",X"D8",X"48",X"CD",X"DE",X"0B",X"CD",
		X"57",X"23",X"92",X"29",X"40",X"66",X"0A",X"C2",X"A6",X"29",X"4D",X"C4",X"89",X"C2",X"A6",X"29",
		X"21",X"20",X"E8",X"39",X"A8",X"48",X"0E",X"68",X"CD",X"81",X"0D",X"21",X"28",X"4B",X"39",X"28",
		X"C6",X"8E",X"08",X"C5",X"A1",X"25",X"4D",X"AA",X"8C",X"43",X"A6",X"29",X"92",X"29",X"40",X"66",
		X"29",X"12",X"2A",X"48",X"20",X"2B",X"12",X"2B",X"E8",X"A7",X"C9",X"12",X"28",X"48",X"E6",X"29",
		X"80",X"2E",X"4D",X"79",X"AA",X"43",X"9C",X"22",X"A1",X"BE",X"9E",X"19",X"52",X"C6",X"4D",X"5E",
		X"0A",X"CD",X"7B",X"AC",X"AE",X"A9",X"81",X"CA",X"38",X"39",X"08",X"60",X"6D",X"4C",X"0A",X"12",
		X"89",X"48",X"EE",X"2A",X"A0",X"34",X"92",X"28",X"48",X"66",X"89",X"A8",X"8E",X"BA",X"8D",X"48",
		X"07",X"20",X"0F",X"39",X"24",X"60",X"81",X"EA",X"38",X"CD",X"EC",X"AA",X"6D",X"BA",X"18",X"EB",
		X"C1",X"30",X"A1",X"6E",X"98",X"19",X"84",X"C0",X"4D",X"4C",X"AA",X"C5",X"BA",X"30",X"6B",X"70",
		X"18",X"21",X"4E",X"98",X"99",X"60",X"C6",X"EB",X"FE",X"AA",X"EF",X"2E",X"28",X"09",X"F6",X"C9",
		X"3F",X"53",X"BA",X"BE",X"2F",X"53",X"BA",X"BE",X"8F",X"53",X"BA",X"17",X"7B",X"33",X"96",X"47",
		X"5B",X"BB",X"1F",X"FB",X"1B",X"16",X"2F",X"FB",X"1B",X"C9",X"81",X"C7",X"E8",X"36",X"2C",X"D3",
		X"F6",X"FE",X"AF",X"28",X"72",X"73",X"49",X"29",X"88",X"48",X"31",X"29",X"48",X"09",X"50",X"27",
		X"96",X"88",X"65",X"B0",X"69",X"21",X"28",X"40",X"B8",X"8B",X"81",X"88",X"C0",X"29",X"D7",X"8E",
		X"B6",X"28",X"55",X"5C",X"33",X"E5",X"B8",X"C1",X"A1",X"58",X"66",X"BA",X"D8",X"48",X"4D",X"B5",
		X"0B",X"F5",X"F0",X"D6",X"30",X"00",X"2D",X"70",X"83",X"36",X"08",X"03",X"51",X"23",X"83",X"77",
		X"A3",X"3E",X"A8",X"C1",X"66",X"2B",X"D6",X"1A",X"A3",X"1B",X"AF",X"BE",X"A8",X"A8",X"8A",X"BE",
		X"09",X"3A",X"9B",X"38",X"F1",X"C9",X"AE",X"A8",X"CE",X"23",X"F6",X"3A",X"83",X"3B",X"07",X"00",
		X"8F",X"F6",X"C8",X"BE",X"A8",X"38",X"89",X"F9",X"32",X"1B",X"30",X"C6",X"49",X"4E",X"96",X"A8",
		X"9A",X"3B",X"B6",X"88",X"9A",X"3B",X"98",X"56",X"69",X"F5",X"45",X"21",X"28",X"80",X"B8",X"8D",
		X"FD",X"65",X"A1",X"28",X"00",X"AB",X"D5",X"34",X"A0",X"D3",X"E9",X"71",X"49",X"19",X"08",X"4B",
		X"21",X"71",X"31",X"56",X"2E",X"28",X"23",X"4E",X"23",X"E5",X"66",X"41",X"0E",X"2D",X"C5",X"B0",
		X"06",X"32",X"C3",X"6A",X"33",X"3E",X"08",X"E5",X"B8",X"61",X"A3",X"BD",X"A0",X"C1",X"26",X"A8",
		X"BF",X"21",X"2D",X"4B",X"39",X"A8",X"28",X"77",X"14",X"19",X"38",X"D3",X"C9",X"F5",X"E6",X"D8",
		X"07",X"8F",X"07",X"8F",X"6E",X"B8",X"67",X"71",X"EE",X"27",X"6E",X"B8",X"49",X"07",X"C7",X"2E",
		X"28",X"29",X"54",X"66",X"09",X"56",X"23",X"66",X"47",X"E5",X"DD",X"E1",X"C9",X"21",X"2A",X"48",
		X"92",X"29",X"40",X"66",X"09",X"A8",X"0B",X"29",X"0B",X"48",X"D6",X"BD",X"06",X"2F",X"A1",X"4C",
		X"C6",X"A7",X"39",X"A8",X"28",X"00",X"2C",X"39",X"28",X"27",X"15",X"73",X"23",X"72",X"23",X"0D",
		X"A0",X"C7",X"49",X"BA",X"08",X"48",X"EE",X"29",X"80",X"2B",X"96",X"29",X"49",X"BA",X"0C",X"48",
		X"E6",X"24",X"0F",X"0F",X"21",X"8B",X"38",X"EB",X"5A",X"22",X"12",X"78",X"E8",X"15",X"6F",X"E6",
		X"8F",X"F6",X"8F",X"F8",X"26",X"28",X"A0",X"2C",X"EE",X"D8",X"26",X"21",X"B8",X"3A",X"58",X"48",
		X"C9",X"12",X"78",X"48",X"D6",X"2A",X"21",X"BB",X"38",X"10",X"2B",X"21",X"12",X"38",X"39",X"4A",
		X"E6",X"C5",X"56",X"22",X"6B",X"80",X"8A",X"29",X"DA",X"38",X"31",X"24",X"E2",X"BA",X"58",X"48",
		X"D6",X"29",X"C8",X"21",X"46",X"38",X"C9",X"21",X"67",X"48",X"36",X"20",X"D3",X"76",X"56",X"A7",
		X"A0",X"D2",X"49",X"29",X"63",X"29",X"92",X"29",X"40",X"66",X"09",X"A8",X"0A",X"E5",X"64",X"2A",
		X"D4",X"C7",X"22",X"E1",X"E8",X"C9",X"21",X"28",X"E9",X"39",X"29",X"49",X"36",X"28",X"29",X"D7",
		X"89",X"E5",X"B8",X"C1",X"92",X"28",X"48",X"66",X"89",X"A8",X"8C",X"BA",X"B1",X"48",X"49",X"BA",
		X"29",X"48",X"6B",X"6F",X"A0",X"A8",X"46",X"08",X"80",X"8C",X"1F",X"DB",X"2C",X"C9",X"1F",X"DB",
		X"88",X"C1",X"92",X"29",X"48",X"E6",X"89",X"3A",X"89",X"48",X"49",X"BA",X"C5",X"48",X"EE",X"F7",
		X"CF",X"12",X"29",X"48",X"46",X"08",X"F0",X"20",X"0A",X"12",X"29",X"48",X"46",X"89",X"F0",X"00",
		X"8A",X"76",X"08",X"53",X"B9",X"3A",X"C5",X"48",X"49",X"3E",X"80",X"2B",X"B6",X"29",X"A3",X"BD",
		X"80",X"57",X"69",X"21",X"D0",X"66",X"AE",X"88",X"B2",X"A8",X"E8",X"EE",X"29",X"27",X"CF",X"E6",
		X"50",X"8F",X"07",X"8F",X"07",X"C5",X"0A",X"30",X"D0",X"66",X"AF",X"43",X"0A",X"30",X"B6",X"28",
		X"83",X"36",X"28",X"23",X"8D",X"EA",X"46",X"AC",X"69",X"21",X"28",X"78",X"99",X"89",X"D8",X"36",
		X"88",X"09",X"77",X"29",X"CD",X"30",X"A1",X"5E",X"98",X"19",X"88",X"52",X"21",X"28",X"8A",X"E5",
		X"10",X"21",X"FE",X"98",X"99",X"88",X"DC",X"29",X"28",X"8A",X"65",X"B0",X"81",X"8C",X"DB",X"36",
		X"88",X"29",X"8C",X"55",X"B6",X"28",X"96",X"D7",X"B2",X"E5",X"48",X"C1",X"92",X"ED",X"48",X"76",
		X"38",X"FB",X"19",X"C9",X"81",X"88",X"E0",X"2E",X"20",X"0E",X"1C",X"1E",X"28",X"16",X"28",X"77",
		X"A3",X"7B",X"A3",X"0D",X"A0",X"D1",X"26",X"A8",X"05",X"28",X"54",X"C1",X"A1",X"5E",X"64",X"0E",
		X"09",X"CD",X"D9",X"AC",X"81",X"DC",X"C4",X"2E",X"0B",X"36",X"20",X"23",X"96",X"88",X"83",X"2D",
		X"6A",X"51",X"AC",X"C1",X"36",X"34",X"21",X"B7",X"88",X"3E",X"89",X"2B",X"B6",X"20",X"01",X"1D",
		X"80",X"57",X"69",X"BF",X"92",X"9B",X"E8",X"12",X"08",X"48",X"76",X"38",X"A0",X"8B",X"4E",X"89",
		X"A7",X"3A",X"88",X"48",X"92",X"30",X"40",X"BC",X"B2",X"30",X"40",X"17",X"B2",X"27",X"40",X"C5",
		X"AD",X"AF",X"21",X"38",X"E8",X"39",X"39",X"48",X"36",X"28",X"29",X"2B",X"28",X"C5",X"B0",X"CD",
		X"A9",X"25",X"A1",X"28",X"08",X"2A",X"9A",X"48",X"49",X"D5",X"ED",X"BE",X"08",X"75",X"4D",X"65",
		X"0B",X"DD",X"56",X"2D",X"2F",X"4F",X"2E",X"28",X"12",X"E7",X"E8",X"E6",X"29",X"00",X"2E",X"21",
		X"63",X"25",X"6B",X"7C",X"8D",X"29",X"73",X"25",X"01",X"65",X"92",X"3C",X"40",X"DF",X"A6",X"38",
		X"CD",X"79",X"6C",X"E9",X"09",X"56",X"CB",X"2F",X"2E",X"28",X"30",X"29",X"2C",X"DD",X"77",X"2F",
		X"5D",X"78",X"88",X"2B",X"D6",X"D5",X"F7",X"21",X"5D",X"3E",X"08",X"98",X"5D",X"3E",X"9A",X"28",
		X"CD",X"6D",X"17",X"CD",X"9B",X"32",X"F1",X"14",X"D6",X"20",X"10",X"99",X"12",X"20",X"E8",X"D6",
		X"0A",X"38",X"8F",X"BA",X"08",X"48",X"EE",X"29",X"A0",X"20",X"92",X"3B",X"40",X"76",X"19",X"3A",
		X"3B",X"48",X"21",X"28",X"EB",X"12",X"3B",X"48",X"29",X"A8",X"28",X"1E",X"08",X"0F",X"30",X"2A",
		X"4B",X"B6",X"01",X"9D",X"A0",X"DF",X"5D",X"61",X"49",X"9A",X"66",X"7F",X"D0",X"1A",X"A3",X"1B",
		X"0D",X"20",X"F6",X"C9",X"12",X"BE",X"E8",X"CD",X"6B",X"37",X"12",X"BE",X"E8",X"14",X"32",X"BE",
		X"40",X"C1",X"06",X"20",X"6B",X"41",X"8D",X"8E",X"89",X"4F",X"EE",X"D8",X"80",X"22",X"07",X"8F",
		X"0F",X"0F",X"EE",X"B8",X"77",X"23",X"71",X"03",X"23",X"23",X"50",X"E6",X"0F",X"EE",X"30",X"77",
		X"A3",X"79",X"49",X"38",X"40",X"A8",X"30",X"B8",X"A0",X"68",X"14",X"78",X"10",X"E8",X"14",X"F8",
		X"A2",X"F0",X"B0",X"68",X"20",X"B0",X"58",X"68",X"88",X"68",X"90",X"48",X"20",X"50",X"7C",X"58",
		X"28",X"58",X"30",X"28",X"B0",X"28",X"E0",X"28",X"38",X"E0",X"D8",X"E8",X"10",X"10",X"D8",X"88",
		X"B0",X"08",X"A8",X"A0",X"48",X"E8",X"88",X"F8",X"18",X"F0",X"84",X"10",X"48",X"40",X"18",X"08",
		X"F0",X"C8",X"10",X"A8",X"F8",X"7C",X"A0",X"78",X"30",X"10",X"F8",X"10",X"28",X"40",X"A0",X"50",
		X"90",X"50",X"A8",X"A0",X"18",X"C8",X"58",X"98",X"90",X"C8",X"A8",X"F0",X"88",X"D0",X"90",X"00",
		X"B8",X"48",X"C0",X"20",X"E8",X"B8",X"10",X"68",X"80",X"68",X"D0",X"08",X"F8",X"08",X"28",X"48",
		X"00",X"58",X"B0",X"D8",X"20",X"30",X"20",X"B0",X"58",X"58",X"58",X"D8",X"88",X"98",X"90",X"08",
		X"30",X"20",X"90",X"B0",X"B8",X"58",X"B8",X"B8",X"E8",X"B8",X"F0",X"08",X"D8",X"08",X"10",X"58",
		X"58",X"10",X"A8",X"08",X"38",X"D8",X"34",X"30",X"34",X"08",X"78",X"C8",X"50",X"80",X"A0",X"48",
		X"F0",X"50",X"00",X"A8",X"B8",X"F8",X"B8",X"D8",X"80",X"40",X"B0",X"30",X"C0",X"E0",X"F8",X"10",
		X"40",X"58",X"80",X"A8",X"10",X"98",X"98",X"A0",X"40",X"E0",X"B8",X"00",X"B8",X"10",X"10",X"60",
		X"E8",X"D8",X"38",X"A0",X"90",X"A8",X"18",X"78",X"E8",X"48",X"D8",X"18",X"D0",X"70",X"20",X"00",
		X"E8",X"48",X"80",X"B0",X"B0",X"C8",X"58",X"E8",X"00",X"08",X"58",X"00",X"80",X"48",X"78",X"40",
		X"A0",X"D8",X"F0",X"20",X"E0",X"30",X"20",X"A8",X"B0",X"70",X"08",X"08",X"E0",X"80",X"08",X"C8",
		X"30",X"40",X"80",X"C8",X"18",X"48",X"18",X"88",X"60",X"D8",X"48",X"D8",X"50",X"08",X"40",X"10",
		X"E8",X"98",X"F0",X"A0",X"D8",X"70",X"A0",X"60",X"48",X"E0",X"1C",X"10",X"1C",X"98",X"A0",X"98",
		X"E8",X"50",X"78",X"90",X"00",X"C8",X"98",X"D8",X"60",X"08",X"20",X"10",X"60",X"48",X"98",X"58",
		X"A8",X"28",X"E8",X"28",X"78",X"A0",X"48",X"60",X"28",X"70",X"F8",X"08",X"68",X"80",X"00",X"90",
		X"20",X"50",X"68",X"30",X"40",X"60",X"18",X"78",X"88",X"78",X"92",X"F8",X"68",X"80",X"92",X"C8",
		X"28",X"C0",X"E8",X"30",X"30",X"B8",X"78",X"70",X"58",X"08",X"80",X"88",X"E8",X"40",X"18",X"40",
		X"60",X"D8",X"60",X"E8",X"38",X"78",X"92",X"08",X"68",X"08",X"88",X"98",X"92",X"28",X"18",X"28",
		X"E8",X"28",X"A0",X"28",X"A0",X"B8",X"00",X"60",X"58",X"18",X"E8",X"18",X"10",X"88",X"40",X"D8",
		X"20",X"C0",X"A8",X"38",X"20",X"B8",X"70",X"B0",X"90",X"E8",X"68",X"F0",X"98",X"10",X"18",X"98",
		X"78",X"40",X"B0",X"24",X"58",X"A8",X"A0",X"B8",X"E8",X"08",X"28",X"08",X"78",X"40",X"E8",X"50",
		X"80",X"C4",X"78",X"B0",X"18",X"30",X"50",X"78",X"78",X"B0",X"90",X"80",X"78",X"40",X"18",X"40",
		X"B0",X"C0",X"F8",X"28",X"E8",X"60",X"E8",X"E8",X"B8",X"E8",X"90",X"0C",X"D8",X"80",X"90",X"98",
		X"10",X"48",X"40",X"A8",X"48",X"A8",X"A8",X"70",X"B0",X"0C",X"68",X"0C",X"A8",X"98",X"B0",X"D8",
		X"48",X"D8",X"00",X"28",X"B8",X"28",X"00",X"B0",X"B0",X"60",X"28",X"E8",X"78",X"90",X"78",X"58",
		X"90",X"50",X"20",X"28",X"78",X"A8",X"88",X"68",X"78",X"E8",X"30",X"08",X"A0",X"88",X"30",X"40",
		X"58",X"50",X"80",X"B0",X"98",X"70",X"D8",X"08",X"D8",X"80",X"D8",X"70",X"20",X"08",X"20",X"80",
		X"A0",X"08",X"18",X"68",X"18",X"68",X"70",X"68",X"90",X"EC",X"58",X"8C",X"58",X"48",X"18",X"48",
		X"B0",X"40",X"78",X"38",X"30",X"B0",X"F8",X"78",X"30",X"E8",X"48",X"F0",X"F8",X"90",X"F8",X"58",
		X"B0",X"D0",X"50",X"B0",X"10",X"B0",X"50",X"08",X"68",X"08",X"70",X"08",X"A0",X"48",X"10",X"C8",
		X"70",X"F0",X"30",X"08",X"60",X"08",X"10",X"4C",X"B0",X"DC",X"80",X"04",X"38",X"04",X"10",X"A4",
		X"88",X"4C",X"B8",X"A8",X"30",X"60",X"00",X"E8",X"68",X"08",X"18",X"88",X"68",X"90",X"00",X"C8",
		X"38",X"08",X"E0",X"28",X"3C",X"BC",X"FC",X"E8",X"3C",X"F8",X"0C",X"10",X"0C",X"20",X"3C",X"C4",
		X"7C",X"C0",X"34",X"2E",X"6B",X"7A",X"6D",X"6C",X"61",X"7C",X"2F",X"6B",X"7A",X"6D",X"6C",X"61",
		X"FC",X"5B",X"AB",X"60",X"C1",X"62",X"AB",X"63",X"C1",X"62",X"AB",X"64",X"C5",X"66",X"2B",X"A9",
		X"28",X"7B",X"6D",X"6F",X"69",X"28",X"B9",X"B1",X"B0",X"BC",X"3B",X"B9",X"28",X"78",X"64",X"69",
		X"79",X"4D",X"FA",X"08",X"FB",X"5C",X"E9",X"5A",X"FC",X"08",X"6F",X"CE",X"6C",X"D9",X"BB",X"39",
		X"28",X"67",X"7A",X"28",X"BA",X"28",X"78",X"64",X"69",X"71",X"6D",X"7A",X"28",X"7B",X"7C",X"69",
		X"FA",X"5C",X"29",X"4F",X"E9",X"CD",X"ED",X"09",X"6F",X"5E",X"ED",X"5A",X"2B",X"C9",X"6E",X"5B",
		X"6D",X"7A",X"7C",X"29",X"6B",X"67",X"61",X"66",X"22",X"7C",X"61",X"65",X"6D",X"28",X"6A",X"67",
		X"6E",X"5D",X"FB",X"0B",X"AC",X"0D",X"AE",X"8E",X"F8",X"CC",X"E9",X"D9",X"ED",X"5A",X"A9",X"39",
		X"29",X"7B",X"7C",X"69",X"7A",X"7C",X"26",X"78",X"64",X"69",X"71",X"6D",X"7A",X"29",X"BA",X"29",
		X"FB",X"5C",X"E9",X"5A",X"FC",X"0C",X"FC",X"C9",X"6D",X"4D",X"2B",X"4A",X"6F",X"CE",X"FD",X"5B",
		X"28",X"7A",X"67",X"7D",X"66",X"6C",X"28",X"28",X"C0",X"28",X"28",X"28",X"28",X"28",X"28",X"D7",
		X"A8",X"B8",X"37",X"40",X"CF",X"F7",X"A8",X"F7",X"A8",X"B8",X"37",X"40",X"CF",X"F7",X"A8",X"35",
		X"83",X"83",X"8C",X"37",X"3E",X"3C",X"28",X"48",X"D7",X"28",X"28",X"28",X"28",X"28",X"28",X"D7",
		X"E0",X"2C",X"AD",X"AE",X"2D",X"A5",X"08",X"BF",X"93",X"E4",X"CA",X"2D",X"F7",X"83",X"08",X"40",
		X"17",X"D8",X"1C",X"AD",X"9B",X"03",X"28",X"13",X"5B",X"8C",X"85",X"9E",X"BC",X"35",X"28",X"D7",
		X"08",X"08",X"08",X"08",X"08",X"0F",X"08",X"F7",X"08",X"08",X"08",X"08",X"08",X"F7",X"08",X"06",
		X"E7",X"D7",X"28",X"28",X"28",X"28",X"28",X"A3",X"03",X"AA",X"22",X"CF",X"D7",X"B7",X"28",X"D0",
		X"AB",X"2B",X"AB",X"AF",X"0E",X"92",X"08",X"08",X"89",X"8A",X"19",X"9A",X"08",X"0A",X"08",X"0F",
		X"D7",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"3A",X"33",X"05",X"BE",X"3B",X"34",X"28",X"D7",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"F7",X"08",X"08",X"08",X"08",X"08",X"08",X"DA",X"F5",
		X"F4",X"C3",X"A0",X"10",X"28",X"2D",X"28",X"DD",X"86",X"84",X"C4",X"8D",X"A3",X"AC",X"28",X"86",
		X"A4",X"A5",X"AD",X"2C",X"0C",X"75",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"28",X"28",X"28",X"28",X"28",X"28",X"5A",X"28",X"3A",X"33",X"05",X"BE",X"3B",X"34",X"28",X"D7",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"F7",X"08",X"08",X"08",X"08",X"08",X"08",X"DA",X"F5",
		X"F4",X"C3",X"A0",X"10",X"28",X"2D",X"28",X"16",X"85",X"8D",X"BD",X"8C",X"30",X"B7",X"28",X"85",
		X"96",X"25",X"AD",X"45",X"7E",X"9B",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"28",X"28",X"28",X"28",X"28",X"28",X"5A",X"28",X"3A",X"33",X"05",X"BE",X"3B",X"34",X"28",X"D7",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"F7",X"08",X"08",X"08",X"08",X"08",X"08",X"DA",X"F5",
		X"F4",X"C3",X"A0",X"10",X"28",X"2D",X"28",X"12",X"A3",X"73",X"25",X"15",X"EE",X"3B",X"28",X"DC",
		X"05",X"23",X"A5",X"9A",X"7B",X"0F",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"08",
		X"28",X"28",X"28",X"28",X"28",X"28",X"72",X"28",X"3A",X"33",X"A5",X"BE",X"3B",X"34",X"28",X"D7",
		X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"F7",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"7A",X"F5",
		X"DC",X"C3",X"88",X"10",X"28",X"2D",X"28",X"28",X"28",X"28",X"28",X"28",X"33",X"3A",X"28",X"AB",
		X"16",X"36",X"D8",X"E0",X"88",X"48",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"08",
		X"28",X"28",X"28",X"28",X"28",X"28",X"72",X"28",X"3A",X"33",X"A5",X"BE",X"3B",X"34",X"28",X"D7",
		X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"F7",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"7A",X"F5",
		X"DC",X"C3",X"88",X"10",X"28",X"2D",X"28",X"B7",X"2F",X"D8",X"48",X"08",X"68",X"D7",X"28",X"2F",
		X"17",X"36",X"D8",X"E0",X"88",X"F7",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"08",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"33",X"C0",X"10",X"B7",X"A6",X"D7",X"C7",X"28",X"D7",
		X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"F7",X"A8",X"08",X"A8",X"08",X"A8",X"08",X"A8",X"65",
		X"B5",X"BB",X"A3",X"C0",X"AC",X"3B",X"28",X"2F",X"DF",X"CD",X"A4",X"BB",X"B3",X"34",X"28",X"CD",
		X"57",X"AB",X"40",X"08",X"A8",X"08",X"58",X"E0",X"A4",X"AD",X"B6",X"60",X"05",X"08",X"A8",X"F7",
		X"C0",X"AC",X"10",X"A7",X"AD",X"85",X"28",X"A3",X"A3",X"AA",X"AA",X"CF",X"D7",X"B7",X"28",X"D0",
		X"23",X"2B",X"23",X"AF",X"AE",X"92",X"A8",X"75",X"06",X"A4",X"44",X"25",X"83",X"2C",X"A8",X"A6",
		X"84",X"85",X"A5",X"AC",X"2C",X"DD",X"28",X"16",X"85",X"8D",X"1D",X"8C",X"B8",X"B7",X"28",X"85",
		X"96",X"25",X"AD",X"45",X"7E",X"9B",X"08",X"92",X"23",X"DB",X"2D",X"95",X"46",X"1B",X"08",X"74",
		X"85",X"8B",X"25",X"32",X"5B",X"2F",X"28",X"28",X"28",X"28",X"28",X"28",X"1B",X"3A",X"28",X"AB",
		X"B6",X"36",X"50",X"E0",X"00",X"48",X"08",X"36",X"A5",X"24",X"A5",X"67",X"F7",X"BF",X"08",X"F0",
		X"B6",X"AB",X"85",X"A7",X"2E",X"12",X"28",X"AD",X"83",X"89",X"1C",X"8A",X"99",X"AC",X"28",X"83",
		X"21",X"A5",X"2E",X"9C",X"0D",X"AD",X"08",X"9D",X"2D",X"9C",X"9B",X"1A",X"28",X"0F",X"08",X"A5",
		X"1F",X"BE",X"30",X"A0",X"3C",X"2F",X"28",X"2C",X"28",X"34",X"3D",X"34",X"25",X"3B",X"28",X"97",
		X"D5",X"08",X"1D",X"AD",X"9C",X"E7",X"08",X"0B",X"0C",X"0D",X"9E",X"0A",X"08",X"08",X"08",X"A5",
		X"F7",X"CF",X"F8",X"C0",X"A8",X"68",X"09",X"6F",X"69",X"65",X"6D",X"28",X"7C",X"61",X"4D",X"6D",
		X"0C",X"CD",X"C9",X"CE",X"DC",X"0C",X"5B",X"4D",X"4B",X"DC",X"3A",X"38",X"38",X"38",X"38",X"08",
		X"78",X"7C",X"7B",X"74",X"31",X"B8",X"30",X"B8",X"30",X"28",X"78",X"7C",X"7B",X"74",X"28",X"BD",
		X"38",X"38",X"38",X"08",X"58",X"5C",X"5B",X"DC",X"08",X"3B",X"38",X"38",X"38",X"08",X"58",X"5C",
		X"7B",X"74",X"28",X"B9",X"30",X"B8",X"30",X"28",X"78",X"7C",X"7B",X"74",X"28",X"66",X"4F",X"28",
		X"4A",X"CF",X"CE",X"5D",X"5B",X"08",X"82",X"1B",X"14",X"1B",X"96",X"1B",X"A0",X"1B",X"32",X"1B",
		X"94",X"3B",X"EF",X"4F",X"7F",X"BF",X"37",X"AF",X"37",X"A7",X"A7",X"8F",X"EF",X"A7",X"27",X"BF",
		X"47",X"47",X"47",X"47",X"9F",X"47",X"9F",X"9F",X"47",X"47",X"5F",X"47",X"47",X"27",X"DF",X"47",
		X"EF",X"4F",X"1F",X"FF",X"1F",X"4F",X"28",X"A7",X"07",X"97",X"1E",X"AE",X"1E",X"AC",X"28",X"A5",
		X"A4",X"9A",X"25",X"2C",X"3A",X"2C",X"A8",X"A5",X"05",X"F7",X"1B",X"24",X"84",X"F7",X"A8",X"67",
		X"CF",X"D7",X"0E",X"0E",X"0E",X"D7",X"28",X"BE",X"A5",X"97",X"A5",X"33",X"AC",X"9F",X"28",X"85",
		X"3B",X"76",X"05",X"08",X"3B",X"23",X"A8",X"38",X"90",X"3D",X"B3",X"98",X"A2",X"2A",X"A8",X"AE",
		X"2C",X"36",X"A6",X"2C",X"36",X"2C",X"28",X"DE",X"C5",X"D6",X"CC",X"8C",X"13",X"DC",X"28",X"BF",
		X"B7",X"2D",X"26",X"9B",X"25",X"9B",X"A8",X"B7",X"80",X"F0",X"90",X"20",X"00",X"BF",X"A8",X"65",
		X"CD",X"D5",X"0C",X"0C",X"0C",X"D5",X"76",X"3C",X"86",X"3C",X"D6",X"3C",X"66",X"3D",X"28",X"28",
		X"38",X"34",X"D1",X"F7",X"38",X"34",X"C2",X"F7",X"38",X"34",X"DB",X"F7",X"38",X"34",X"F4",X"0A",
		X"C0",X"9C",X"0B",X"2A",X"C0",X"9C",X"1A",X"2A",X"C0",X"9C",X"89",X"2A",X"C0",X"9C",X"30",X"D7",
		X"38",X"35",X"29",X"F7",X"38",X"35",X"52",X"F6",X"38",X"35",X"43",X"F6",X"38",X"35",X"7C",X"0B",
		X"C0",X"9B",X"E3",X"2B",X"C0",X"9B",X"F2",X"2B",X"C0",X"9B",X"01",X"2B",X"C0",X"9B",X"B8",X"D6",
		X"38",X"34",X"A1",X"F6",X"38",X"34",X"BA",X"F6",X"38",X"34",X"AB",X"F6",X"38",X"34",X"A8",X"08",
		X"30",X"9C",X"D9",X"D7",X"3C",X"9C",X"CA",X"D7",X"38",X"9C",X"5B",X"D7",X"24",X"9C",X"FC",X"2A",
		X"40",X"34",X"8B",X"0A",X"44",X"34",X"9A",X"0A",X"D0",X"34",X"81",X"0A",X"D4",X"34",X"38",X"F7",
		X"30",X"9D",X"21",X"D7",X"3C",X"9D",X"D2",X"D6",X"38",X"9D",X"C3",X"D6",X"24",X"9D",X"74",X"2B",
		X"40",X"33",X"63",X"0B",X"44",X"33",X"72",X"0B",X"D0",X"33",X"09",X"0B",X"D4",X"33",X"B0",X"F6",
		X"30",X"9C",X"A9",X"D6",X"3C",X"9C",X"3A",X"D6",X"38",X"9C",X"2B",X"D6",X"24",X"9C",X"28",X"28",
		X"98",X"34",X"71",X"F7",X"98",X"B0",X"62",X"F7",X"98",X"B4",X"53",X"F7",X"98",X"40",X"7C",X"0A",
		X"C0",X"9C",X"AB",X"2A",X"C0",X"90",X"BA",X"2A",X"C0",X"94",X"A1",X"2A",X"C0",X"48",X"18",X"D7",
		X"98",X"34",X"89",X"F7",X"98",X"B0",X"F2",X"F6",X"98",X"B4",X"E3",X"F6",X"98",X"40",X"DC",X"0B",
		X"C0",X"9C",X"43",X"2B",X"C0",X"90",X"52",X"2B",X"C0",X"94",X"89",X"2B",X"C0",X"48",X"30",X"D6",
		X"98",X"34",X"29",X"F6",X"98",X"B0",X"1A",X"F6",X"98",X"B4",X"0B",X"F6",X"98",X"40",X"08",X"08",
		X"3A",X"9C",X"F1",X"D7",X"3A",X"9C",X"E2",X"D7",X"3A",X"9C",X"FB",X"D7",X"3A",X"9C",X"28",X"2A",
		X"E6",X"34",X"8F",X"0A",X"E6",X"34",X"9E",X"0A",X"E6",X"34",X"AD",X"0A",X"E6",X"34",X"98",X"F7",
		X"3A",X"9D",X"09",X"D7",X"3A",X"9D",X"D2",X"D6",X"3A",X"9D",X"C3",X"D6",X"3A",X"9D",X"C0",X"2A",
		X"E6",X"33",X"77",X"0A",X"E6",X"33",X"0E",X"0B",X"E6",X"33",X"1D",X"0B",X"E6",X"33",X"38",X"F6",
		X"0B",X"9C",X"21",X"D6",X"38",X"9C",X"3A",X"D6",X"3D",X"9C",X"2B",X"D6",X"1A",X"9C",X"B6",X"3D",
		X"36",X"1D",X"36",X"1D",X"36",X"1D",X"37",X"1D",X"41",X"1D",X"C6",X"1D",X"D0",X"1D",X"65",X"1D",
		X"C7",X"3D",X"F6",X"3D",X"28",X"3E",X"D7",X"29",X"38",X"B8",X"38",X"D6",X"E0",X"60",X"29",X"A8",
		X"F7",X"0A",X"F7",X"08",X"48",X"0A",X"28",X"78",X"F4",X"60",X"14",X"0A",X"38",X"F7",X"0C",X"09",
		X"20",X"08",X"D7",X"28",X"B0",X"58",X"B8",X"D7",X"2A",X"D7",X"28",X"68",X"2C",X"F8",X"A8",X"D0",
		X"10",X"B0",X"0A",X"70",X"F7",X"00",X"F0",X"20",X"20",X"18",X"38",X"40",X"F7",X"08",X"F7",X"0A",
		X"F8",X"58",X"18",X"2A",X"10",X"D7",X"2C",X"B8",X"70",X"38",X"D6",X"58",X"A8",X"2A",X"20",X"D7",
		X"AC",X"F7",X"A8",X"48",X"A9",X"78",X"57",X"1D",X"34",X"08",X"B2",X"3D",X"B0",X"08",X"F8",X"5C",
		X"7B",X"74",X"B6",X"28",X"28",X"B8",X"B8",X"B8",X"28",X"78",X"7C",X"7B",X"74",X"25",X"78",X"6D",
		X"FA",X"4E",X"ED",X"4B",X"FC",X"08",X"EA",X"CF",X"6E",X"5D",X"FB",X"8A",X"B1",X"38",X"B0",X"38",
		X"B8",X"28",X"78",X"7C",X"7B",X"74",X"2C",X"7A",X"6C",X"74",X"29",X"39",X"6F",X"69",X"7C",X"60",
		X"ED",X"5A",X"A8",X"5D",X"F8",X"08",X"F8",X"C9",X"6F",X"58",X"69",X"CF",X"E8",X"19",X"EC",X"4D",
		X"6E",X"6D",X"69",X"7C",X"28",X"66",X"71",X"69",X"66",X"66",X"71",X"69",X"66",X"68",X"28",X"39",
		X"FC",X"49",X"6B",X"4D",X"A8",X"58",X"69",X"CF",X"F8",X"C9",X"6F",X"08",X"68",X"CF",X"6D",X"4D",
		X"68",X"28",X"A8",X"28",X"38",X"28",X"2D",X"28",X"2B",X"28",X"29",X"28",X"28",X"A3",X"84",X"8D",
		X"E8",X"A5",X"A8",X"A5",X"81",X"9C",X"BD",X"0B",X"A8",X"08",X"A5",X"58",X"F5",X"D5",X"92",X"6E",
		X"48",X"87",X"00",X"2B",X"F1",X"53",X"C9",X"32",X"EF",X"48",X"A7",X"CA",X"E0",X"3F",X"ED",X"DD",
		X"ED",X"A1",X"A8",X"41",X"31",X"08",X"D8",X"AE",X"A8",X"36",X"3F",X"2E",X"28",X"4B",X"D6",X"CA",
		X"93",X"3E",X"C3",X"29",X"09",X"43",X"0C",X"29",X"EB",X"4B",X"3E",X"A3",X"C5",X"90",X"C3",X"2E",
		X"28",X"29",X"CB",X"35",X"6A",X"A3",X"BE",X"22",X"61",X"40",X"A2",X"F4",X"47",X"A6",X"CF",X"BE",
		X"50",X"32",X"4C",X"48",X"E6",X"2F",X"CB",X"2F",X"CB",X"2F",X"5F",X"C6",X"29",X"4A",X"CC",X"3E",
		X"4B",X"8B",X"A4",X"BC",X"C3",X"A9",X"E8",X"08",X"CD",X"90",X"92",X"3F",X"C8",X"B2",X"B6",X"D4",
		X"32",X"79",X"52",X"22",X"BB",X"48",X"22",X"6E",X"54",X"32",X"E5",X"48",X"32",X"61",X"52",X"32",
		X"D0",X"40",X"AF",X"32",X"6D",X"40",X"4A",X"8E",X"1F",X"D6",X"18",X"CB",X"18",X"1F",X"EE",X"E7",
		X"32",X"ED",X"E8",X"4D",X"6B",X"24",X"21",X"4C",X"E8",X"B4",X"21",X"E0",X"E8",X"B4",X"12",X"48",
		X"40",X"CE",X"09",X"56",X"BC",X"30",X"3D",X"32",X"18",X"40",X"6E",X"09",X"A7",X"56",X"68",X"30",
		X"0A",X"92",X"39",X"48",X"EE",X"29",X"27",X"B2",X"39",X"48",X"BF",X"B2",X"38",X"48",X"12",X"22",
		X"40",X"CE",X"09",X"A7",X"DE",X"68",X"90",X"18",X"92",X"8B",X"40",X"CE",X"09",X"A7",X"DE",X"68",
		X"10",X"2A",X"16",X"E8",X"32",X"23",X"E8",X"3F",X"32",X"22",X"E8",X"3F",X"32",X"48",X"E8",X"4D",
		X"26",X"98",X"E9",X"D9",X"69",X"D1",X"DB",X"49",X"6D",X"DD",X"ED",X"A1",X"6F",X"40",X"B5",X"76",
		X"21",X"28",X"F8",X"2C",X"67",X"3F",X"6F",X"F7",X"23",X"30",X"D4",X"E9",X"F9",X"69",X"F1",X"DB",
		X"49",X"C5",X"A1",X"F7",X"F7",X"25",X"A0",X"F5",X"A5",X"A0",X"F2",X"C1",X"49",X"EF",X"92",X"08",
		X"E8",X"EE",X"29",X"68",X"50",X"EE",X"0F",X"27",X"4F",X"26",X"28",X"A1",X"55",X"32",X"09",X"46",
		X"A3",X"EE",X"4D",X"8D",X"98",X"71",X"2E",X"A7",X"F7",X"23",X"D0",X"0E",X"A7",X"F7",X"83",X"36",
		X"28",X"0E",X"27",X"DE",X"99",X"B0",X"29",X"F7",X"E6",X"27",X"2F",X"27",X"2F",X"27",X"5F",X"A3",
		X"D6",X"C6",X"70",X"2F",X"07",X"2F",X"07",X"93",X"57",X"A1",X"ED",X"9A",X"92",X"0C",X"40",X"C6",
		X"30",X"07",X"0F",X"47",X"2E",X"28",X"09",X"92",X"0E",X"48",X"4F",X"01",X"56",X"9B",X"00",X"2A",
		X"B0",X"28",X"92",X"8E",X"40",X"34",X"B2",X"8E",X"40",X"36",X"09",X"B2",X"8D",X"40",X"A1",X"0A",
		X"E8",X"92",X"29",X"48",X"E6",X"29",X"00",X"29",X"04",X"B4",X"CD",X"E2",X"0B",X"96",X"B8",X"4D",
		X"B5",X"4D",X"92",X"09",X"C8",X"C6",X"A9",X"CA",X"78",X"98",X"6B",X"9A",X"38",X"A1",X"D9",X"40",
		X"12",X"29",X"48",X"C6",X"29",X"48",X"21",X"5C",X"48",X"49",X"21",X"26",X"C0",X"B9",X"47",X"48",
		X"4D",X"6F",X"38",X"32",X"A9",X"40",X"EE",X"0A",X"68",X"22",X"DD",X"40",X"75",X"7C",X"82",X"C7",
		X"48",X"75",X"44",X"E7",X"B7",X"45",X"7A",X"58",X"20",X"22",X"12",X"5F",X"48",X"7F",X"12",X"59",
		X"C8",X"13",X"48",X"58",X"31",X"55",X"C8",X"A1",X"4F",X"40",X"21",X"0B",X"A8",X"45",X"B8",X"B9",
		X"47",X"48",X"21",X"A2",X"C0",X"CB",X"EF",X"30",X"21",X"A2",X"C0",X"B9",X"5A",X"48",X"EB",X"EF",
		X"38",X"A1",X"22",X"E0",X"31",X"55",X"C8",X"AE",X"AB",X"2E",X"A8",X"C5",X"4D",X"F2",X"39",X"B6",
		X"B8",X"24",X"36",X"20",X"E1",X"71",X"A7",X"C8",X"FD",X"B9",X"71",X"32",X"C3",X"4D",X"5E",X"22",
		X"79",X"49",X"6E",X"38",X"05",X"2E",X"A9",X"4A",X"9F",X"98",X"DE",X"38",X"A0",X"89",X"06",X"08",
		X"36",X"A8",X"23",X"B6",X"20",X"38",X"2C",X"F7",X"23",X"B6",X"20",X"A3",X"C9",X"8A",X"27",X"FF",
		X"D3",X"4E",X"A8",X"A7",X"57",X"49",X"92",X"D1",X"C8",X"87",X"68",X"9F",X"5B",X"88",X"67",X"32",
		X"79",X"48",X"4F",X"4B",X"58",X"20",X"32",X"4B",X"59",X"20",X"30",X"4B",X"99",X"A1",X"78",X"48",
		X"D6",X"56",X"29",X"30",X"AD",X"36",X"29",X"CB",X"4D",X"98",X"6E",X"09",X"A7",X"F7",X"6B",X"53",
		X"30",X"4B",X"D9",X"A1",X"7A",X"48",X"39",X"72",X"48",X"4B",X"68",X"20",X"24",X"4B",X"69",X"20",
		X"2A",X"4B",X"29",X"4D",X"A1",X"99",X"6B",X"E3",X"38",X"4B",X"69",X"76",X"6D",X"EF",X"92",X"5D",
		X"48",X"10",X"00",X"2E",X"21",X"7D",X"48",X"B9",X"74",X"48",X"E9",X"4B",X"48",X"20",X"24",X"4B",
		X"41",X"20",X"8A",X"4B",X"09",X"4D",X"29",X"99",X"6B",X"8D",X"99",X"4B",X"49",X"71",X"B2",X"59",
		X"E8",X"A1",X"5A",X"48",X"0E",X"29",X"CD",X"9C",X"19",X"A1",X"5C",X"48",X"0E",X"2A",X"EB",X"9C",
		X"99",X"CD",X"ED",X"DD",X"D6",X"AF",X"DE",X"1C",X"B0",X"4E",X"47",X"AE",X"08",X"43",X"33",X"A1",
		X"3A",X"32",X"09",X"D6",X"23",X"E6",X"47",X"3F",X"C1",X"94",X"14",X"94",X"14",X"94",X"14",X"4D",
		X"17",X"99",X"10",X"CC",X"12",X"56",X"09",X"B0",X"99",X"38",X"1B",X"3A",X"DE",X"0A",X"B0",X"1A",
		X"18",X"24",X"1A",X"DE",X"2B",X"B0",X"0B",X"10",X"2D",X"12",X"D6",X"29",X"30",X"24",X"14",X"32",
		X"10",X"AE",X"3F",X"BA",X"94",X"4D",X"17",X"99",X"10",X"2E",X"3F",X"BA",X"94",X"34",X"10",X"74",
		X"FE",X"3C",X"4F",X"26",X"28",X"CB",X"3B",X"33",X"21",X"AE",X"1A",X"01",X"56",X"A3",X"66",X"C7",
		X"12",X"34",X"47",X"16",X"90",X"09",X"3F",X"BA",X"26",X"08",X"01",X"76",X"AF",X"CC",X"17",X"99",
		X"F9",X"E9",X"E9",X"12",X"14",X"32",X"C9",X"77",X"12",X"78",X"E8",X"2A",X"27",X"77",X"D6",X"21",
		X"90",X"0D",X"96",X"89",X"6B",X"30",X"99",X"4D",X"AA",X"4D",X"96",X"87",X"4D",X"BD",X"4D",X"72",
		X"32",X"78",X"E8",X"49",X"56",X"AF",X"C8",X"4B",X"57",X"6A",X"FB",X"31",X"23",X"D6",X"A7",X"6A",
		X"C0",X"99",X"4D",X"D5",X"99",X"B6",X"0E",X"49",X"B5",X"C8",X"4D",X"E1",X"99",X"B6",X"0E",X"23",
		X"CB",X"DE",X"C9",X"A3",X"35",X"68",X"03",X"D6",X"E6",X"F7",X"15",X"F7",X"C9",X"ED",X"12",X"ED",
		X"40",X"91",X"B2",X"6D",X"40",X"DB",X"99",X"C1",X"49",X"C5",X"6D",X"71",X"87",X"6F",X"92",X"6D",
		X"E8",X"A9",X"32",X"ED",X"E8",X"7B",X"19",X"69",X"E1",X"49",X"1A",X"4B",X"17",X"4B",X"17",X"4B",
		X"97",X"4B",X"97",X"4D",X"8A",X"98",X"12",X"C6",X"2F",X"4D",X"8A",X"98",X"25",X"48",X"33",X"CB",
		X"D2",X"31",X"B6",X"31",X"B5",X"31",X"B4",X"31",X"B3",X"31",X"B2",X"31",X"B1",X"31",X"6C",X"31",
		X"6B",X"99",X"FA",X"99",X"79",X"99",X"B4",X"9A",X"33",X"9A",X"E8",X"9A",X"EE",X"9A",X"6B",X"9A",
		X"66",X"32",X"7C",X"32",X"2E",X"28",X"29",X"28",X"29",X"29",X"29",X"2C",X"28",X"29",X"28",X"2A",
		X"AD",X"09",X"A9",X"09",X"A9",X"0A",X"AC",X"09",X"A9",X"09",X"AA",X"0A",X"A9",X"0A",X"AD",X"0A",
		X"2A",X"2A",X"2A",X"2B",X"2C",X"2A",X"2A",X"2A",X"2B",X"2F",X"28",X"28",X"28",X"28",X"28",X"28",
		X"B0",X"8F",X"2E",X"8D",X"2C",X"8B",X"2A",X"89",X"2A",X"8B",X"2C",X"8D",X"2E",X"0B",X"28",X"1E",
		X"D7",X"2B",X"38",X"A8",X"D7",X"2C",X"3A",X"AC",X"D7",X"2C",X"3C",X"A0",X"D7",X"28",X"28",X"29",
		X"A8",X"0A",X"A8",X"0B",X"A8",X"0D",X"A8",X"18",X"A8",X"28",X"A8",X"38",X"A8",X"48",X"A8",X"58",
		X"28",X"08",X"28",X"28",X"29",X"28",X"2A",X"28",X"2B",X"28",X"2D",X"4D",X"9B",X"32",X"DD",X"7E",
		X"A9",X"5D",X"76",X"0A",X"CB",X"A9",X"AC",X"08",X"01",X"76",X"A3",X"E6",X"C7",X"A9",X"2F",X"08",
		X"C5",X"90",X"C9",X"A1",X"28",X"4F",X"DD",X"76",X"2D",X"4B",X"67",X"20",X"29",X"A4",X"E6",X"27",
		X"27",X"AF",X"27",X"AF",X"C7",X"49",X"92",X"4C",X"C8",X"87",X"68",X"32",X"A8",X"40",X"EE",X"09",
		X"CA",X"68",X"33",X"32",X"4C",X"48",X"E6",X"27",X"EA",X"68",X"33",X"A1",X"05",X"B8",X"12",X"E7",
		X"C8",X"87",X"80",X"18",X"DE",X"09",X"80",X"99",X"92",X"4D",X"C8",X"87",X"A0",X"5A",X"A1",X"30",
		X"B8",X"CB",X"29",X"33",X"21",X"22",X"B8",X"32",X"E6",X"48",X"E6",X"29",X"20",X"2B",X"21",X"6A",
		X"38",X"32",X"B8",X"40",X"47",X"AE",X"08",X"29",X"DE",X"58",X"B0",X"3C",X"D6",X"B2",X"B9",X"40",
		X"51",X"94",X"32",X"B0",X"E8",X"92",X"47",X"48",X"D6",X"29",X"20",X"AC",X"12",X"B0",X"E8",X"A1",
		X"BB",X"1E",X"31",X"50",X"E3",X"56",X"09",X"20",X"1C",X"A1",X"CD",X"1E",X"31",X"50",X"E3",X"56",
		X"0D",X"80",X"0A",X"DE",X"3C",X"A0",X"09",X"A1",X"5F",X"3E",X"39",X"58",X"C3",X"4D",X"EC",X"22",
		X"3F",X"5B",X"88",X"4B",X"77",X"A0",X"0D",X"36",X"09",X"B2",X"D1",X"40",X"92",X"AC",X"40",X"87",
		X"EA",X"4A",X"1D",X"92",X"47",X"48",X"D6",X"2A",X"CA",X"4A",X"1D",X"92",X"EC",X"48",X"E6",X"24",
		X"07",X"2F",X"47",X"AE",X"08",X"A1",X"0E",X"38",X"01",X"76",X"B2",X"3F",X"40",X"32",X"40",X"40",
		X"E6",X"29",X"20",X"A8",X"12",X"BE",X"E8",X"AF",X"00",X"32",X"D6",X"2F",X"20",X"27",X"12",X"3B",
		X"40",X"56",X"F7",X"20",X"0E",X"32",X"A8",X"40",X"AF",X"A0",X"89",X"36",X"0F",X"35",X"B2",X"3E",
		X"E8",X"4D",X"6B",X"37",X"29",X"28",X"28",X"92",X"00",X"48",X"A7",X"6A",X"BB",X"36",X"12",X"28",
		X"44",X"C6",X"0C",X"CA",X"DF",X"9C",X"92",X"08",X"46",X"C6",X"28",X"CA",X"DF",X"9C",X"92",X"49",
		X"E8",X"DE",X"2E",X"B0",X"2B",X"AF",X"20",X"67",X"CD",X"2C",X"0C",X"DE",X"D7",X"80",X"3B",X"DE",
		X"F3",X"20",X"8F",X"56",X"F5",X"20",X"8B",X"56",X"F1",X"20",X"0F",X"9F",X"B2",X"4E",X"40",X"CB",
		X"DD",X"33",X"12",X"6E",X"E8",X"94",X"32",X"6E",X"E8",X"DE",X"D7",X"80",X"32",X"92",X"0B",X"48",
		X"AF",X"A0",X"1D",X"32",X"0C",X"40",X"EE",X"48",X"4A",X"DF",X"9C",X"32",X"8A",X"40",X"DE",X"48",
		X"DA",X"77",X"1C",X"26",X"0F",X"6B",X"2B",X"34",X"2E",X"2F",X"12",X"22",X"E8",X"DE",X"20",X"90",
		X"AA",X"AE",X"AB",X"80",X"6A",X"DF",X"3C",X"32",X"C8",X"40",X"EE",X"0B",X"6A",X"DF",X"3C",X"A1",
		X"50",X"B8",X"12",X"69",X"48",X"56",X"2E",X"DA",X"B6",X"34",X"2F",X"6F",X"2E",X"28",X"2F",X"89",
		X"47",X"29",X"55",X"FC",X"82",X"BF",X"C8",X"A9",X"35",X"08",X"4D",X"A7",X"3D",X"4D",X"07",X"9D",
		X"CD",X"87",X"35",X"32",X"69",X"48",X"14",X"B2",X"69",X"48",X"D6",X"2E",X"20",X"A9",X"02",X"B7",
		X"C8",X"6D",X"64",X"4D",X"7E",X"2F",X"21",X"0B",X"A8",X"97",X"CD",X"EA",X"A2",X"0F",X"CE",X"C6",
		X"D0",X"CE",X"22",X"B2",X"21",X"4E",X"16",X"98",X"32",X"28",X"4E",X"9F",X"32",X"2E",X"4E",X"32",
		X"CC",X"40",X"EE",X"0F",X"A0",X"C9",X"92",X"08",X"CC",X"C6",X"AC",X"A0",X"EA",X"32",X"B1",X"40",
		X"A7",X"20",X"33",X"56",X"39",X"30",X"21",X"9F",X"32",X"B9",X"48",X"2E",X"28",X"CB",X"7E",X"35",
		X"DD",X"A1",X"25",X"40",X"4D",X"EF",X"A0",X"32",X"B1",X"40",X"94",X"B2",X"B1",X"40",X"92",X"3A",
		X"48",X"87",X"00",X"33",X"D6",X"39",X"10",X"21",X"BF",X"B2",X"BA",X"48",X"0E",X"29",X"EB",X"7E",
		X"3D",X"55",X"A1",X"AF",X"C8",X"4D",X"67",X"28",X"92",X"3A",X"C8",X"34",X"B2",X"3A",X"C8",X"2E",
		X"28",X"32",X"B9",X"48",X"D6",X"2D",X"10",X"2C",X"D6",X"38",X"20",X"23",X"12",X"BA",X"48",X"56",
		X"AD",X"30",X"29",X"56",X"B8",X"20",X"AD",X"DE",X"AC",X"C6",X"AB",X"6F",X"4B",X"A9",X"26",X"08",
		X"21",X"D6",X"A7",X"29",X"56",X"B2",X"BB",X"48",X"23",X"76",X"32",X"BC",X"48",X"3E",X"28",X"32",
		X"A0",X"44",X"EE",X"00",X"80",X"09",X"14",X"32",X"E8",X"44",X"EE",X"00",X"80",X"09",X"14",X"73",
		X"D6",X"2A",X"20",X"3B",X"12",X"E8",X"4C",X"C6",X"08",X"CA",X"8B",X"35",X"12",X"30",X"48",X"56",
		X"89",X"5A",X"23",X"9D",X"6B",X"8A",X"9D",X"87",X"80",X"3F",X"92",X"44",X"40",X"C6",X"FF",X"CA",
		X"1C",X"35",X"12",X"AF",X"E8",X"94",X"A7",X"80",X"2B",X"B2",X"27",X"48",X"12",X"48",X"E8",X"AF",
		X"6A",X"23",X"9D",X"32",X"F3",X"46",X"94",X"B2",X"F3",X"46",X"92",X"88",X"40",X"56",X"88",X"30",
		X"2A",X"96",X"2F",X"47",X"2E",X"28",X"21",X"2E",X"00",X"01",X"6E",X"92",X"D3",X"4E",X"90",X"90",
		X"6A",X"A1",X"39",X"40",X"92",X"28",X"44",X"C6",X"00",X"20",X"09",X"A3",X"D6",X"87",X"6A",X"23",
		X"1D",X"B6",X"29",X"6B",X"A3",X"35",X"BF",X"B2",X"D3",X"4E",X"DD",X"ED",X"51",X"5D",X"21",X"A8",
		X"44",X"87",X"80",X"8E",X"5D",X"A1",X"48",X"44",X"5D",X"4B",X"08",X"FE",X"80",X"0C",X"5D",X"A1",
		X"60",X"4C",X"DD",X"D6",X"2D",X"DE",X"0B",X"A0",X"09",X"4D",X"36",X"AF",X"CD",X"92",X"64",X"6B",
		X"21",X"9D",X"4D",X"3E",X"2F",X"4D",X"3D",X"6C",X"92",X"19",X"40",X"87",X"A1",X"6D",X"C8",X"A0",
		X"0A",X"92",X"38",X"48",X"D6",X"B8",X"30",X"2B",X"21",X"9D",X"48",X"5D",X"75",X"2B",X"DD",X"F4",
		X"0C",X"5D",X"E9",X"32",X"08",X"44",X"EE",X"0C",X"80",X"98",X"3F",X"B2",X"72",X"46",X"49",X"3A",
		X"77",X"84",X"56",X"FE",X"2F",X"F7",X"3B",X"12",X"04",X"F7",X"04",X"D6",X"F6",X"2F",X"77",X"33",
		X"01",X"49",X"4D",X"0C",X"8C",X"4B",X"D7",X"CA",X"64",X"9D",X"5D",X"76",X"8B",X"87",X"80",X"0D",
		X"E6",X"08",X"CA",X"34",X"1E",X"5D",X"CB",X"28",X"9E",X"5D",X"36",X"23",X"30",X"5D",X"36",X"24",
		X"0B",X"CB",X"9C",X"9E",X"4B",X"F7",X"A0",X"1E",X"5D",X"4B",X"8B",X"FE",X"6A",X"9C",X"9E",X"5D",
		X"CB",X"28",X"9E",X"5D",X"36",X"23",X"F8",X"5D",X"36",X"24",X"D5",X"6B",X"1C",X"36",X"12",X"A9",
		X"C8",X"87",X"80",X"29",X"92",X"72",X"CE",X"87",X"48",X"5D",X"B6",X"8B",X"A8",X"C6",X"88",X"36",
		X"29",X"A0",X"2A",X"45",X"6C",X"B2",X"C4",X"4E",X"DD",X"4B",X"28",X"16",X"DD",X"4B",X"28",X"76",
		X"A0",X"0B",X"4D",X"BF",X"F3",X"32",X"D3",X"46",X"5D",X"EE",X"BA",X"88",X"67",X"C6",X"2F",X"B2",
		X"DB",X"4E",X"50",X"AE",X"28",X"C6",X"D8",X"2F",X"0F",X"2F",X"0F",X"4B",X"5F",X"20",X"2B",X"D6",
		X"D0",X"AD",X"47",X"32",X"24",X"40",X"AF",X"A0",X"BA",X"32",X"67",X"40",X"DE",X"0A",X"A0",X"2D",
		X"41",X"E0",X"22",X"3E",X"48",X"32",X"6D",X"48",X"A7",X"A0",X"25",X"22",X"2F",X"4C",X"B7",X"45",
		X"62",X"74",X"EE",X"09",X"E7",X"A2",X"AF",X"44",X"21",X"08",X"A8",X"32",X"67",X"40",X"DE",X"0A",
		X"00",X"AE",X"EB",X"1B",X"36",X"36",X"28",X"A1",X"2F",X"4B",X"D6",X"20",X"00",X"21",X"5E",X"A3",
		X"76",X"43",X"01",X"43",X"F2",X"23",X"F3",X"34",X"DE",X"9B",X"B0",X"0F",X"31",X"28",X"A8",X"39",
		X"EB",X"F2",X"36",X"61",X"60",X"A2",X"3E",X"48",X"02",X"32",X"48",X"29",X"22",X"32",X"48",X"22",
		X"3A",X"40",X"92",X"09",X"C8",X"4B",X"67",X"20",X"2B",X"C6",X"88",X"A0",X"AF",X"A9",X"BA",X"08",
		X"09",X"CB",X"92",X"36",X"29",X"34",X"28",X"97",X"C5",X"EA",X"22",X"E1",X"48",X"49",X"12",X"AD",
		X"C8",X"67",X"A6",X"42",X"92",X"89",X"CC",X"F7",X"85",X"75",X"DE",X"48",X"B0",X"0A",X"96",X"6F",
		X"32",X"AD",X"48",X"32",X"AE",X"48",X"3E",X"4A",X"5F",X"22",X"3E",X"48",X"54",X"BA",X"1D",X"75",
		X"32",X"3D",X"D3",X"56",X"88",X"B0",X"AA",X"36",X"4F",X"B2",X"A6",X"40",X"92",X"1D",X"C8",X"87",
		X"C8",X"EF",X"D5",X"A1",X"C8",X"4A",X"02",X"2F",X"4C",X"2E",X"2D",X"CD",X"1C",X"73",X"D6",X"58",
		X"90",X"0A",X"16",X"00",X"12",X"6F",X"14",X"3A",X"67",X"29",X"69",X"2D",X"A0",X"E5",X"DD",X"F5",
		X"28",X"DD",X"74",X"29",X"2D",X"48",X"D5",X"A3",X"D5",X"A3",X"EB",X"D1",X"1E",X"49",X"BF",X"B2",
		X"3D",X"40",X"4D",X"12",X"9F",X"B6",X"40",X"24",X"D6",X"C6",X"F0",X"F7",X"84",X"B6",X"41",X"24",
		X"56",X"EE",X"D0",X"F7",X"04",X"B6",X"EA",X"84",X"56",X"EE",X"D0",X"B6",X"28",X"92",X"35",X"48",
		X"6B",X"CE",X"9F",X"A1",X"61",X"9F",X"47",X"AE",X"08",X"29",X"D6",X"B2",X"3D",X"40",X"47",X"AF",
		X"2F",X"27",X"A9",X"47",X"2E",X"28",X"21",X"8A",X"1F",X"01",X"5D",X"74",X"CD",X"1A",X"1F",X"21",
		X"48",X"08",X"01",X"A9",X"BB",X"08",X"4D",X"EC",X"9F",X"4D",X"EC",X"9F",X"12",X"F7",X"A3",X"76",
		X"E6",X"D0",X"77",X"A3",X"3B",X"12",X"77",X"A3",X"56",X"EE",X"D0",X"F7",X"23",X"33",X"1A",X"F7",
		X"A3",X"76",X"EE",X"F0",X"F7",X"29",X"33",X"49",X"A1",X"45",X"28",X"32",X"1C",X"40",X"27",X"CB",
		X"98",X"37",X"21",X"C7",X"1F",X"92",X"3C",X"48",X"2F",X"47",X"2E",X"28",X"09",X"D6",X"23",X"E6",
		X"C7",X"49",X"43",X"46",X"C1",X"44",X"47",X"C2",X"45",X"C0",X"C3",X"C4",X"D0",X"C7",X"C5",X"60",
		X"F8",X"46",X"E1",X"59",X"FA",X"CA",X"FD",X"5B",X"E3",X"5E",X"FC",X"CC",X"FF",X"CD",X"C0",X"C3",
		X"66",X"E1",X"E4",X"67",X"E2",X"E5",X"E6",X"E0",X"71",X"E7",X"E1",X"72",X"70",X"E2",X"73",X"74",
		X"C0",X"DF",X"F5",X"C1",X"D0",X"DE",X"C2",X"D1",X"D2",X"C0",X"D5",X"D3",X"C1",X"D6",X"D4",X"C2",
		X"F7",X"08",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"96",
		X"E5",X"16",X"E5",X"36",X"E2",X"36",X"E1",X"36",X"E1",X"16",X"E0",X"36",X"E1",X"56",X"E0",X"16",
		X"44",X"16",X"44",X"16",X"45",X"56",X"40",X"16",X"40",X"36",X"41",X"16",X"45",X"16",X"45",X"16",
		X"E5",X"3E",X"E5",X"FE",X"E0",X"3E",X"E5",X"FE",X"E0",X"FE",X"E0",X"3E",X"E5",X"3E",X"E5",X"BE",
		X"42",X"16",X"45",X"16",X"45",X"16",X"44",X"76",X"42",X"16",X"45",X"16",X"45",X"16",X"45",X"76",
		X"E0",X"BE",X"E3",X"FE",X"E0",X"3E",X"E5",X"12",X"47",X"48",X"81",X"49",X"20",X"A7",X"80",X"AC",
		X"92",X"3C",X"48",X"0F",X"27",X"CF",X"26",X"28",X"A1",X"4D",X"80",X"89",X"56",X"2B",X"76",X"E3",
		X"82",X"A5",X"E8",X"D5",X"81",X"A5",X"E8",X"12",X"31",X"48",X"5D",X"CD",X"47",X"80",X"59",X"3B",
		X"CB",X"CE",X"A3",X"6E",X"C1",X"2A",X"A7",X"48",X"DD",X"29",X"A7",X"48",X"92",X"BA",X"48",X"29",
		X"81",X"80",X"76",X"8D",X"B0",X"A8",X"76",X"98",X"B6",X"88",X"A0",X"8A",X"B6",X"8C",X"8F",X"2F",
		X"47",X"0E",X"88",X"89",X"55",X"5C",X"DD",X"EE",X"88",X"F5",X"E6",X"29",X"4D",X"1C",X"80",X"09",
		X"15",X"88",X"A9",X"3B",X"BA",X"77",X"83",X"56",X"46",X"50",X"56",X"89",X"D7",X"23",X"9B",X"1A",
		X"F7",X"2B",X"D6",X"66",X"50",X"76",X"89",X"7F",X"49",X"28",X"8A",X"29",X"8B",X"2C",X"8A",X"2D",
		X"2B",X"8E",X"08",X"8F",X"09",X"AA",X"0C",X"AB",X"0D",X"AE",X"38",X"AF",X"39",X"88",X"2A",X"89",
		X"8B",X"AE",X"46",X"AE",X"46",X"9E",X"41",X"A4",X"46",X"56",X"42",X"76",X"41",X"20",X"41",X"36",
		X"E6",X"32",X"E1",X"A2",X"E6",X"14",X"E0",X"94",X"E6",X"AE",X"E2",X"A6",X"E4",X"2E",X"E1",X"24",
		X"44",X"28",X"42",X"AA",X"46",X"2E",X"46",X"DA",X"41",X"C0",X"41",X"20",X"46",X"3A",X"42",X"9E",
		X"E3",X"54",X"E0",X"78",X"E3",X"8E",X"E2",X"A6",X"E6",X"1C",X"E0",X"A0",X"E6",X"94",X"E1",X"AE",
		X"66",X"16",X"61",X"A6",X"66",X"D4",X"60",X"22",X"66",X"CE",X"60",X"2E",X"66",X"56",X"62",X"36",
		X"E6",X"58",X"E0",X"24",X"E6",X"56",X"E2",X"36",X"E6",X"A2",X"E2",X"32",X"E6",X"18",X"E0",X"98",
		X"60",X"46",X"60",X"56",X"64",X"DC",X"60",X"60",X"64",X"FE",X"61",X"2E",X"66",X"D0",X"60",X"38",
		X"E6",X"88",X"E0",X"B4",X"E6",X"3A",X"E6",X"82",X"E4",X"1E",X"E1",X"5E",X"E3",X"06",X"E2",X"86",
		X"62",X"50",X"60",X"D0",X"60",X"6E",X"64",X"AE",X"66",X"78",X"62",X"BE",X"66",X"02",X"62",X"BA",
		X"E6",X"88",X"E2",X"68",X"E4",X"12",X"3C",X"48",X"2F",X"4F",X"2E",X"28",X"21",X"E6",X"21",X"09",
		X"46",X"2B",X"E6",X"E9",X"A2",X"B7",X"40",X"1E",X"60",X"9E",X"0F",X"43",X"71",X"A9",X"E0",X"C8",
		X"E6",X"C8",X"26",X"CD",X"98",X"CD",X"2A",X"CA",X"AA",X"CD",X"0C",X"CC",X"9A",X"CD",X"90",X"CB",
		X"36",X"CD",X"68",X"CC",X"36",X"CD",X"12",X"CD",X"B2",X"CD",X"80",X"C8",X"40",X"CA",X"F8",X"CB",
		X"14",X"C9",X"14",X"CC",X"6C",X"CB",X"90",X"CD",X"34",X"CB",X"94",X"CD",X"EA",X"CC",X"EA",X"CA",
		X"00",X"CD",X"0C",X"CA",X"D6",X"CD",X"9E",X"CC",X"96",X"CB",X"DE",X"CA",X"16",X"CA",X"00",X"C9",
		X"34",X"C9",X"DE",X"C9",X"20",X"C9",X"12",X"3C",X"E8",X"2F",X"4F",X"2E",X"28",X"21",X"6D",X"A6",
		X"01",X"CE",X"A3",X"6E",X"C1",X"FE",X"AF",X"C0",X"A3",X"DE",X"A3",X"5E",X"CB",X"75",X"92",X"30",
		X"E8",X"E6",X"1C",X"0F",X"0F",X"D6",X"2D",X"10",X"2A",X"FE",X"2D",X"2F",X"4F",X"2F",X"A9",X"EE",
		X"20",X"55",X"77",X"9E",X"08",X"C5",X"71",X"A9",X"79",X"71",X"95",X"C0",X"CB",X"2B",X"6B",X"41",
		X"21",X"72",X"04",X"73",X"29",X"B7",X"28",X"09",X"3C",X"72",X"04",X"73",X"09",X"3C",X"72",X"04",
		X"F3",X"AB",X"4D",X"DD",X"B2",X"FA",X"6E",X"2B",X"77",X"7A",X"84",X"7B",X"BF",X"09",X"C9",X"28",
		X"65",X"6A",X"9D",X"72",X"A4",X"73",X"17",X"C5",X"CA",X"3D",X"D2",X"04",X"D3",X"C9",X"B2",X"9C",
		X"48",X"0F",X"47",X"0E",X"88",X"29",X"F9",X"AA",X"01",X"CE",X"A3",X"6E",X"C1",X"FE",X"AF",X"C0",
		X"83",X"5E",X"83",X"7E",X"83",X"C3",X"55",X"FD",X"B2",X"B2",X"E8",X"1E",X"AD",X"3E",X"2B",X"E5",
		X"06",X"2E",X"F3",X"2B",X"F7",X"2B",X"14",X"8D",X"A0",X"D0",X"E9",X"09",X"C8",X"28",X"01",X"1D",
		X"80",X"65",X"41",X"F1",X"B5",X"C8",X"4B",X"91",X"22",X"01",X"22",X"02",X"22",X"05",X"22",X"30",
		X"82",X"91",X"82",X"94",X"82",X"95",X"82",X"96",X"82",X"97",X"82",X"4A",X"82",X"4D",X"82",X"42",
		X"22",X"6A",X"22",X"6B",X"22",X"58",X"22",X"5D",X"22",X"7E",X"22",X"61",X"22",X"64",X"22",X"65",
		X"82",X"D8",X"82",X"D9",X"82",X"DA",X"82",X"DB",X"82",X"DE",X"82",X"D1",X"82",X"D1",X"82",X"D2",
		X"22",X"75",X"22",X"76",X"22",X"89",X"23",X"8E",X"23",X"8F",X"23",X"9E",X"23",X"81",X"23",X"A0",
		X"83",X"28",X"89",X"46",X"40",X"21",X"48",X"C8",X"58",X"C8",X"7C",X"C8",X"50",X"C8",X"A8",X"CA",
		X"34",X"42",X"8A",X"43",X"E2",X"43",X"46",X"45",X"28",X"89",X"6C",X"41",X"28",X"88",X"28",X"89",
		X"10",X"CC",X"89",X"6E",X"45",X"2A",X"6C",X"CD",X"A0",X"CD",X"88",X"2A",X"3A",X"CA",X"FA",X"CB",
		X"2A",X"AA",X"E2",X"50",X"E5",X"8C",X"CC",X"40",X"02",X"41",X"EC",X"42",X"C6",X"41",X"2D",X"88",
		X"43",X"24",X"43",X"42",X"44",X"5A",X"45",X"EE",X"43",X"29",X"C8",X"C9",X"88",X"29",X"CE",X"CA",
		X"28",X"88",X"28",X"89",X"C0",X"41",X"29",X"28",X"E5",X"88",X"29",X"08",X"E5",X"88",X"29",X"4E",
		X"64",X"2A",X"50",X"CD",X"64",X"CD",X"08",X"2F",X"18",X"CA",X"C4",X"CA",X"06",X"CB",X"56",X"CC",
		X"04",X"C9",X"B0",X"CB",X"F2",X"CD",X"2D",X"4A",X"E2",X"0E",X"E5",X"1A",X"E1",X"CE",X"E0",X"D8",
		X"61",X"2B",X"42",X"C9",X"72",X"C8",X"34",X"C9",X"08",X"BA",X"EF",X"48",X"AF",X"40",X"4D",X"36",
		X"22",X"12",X"3C",X"48",X"D6",X"30",X"F8",X"2F",X"4F",X"2E",X"28",X"21",X"AD",X"AB",X"09",X"4E",
		X"A3",X"6E",X"C1",X"FE",X"AF",X"C0",X"A3",X"DE",X"A3",X"5E",X"A3",X"65",X"C3",X"6A",X"FD",X"BA",
		X"12",X"48",X"7F",X"1E",X"B0",X"E5",X"CD",X"F0",X"23",X"E1",X"29",X"68",X"28",X"09",X"E5",X"CD",
		X"F8",X"AB",X"E9",X"8E",X"48",X"89",X"ED",X"C5",X"F8",X"AB",X"E9",X"8E",X"48",X"89",X"4D",X"F0",
		X"23",X"F1",X"E1",X"15",X"C8",X"EB",X"6F",X"AB",X"0E",X"2C",X"73",X"04",X"72",X"1C",X"CD",X"91",
		X"2F",X"8D",X"A0",X"DE",X"49",X"45",X"2B",X"45",X"2B",X"46",X"2B",X"45",X"2B",X"45",X"2B",X"45",
		X"23",X"5F",X"23",X"52",X"23",X"55",X"23",X"CA",X"23",X"CF",X"23",X"C6",X"23",X"D9",X"23",X"DE",
		X"2B",X"45",X"2B",X"D1",X"2B",X"28",X"2C",X"45",X"2B",X"2D",X"2C",X"45",X"2B",X"45",X"2B",X"45",
		X"23",X"45",X"23",X"45",X"23",X"45",X"23",X"20",X"24",X"23",X"24",X"26",X"24",X"3B",X"24",X"45",
		X"2B",X"45",X"2B",X"32",X"2C",X"37",X"2C",X"AC",X"2C",X"A1",X"2C",X"A6",X"2C",X"28",X"0C",X"66",
		X"E4",X"3C",X"E2",X"86",X"E3",X"DE",X"E2",X"29",X"9C",X"CA",X"29",X"06",X"E5",X"2A",X"28",X"CC",
		X"8A",X"CB",X"0A",X"48",X"62",X"C6",X"60",X"2B",X"08",X"C9",X"72",X"C8",X"B0",X"CA",X"09",X"02",
		X"E2",X"2A",X"C4",X"C8",X"28",X"CB",X"29",X"48",X"E4",X"2B",X"EA",X"C9",X"8A",X"C9",X"10",X"CB",
		X"8A",X"54",X"40",X"16",X"43",X"29",X"70",X"CA",X"89",X"FC",X"45",X"29",X"BC",X"CA",X"8A",X"28",
		X"E1",X"B0",X"E2",X"8B",X"CC",X"40",X"42",X"41",X"9C",X"45",X"2A",X"28",X"E3",X"E6",X"E5",X"8A",
		X"0C",X"CA",X"42",X"CC",X"8A",X"4E",X"40",X"12",X"44",X"2A",X"48",X"C8",X"6E",X"CB",X"89",X"3E",
		X"E5",X"12",X"47",X"48",X"76",X"8A",X"80",X"F4",X"81",X"88",X"E0",X"1E",X"3A",X"2E",X"2A",X"0E",
		X"88",X"C5",X"61",X"AF",X"31",X"8F",X"FF",X"F5",X"A1",X"9E",X"FF",X"0E",X"8B",X"8E",X"8D",X"BE",
		X"2F",X"CD",X"AB",X"84",X"99",X"4C",X"5F",X"D5",X"81",X"7C",X"5F",X"2E",X"2C",X"0E",X"2D",X"16",
		X"A8",X"C5",X"0B",X"AC",X"31",X"C4",X"FF",X"F5",X"A1",X"9A",X"84",X"0E",X"AB",X"8E",X"8D",X"BE",
		X"29",X"CD",X"AB",X"84",X"81",X"09",X"E6",X"2E",X"68",X"56",X"56",X"90",X"D7",X"23",X"83",X"2D",
		X"A0",X"DF",X"49",X"55",X"FD",X"45",X"DD",X"EE",X"88",X"F5",X"A3",X"F5",X"E6",X"28",X"DD",X"2B",
		X"4D",X"E5",X"BA",X"77",X"83",X"3B",X"96",X"8F",X"83",X"2D",X"80",X"56",X"41",X"E9",X"AD",X"00",
		X"A9",X"45",X"21",X"68",X"88",X"89",X"69",X"43",X"18",X"AC",X"69",X"71",X"79",X"BD",X"48",X"43",
		X"AB",X"84",X"9E",X"44",X"81",X"08",X"E0",X"1E",X"18",X"12",X"28",X"48",X"46",X"89",X"A0",X"AE",
		X"92",X"E6",X"48",X"66",X"89",X"BE",X"A8",X"A8",X"A8",X"BE",X"8C",X"43",X"59",X"AC",X"92",X"30",
		X"E8",X"14",X"46",X"74",X"AF",X"0F",X"76",X"8E",X"B0",X"8D",X"5E",X"8E",X"4B",X"5E",X"24",X"14",
		X"B2",X"B2",X"48",X"CF",X"26",X"08",X"92",X"A4",X"48",X"27",X"A0",X"2E",X"92",X"E7",X"48",X"27",
		X"A0",X"8C",X"8E",X"88",X"AE",X"88",X"6D",X"61",X"27",X"12",X"12",X"48",X"AE",X"00",X"56",X"90",
		X"67",X"29",X"08",X"C8",X"4D",X"5E",X"2F",X"8E",X"24",X"29",X"48",X"C8",X"4D",X"5A",X"2F",X"BA",
		X"47",X"48",X"A7",X"EA",X"76",X"AE",X"12",X"A4",X"E8",X"A7",X"20",X"39",X"21",X"08",X"E0",X"0E",
		X"02",X"9E",X"28",X"BA",X"BA",X"48",X"F1",X"AC",X"F7",X"AC",X"15",X"28",X"F1",X"BA",X"AC",X"48",
		X"A7",X"00",X"39",X"21",X"68",X"CD",X"1E",X"A8",X"36",X"EB",X"23",X"36",X"38",X"23",X"1D",X"20",
		X"77",X"43",X"7E",X"AE",X"92",X"3C",X"40",X"0F",X"47",X"0E",X"08",X"29",X"8F",X"A0",X"01",X"CE",
		X"23",X"66",X"41",X"56",X"A7",X"00",X"7F",X"4F",X"23",X"5E",X"23",X"7E",X"23",X"6E",X"C3",X"ED",
		X"ED",X"3E",X"EA",X"AC",X"B6",X"38",X"4D",X"91",X"2F",X"0D",X"B6",X"EB",X"84",X"3E",X"18",X"0D",
		X"00",X"2E",X"CD",X"91",X"27",X"EB",X"42",X"AD",X"05",X"36",X"43",X"04",X"CD",X"91",X"27",X"36",
		X"03",X"AC",X"92",X"B2",X"40",X"7F",X"E9",X"55",X"31",X"68",X"08",X"99",X"79",X"41",X"B6",X"09",
		X"04",X"77",X"CD",X"91",X"27",X"2D",X"36",X"0A",X"04",X"12",X"12",X"48",X"77",X"CD",X"91",X"AF",
		X"25",X"28",X"73",X"3E",X"04",X"AC",X"92",X"B2",X"40",X"7F",X"CB",X"8D",X"A0",X"82",X"92",X"3C",
		X"E8",X"2F",X"4F",X"2E",X"28",X"21",X"7F",X"A0",X"09",X"4E",X"23",X"66",X"41",X"56",X"A7",X"CA",
		X"7E",X"AE",X"A3",X"75",X"56",X"2B",X"76",X"2B",X"46",X"2B",X"CB",X"55",X"ED",X"49",X"6D",X"0E",
		X"28",X"5D",X"7C",X"CD",X"EB",X"AF",X"56",X"E6",X"F0",X"D6",X"60",X"20",X"29",X"2C",X"43",X"62",
		X"84",X"C5",X"B1",X"AF",X"D6",X"66",X"70",X"F6",X"68",X"28",X"0A",X"C3",X"48",X"EB",X"E2",X"19",
		X"68",X"28",X"B7",X"C5",X"7A",X"56",X"E6",X"D8",X"D6",X"E8",X"20",X"2A",X"CB",X"F8",X"0D",X"00",
		X"8A",X"C3",X"58",X"8C",X"11",X"65",X"50",X"1E",X"88",X"29",X"56",X"AF",X"11",X"DE",X"E9",X"FE",
		X"46",X"50",X"76",X"00",X"80",X"8E",X"A4",X"CB",X"46",X"EB",X"21",X"86",X"D3",X"04",X"96",X"98",
		X"D3",X"19",X"B7",X"28",X"11",X"41",X"05",X"42",X"6E",X"AD",X"06",X"0A",X"DE",X"EE",X"80",X"2E",
		X"76",X"C7",X"A0",X"8A",X"AE",X"09",X"D1",X"04",X"B2",X"B2",X"E8",X"77",X"41",X"ED",X"A4",X"CD",
		X"31",X"AF",X"31",X"68",X"88",X"FE",X"EE",X"D8",X"DE",X"E8",X"80",X"24",X"DE",X"88",X"80",X"20",
		X"96",X"0B",X"83",X"12",X"12",X"48",X"D7",X"03",X"B9",X"56",X"76",X"0A",X"A0",X"AE",X"46",X"50",
		X"DE",X"E8",X"80",X"20",X"B6",X"0C",X"84",X"BA",X"B2",X"48",X"F7",X"AD",X"25",X"28",X"61",X"41",
		X"41",X"F1",X"B5",X"EA",X"EB",X"85",X"81",X"08",X"E6",X"0E",X"80",X"12",X"12",X"48",X"56",X"90",
		X"67",X"C5",X"5E",X"AF",X"A1",X"48",X"46",X"8E",X"24",X"C5",X"5E",X"AF",X"92",X"A4",X"48",X"27",
		X"48",X"12",X"47",X"48",X"07",X"20",X"69",X"12",X"3C",X"48",X"76",X"BA",X"81",X"74",X"30",X"00",
		X"AE",X"29",X"9D",X"B9",X"DE",X"A9",X"80",X"2F",X"DE",X"AB",X"A0",X"AE",X"A1",X"BA",X"91",X"FE",
		X"83",X"5E",X"83",X"7E",X"83",X"3B",X"EE",X"23",X"CE",X"23",X"63",X"FD",X"99",X"C8",X"28",X"E5",
		X"6D",X"C3",X"EE",X"2B",X"A3",X"8D",X"A0",X"D1",X"69",X"61",X"11",X"0D",X"A0",X"D9",X"E9",X"BD",
		X"80",X"7F",X"6D",X"16",X"21",X"CD",X"7D",X"81",X"6D",X"BE",X"1F",X"CD",X"37",X"80",X"6D",X"A1",
		X"83",X"29",X"D8",X"E2",X"16",X"A8",X"4D",X"DE",X"86",X"29",X"38",X"E2",X"16",X"68",X"4D",X"DE",
		X"26",X"21",X"8E",X"E6",X"BE",X"08",X"B2",X"9C",X"E8",X"2F",X"EF",X"2E",X"28",X"09",X"EE",X"23",
		X"E6",X"E9",X"D6",X"27",X"48",X"5F",X"A3",X"CE",X"A3",X"4E",X"23",X"8A",X"BB",X"0A",X"35",X"28",
		X"F5",X"C9",X"21",X"28",X"EB",X"1E",X"08",X"29",X"20",X"28",X"CB",X"56",X"00",X"3B",X"29",X"32",
		X"08",X"89",X"4B",X"CE",X"A0",X"2E",X"4B",X"C6",X"3F",X"3A",X"F3",X"4E",X"35",X"C0",X"21",X"2E",
		X"28",X"09",X"1D",X"20",X"E5",X"C9",X"12",X"E7",X"E8",X"A7",X"00",X"2E",X"21",X"49",X"20",X"EB",
		X"CE",X"AF",X"92",X"3C",X"40",X"0F",X"27",X"CF",X"26",X"28",X"A1",X"4D",X"28",X"89",X"5D",X"FE",
		X"2D",X"D6",X"0B",X"00",X"2C",X"E6",X"29",X"20",X"2A",X"23",X"23",X"4E",X"23",X"6E",X"51",X"E6",
		X"F0",X"8F",X"07",X"8F",X"57",X"F8",X"EE",X"2F",X"07",X"8F",X"07",X"33",X"67",X"F9",X"6E",X"2A",
		X"E6",X"B7",X"2F",X"2F",X"2F",X"3E",X"28",X"30",X"29",X"3C",X"5F",X"02",X"1A",X"48",X"19",X"54",
		X"EE",X"29",X"E7",X"F8",X"49",X"BA",X"98",X"48",X"DE",X"B8",X"90",X"2D",X"7E",X"B8",X"6B",X"00",
		X"27",X"21",X"CA",X"A7",X"4F",X"2E",X"28",X"09",X"56",X"32",X"3C",X"48",X"C9",X"7F",X"0E",X"29",
		X"EE",X"D8",X"07",X"8F",X"07",X"8F",X"AF",X"28",X"0F",X"3E",X"08",X"2B",X"A3",X"43",X"33",X"AF",
		X"CD",X"0A",X"18",X"52",X"E6",X"27",X"EB",X"0A",X"18",X"04",X"55",X"E6",X"17",X"E8",X"55",X"FE",
		X"48",X"EF",X"49",X"FD",X"EE",X"B7",X"A0",X"2F",X"D5",X"66",X"40",X"76",X"BE",X"EF",X"49",X"AD",
		X"05",X"C9",X"12",X"B2",X"E8",X"6F",X"3E",X"28",X"1E",X"A8",X"51",X"AA",X"77",X"04",X"70",X"04",
		X"34",X"FA",X"EE",X"2B",X"77",X"9D",X"A0",X"DA",X"49",X"1E",X"28",X"78",X"84",X"79",X"A3",X"1D",
		X"20",X"D1",X"1D",X"20",X"F4",X"C9",X"41",X"E3",X"42",X"EB",X"41",X"EF",X"65",X"EE",X"40",X"EA",
		X"C0",X"E9",X"C4",X"E5",X"E4",X"E4",X"8F",X"2E",X"8D",X"2C",X"8B",X"2A",X"8A",X"29",X"89",X"17",
		X"00",X"22",X"00",X"49",X"00",X"7E",X"00",X"8C",X"01",X"A2",X"01",X"C9",X"01",X"EC",X"01",X"0C",
		X"A1",X"1D",X"A1",X"4F",X"A1",X"53",X"A1",X"2C",X"A2",X"B8",X"A2",X"71",X"A2",X"F7",X"A2",X"18",
		X"02",X"4D",X"02",X"75",X"02",X"80",X"03",X"E9",X"03",X"FA",X"03",X"E3",X"03",X"3D",X"03",X"35",
		X"A3",X"40",X"A3",X"28",X"A4",X"B3",X"A4",X"EF",X"A4",X"FD",X"A4",X"07",X"A4",X"45",X"A4",X"3F",
		X"05",X"82",X"05",X"F3",X"05",X"31",X"05",X"21",X"00",X"48",X"00",X"7A",X"00",X"51",X"00",X"BA",
		X"A1",X"68",X"A1",X"63",X"A1",X"FC",X"A1",X"1C",X"A1",X"92",X"A1",X"52",X"A1",X"DF",X"A1",X"A7",
		X"02",X"EC",X"02",X"D2",X"02",X"2F",X"02",X"12",X"02",X"44",X"02",X"9B",X"03",X"96",X"03",X"F9",
		X"A3",X"EF",X"A3",X"0C",X"A3",X"9B",X"A3",X"4F",X"A3",X"DB",X"A3",X"31",X"A4",X"7F",X"A4",X"FC",
		X"04",X"0D",X"04",X"6C",X"04",X"52",X"04",X"81",X"05",X"D8",X"05",X"1F",X"05",X"77",X"05",X"8B",
		X"86",X"CA",X"BA",X"8E",X"43",X"32",X"86",X"CD",X"BA",X"28",X"8F",X"BC",X"41",X"24",X"14",X"CA",
		X"0C",X"94",X"E4",X"AC",X"B4",X"45",X"0C",X"5C",X"E1",X"AC",X"7C",X"43",X"0C",X"5C",X"E4",X"AC",
		X"88",X"20",X"36",X"C9",X"AE",X"8E",X"41",X"2F",X"B6",X"CB",X"BB",X"96",X"44",X"2F",X"38",X"CC",
		X"0E",X"34",X"E5",X"AF",X"24",X"46",X"2C",X"C4",X"E6",X"8C",X"29",X"B8",X"E3",X"AB",X"2E",X"9E",
		X"42",X"23",X"96",X"CA",X"AC",X"08",X"43",X"24",X"00",X"CB",X"AC",X"22",X"45",X"24",X"A2",X"CD",
		X"0C",X"8E",X"4C",X"40",X"08",X"9E",X"E2",X"8F",X"36",X"42",X"2F",X"08",X"E3",X"8F",X"A0",X"43",
		X"0F",X"22",X"65",X"2F",X"0F",X"A6",X"61",X"2F",X"1E",X"CA",X"1C",X"B4",X"63",X"2F",X"16",X"CB",
		X"0B",X"3E",X"E5",X"2F",X"36",X"CC",X"0A",X"A4",X"E5",X"39",X"2D",X"20",X"E3",X"2D",X"0C",X"CD",
		X"0E",X"1E",X"63",X"2F",X"AE",X"C9",X"0D",X"B4",X"62",X"2D",X"0F",X"00",X"62",X"20",X"80",X"CC",
		X"08",X"10",X"E1",X"20",X"98",X"CD",X"08",X"80",X"E2",X"20",X"80",X"CC",X"08",X"90",X"E3",X"20",
		X"08",X"2B",X"0E",X"CA",X"9A",X"8E",X"63",X"32",X"0E",X"CD",X"9A",X"28",X"8D",X"0E",X"61",X"2D",
		X"2E",X"CB",X"2D",X"0E",X"E4",X"2D",X"D8",X"C9",X"08",X"70",X"E3",X"20",X"D8",X"CC",X"08",X"B0",
		X"61",X"20",X"3A",X"CA",X"0C",X"90",X"62",X"20",X"30",X"CB",X"0C",X"BE",X"64",X"21",X"38",X"CD",
		X"2C",X"9E",X"E5",X"21",X"2D",X"2E",X"E1",X"2B",X"AE",X"CA",X"2B",X"2E",X"E4",X"2B",X"10",X"C9",
		X"0F",X"9E",X"63",X"21",X"0D",X"2E",X"61",X"32",X"6C",X"CA",X"9C",X"74",X"63",X"2C",X"D8",X"CC",
		X"08",X"1C",X"E5",X"24",X"28",X"24",X"CC",X"C9",X"2D",X"7C",X"E1",X"20",X"62",X"CA",X"2D",X"D0",
		X"61",X"2E",X"CC",X"CB",X"0C",X"E4",X"63",X"2C",X"4C",X"CC",X"0C",X"7A",X"64",X"2D",X"6C",X"CC",
		X"2D",X"FC",X"E4",X"2C",X"BC",X"CD",X"0C",X"F4",X"E5",X"2C",X"2C",X"7C",X"E1",X"2B",X"62",X"C9",
		X"0D",X"7A",X"63",X"2D",X"EC",X"CB",X"0D",X"2E",X"D8",X"C9",X"88",X"06",X"62",X"2E",X"26",X"CA",
		X"2E",X"2C",X"E4",X"2E",X"30",X"CC",X"2E",X"92",X"E5",X"2E",X"28",X"21",X"78",X"C9",X"2D",X"50",
		X"61",X"25",X"78",X"C9",X"0C",X"50",X"62",X"21",X"F0",X"CA",X"88",X"78",X"64",X"20",X"E8",X"CC",
		X"08",X"74",X"E5",X"2F",X"A8",X"CD",X"09",X"2C",X"58",X"C9",X"2B",X"F8",X"E1",X"2B",X"C0",X"CA",
		X"AB",X"78",X"44",X"2E",X"AE",X"14",X"41",X"2C",X"34",X"C9",X"8C",X"0C",X"42",X"2C",X"1C",X"CA",
		X"2C",X"04",X"E2",X"8C",X"B4",X"42",X"2C",X"2C",X"E3",X"8C",X"84",X"43",X"2C",X"0C",X"E4",X"8C",
		X"1C",X"CC",X"8C",X"8C",X"44",X"2C",X"14",X"CC",X"8C",X"14",X"45",X"2C",X"34",X"CD",X"8C",X"28",
		X"09",X"BC",X"E2",X"8C",X"0E",X"41",X"2E",X"86",X"E1",X"8E",X"AC",X"42",X"2E",X"10",X"E2",X"8E",
		X"8C",X"CC",X"8E",X"B8",X"44",X"2E",X"2E",X"CD",X"8E",X"8E",X"45",X"2E",X"8C",X"26",X"41",X"2F",
		X"0E",X"44",X"2F",X"90",X"E1",X"8F",X"30",X"44",X"2F",X"A8",X"AC",X"41",X"0C",X"04",X"E1",X"AC",
		X"8C",X"CC",X"8E",X"58",X"42",X"2E",X"44",X"CA",X"8E",X"B8",X"44",X"2E",X"CC",X"CD",X"AC",X"EC",
		X"E5",X"AC",X"2C",X"0C",X"E1",X"AB",X"DA",X"42",X"0B",X"44",X"E2",X"AB",X"92",X"41",X"0B",X"8D",
		X"BC",X"C9",X"8C",X"30",X"42",X"20",X"9A",X"CB",X"AE",X"24",X"44",X"3C",X"CE",X"CD",X"BA",X"28",
		X"0B",X"98",X"E1",X"8D",X"26",X"41",X"2D",X"F4",X"E1",X"8C",X"AE",X"42",X"2D",X"10",X"E2",X"8D",
		X"98",X"CC",X"8D",X"AE",X"44",X"2D",X"F0",X"CC",X"A8",X"70",X"45",X"20",X"0E",X"CD",X"8D",X"98",
		X"E5",X"8D",X"2E",X"B8",X"E1",X"8E",X"26",X"41",X"2E",X"CE",X"E4",X"8E",X"18",X"44",X"2E",X"86",
		X"44",X"2E",X"F0",X"CC",X"8E",X"22",X"8C",X"CD",X"8C",X"42",X"43",X"2C",X"18",X"CA",X"8C",X"7E",
		X"E1",X"8B",X"BC",X"45",X"2C",X"04",X"E5",X"8C",X"64",X"41",X"2B",X"20",X"E2",X"8C",X"C6",X"43",
		X"8C",X"BC",X"45",X"2C",X"A8",X"42",X"43",X"2E",X"18",X"CA",X"8E",X"7E",X"41",X"2E",X"FA",X"C9",
		X"3A",X"C4",X"E1",X"9A",X"40",X"41",X"2E",X"26",X"E2",X"8E",X"F4",X"43",X"2E",X"8F",X"6C",X"41",
		X"1C",X"E2",X"62",X"2D",X"FC",X"CA",X"8C",X"64",X"63",X"3C",X"4A",X"CC",X"0E",X"E8",X"64",X"24",
		X"6C",X"CD",X"1C",X"2C",X"42",X"C9",X"2D",X"FA",X"E2",X"2D",X"4C",X"CB",X"2D",X"6C",X"E4",X"2D",
		X"0F",X"68",X"61",X"3A",X"EC",X"C9",X"0E",X"EA",X"62",X"2E",X"DA",X"CB",X"0D",X"7A",X"64",X"2D",
		X"64",X"CC",X"2D",X"62",X"E5",X"3A",X"2E",X"68",X"E0",X"32",X"76",X"C9",X"39",X"EA",X"E2",X"2D",
		X"DA",X"CB",X"0D",X"7A",X"64",X"2D",X"EC",X"CA",X"89",X"2D",X"C8",X"C9",X"98",X"EE",X"62",X"32",
		X"48",X"CB",X"18",X"EE",X"E4",X"32",X"48",X"CD",X"18",X"28",X"2C",X"6E",X"E1",X"30",X"98",X"CA",
		X"1C",X"58",X"63",X"39",X"4E",X"CD",X"9A",X"29",X"4E",X"C9",X"19",X"20",X"8C",X"C9",X"0E",X"68",
		X"E2",X"2F",X"04",X"C9",X"2E",X"E8",X"E2",X"2F",X"FC",X"CB",X"2F",X"20",X"E5",X"2F",X"F4",X"CB",
		X"0F",X"A0",X"65",X"2F",X"88",X"68",X"62",X"2F",X"8C",X"C9",X"0E",X"A4",X"61",X"2E",X"68",X"CA",
		X"2F",X"5C",X"E3",X"2E",X"08",X"CD",X"2F",X"DC",X"E3",X"2E",X"00",X"CD",X"2F",X"2F",X"6E",X"C9",
		X"89",X"EE",X"61",X"21",X"06",X"CA",X"8A",X"8C",X"62",X"22",X"0E",X"CC",X"8A",X"AC",X"64",X"22",
		X"78",X"CD",X"0F",X"2B",X"6E",X"C9",X"0C",X"FE",X"E1",X"24",X"56",X"C8",X"1A",X"2B",X"64",X"C9",
		X"9C",X"34",X"63",X"2C",X"64",X"CC",X"9C",X"28",X"8E",X"4C",X"61",X"2D",X"4C",X"CB",X"0D",X"4C",
		X"E4",X"2D",X"3C",X"C9",X"2D",X"1C",X"E2",X"2D",X"3C",X"CC",X"2D",X"1C",X"E5",X"2D",X"24",X"C9",
		X"0D",X"8C",X"62",X"2D",X"2C",X"CC",X"0D",X"8C",X"65",X"2D",X"74",X"C9",X"0D",X"FC",X"63",X"2D",
		X"F4",X"CC",X"2D",X"2C",X"EC",X"C9",X"0D",X"34",X"E1",X"3B",X"24",X"C9",X"3B",X"D4",X"E1",X"25",
		X"A8",X"EC",X"41",X"35",X"84",X"CB",X"BD",X"66",X"42",X"2C",X"E4",X"CA",X"8C",X"26",X"44",X"2C",
		X"04",X"44",X"2C",X"44",X"E4",X"BD",X"F4",X"45",X"0D",X"AB",X"68",X"41",X"0F",X"EE",X"E2",X"8C",
		X"DC",X"CA",X"8C",X"E4",X"42",X"2C",X"D2",X"CA",X"8C",X"26",X"44",X"2C",X"9C",X"CC",X"8C",X"A4",
		X"E4",X"8C",X"32",X"44",X"2C",X"6C",X"E5",X"8C",X"F4",X"45",X"2C",X"A9",X"18",X"41",X"09",X"AC",
		X"42",X"22",X"A0",X"CA",X"8E",X"2E",X"43",X"2C",X"80",X"CB",X"8C",X"BA",X"43",X"2E",X"4A",X"CC",
		X"0B",X"60",X"E4",X"A9",X"BE",X"45",X"0A",X"8D",X"00",X"41",X"2D",X"AC",X"E2",X"AC",X"FE",X"44",
		X"8C",X"C0",X"44",X"2C",X"92",X"CA",X"AC",X"2C",X"FC",X"CB",X"8C",X"38",X"45",X"2C",X"A0",X"CD",
		X"2C",X"B4",X"E5",X"8C",X"28",X"8D",X"1C",X"41",X"1B",X"A4",X"E2",X"B8",X"64",X"43",X"18",X"E6",
		X"44",X"3F",X"04",X"CD",X"9F",X"2B",X"84",X"C9",X"9B",X"32",X"42",X"2D",X"FA",X"CC",X"AA",X"3C",
		X"0C",X"41",X"2D",X"BC",X"E1",X"8D",X"04",X"41",X"2D",X"B4",X"E1",X"8D",X"2C",X"42",X"2D",X"9C",
		X"42",X"2D",X"84",X"CA",X"8D",X"BC",X"42",X"2D",X"AC",X"CB",X"8D",X"34",X"43",X"2D",X"A4",X"CB",
		X"2D",X"B4",X"E3",X"8D",X"2C",X"44",X"2D",X"9C",X"E4",X"8D",X"24",X"44",X"2D",X"94",X"E4",X"8D",
		X"AC",X"CD",X"8D",X"34",X"45",X"2D",X"A4",X"CD",X"8D",X"B4",X"45",X"2D",X"88",X"24",X"CE",X"C9",
		X"2C",X"DE",X"E1",X"8C",X"66",X"41",X"2C",X"D6",X"E1",X"8C",X"0C",X"43",X"2C",X"BC",X"E3",X"8C",
		X"A4",X"CB",X"8C",X"B4",X"43",X"2C",X"4A",X"CC",X"8C",X"5A",X"44",X"2C",X"42",X"CC",X"8C",X"DA",
		X"E4",X"8C",X"0C",X"EC",X"E1",X"A8",X"5C",X"41",X"08",X"E4",X"E1",X"A8",X"54",X"41",X"08",X"8A",
		X"63",X"20",X"1A",X"CB",X"88",X"AA",X"63",X"20",X"3A",X"CB",X"88",X"40",X"64",X"20",X"D0",X"CC",
		X"08",X"C0",X"E4",X"20",X"D0",X"CC",X"08",X"2B",X"5C",X"C9",X"2C",X"A4",X"E3",X"2E",X"E8",X"CC",
		X"88",X"28",X"8F",X"76",X"61",X"2B",X"FE",X"C9",X"0B",X"36",X"62",X"2B",X"BE",X"CA",X"0B",X"46",
		X"E2",X"2B",X"8E",X"CB",X"2B",X"C6",X"E2",X"2B",X"86",X"CB",X"2B",X"F6",X"E4",X"2B",X"16",X"CD",
		X"0B",X"1C",X"65",X"2B",X"5C",X"CE",X"0B",X"80",X"65",X"2B",X"E8",X"CE",X"0B",X"34",X"64",X"2D",
		X"0E",X"6A",X"E1",X"2C",X"56",X"C9",X"2C",X"76",X"E1",X"2C",X"62",X"C9",X"2C",X"46",X"E2",X"2C",
		X"52",X"CA",X"0C",X"C6",X"62",X"2C",X"72",X"CA",X"0C",X"6A",X"64",X"2C",X"FE",X"CC",X"0C",X"1C",
		X"E5",X"2C",X"98",X"CD",X"2C",X"80",X"E5",X"2C",X"84",X"CD",X"2C",X"21",X"78",X"C9",X"38",X"16",
		X"62",X"2A",X"8A",X"CB",X"0C",X"A6",X"63",X"2C",X"D0",X"CB",X"88",X"4C",X"64",X"2C",X"74",X"CC",
		X"2C",X"1A",X"E5",X"2C",X"A0",X"CD",X"2F",X"23",X"EC",X"CC",X"2C",X"22",X"E3",X"20",X"78",X"C9",
		X"88",X"1A",X"65",X"2D",X"D0",X"CB",X"88",X"16",X"62",X"2E",X"20",X"CA",X"0E",X"CE",X"63",X"20",
		X"46",X"C9",X"08",X"BC",X"E3",X"20",X"D2",X"CC",X"08",X"3F",X"6E",X"C9",X"2B",X"7E",X"E1",X"2B",
		X"0E",X"CA",X"8B",X"EE",X"61",X"2B",X"7E",X"C9",X"0B",X"AE",X"62",X"23",X"1C",X"CB",X"8D",X"5C",
		X"E3",X"25",X"10",X"CB",X"09",X"D0",X"E3",X"21",X"C6",X"CC",X"3B",X"6A",X"E5",X"2B",X"6A",X"CE",
		X"0B",X"62",X"65",X"2B",X"C2",X"CD",X"0B",X"56",X"64",X"2B",X"DE",X"CD",X"0B",X"FA",X"65",X"2B",
		X"F2",X"CD",X"2B",X"FA",X"E6",X"2B",X"52",X"CD",X"2B",X"D2",X"E5",X"2B",X"52",X"CE",X"2B",X"3F",
		X"2A",X"C8",X"8C",X"1E",X"40",X"2C",X"CE",X"C9",X"8C",X"72",X"41",X"2C",X"22",X"C8",X"8C",X"9E",
		X"E0",X"8C",X"66",X"41",X"2C",X"F2",X"E1",X"8C",X"08",X"43",X"2C",X"9C",X"E3",X"8C",X"04",X"43",
		X"8C",X"B0",X"43",X"2C",X"CA",X"CD",X"8D",X"4E",X"45",X"2B",X"EA",X"CD",X"8D",X"66",X"45",X"2D",
		X"FA",X"44",X"2F",X"7E",X"E4",X"8B",X"E2",X"44",X"2B",X"66",X"E4",X"8F",X"72",X"45",X"2B",X"56",
		X"45",X"2B",X"F2",X"CD",X"8D",X"05",X"A6",X"9C",X"A6",X"4D",X"A6",X"4E",X"A6",X"59",X"A6",X"50",
		X"06",X"41",X"06",X"62",X"06",X"51",X"06",X"54",X"06",X"73",X"06",X"88",X"07",X"8F",X"07",X"98",
		X"A7",X"3D",X"A7",X"AA",X"A7",X"AB",X"A7",X"AC",X"A7",X"BD",X"A7",X"B6",X"A7",X"6F",X"A7",X"70",
		X"07",X"C3",X"07",X"F0",X"07",X"09",X"07",X"2A",X"07",X"1B",X"07",X"3C",X"07",X"05",X"07",X"26",
		X"A7",X"9F",X"A7",X"48",X"A7",X"41",X"A7",X"41",X"A7",X"41",X"A7",X"41",X"A7",X"3B",X"8A",X"C9",
		X"2E",X"41",X"0E",X"41",X"12",X"41",X"8E",X"42",X"BA",X"42",X"82",X"42",X"86",X"42",X"B6",X"42",
		X"32",X"CA",X"8A",X"CC",X"8E",X"CC",X"AE",X"CC",X"A2",X"CC",X"08",X"CD",X"0E",X"CD",X"2A",X"CD",
		X"B6",X"45",X"92",X"45",X"08",X"08",X"E1",X"88",X"E3",X"08",X"E4",X"7C",X"E3",X"40",X"E3",X"34",
		X"41",X"B4",X"43",X"94",X"44",X"28",X"8D",X"26",X"44",X"3A",X"44",X"30",X"41",X"36",X"41",X"AE",
		X"E1",X"8B",X"9A",X"42",X"9E",X"42",X"84",X"45",X"2C",X"2C",X"E3",X"18",X"E3",X"3C",X"E4",X"00",
		X"44",X"2C",X"1A",X"CA",X"1A",X"CD",X"30",X"CA",X"10",X"CD",X"8B",X"02",X"43",X"56",X"43",X"B8",
		X"E4",X"89",X"B4",X"45",X"2B",X"DE",X"E3",X"C6",X"E3",X"D6",X"E3",X"8A",X"08",X"43",X"84",X"41",
		X"0B",X"0C",X"64",X"E6",X"63",X"FA",X"63",X"2C",X"16",X"C9",X"16",X"CB",X"26",X"C9",X"26",X"CB",
		X"2A",X"00",X"E1",X"9C",X"E1",X"2E",X"BA",X"C8",X"BE",X"C8",X"08",X"CB",X"34",X"CB",X"7C",X"CC",
		X"EA",X"CC",X"08",X"28",X"88",X"18",X"61",X"42",X"62",X"2C",X"64",X"1C",X"64",X"80",X"64",X"84",
		X"E1",X"DA",X"E2",X"B0",X"E4",X"2C",X"58",X"CA",X"64",X"CA",X"7C",X"CC",X"58",X"CC",X"2C",X"EE",
		X"61",X"74",X"62",X"7C",X"63",X"64",X"64",X"20",X"48",X"C9",X"48",X"CB",X"00",X"CD",X"DC",X"CC",
		X"60",X"CC",X"54",X"C9",X"54",X"CB",X"94",X"CD",X"2D",X"5A",X"E2",X"7E",X"E4",X"72",X"E4",X"EC",
		X"64",X"E0",X"64",X"22",X"6A",X"C9",X"6E",X"C9",X"56",X"CA",X"D2",X"CA",X"8A",X"CC",X"8E",X"CC",
		X"02",X"CC",X"06",X"CC",X"D0",X"CA",X"D4",X"CA",X"2C",X"3C",X"E3",X"AE",X"E3",X"00",X"E5",X"9A",
		X"65",X"2C",X"52",X"CB",X"56",X"CB",X"E0",X"CB",X"E4",X"CB",X"0C",X"60",X"62",X"40",X"63",X"FE",
		X"E2",X"DE",X"E3",X"2C",X"18",X"CA",X"D8",X"CB",X"26",X"CA",X"E6",X"CB",X"2C",X"58",X"E3",X"5C",
		X"63",X"C0",X"63",X"C4",X"63",X"2C",X"06",X"CA",X"82",X"CA",X"32",X"CA",X"36",X"CA",X"0C",X"E6",
		X"E2",X"FA",X"E2",X"86",X"E4",X"9A",X"E4",X"2C",X"AE",X"CD",X"8A",X"CD",X"B2",X"CD",X"B6",X"CD",
		X"0C",X"48",X"61",X"4C",X"61",X"C8",X"61",X"CC",X"61",X"28",X"09",X"2E",X"08",X"28",X"0D",X"2B",
		X"28",X"2C",X"0E",X"2F",X"28",X"20",X"09",X"22",X"28",X"23",X"0C",X"25",X"28",X"2A",X"0F",X"38",
		X"08",X"39",X"1A",X"3B",X"08",X"3C",X"1D",X"3E",X"08",X"3F",X"98",X"31",X"08",X"32",X"9B",X"34",
		X"28",X"35",X"1E",X"37",X"28",X"A8",X"21",X"AA",X"28",X"AB",X"0E",X"22",X"08",X"2C",X"BC",X"35",
		X"1B",X"AF",X"19",X"B7",X"84",X"F7",X"57",X"0F",X"AB",X"0F",X"57",X"F7",X"57",X"F7",X"73",X"FF",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"97",X"97",X"97",X"97",X"97",X"F7",X"F7",X"F7",X"97",X"97",X"97",
		X"15",X"B7",X"17",X"F7",X"17",X"FF",X"75",X"FF",X"77",X"F7",X"17",X"B7",X"17",X"F7",X"57",X"FD",
		X"F7",X"D7",X"F1",X"F7",X"F1",X"F7",X"F7",X"91",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"97",X"97",
		X"17",X"B7",X"A8",X"F7",X"57",X"F7",X"77",X"FF",X"17",X"FF",X"77",X"FF",X"17",X"B5",X"77",X"FF",
		X"D7",X"F7",X"F7",X"F5",X"F7",X"F7",X"F7",X"F7",X"F7",X"97",X"97",X"D5",X"D7",X"F7",X"97",X"97",
		X"77",X"FF",X"17",X"B5",X"77",X"F7",X"17",X"B7",X"57",X"F7",X"75",X"B7",X"17",X"B7",X"77",X"FD",
		X"F7",X"F7",X"D7",X"97",X"97",X"97",X"97",X"D7",X"D7",X"F7",X"F7",X"D7",X"97",X"F7",X"D7",X"97",
		X"17",X"B3",X"57",X"B7",X"17",X"B7",X"13",X"B3",X"17",X"B7",X"17",X"B7",X"17",X"F7",X"57",X"F7",
		X"F7",X"D1",X"F7",X"D7",X"D7",X"F7",X"D7",X"D7",X"D7",X"97",X"97",X"97",X"97",X"F7",X"F7",X"F1",
		X"77",X"F7",X"57",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",
		X"D7",X"D7",X"97",X"91",X"F7",X"D7",X"D7",X"97",X"D7",X"97",X"F1",X"F7",X"F7",X"97",X"97",X"97",
		X"57",X"B1",X"57",X"F7",X"77",X"FF",X"71",X"B7",X"17",X"B7",X"77",X"B7",X"77",X"F9",X"77",X"FF",
		X"F1",X"F7",X"F7",X"F7",X"D7",X"D7",X"D7",X"D7",X"C8",X"CB",X"C9",X"CC",X"CA",X"CD",X"C8",X"CB",
		X"C6",X"E0",X"C7",X"E1",X"C0",X"E4",X"42",X"E5",X"43",X"E6",X"C0",X"71",X"47",X"72",X"D0",X"73",
		X"C8",X"DE",X"DC",X"DF",X"DD",X"D0",X"C8",X"D3",X"D1",X"D4",X"D2",X"D5",X"2E",X"18",X"CA",X"2A",
		X"0A",X"A6",X"62",X"0A",X"0A",X"58",X"64",X"0A",X"0A",X"EE",X"64",X"0A",X"0A",X"08",X"66",X"0E",
		X"2A",X"BE",X"E6",X"2D",X"2A",X"2F",X"A8",X"C9",X"29",X"2A",X"A8",X"CC",X"29",X"2A",X"38",X"CB",
		X"09",X"0A",X"56",X"65",X"09",X"0A",X"20",X"61",X"09",X"0A",X"E2",X"65",X"09",X"0A",X"38",X"63",
		X"29",X"2A",X"09",X"68",X"E3",X"2C",X"2A",X"7E",X"E3",X"23",X"2A",X"F2",X"E3",X"2B",X"2A",X"28",
		X"65",X"89",X"0E",X"38",X"65",X"88",X"0E",X"CA",X"60",X"0F",X"0D",X"EA",X"60",X"0F",X"0D",X"80",
		X"E1",X"21",X"2A",X"80",X"E1",X"21",X"2A",X"28",X"28",X"A8",X"6A",X"BA",X"6A",X"BA",X"6A",X"BA",
		X"4A",X"3A",X"4A",X"3A",X"4A",X"3A",X"4A",X"3A",X"4A",X"3A",X"59",X"3A",X"AE",X"3A",X"AE",X"3A",
		X"15",X"BA",X"01",X"BA",X"01",X"BA",X"01",X"BA",X"01",X"BA",X"01",X"BA",X"01",X"BA",X"B2",X"67",
		X"32",X"CF",X"C8",X"58",X"C8",X"58",X"C8",X"58",X"C8",X"58",X"3B",X"3A",X"68",X"5A",X"68",X"5A",
		X"7E",X"BA",X"7E",X"BA",X"7E",X"BA",X"7E",X"BA",X"5B",X"BA",X"10",X"BA",X"10",X"BA",X"09",X"7B",
		X"89",X"5B",X"5E",X"3A",X"5E",X"3A",X"5E",X"3A",X"5E",X"3A",X"59",X"3A",X"CC",X"3A",X"CC",X"3A",
		X"4C",X"BA",X"4C",X"BA",X"4C",X"BA",X"4C",X"BA",X"4C",X"BA",X"4C",X"BA",X"4C",X"BA",X"4C",X"BA",
		X"CC",X"3A",X"CC",X"3A",X"CC",X"3A",X"CC",X"3A",X"CC",X"3A",X"CC",X"3A",X"CC",X"3A",X"CC",X"3A",
		X"4C",X"BA",X"4C",X"BA",X"7E",X"BA",X"6F",X"BA",X"5B",X"BA",X"64",X"76",X"1A",X"BA",X"1F",X"BA",
		X"9F",X"3A",X"9F",X"3A",X"9F",X"3A",X"9F",X"3A",X"9F",X"3A",X"2C",X"3A",X"E9",X"DE",X"EE",X"DE",
		X"46",X"76",X"46",X"76",X"46",X"76",X"46",X"76",X"46",X"76",X"50",X"76",X"73",X"76",X"55",X"76",
		X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",
		X"7E",X"BA",X"7E",X"BA",X"7E",X"BA",X"7E",X"BA",X"73",X"BA",X"98",X"E8",X"BA",X"80",X"BC",X"99",
		X"1E",X"3B",X"F1",X"BB",X"91",X"08",X"B4",X"D3",X"B4",X"30",X"E9",X"3C",X"4D",X"4D",X"A8",X"4A",
		X"E0",X"9D",X"60",X"08",X"F7",X"BA",X"60",X"6A",X"98",X"64",X"BB",X"DC",X"69",X"28",X"28",X"28",
		X"2E",X"5B",X"90",X"B7",X"B3",X"79",X"33",X"30",X"63",X"3B",X"FA",X"49",X"88",X"34",X"B3",X"68",
		X"68",X"08",X"BC",X"BC",X"BF",X"BD",X"08",X"6B",X"BB",X"8F",X"BC",X"08",X"6B",X"BB",X"4E",X"32",
		X"29",X"8B",X"78",X"08",X"67",X"3A",X"AC",X"E9",X"B9",X"C8",X"3F",X"C6",X"26",X"39",X"27",X"3B",
		X"D8",X"C8",X"48",X"B7",X"A6",X"AD",X"C7",X"28",X"85",X"D7",X"96",X"84",X"33",X"2F",X"AA",X"2C",
		X"28",X"98",X"A8",X"3B",X"B3",X"09",X"F0",X"48",X"28",X"88",X"30",X"08",X"B3",X"3B",X"A9",X"10",
		X"68",X"24",X"20",X"70",X"28",X"BB",X"BB",X"29",X"58",X"68",X"26",X"20",X"E0",X"28",X"BB",X"BB",
		X"A9",X"38",X"E9",X"1D",X"2A",X"C0",X"A8",X"3B",X"B3",X"09",X"80",X"49",X"38",X"8A",X"C6",X"08",
		X"BB",X"BB",X"29",X"FA",X"6A",X"32",X"22",X"D2",X"28",X"BB",X"BB",X"29",X"EA",X"6B",X"32",X"22",
		X"52",X"08",X"B3",X"3B",X"A9",X"6E",X"EC",X"9A",X"2A",X"F2",X"A8",X"3B",X"B3",X"09",X"62",X"4D",
		X"32",X"22",X"D2",X"28",X"BB",X"BB",X"29",X"E6",X"6E",X"31",X"23",X"20",X"29",X"BB",X"BB",X"29",
		X"F2",X"4F",X"BF",X"8C",X"28",X"09",X"B3",X"3B",X"A9",X"05",X"68",X"99",X"2A",X"70",X"A8",X"3B",
		X"BB",X"29",X"11",X"61",X"32",X"22",X"D2",X"28",X"BB",X"BB",X"29",X"1B",X"62",X"32",X"21",X"C9",
		X"08",X"3B",X"3B",X"09",X"17",X"CB",X"9C",X"89",X"73",X"08",X"3B",X"3B",X"09",X"01",X"CC",X"9A",
		X"0A",X"D2",X"28",X"BB",X"33",X"29",X"55",X"65",X"1A",X"22",X"D2",X"28",X"33",X"BB",X"29",X"09",
		X"CE",X"9A",X"8A",X"F2",X"08",X"3B",X"3B",X"09",X"05",X"CF",X"99",X"8A",X"70",X"08",X"3B",X"3B",
		X"29",X"01",X"78",X"9C",X"28",X"3C",X"1D",X"AE",X"07",X"BF",X"17",X"D7",X"2D",X"AD",X"05",X"BD",
		X"A5",X"B7",X"74",X"8E",X"0F",X"DB",X"08",X"5F",X"3C",X"09",X"08",X"08",X"18",X"19",X"F7",X"08",
		X"5B",X"BB",X"2C",X"51",X"0C",X"C1",X"0D",X"D1",X"0E",X"C1",X"0D",X"A0",X"28",X"2C",X"24",X"2F",
		X"6F",X"27",X"67",X"E7",X"F7",X"24",X"E4",X"50",X"65",X"00",X"24",X"8C",X"89",X"6B",X"08",X"70",
		X"33",X"29",X"D2",X"23",X"0A",X"21",X"79",X"28",X"F0",X"BB",X"29",X"EE",X"0C",X"24",X"2E",X"6A",
		X"08",X"60",X"3B",X"0A",X"6B",X"1B",X"32",X"9F",X"8C",X"0E",X"4A",X"08",X"60",X"3B",X"0A",X"A3",
		X"3B",X"D2",X"1F",X"23",X"2E",X"B4",X"28",X"C8",X"33",X"2A",X"F3",X"3B",X"6A",X"A8",X"0B",X"2E",
		X"BC",X"08",X"60",X"3B",X"0A",X"3D",X"1C",X"04",X"28",X"8A",X"0E",X"3E",X"08",X"60",X"3B",X"0A",
		X"77",X"3C",X"EE",X"A8",X"0B",X"2E",X"14",X"28",X"E0",X"BB",X"2A",X"7D",X"3D",X"2A",X"21",X"22",
		X"0D",X"AD",X"08",X"60",X"3B",X"0A",X"17",X"1D",X"4C",X"29",X"8C",X"0D",X"3F",X"08",X"60",X"3B",
		X"2A",X"41",X"3D",X"FE",X"21",X"24",X"2D",X"BF",X"28",X"C8",X"33",X"2A",X"2D",X"3E",X"B2",X"A9",
		X"08",X"F7",X"B7",X"BF",X"3E",X"AD",X"2C",X"08",X"3F",X"AF",X"2E",X"A5",X"A4",X"23",X"08",X"B8",
		X"28",X"D5",X"24",X"2F",X"05",X"D7",X"76",X"8D",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"BA",X"0E",X"E6",X"08",X"FF",X"3C",X"A9",X"14",X"27",X"19",X"AE",X"68",X"A8",X"5F",X"B4",X"09",
		X"28",X"B8",X"38",X"2E",X"72",X"28",X"7F",X"BC",X"29",X"EE",X"B8",X"39",X"2E",X"E8",X"28",X"7F",
		X"B4",X"09",X"CE",X"38",X"A8",X"3C",X"29",X"3C",X"BA",X"3C",X"3B",X"3C",X"3B",X"3C",X"BA",X"3C",
		X"21",X"BC",X"28",X"BC",X"3A",X"2E",X"EE",X"28",X"7F",X"BC",X"2B",X"28",X"28",X"28",X"28",X"99",
		X"33",X"1A",X"AE",X"6E",X"A8",X"6F",X"B4",X"0A",X"A8",X"08",X"A8",X"08",X"BA",X"0E",X"E6",X"08",
		X"7F",X"BC",X"2A",X"04",X"29",X"D0",X"29",X"28",X"D8",X"C8",X"48",X"B7",X"A6",X"AD",X"C7",X"68",
		X"56",X"F7",X"16",X"A4",X"3B",X"0F",X"A2",X"08",X"57",X"7F",X"F7",X"7E",X"F7",X"7F",X"47",X"2D",
		X"84",X"9D",X"96",X"CD",X"88",X"2F",X"AA",X"26",X"22",X"0A",X"28",X"7F",X"BC",X"2A",X"EC",X"2A",
		X"D0",X"0A",X"BA",X"8A",X"02",X"08",X"FF",X"3C",X"AA",X"DC",X"AD",X"DC",X"AD",X"18",X"AE",X"DA",
		X"28",X"7F",X"BC",X"2A",X"44",X"28",X"A4",X"29",X"38",X"2E",X"72",X"28",X"7F",X"BC",X"2C",X"38",
		X"AE",X"78",X"AE",X"50",X"AE",X"38",X"AF",X"49",X"5D",X"76",X"BE",X"34",X"5D",X"F7",X"BE",X"C6",
		X"2B",X"A0",X"21",X"5D",X"56",X"25",X"14",X"C6",X"2B",X"5D",X"77",X"25",X"12",X"28",X"4C",X"C6",
		X"A9",X"EF",X"5D",X"76",X"A8",X"C6",X"56",X"90",X"5D",X"F7",X"A8",X"22",X"AF",X"44",X"5D",X"F5",
		X"2F",X"5D",X"74",X"20",X"54",X"56",X"2A",X"D8",X"EB",X"8C",X"6B",X"5D",X"34",X"3E",X"DD",X"76",
		X"BE",X"C6",X"AF",X"A0",X"29",X"5D",X"D6",X"1F",X"94",X"C6",X"AF",X"5D",X"F7",X"1F",X"4D",X"D4",
		X"FA",X"A1",X"AC",X"BC",X"CD",X"66",X"68",X"32",X"20",X"4C",X"D6",X"2A",X"F8",X"4D",X"8C",X"6B",
		X"92",X"88",X"44",X"87",X"68",X"32",X"0F",X"44",X"DE",X"28",X"78",X"A1",X"3F",X"3D",X"A2",X"0B",
		X"EC",X"3F",X"32",X"6D",X"E8",X"B2",X"3A",X"4C",X"32",X"DA",X"EE",X"49",X"DD",X"B4",X"3E",X"5D",
		X"D6",X"1E",X"EE",X"0F",X"6A",X"24",X"4B",X"5D",X"D6",X"8D",X"94",X"56",X"0B",X"30",X"0A",X"36",
		X"29",X"5D",X"77",X"25",X"EB",X"8C",X"6B",X"5D",X"CB",X"28",X"7E",X"4A",X"CA",X"BD",X"12",X"A9",
		X"40",X"87",X"4A",X"C2",X"3D",X"32",X"1E",X"44",X"94",X"B2",X"1E",X"44",X"EE",X"0B",X"68",X"32",
		X"3F",X"4C",X"14",X"B2",X"3F",X"4C",X"D6",X"30",X"30",X"EC",X"D6",X"2B",X"20",X"60",X"DD",X"ED",
		X"5D",X"A1",X"28",X"44",X"4D",X"AA",X"4C",X"5D",X"4B",X"08",X"B6",X"5D",X"A1",X"48",X"44",X"4D",
		X"02",X"6C",X"DD",X"4B",X"28",X"96",X"DD",X"A1",X"60",X"4C",X"CD",X"A2",X"6C",X"5D",X"CB",X"28",
		X"B6",X"5D",X"A1",X"08",X"46",X"4D",X"AA",X"4C",X"5D",X"4B",X"08",X"A6",X"5D",X"A1",X"28",X"46",
		X"CD",X"A2",X"6C",X"5D",X"CB",X"28",X"96",X"5D",X"21",X"68",X"EE",X"4D",X"02",X"6C",X"DD",X"4B",
		X"08",X"B6",X"5D",X"C1",X"96",X"0F",X"EE",X"0F",X"A1",X"36",X"3D",X"6F",X"26",X"08",X"01",X"76",
		X"32",X"25",X"EC",X"6B",X"A4",X"6B",X"28",X"28",X"29",X"2A",X"2B",X"2A",X"2B",X"2A",X"DD",X"4B",
		X"08",X"16",X"96",X"F7",X"B2",X"3F",X"40",X"CB",X"AE",X"89",X"4D",X"48",X"4D",X"CA",X"E0",X"3D",
		X"12",X"AC",X"E8",X"DE",X"29",X"B0",X"2F",X"94",X"32",X"AC",X"E8",X"6B",X"C4",X"BD",X"BF",X"B2",
		X"29",X"40",X"B2",X"28",X"40",X"CB",X"1E",X"B8",X"3F",X"B2",X"2C",X"40",X"92",X"0E",X"44",X"56",
		X"2B",X"80",X"0B",X"AF",X"00",X"20",X"12",X"21",X"EC",X"7E",X"08",X"6B",X"29",X"BE",X"12",X"21",
		X"CC",X"4D",X"97",X"BF",X"21",X"48",X"A8",X"BE",X"AB",X"78",X"4B",X"E6",X"4A",X"18",X"B6",X"3C",
		X"CB",X"AB",X"3D",X"20",X"2C",X"29",X"EB",X"22",X"BE",X"4D",X"DD",X"B2",X"CB",X"E6",X"CA",X"AA",
		X"B6",X"3C",X"4B",X"AB",X"BF",X"2E",X"88",X"32",X"BD",X"40",X"AF",X"20",X"7A",X"2E",X"E9",X"97",
		X"C5",X"EA",X"56",X"A3",X"0E",X"68",X"E6",X"D8",X"D6",X"48",X"20",X"63",X"12",X"A9",X"48",X"87",
		X"4A",X"07",X"B6",X"32",X"20",X"40",X"AF",X"A0",X"36",X"C5",X"7D",X"2E",X"A0",X"BE",X"28",X"A1",
		X"32",X"4B",X"CB",X"EE",X"00",X"26",X"0E",X"32",X"B7",X"45",X"6A",X"4B",X"56",X"20",X"2A",X"4B",
		X"7E",X"29",X"06",X"28",X"35",X"20",X"AC",X"29",X"6B",X"5A",X"B6",X"36",X"A9",X"B2",X"20",X"40",
		X"32",X"A1",X"48",X"9F",X"32",X"A3",X"48",X"32",X"BE",X"48",X"A7",X"A0",X"2D",X"36",X"25",X"B2",
		X"B6",X"40",X"79",X"C1",X"21",X"48",X"A8",X"97",X"CD",X"EA",X"4B",X"E6",X"4A",X"10",X"B6",X"3C",
		X"CB",X"AB",X"CD",X"DD",X"B2",X"2E",X"68",X"BE",X"2B",X"4B",X"66",X"4A",X"17",X"BE",X"1C",X"BD",
		X"4A",X"A1",X"B6",X"4B",X"23",X"29",X"6B",X"91",X"B6",X"9F",X"B2",X"2A",X"C8",X"73",X"EE",X"70",
		X"D6",X"48",X"30",X"20",X"D6",X"F8",X"00",X"2C",X"D6",X"E8",X"20",X"AB",X"12",X"A9",X"48",X"87",
		X"80",X"8D",X"92",X"9A",X"C8",X"C6",X"2E",X"56",X"2C",X"B0",X"BC",X"56",X"28",X"30",X"B8",X"32",
		X"DA",X"4E",X"CB",X"77",X"20",X"67",X"3E",X"58",X"EE",X"20",X"C5",X"EC",X"EB",X"3E",X"BF",X"73",
		X"EE",X"98",X"DE",X"98",X"80",X"18",X"D3",X"C6",X"2F",X"56",X"AB",X"20",X"29",X"56",X"AE",X"20",
		X"2D",X"56",X"2F",X"CA",X"A2",X"BF",X"12",X"A9",X"48",X"87",X"00",X"25",X"12",X"32",X"48",X"C6",
		X"8E",X"56",X"88",X"B0",X"2D",X"56",X"0C",X"30",X"29",X"32",X"72",X"46",X"4B",X"77",X"80",X"1D",
		X"C5",X"64",X"EE",X"20",X"3E",X"B8",X"32",X"DA",X"EE",X"D2",X"32",X"C3",X"EE",X"92",X"E0",X"4E",
		X"4B",X"1F",X"B2",X"60",X"46",X"36",X"09",X"B2",X"2A",X"40",X"D3",X"C6",X"39",X"56",X"39",X"4A",
		X"C3",X"BF",X"D6",X"B8",X"CA",X"C3",X"37",X"DE",X"39",X"4A",X"C3",X"BF",X"D6",X"A8",X"20",X"22",
		X"92",X"0E",X"44",X"87",X"4A",X"E3",X"3F",X"CB",X"5D",X"3F",X"DE",X"09",X"A0",X"0F",X"92",X"0E",
		X"EC",X"AF",X"CA",X"C3",X"37",X"3F",X"32",X"A9",X"E8",X"D3",X"E6",X"04",X"D6",X"04",X"00",X"EB",
		X"DE",X"80",X"80",X"DF",X"DE",X"8C",X"80",X"DB",X"92",X"28",X"40",X"87",X"6A",X"1E",X"B8",X"32",
		X"21",X"48",X"A7",X"6A",X"3E",X"B0",X"53",X"EE",X"6A",X"4A",X"B1",X"BF",X"D6",X"6A",X"00",X"B3",
		X"92",X"2A",X"40",X"87",X"A0",X"AB",X"26",X"08",X"D3",X"56",X"48",X"20",X"0D",X"AC",X"DE",X"0A",
		X"20",X"A1",X"12",X"2E",X"EC",X"DE",X"2A",X"B0",X"22",X"96",X"18",X"4B",X"68",X"A0",X"2A",X"CD",
		X"64",X"B2",X"72",X"46",X"92",X"60",X"46",X"4B",X"1F",X"B2",X"60",X"46",X"96",X"00",X"B2",X"2A",
		X"E8",X"3F",X"32",X"A8",X"E8",X"B2",X"21",X"48",X"EB",X"3E",X"10",X"92",X"3C",X"4C",X"CB",X"D7",
		X"4A",X"E3",X"3F",X"32",X"28",X"40",X"AF",X"CA",X"1E",X"B8",X"96",X"09",X"B2",X"28",X"40",X"AE",
		X"2B",X"D3",X"E6",X"6A",X"00",X"2A",X"2E",X"23",X"12",X"2E",X"EC",X"DE",X"2A",X"B0",X"2B",X"24",
		X"24",X"AC",X"92",X"89",X"44",X"C6",X"F0",X"88",X"6B",X"18",X"B8",X"32",X"29",X"40",X"AF",X"CA",
		X"3E",X"B0",X"16",X"29",X"32",X"A9",X"E8",X"06",X"29",X"92",X"2E",X"4C",X"D6",X"2A",X"20",X"2F",
		X"D3",X"C6",X"EA",X"20",X"AA",X"2E",X"29",X"32",X"29",X"44",X"EE",X"F0",X"4A",X"1E",X"30",X"99",
		X"32",X"21",X"4C",X"4D",X"29",X"B3",X"12",X"A0",X"48",X"87",X"00",X"22",X"12",X"A9",X"48",X"87",
		X"6A",X"23",X"30",X"CB",X"2E",X"B9",X"3F",X"B2",X"A3",X"40",X"4D",X"0C",X"2C",X"27",X"B2",X"BE",
		X"48",X"C6",X"2E",X"A0",X"20",X"32",X"32",X"4C",X"E6",X"F6",X"32",X"32",X"4C",X"32",X"A9",X"48",
		X"AF",X"4A",X"15",X"B8",X"4D",X"09",X"33",X"5D",X"4B",X"08",X"FE",X"CA",X"5E",X"BA",X"92",X"BE",
		X"48",X"C6",X"2E",X"20",X"A6",X"32",X"32",X"4C",X"CB",X"EF",X"20",X"3B",X"F6",X"29",X"32",X"32",
		X"CC",X"36",X"DF",X"B2",X"BC",X"44",X"3F",X"B2",X"A1",X"40",X"96",X"04",X"4D",X"3D",X"ED",X"32",
		X"32",X"4C",X"CB",X"77",X"20",X"25",X"F6",X"08",X"32",X"32",X"4C",X"36",X"29",X"B2",X"AB",X"48",
		X"6B",X"B5",X"30",X"32",X"A2",X"40",X"EE",X"09",X"A0",X"1B",X"92",X"72",X"CE",X"87",X"80",X"8D",
		X"6F",X"32",X"C4",X"4E",X"E6",X"08",X"50",X"20",X"30",X"C6",X"08",X"20",X"30",X"32",X"DA",X"4E",
		X"AF",X"A0",X"AF",X"9F",X"A1",X"3C",X"B4",X"CB",X"3B",X"B9",X"3F",X"A1",X"6C",X"3C",X"6B",X"9B",
		X"B1",X"C6",X"08",X"20",X"C0",X"36",X"2B",X"A1",X"0A",X"BC",X"EB",X"33",X"B1",X"4D",X"92",X"FB",
		X"26",X"08",X"4D",X"D4",X"F2",X"32",X"29",X"44",X"DE",X"C3",X"5A",X"C7",X"30",X"36",X"4B",X"56",
		X"25",X"B0",X"2A",X"36",X"25",X"B2",X"21",X"4C",X"DD",X"4B",X"28",X"7E",X"00",X"22",X"16",X"29",
		X"A1",X"90",X"B4",X"AE",X"AB",X"CB",X"3D",X"B9",X"92",X"2A",X"C8",X"C6",X"88",X"A0",X"3F",X"32",
		X"B6",X"48",X"E6",X"2E",X"00",X"39",X"12",X"32",X"4C",X"4B",X"57",X"A0",X"22",X"D6",X"08",X"B2",
		X"9A",X"44",X"96",X"09",X"B2",X"2B",X"40",X"32",X"72",X"46",X"EE",X"F0",X"A0",X"88",X"96",X"09",
		X"21",X"05",X"34",X"6B",X"1B",X"B1",X"16",X"2A",X"21",X"FF",X"34",X"26",X"29",X"A2",X"29",X"4C",
		X"B2",X"0E",X"44",X"32",X"1E",X"44",X"AF",X"4A",X"39",X"B9",X"95",X"B2",X"1E",X"44",X"6B",X"BE",
		X"11",X"96",X"2A",X"B2",X"3E",X"4C",X"12",X"25",X"EC",X"94",X"A0",X"B2",X"0D",X"4C",X"12",X"DA",
		X"46",X"87",X"80",X"8F",X"5D",X"4B",X"08",X"06",X"92",X"72",X"46",X"C6",X"00",X"A0",X"0C",X"5D",
		X"CB",X"28",X"EE",X"92",X"23",X"48",X"A7",X"A0",X"38",X"92",X"3C",X"4C",X"CB",X"D7",X"00",X"A0",
		X"DE",X"E0",X"B0",X"2C",X"96",X"09",X"B2",X"2B",X"40",X"32",X"9A",X"44",X"4B",X"F7",X"80",X"98",
		X"E6",X"97",X"32",X"32",X"EC",X"96",X"8A",X"4D",X"35",X"6D",X"21",X"12",X"EC",X"21",X"20",X"28",
		X"36",X"0E",X"4B",X"16",X"01",X"BD",X"A0",X"F2",X"4D",X"B6",X"9E",X"32",X"AC",X"40",X"AF",X"A0",
		X"27",X"92",X"00",X"D3",X"E6",X"29",X"16",X"28",X"32",X"A0",X"D3",X"6A",X"C9",X"B2",X"12",X"60",
		X"F3",X"C6",X"09",X"36",X"08",X"B2",X"C8",X"F3",X"6A",X"C1",X"BA",X"32",X"88",X"F3",X"EE",X"09",
		X"16",X"28",X"32",X"20",X"D3",X"6A",X"C9",X"B2",X"12",X"A0",X"E8",X"AF",X"20",X"22",X"CD",X"75",
		X"4C",X"32",X"38",X"42",X"DE",X"F7",X"A0",X"9A",X"92",X"0E",X"44",X"56",X"0B",X"CA",X"24",X"4B",
		X"12",X"21",X"EC",X"94",X"32",X"21",X"EC",X"4D",X"A4",X"6B",X"12",X"21",X"EC",X"95",X"32",X"21",
		X"44",X"49",X"92",X"AC",X"40",X"87",X"92",X"38",X"42",X"A0",X"D5",X"B9",X"38",X"42",X"A1",X"2E",
		X"EC",X"DE",X"09",X"4A",X"88",X"B2",X"D6",X"22",X"CA",X"00",X"12",X"A1",X"40",X"4C",X"D6",X"23",
		X"4A",X"17",X"32",X"56",X"BA",X"20",X"3A",X"56",X"BB",X"A0",X"36",X"32",X"E0",X"45",X"4B",X"67",
		X"CA",X"40",X"B1",X"C6",X"57",X"B2",X"E8",X"4D",X"02",X"EF",X"4D",X"32",X"E1",X"4D",X"EB",X"BC",
		X"32",X"32",X"E8",X"45",X"4B",X"67",X"4A",X"C0",X"31",X"C6",X"5F",X"B2",X"E8",X"45",X"82",X"4F",
		X"4D",X"32",X"61",X"4D",X"FE",X"22",X"4F",X"32",X"3D",X"48",X"EE",X"2D",X"2E",X"A8",X"CD",X"41",
		X"6E",X"36",X"99",X"4D",X"B5",X"4D",X"6B",X"C0",X"31",X"EF",X"92",X"2B",X"C8",X"87",X"A0",X"AE",
		X"12",X"32",X"4C",X"C6",X"68",X"70",X"20",X"AE",X"21",X"08",X"4C",X"DE",X"24",X"2F",X"0F",X"2F",
		X"26",X"08",X"47",X"29",X"4B",X"66",X"80",X"1E",X"06",X"9A",X"01",X"4B",X"F6",X"A0",X"2F",X"4B",
		X"D6",X"32",X"32",X"4C",X"F6",X"68",X"32",X"32",X"4C",X"36",X"00",X"4D",X"BD",X"6D",X"3B",X"3A",
		X"DE",X"F7",X"4A",X"C0",X"31",X"CB",X"46",X"B9",X"7E",X"89",X"07",X"2F",X"07",X"6F",X"26",X"08",
		X"09",X"76",X"A7",X"A0",X"C1",X"A3",X"23",X"76",X"03",X"C6",X"29",X"76",X"20",X"2F",X"D6",X"D1",
		X"90",X"D4",X"6B",X"A1",X"32",X"56",X"AF",X"B0",X"DD",X"A3",X"A3",X"76",X"5D",X"EE",X"29",X"10",
		X"30",X"20",X"EE",X"24",X"90",X"30",X"4F",X"CB",X"48",X"B2",X"FE",X"24",X"90",X"DA",X"F6",X"B2",
		X"21",X"19",X"A8",X"29",X"4B",X"E6",X"6A",X"24",X"EB",X"5D",X"4B",X"08",X"FE",X"CA",X"84",X"4B",
		X"DD",X"4B",X"28",X"5E",X"16",X"0E",X"CD",X"BD",X"6D",X"36",X"29",X"B2",X"A1",X"48",X"BF",X"B2",
		X"BE",X"44",X"B2",X"8D",X"CC",X"B2",X"BF",X"44",X"A1",X"90",X"B4",X"A2",X"A9",X"44",X"94",X"B2",
		X"2E",X"4C",X"EB",X"8C",X"6B",X"75",X"E6",X"48",X"4F",X"75",X"14",X"34",X"E6",X"B7",X"B1",X"67",
		X"49",X"5D",X"4B",X"08",X"96",X"32",X"28",X"40",X"AF",X"20",X"8B",X"32",X"1C",X"44",X"4B",X"77",
		X"C8",X"3F",X"32",X"3C",X"EC",X"49",X"12",X"3C",X"EC",X"4B",X"57",X"68",X"BF",X"B2",X"3C",X"4C",
		X"49",X"9F",X"B2",X"8D",X"44",X"32",X"1E",X"44",X"94",X"C6",X"0B",X"B2",X"1E",X"44",X"A0",X"8B",
		X"12",X"3F",X"EC",X"94",X"E6",X"2B",X"F6",X"08",X"32",X"3F",X"EC",X"92",X"3F",X"4C",X"E6",X"2B",
		X"27",X"6F",X"26",X"08",X"A1",X"2C",X"3C",X"29",X"D6",X"B2",X"09",X"44",X"A3",X"76",X"B2",X"0A",
		X"EC",X"6B",X"16",X"B1",X"DD",X"D6",X"3E",X"94",X"E6",X"2B",X"DD",X"F7",X"3E",X"A0",X"09",X"5D",
		X"D6",X"1F",X"94",X"C6",X"0B",X"5D",X"F7",X"1F",X"A1",X"69",X"BD",X"4D",X"CE",X"48",X"6B",X"24",
		X"6B",X"5D",X"34",X"3E",X"DD",X"D6",X"3E",X"EE",X"2B",X"A0",X"09",X"5D",X"56",X"3F",X"14",X"EE",
		X"0B",X"5D",X"F7",X"1F",X"5D",X"4B",X"9A",X"4E",X"4A",X"7F",X"BD",X"32",X"08",X"44",X"EE",X"0C",
		X"20",X"B9",X"12",X"A0",X"E8",X"AF",X"EA",X"20",X"14",X"92",X"12",X"4C",X"CB",X"E7",X"20",X"26",
		X"A1",X"28",X"F1",X"5D",X"D6",X"0D",X"BD",X"67",X"4B",X"EE",X"B6",X"08",X"A0",X"1D",X"92",X"DA",
		X"EC",X"4B",X"67",X"A0",X"7B",X"A1",X"68",X"D1",X"DD",X"D6",X"2D",X"BD",X"47",X"4B",X"6E",X"B6",
		X"08",X"20",X"4D",X"5D",X"4B",X"9A",X"06",X"5D",X"4B",X"9A",X"C6",X"5D",X"56",X"9C",X"92",X"1D",
		X"E8",X"9B",X"10",X"BC",X"53",X"B2",X"3D",X"48",X"21",X"32",X"EB",X"36",X"08",X"26",X"28",X"06",
		X"28",X"4B",X"66",X"20",X"9C",X"2E",X"0A",X"29",X"D6",X"13",X"B0",X"0D",X"06",X"9E",X"6B",X"09",
		X"14",X"BF",X"C5",X"62",X"CB",X"2E",X"CB",X"4E",X"0E",X"2E",X"B7",X"CD",X"6A",X"B6",X"28",X"06",
		X"A6",X"BD",X"80",X"0C",X"01",X"CB",X"5F",X"BB",X"5D",X"76",X"3C",X"6F",X"27",X"AF",X"29",X"6F",
		X"2E",X"28",X"12",X"AD",X"48",X"34",X"47",X"A6",X"4A",X"29",X"55",X"56",X"E0",X"30",X"2B",X"DE",
		X"20",X"67",X"D6",X"5D",X"F7",X"89",X"A1",X"60",X"CA",X"5D",X"46",X"9C",X"4B",X"A9",X"01",X"76",
		X"DD",X"F7",X"2F",X"6F",X"23",X"76",X"DD",X"F7",X"20",X"EF",X"12",X"E7",X"48",X"56",X"2A",X"70",
		X"A0",X"38",X"82",X"0F",X"CC",X"97",X"CD",X"EA",X"D5",X"B0",X"29",X"5D",X"4B",X"08",X"CE",X"45",
		X"6C",X"CB",X"73",X"B4",X"A7",X"20",X"2C",X"5D",X"CB",X"28",X"0E",X"D5",X"CD",X"68",X"6D",X"D1",
		X"A1",X"D9",X"35",X"A0",X"ED",X"56",X"2C",X"A1",X"E1",X"BD",X"B0",X"BE",X"A1",X"E9",X"35",X"CB",
		X"82",X"B4",X"E6",X"29",X"20",X"2F",X"DD",X"4B",X"28",X"0E",X"EB",X"0D",X"B4",X"71",X"A7",X"20",
		X"AC",X"5D",X"4B",X"08",X"CE",X"4D",X"E8",X"4D",X"80",X"0E",X"A1",X"D9",X"35",X"CB",X"02",X"BC",
		X"21",X"E9",X"B5",X"5D",X"CB",X"20",X"6E",X"5D",X"56",X"2F",X"20",X"2F",X"D6",X"DC",X"10",X"22",
		X"6B",X"27",X"34",X"56",X"2C",X"B0",X"AB",X"A1",X"61",X"BD",X"4D",X"CE",X"E8",X"5D",X"D6",X"89",
		X"EE",X"2B",X"DD",X"F7",X"21",X"4D",X"8C",X"6B",X"DD",X"76",X"21",X"DE",X"2B",X"5D",X"77",X"21",
		X"5D",X"4B",X"A8",X"5E",X"48",X"32",X"20",X"40",X"AF",X"48",X"92",X"AB",X"C8",X"5D",X"66",X"9C",
		X"90",X"C8",X"12",X"21",X"4C",X"5D",X"6E",X"21",X"90",X"C8",X"DD",X"76",X"2F",X"87",X"E8",X"4D",
		X"B1",X"48",X"5D",X"4B",X"A8",X"B6",X"4D",X"AA",X"EC",X"36",X"8D",X"4D",X"B5",X"4D",X"4D",X"F1",
		X"22",X"32",X"A3",X"48",X"4F",X"34",X"32",X"A3",X"48",X"AE",X"28",X"A1",X"6E",X"68",X"09",X"76",
		X"FD",X"32",X"AB",X"40",X"27",X"AF",X"27",X"6F",X"92",X"89",X"44",X"56",X"00",X"B0",X"0E",X"CE",
		X"09",X"29",X"EB",X"30",X"15",X"7E",X"09",X"39",X"4F",X"A1",X"28",X"29",X"F1",X"26",X"20",X"4D",
		X"C1",X"CE",X"92",X"AB",X"40",X"EF",X"92",X"1D",X"40",X"10",X"68",X"32",X"1B",X"40",X"DE",X"F7",
		X"20",X"2C",X"BF",X"6B",X"49",X"B5",X"BF",X"B2",X"00",X"48",X"12",X"30",X"E8",X"94",X"E6",X"2B",
		X"DE",X"0B",X"96",X"08",X"80",X"0B",X"B2",X"A9",X"40",X"B2",X"1D",X"40",X"B2",X"72",X"46",X"B2",
		X"F3",X"4E",X"32",X"C4",X"EE",X"B2",X"C3",X"4E",X"C9",X"F5",X"33",X"00",X"33",X"1B",X"33",X"00",
		X"3B",X"96",X"3B",X"A1",X"3B",X"96",X"3B",X"A1",X"3B",X"34",X"3B",X"B7",X"3B",X"34",X"3B",X"B7",
		X"33",X"42",X"33",X"5D",X"33",X"42",X"33",X"92",X"47",X"48",X"D6",X"2A",X"20",X"2E",X"DD",X"D6",
		X"9A",X"87",X"80",X"2C",X"5D",X"76",X"88",X"C6",X"09",X"5D",X"F7",X"88",X"4D",X"25",X"4C",X"32",
		X"00",X"48",X"A7",X"A0",X"3B",X"92",X"28",X"4C",X"E6",X"2C",X"20",X"24",X"26",X"D1",X"DD",X"C6",
		X"0D",X"4B",X"66",X"B6",X"08",X"CA",X"11",X"BF",X"5D",X"4B",X"9A",X"CE",X"6A",X"59",X"BE",X"32",
		X"47",X"48",X"D6",X"2A",X"EA",X"D5",X"15",X"A1",X"6F",X"4C",X"DD",X"D6",X"2D",X"7E",X"2A",X"07",
		X"07",X"2F",X"47",X"AE",X"08",X"29",X"D6",X"5D",X"F7",X"0F",X"A3",X"76",X"5D",X"F7",X"88",X"87",
		X"00",X"2B",X"D6",X"29",X"E8",X"A3",X"56",X"6E",X"19",X"5D",X"77",X"21",X"29",X"2B",X"28",X"BF",
		X"CD",X"EA",X"D6",X"87",X"4A",X"35",X"48",X"5D",X"4B",X"9A",X"C6",X"A9",X"8C",X"08",X"01",X"76",
		X"DD",X"F7",X"3A",X"A6",X"D1",X"5D",X"46",X"2D",X"36",X"28",X"EB",X"B2",X"69",X"A1",X"41",X"B5",
		X"4D",X"CE",X"E8",X"5D",X"D6",X"1E",X"EE",X"9F",X"6A",X"1B",X"36",X"5D",X"D6",X"08",X"CE",X"09",
		X"DD",X"F7",X"28",X"5D",X"56",X"38",X"2E",X"2C",X"D6",X"68",X"10",X"2E",X"D6",X"48",X"30",X"2A",
		X"26",X"0B",X"28",X"5D",X"F7",X"18",X"27",X"67",X"A6",X"08",X"B0",X"09",X"A4",X"4D",X"41",X"4C",
		X"55",X"C6",X"48",X"AF",X"2F",X"4B",X"54",X"20",X"2A",X"45",X"6C",X"5D",X"46",X"21",X"F5",X"8D",
		X"5D",X"F7",X"29",X"4D",X"84",X"4B",X"F9",X"45",X"64",X"5D",X"C6",X"89",X"2D",X"5D",X"F7",X"89",
		X"C9",X"5D",X"56",X"21",X"CD",X"CF",X"B7",X"BE",X"28",X"4B",X"66",X"20",X"29",X"BC",X"29",X"68",
		X"A8",X"29",X"4B",X"E6",X"80",X"0A",X"4B",X"4A",X"4D",X"75",X"32",X"4B",X"E6",X"20",X"AA",X"4B",
		X"FA",X"A9",X"68",X"28",X"B7",X"45",X"6A",X"4B",X"66",X"20",X"2A",X"4B",X"DA",X"72",X"A7",X"4A",
		X"F6",X"BF",X"DE",X"89",X"A0",X"8A",X"5D",X"76",X"29",X"C6",X"50",X"DE",X"AF",X"CB",X"DC",X"BE",
		X"CB",X"EA",X"00",X"3C",X"DD",X"4B",X"3A",X"F6",X"00",X"AE",X"DD",X"76",X"3A",X"45",X"6C",X"5D",
		X"F7",X"1A",X"4D",X"6C",X"37",X"CB",X"46",X"BE",X"4B",X"7F",X"80",X"1C",X"5D",X"4B",X"BA",X"FE",
		X"20",X"26",X"DD",X"76",X"3A",X"45",X"6C",X"5D",X"77",X"3A",X"CD",X"78",X"B7",X"CB",X"C6",X"B6",
		X"5D",X"4B",X"3A",X"5E",X"A0",X"0F",X"5D",X"4B",X"3A",X"56",X"4D",X"CA",X"37",X"5D",X"D6",X"89",
		X"E6",X"D0",X"EE",X"2A",X"DD",X"F7",X"21",X"5D",X"36",X"3C",X"28",X"5D",X"CB",X"28",X"76",X"CC",
		X"ED",X"BF",X"5D",X"4B",X"3A",X"DE",X"A0",X"1A",X"5D",X"76",X"BA",X"87",X"A0",X"4A",X"5D",X"4B",
		X"32",X"56",X"DD",X"B6",X"2E",X"28",X"DD",X"B6",X"3E",X"28",X"DD",X"76",X"3E",X"C6",X"27",X"A0",
		X"2B",X"5D",X"B4",X"0E",X"5D",X"76",X"0E",X"56",X"0A",X"A0",X"8E",X"5D",X"4B",X"08",X"06",X"5D",
		X"CB",X"23",X"56",X"80",X"2C",X"5D",X"CB",X"28",X"EE",X"DE",X"2B",X"90",X"2F",X"5D",X"CB",X"32",
		X"96",X"CB",X"38",X"BF",X"A1",X"79",X"BD",X"5D",X"46",X"0E",X"4D",X"59",X"48",X"CB",X"24",X"4B",
		X"DD",X"4B",X"28",X"76",X"20",X"2B",X"CD",X"B7",X"73",X"4D",X"DC",X"FA",X"21",X"71",X"15",X"4D",
		X"CE",X"48",X"6B",X"24",X"4B",X"5D",X"4B",X"8D",X"4E",X"C8",X"5D",X"4B",X"1A",X"FE",X"A0",X"1C",
		X"DD",X"D6",X"2D",X"27",X"C5",X"64",X"EE",X"C4",X"DD",X"F7",X"0B",X"5D",X"36",X"24",X"D7",X"5D",
		X"4B",X"08",X"96",X"49",X"5D",X"76",X"0D",X"AF",X"6E",X"1C",X"5D",X"F7",X"8B",X"5D",X"B6",X"8C",
		X"29",X"5D",X"CB",X"28",X"9E",X"49",X"DD",X"D6",X"3E",X"AF",X"16",X"04",X"CC",X"BD",X"6D",X"5D",
		X"B4",X"1E",X"4D",X"B2",X"7B",X"4D",X"D4",X"7A",X"A1",X"69",X"BD",X"4D",X"CE",X"48",X"6B",X"24",
		X"6B",X"96",X"8B",X"4D",X"35",X"6D",X"12",X"3D",X"E8",X"5D",X"77",X"34",X"14",X"B2",X"3D",X"48",
		X"5D",X"4B",X"9A",X"16",X"5D",X"4B",X"9A",X"46",X"5D",X"4B",X"9A",X"CE",X"6A",X"24",X"4B",X"36",
		X"29",X"4D",X"8D",X"3F",X"EB",X"8C",X"6B",X"67",X"E6",X"30",X"2F",X"27",X"2F",X"47",X"50",X"EE",
		X"60",X"AF",X"27",X"AF",X"FE",X"60",X"67",X"22",X"9A",X"40",X"55",X"FC",X"A1",X"08",X"0A",X"97",
		X"C5",X"72",X"55",X"EE",X"F0",X"07",X"0F",X"07",X"CB",X"64",X"00",X"2A",X"F6",X"A8",X"EE",X"37",
		X"EE",X"BF",X"C7",X"A6",X"08",X"29",X"49",X"EF",X"EE",X"98",X"27",X"AF",X"27",X"6F",X"D0",X"C6",
		X"E0",X"27",X"2F",X"27",X"F6",X"C8",X"6F",X"82",X"1A",X"48",X"5D",X"74",X"21",X"28",X"2A",X"BF",
		X"CD",X"5A",X"D5",X"66",X"50",X"8F",X"07",X"8F",X"4B",X"4C",X"80",X"2A",X"FE",X"A8",X"C7",X"D5",
		X"F6",X"8F",X"46",X"70",X"AF",X"0F",X"AF",X"DD",X"6B",X"A8",X"6E",X"00",X"2A",X"F6",X"20",X"AD",
		X"EE",X"B7",X"FE",X"29",X"C7",X"2E",X"88",X"89",X"49",X"29",X"8A",X"2C",X"A8",X"38",X"80",X"68",
		X"A8",X"DD",X"F6",X"8D",X"5E",X"88",X"EF",X"2E",X"28",X"21",X"01",X"C8",X"A9",X"6E",X"B2",X"9B",
		X"48",X"30",X"B2",X"3B",X"48",X"C1",X"8D",X"2E",X"8F",X"20",X"A9",X"23",X"AC",X"26",X"5D",X"CE",
		X"3F",X"CB",X"89",X"2E",X"28",X"09",X"F6",X"DD",X"D7",X"89",X"83",X"56",X"7D",X"77",X"2A",X"C9",
		X"5D",X"C3",X"88",X"7E",X"68",X"D5",X"B4",X"3E",X"5D",X"FE",X"9E",X"66",X"8B",X"28",X"A9",X"D5",
		X"F6",X"9F",X"B4",X"E6",X"2B",X"DD",X"D7",X"9F",X"7D",X"CB",X"1A",X"CE",X"4A",X"36",X"68",X"DD",
		X"4B",X"3A",X"F6",X"09",X"89",X"28",X"80",X"2B",X"21",X"D7",X"77",X"D5",X"C6",X"2F",X"5D",X"6E",
		X"08",X"09",X"7D",X"75",X"2F",X"DD",X"D4",X"A8",X"F4",X"A7",X"A0",X"8B",X"76",X"89",X"48",X"DD",
		X"4B",X"3A",X"F6",X"FD",X"80",X"2F",X"DE",X"88",X"B0",X"23",X"6B",X"99",X"C8",X"F6",X"08",X"B8",
		X"2C",X"DD",X"96",X"BA",X"29",X"21",X"61",X"B5",X"6D",X"EE",X"68",X"EB",X"A4",X"CB",X"A2",X"CA",
		X"48",X"D5",X"D6",X"2E",X"47",X"0F",X"29",X"CF",X"26",X"28",X"01",X"CE",X"5D",X"FE",X"98",X"BC",
		X"76",X"77",X"A0",X"A1",X"7D",X"77",X"38",X"91",X"80",X"83",X"7D",X"34",X"2E",X"23",X"F6",X"DD",
		X"4B",X"34",X"CE",X"A8",X"AC",X"E5",X"64",X"D5",X"F7",X"24",X"A3",X"FE",X"CD",X"4C",X"6B",X"DE",
		X"68",X"DD",X"D7",X"AC",X"83",X"56",X"7D",X"77",X"0B",X"DD",X"6B",X"88",X"9E",X"DD",X"F6",X"9C",
		X"EE",X"08",X"A0",X"2F",X"5D",X"FE",X"1E",X"66",X"09",X"28",X"A8",X"C5",X"B2",X"FB",X"4D",X"B7",
		X"73",X"CD",X"DC",X"FA",X"DD",X"CB",X"28",X"76",X"00",X"2C",X"DD",X"36",X"0C",X"28",X"DD",X"56",
		X"89",X"F6",X"70",X"B8",X"8E",X"D5",X"4B",X"28",X"56",X"BA",X"BB",X"48",X"94",X"3A",X"BB",X"48",
		X"EB",X"A2",X"6C",X"DD",X"CB",X"3C",X"56",X"EA",X"B5",X"68",X"21",X"E1",X"15",X"DD",X"56",X"3E",
		X"EE",X"37",X"A0",X"20",X"5D",X"FE",X"08",X"E6",X"09",X"D5",X"F7",X"28",X"4D",X"66",X"48",X"43",
		X"A4",X"6B",X"29",X"38",X"28",X"02",X"2F",X"4C",X"12",X"28",X"EC",X"E6",X"29",X"00",X"0A",X"B7",
		X"CD",X"4A",X"5D",X"C3",X"08",X"0E",X"6B",X"E6",X"49",X"89",X"5D",X"C3",X"08",X"4E",X"5D",X"7D",
		X"2F",X"DD",X"74",X"20",X"12",X"21",X"EC",X"EE",X"2F",X"DD",X"77",X"21",X"12",X"DA",X"EE",X"A7",
		X"A1",X"E3",X"3B",X"A8",X"0B",X"29",X"7C",X"BB",X"5D",X"7D",X"09",X"D5",X"F4",X"2A",X"3F",X"29",
		X"E8",X"D3",X"29",X"21",X"28",X"09",X"CB",X"6E",X"36",X"28",X"20",X"21",X"23",X"14",X"D6",X"3C",
		X"90",X"DC",X"6B",X"8C",X"4B",X"46",X"89",X"D5",X"ED",X"C5",X"CD",X"23",X"5D",X"C3",X"08",X"7E",
		X"20",X"B5",X"DD",X"56",X"3C",X"A7",X"00",X"BF",X"E6",X"08",X"20",X"BB",X"16",X"03",X"CD",X"BD",
		X"4D",X"D5",X"4B",X"28",X"56",X"C5",X"AA",X"6C",X"92",X"B3",X"40",X"BC",X"B2",X"B3",X"40",X"BA",
		X"15",X"48",X"21",X"66",X"C1",X"2F",X"4F",X"2E",X"28",X"09",X"36",X"A7",X"04",X"36",X"08",X"12",
		X"BD",X"48",X"94",X"3A",X"BD",X"48",X"92",X"B4",X"40",X"46",X"09",X"2F",X"B2",X"B4",X"40",X"D5",
		X"E1",X"EB",X"A4",X"6B",X"DD",X"34",X"3E",X"DD",X"56",X"3E",X"E6",X"2F",X"E8",X"DD",X"56",X"2E",
		X"94",X"66",X"8F",X"D5",X"F7",X"2E",X"27",X"CF",X"26",X"28",X"A1",X"B0",X"CA",X"89",X"56",X"D5",
		X"F6",X"88",X"46",X"76",X"13",X"DD",X"6B",X"8D",X"6E",X"00",X"2A",X"C6",X"29",X"DD",X"D7",X"88",
		X"A3",X"FE",X"5D",X"7F",X"9F",X"F6",X"8A",X"8E",X"88",X"A8",X"8F",X"66",X"89",X"8E",X"89",X"28",
		X"29",X"0C",X"7D",X"71",X"0D",X"EB",X"A4",X"CB",X"28",X"88",X"28",X"89",X"28",X"8A",X"29",X"8B",
		X"89",X"2C",X"89",X"2B",X"88",X"2A",X"88",X"29",X"5D",X"C3",X"88",X"E6",X"48",X"BA",X"A0",X"48",
		X"07",X"EA",X"2E",X"CB",X"7D",X"56",X"38",X"14",X"B0",X"8B",X"7D",X"77",X"38",X"12",X"3E",X"4E",
		X"94",X"3A",X"9E",X"4E",X"EE",X"2B",X"6A",X"2E",X"CB",X"BA",X"8E",X"4E",X"5D",X"C3",X"BA",X"6E",
		X"A0",X"98",X"B5",X"D6",X"D7",X"20",X"7F",X"DD",X"96",X"BA",X"28",X"DD",X"6B",X"88",X"86",X"EB",
		X"A2",X"6C",X"94",X"F6",X"AC",X"B8",X"CF",X"D5",X"4B",X"32",X"4E",X"D5",X"D6",X"38",X"DE",X"30",
		X"B0",X"B2",X"B2",X"AB",X"E8",X"A7",X"80",X"8F",X"B2",X"AA",X"E8",X"D6",X"0A",X"10",X"05",X"12",
		X"80",X"4E",X"EE",X"08",X"A0",X"21",X"5D",X"65",X"5D",X"29",X"80",X"4E",X"6B",X"94",X"CA",X"BA",
		X"68",X"4E",X"46",X"08",X"80",X"9E",X"7D",X"E5",X"7D",X"21",X"68",X"4E",X"A2",X"8F",X"EE",X"12",
		X"A9",X"4E",X"47",X"C5",X"6B",X"78",X"5D",X"61",X"5D",X"3E",X"98",X"28",X"96",X"23",X"B2",X"2E",
		X"EE",X"D6",X"08",X"10",X"22",X"20",X"2F",X"DD",X"6B",X"BA",X"6E",X"CC",X"03",X"CB",X"B2",X"9F",
		X"4E",X"66",X"8B",X"0F",X"47",X"0E",X"88",X"29",X"D0",X"6B",X"01",X"CE",X"A3",X"6E",X"C1",X"BA",
		X"2E",X"4E",X"5E",X"A8",X"4B",X"72",X"6A",X"21",X"50",X"CB",X"8F",X"4F",X"8E",X"88",X"A9",X"4E",
		X"A3",X"6E",X"C1",X"2A",X"09",X"4E",X"92",X"2E",X"46",X"F6",X"0E",X"B8",X"0A",X"BE",X"0E",X"29",
		X"41",X"6B",X"2E",X"28",X"4F",X"09",X"6E",X"12",X"09",X"4E",X"ED",X"A8",X"32",X"21",X"EE",X"CD",
		X"D2",X"76",X"69",X"BA",X"89",X"4E",X"38",X"3A",X"89",X"4E",X"49",X"BA",X"08",X"4E",X"EE",X"D6",
		X"32",X"28",X"EE",X"12",X"09",X"4C",X"6F",X"0E",X"28",X"12",X"09",X"4E",X"FE",X"B8",X"10",X"2B",
		X"98",X"38",X"1E",X"46",X"68",X"F6",X"60",X"38",X"0D",X"B0",X"06",X"2A",X"90",X"23",X"92",X"20",
		X"EE",X"E6",X"29",X"0E",X"2B",X"20",X"2A",X"0E",X"29",X"51",X"32",X"3F",X"EE",X"D6",X"2B",X"E8",
		X"92",X"28",X"46",X"76",X"09",X"3A",X"08",X"4E",X"49",X"22",X"88",X"2E",X"0D",X"2B",X"0A",X"29",
		X"B8",X"6B",X"88",X"6B",X"98",X"6B",X"88",X"6B",X"57",X"BA",X"88",X"BA",X"B9",X"BA",X"9A",X"BA",
		X"23",X"BA",X"A4",X"BA",X"35",X"BA",X"B6",X"BA",X"47",X"BA",X"50",X"BA",X"D1",X"BA",X"62",X"BA",
		X"C3",X"BA",X"F4",X"BA",X"D5",X"BA",X"2E",X"BB",X"0F",X"BB",X"18",X"BB",X"21",X"BB",X"02",X"BB",
		X"08",X"29",X"0A",X"29",X"5D",X"EE",X"09",X"D5",X"E6",X"2A",X"ED",X"F5",X"E9",X"D1",X"DD",X"DE",
		X"28",X"7B",X"CB",X"13",X"12",X"ED",X"E8",X"E6",X"A8",X"DD",X"56",X"21",X"00",X"2A",X"EE",X"2A",
		X"3B",X"3A",X"28",X"4A",X"2A",X"3A",X"29",X"4A",X"36",X"28",X"DD",X"DE",X"09",X"9D",X"4B",X"2B",
		X"DD",X"46",X"2F",X"DD",X"66",X"20",X"C5",X"7A",X"22",X"AA",X"EA",X"D9",X"DD",X"56",X"0D",X"AF",
		X"6E",X"2F",X"57",X"1E",X"08",X"99",X"D6",X"2B",X"E6",X"EF",X"92",X"ED",X"40",X"66",X"00",X"D5",
		X"56",X"28",X"00",X"2A",X"C6",X"2A",X"1F",X"30",X"08",X"D5",X"5E",X"29",X"1D",X"1D",X"19",X"CB",
		X"DC",X"66",X"89",X"A8",X"8F",X"F5",X"46",X"2A",X"DD",X"4E",X"8B",X"89",X"A2",X"AE",X"4A",X"F5",
		X"E6",X"89",X"C2",X"B7",X"A0",X"8C",X"FA",X"C3",X"65",X"7A",X"82",X"84",X"EA",X"C3",X"A2",X"86",
		X"4A",X"37",X"CD",X"5A",X"A2",X"AE",X"4A",X"43",X"92",X"6C",X"96",X"C8",X"B2",X"A8",X"4A",X"3A",
		X"21",X"4A",X"7D",X"56",X"2D",X"5F",X"0F",X"AF",X"0F",X"AB",X"E7",X"16",X"E9",X"CE",X"28",X"67",
		X"ED",X"3E",X"F6",X"E3",X"A1",X"A8",X"4A",X"1B",X"21",X"20",X"88",X"E5",X"B8",X"61",X"B6",X"D6",
		X"69",X"3E",X"28",X"42",X"8E",X"A8",X"A1",X"30",X"29",X"19",X"98",X"72",X"69",X"21",X"00",X"71",
		X"21",X"A8",X"88",X"BE",X"A9",X"19",X"90",X"4A",X"4B",X"4E",X"B6",X"28",X"80",X"2A",X"32",X"1B",
		X"76",X"9C",X"A0",X"8D",X"B4",X"09",X"4B",X"E0",X"6C",X"16",X"D7",X"3A",X"69",X"CD",X"AB",X"CC",
		X"B6",X"28",X"49",X"2E",X"70",X"D5",X"D6",X"2D",X"DE",X"20",X"90",X"3A",X"27",X"0F",X"27",X"C3",
		X"87",X"30",X"2A",X"CB",X"6C",X"CB",X"87",X"30",X"29",X"24",X"56",X"A8",X"E7",X"C9",X"81",X"88",
		X"71",X"35",X"C7",X"3E",X"88",X"29",X"80",X"D1",X"5D",X"FE",X"8D",X"35",X"C7",X"3E",X"88",X"29",
		X"68",X"71",X"7D",X"56",X"2D",X"B5",X"E7",X"36",X"28",X"C9",X"81",X"48",X"D3",X"16",X"09",X"B5",
		X"C7",X"BE",X"AA",X"3E",X"88",X"2B",X"95",X"28",X"72",X"C1",X"ED",X"AA",X"49",X"48",X"D4",X"8F",
		X"AF",X"84",X"AF",X"85",X"AF",X"0F",X"AF",X"0F",X"25",X"1F",X"65",X"42",X"80",X"8B",X"81",X"B4",
		X"D3",X"E5",X"57",X"A5",X"A2",X"49",X"48",X"61",X"49",X"C3",X"D5",X"A8",X"A9",X"FD",X"CD",X"4C",
		X"52",X"55",X"6C",X"16",X"57",X"47",X"F4",X"26",X"28",X"29",X"4D",X"CD",X"A9",X"E6",X"29",X"46",
		X"A0",X"2B",X"A6",X"28",X"49",X"2E",X"00",X"C1",X"26",X"20",X"CD",X"EA",X"D4",X"D2",X"1C",X"6D",
		X"93",X"DA",X"3F",X"6D",X"BB",X"67",X"B7",X"38",X"F1",X"55",X"3F",X"07",X"C9",X"BF",X"FB",X"30",
		X"49",X"BA",X"08",X"48",X"EE",X"29",X"68",X"17",X"7B",X"30",X"92",X"ED",X"40",X"66",X"77",X"3A",
		X"65",X"48",X"FB",X"31",X"C9",X"6F",X"12",X"28",X"E8",X"E6",X"29",X"E8",X"50",X"FB",X"18",X"C9",
		X"5D",X"FE",X"0D",X"2E",X"70",X"76",X"28",X"EF",X"4B",X"4E",X"B6",X"28",X"49",X"28",X"0B",X"2E",
		X"09",X"25",X"38",X"3B",X"3E",X"31",X"1C",X"37",X"22",X"AD",X"01",X"A4",X"07",X"BA",X"35",X"B0",
		X"BB",X"B6",X"49",X"6C",X"4F",X"62",X"CD",X"78",X"5B",X"7E",X"D9",X"74",X"DF",X"EA",X"6C",X"EF",
		X"42",X"E5",X"70",X"FB",X"75",X"F0",X"53",X"F6",X"A8",X"0B",X"AE",X"00",X"8B",X"06",X"B8",X"1B",
		X"15",X"10",X"92",X"15",X"97",X"8A",X"24",X"8F",X"A1",X"83",X"A6",X"98",X"32",X"9C",X"37",X"91",
		X"93",X"95",X"97",X"49",X"EB",X"4D",X"EF",X"41",X"CB",X"45",X"CF",X"58",X"FA",X"5C",X"FE",X"5F",
		X"D1",X"53",X"D4",X"56",X"D7",X"C9",X"62",X"CC",X"65",X"CF",X"E0",X"C1",X"E2",X"C4",X"E5",X"C6",
		X"C7",X"D8",X"F1",X"DA",X"F3",X"DC",X"F5",X"DE",X"F7",X"DF",X"D0",X"D1",X"D1",X"D2",X"D3",X"D3",
		X"F4",X"D4",X"F5",X"D5",X"F5",X"D6",X"F6",X"D6",X"F7",X"D7",X"F7",X"D7",X"F7",X"D5",X"4B",X"28",
		X"46",X"20",X"2D",X"DD",X"36",X"28",X"28",X"C9",X"12",X"A1",X"E8",X"B7",X"EA",X"01",X"6F",X"DD",
		X"46",X"32",X"4B",X"F9",X"6A",X"98",X"4E",X"C3",X"F1",X"42",X"28",X"6E",X"4B",X"E9",X"4A",X"0A",
		X"6F",X"51",X"F6",X"68",X"E6",X"57",X"DD",X"77",X"1A",X"CD",X"EA",X"FA",X"12",X"28",X"EC",X"0F",
		X"90",X"23",X"5D",X"3E",X"9A",X"F8",X"5D",X"3E",X"AC",X"D7",X"6B",X"3D",X"CE",X"D5",X"B6",X"3A",
		X"B8",X"DD",X"96",X"AC",X"29",X"DD",X"96",X"AB",X"28",X"DD",X"96",X"BB",X"2C",X"EB",X"23",X"CE",
		X"4D",X"5F",X"EC",X"D5",X"4B",X"32",X"DE",X"42",X"96",X"6E",X"4D",X"B7",X"D3",X"38",X"8F",X"D5",
		X"6B",X"88",X"86",X"EB",X"02",X"CC",X"7D",X"56",X"08",X"E6",X"29",X"20",X"2F",X"DD",X"F6",X"8F",
		X"DE",X"20",X"90",X"C3",X"4D",X"1D",X"D2",X"C2",X"F7",X"6F",X"59",X"D5",X"E6",X"3A",X"5D",X"EE",
		X"3C",X"DD",X"DE",X"AC",X"79",X"21",X"30",X"4A",X"F6",X"4F",X"6D",X"1C",X"6F",X"51",X"55",X"D5",
		X"4B",X"32",X"C6",X"28",X"95",X"D1",X"DD",X"7C",X"9A",X"F5",X"F5",X"3C",X"DD",X"7A",X"AC",X"F5",
		X"96",X"AB",X"28",X"D5",X"6B",X"BA",X"D6",X"DD",X"F6",X"BB",X"4E",X"8A",X"7D",X"77",X"1B",X"D9",
		X"ED",X"75",X"5D",X"EE",X"8F",X"D5",X"E6",X"20",X"5D",X"FE",X"A9",X"56",X"A8",X"CF",X"F9",X"0E",
		X"14",X"CD",X"C9",X"EE",X"B6",X"29",X"6D",X"95",X"6D",X"E1",X"83",X"F1",X"CF",X"56",X"76",X"77",
		X"4A",X"F7",X"CF",X"CF",X"31",X"A8",X"88",X"10",X"67",X"F5",X"11",X"18",X"74",X"43",X"FD",X"6E",
		X"7D",X"CB",X"1A",X"66",X"B2",X"88",X"EC",X"4F",X"B2",X"8E",X"EC",X"AF",X"4E",X"6C",X"E7",X"16",
		X"CE",X"C6",X"88",X"6F",X"CD",X"DB",X"8F",X"4C",X"92",X"21",X"4C",X"E1",X"10",X"2E",X"10",X"64",
		X"B8",X"EA",X"B8",X"88",X"6B",X"69",X"80",X"82",X"6D",X"DF",X"6F",X"E5",X"4D",X"09",X"7D",X"75",
		X"8F",X"D5",X"F4",X"20",X"4D",X"58",X"D1",X"C3",X"61",X"41",X"E9",X"C2",X"0A",X"6F",X"BF",X"E5",
		X"CA",X"DD",X"D5",X"8F",X"7D",X"74",X"08",X"EB",X"AA",X"CF",X"6D",X"DF",X"6F",X"E5",X"4D",X"B7",
		X"CD",X"4A",X"5D",X"7D",X"0F",X"D5",X"F4",X"20",X"4D",X"8D",X"79",X"C3",X"71",X"41",X"E9",X"C2",
		X"AA",X"6F",X"09",X"DD",X"75",X"2F",X"DD",X"74",X"08",X"EB",X"AA",X"6F",X"DD",X"73",X"2F",X"DD",
		X"F2",X"20",X"82",X"29",X"44",X"CE",X"4B",X"B9",X"29",X"D5",X"C6",X"29",X"5D",X"6E",X"0A",X"CE",
		X"CB",X"11",X"ED",X"F5",X"CD",X"78",X"72",X"F1",X"E9",X"CB",X"66",X"20",X"39",X"39",X"68",X"28",
		X"11",X"C3",X"E6",X"28",X"0F",X"01",X"5D",X"7F",X"89",X"43",X"02",X"6F",X"6E",X"20",X"EE",X"D0",
		X"B9",X"DD",X"77",X"21",X"EB",X"0A",X"6F",X"F5",X"C3",X"C5",X"5B",X"29",X"EC",X"1A",X"4F",X"CB",
		X"91",X"1B",X"12",X"4F",X"5D",X"DE",X"09",X"D5",X"76",X"2A",X"F9",X"01",X"47",X"9A",X"4B",X"BF",
		X"FD",X"5F",X"51",X"BB",X"DD",X"77",X"09",X"F9",X"3B",X"1A",X"A8",X"4F",X"2E",X"28",X"C9",X"CD",
		X"D4",X"FA",X"5D",X"C3",X"9A",X"FE",X"6C",X"8D",X"4F",X"D5",X"D6",X"20",X"EE",X"29",X"5D",X"7F",
		X"08",X"EB",X"A4",X"6B",X"E5",X"AF",X"47",X"26",X"28",X"39",X"54",X"66",X"19",X"56",X"23",X"66",
		X"C7",X"63",X"DD",X"61",X"49",X"D5",X"B5",X"3E",X"68",X"D5",X"B6",X"3E",X"09",X"D5",X"4B",X"3A",
		X"56",X"DD",X"56",X"2E",X"00",X"2C",X"14",X"EB",X"93",X"6F",X"15",X"E6",X"2F",X"DD",X"77",X"2E",
		X"57",X"1E",X"08",X"29",X"6C",X"EF",X"11",X"D5",X"D6",X"28",X"EE",X"D4",X"BE",X"D5",X"F7",X"28",
		X"21",X"E4",X"67",X"19",X"56",X"DD",X"77",X"25",X"C9",X"DD",X"CB",X"28",X"46",X"20",X"2D",X"DD",
		X"4B",X"28",X"B6",X"C1",X"92",X"A1",X"40",X"37",X"6A",X"14",X"C9",X"D5",X"D6",X"32",X"4B",X"6F",
		X"EA",X"48",X"49",X"DD",X"56",X"2E",X"B7",X"EA",X"51",X"62",X"CB",X"57",X"EA",X"8F",X"49",X"CD",
		X"5F",X"64",X"5D",X"FE",X"BA",X"C3",X"77",X"42",X"E1",X"61",X"4B",X"CF",X"6A",X"70",X"EA",X"C3",
		X"FF",X"EA",X"3F",X"E9",X"B2",X"A9",X"EC",X"EE",X"08",X"DD",X"36",X"A9",X"7C",X"6F",X"4A",X"DD",
		X"D6",X"32",X"4B",X"CF",X"6A",X"70",X"EA",X"C3",X"F7",X"42",X"9F",X"61",X"4D",X"C5",X"EA",X"D5",
		X"6B",X"BA",X"76",X"EA",X"3F",X"E9",X"7D",X"34",X"3F",X"EA",X"5B",X"E9",X"7D",X"56",X"3A",X"C5",
		X"64",X"D5",X"F7",X"30",X"5D",X"3E",X"AB",X"28",X"5D",X"3E",X"98",X"28",X"DA",X"7E",X"E8",X"D5",
		X"96",X"AC",X"08",X"EB",X"5A",X"E8",X"7D",X"36",X"0C",X"70",X"7D",X"56",X"1A",X"F6",X"48",X"DD",
		X"F7",X"32",X"6B",X"3F",X"E9",X"D5",X"4B",X"28",X"E6",X"28",X"8D",X"D5",X"4B",X"28",X"36",X"C1",
		X"B2",X"A1",X"E8",X"B7",X"4A",X"3C",X"49",X"DD",X"F6",X"BA",X"6B",X"67",X"4A",X"48",X"49",X"CB",
		X"D7",X"42",X"07",X"61",X"5D",X"FE",X"8E",X"37",X"6A",X"F1",X"EA",X"C5",X"5F",X"64",X"5D",X"FE",
		X"1A",X"CB",X"DF",X"EA",X"41",X"E9",X"6B",X"4F",X"4A",X"F8",X"4A",X"CB",X"FF",X"EA",X"3F",X"E9",
		X"92",X"21",X"4C",X"46",X"A8",X"D5",X"9E",X"21",X"5C",X"47",X"EA",X"D5",X"4B",X"32",X"EE",X"42",
		X"58",X"EA",X"4B",X"8F",X"49",X"DD",X"6B",X"88",X"46",X"20",X"2D",X"DD",X"6B",X"88",X"96",X"C9",
		X"92",X"A1",X"48",X"37",X"6A",X"14",X"E9",X"D5",X"D6",X"32",X"4B",X"6F",X"6A",X"48",X"E9",X"C3",
		X"F7",X"EA",X"A7",X"E9",X"7D",X"56",X"2E",X"B7",X"4A",X"F1",X"4A",X"CD",X"FF",X"EC",X"7D",X"56",
		X"BA",X"C3",X"77",X"42",X"E1",X"61",X"4B",X"CF",X"6A",X"70",X"EA",X"C3",X"57",X"42",X"9F",X"61",
		X"B2",X"A9",X"EC",X"EE",X"08",X"DD",X"36",X"A9",X"7C",X"6F",X"4A",X"DD",X"F6",X"BA",X"6B",X"4F",
		X"6A",X"70",X"CA",X"C3",X"67",X"A8",X"89",X"D5",X"4B",X"32",X"7E",X"28",X"8A",X"C5",X"E5",X"62",
		X"DD",X"CB",X"1A",X"FE",X"CA",X"73",X"49",X"CD",X"17",X"FB",X"30",X"B1",X"DD",X"CB",X"1A",X"76",
		X"A0",X"2F",X"5D",X"C3",X"9A",X"9E",X"6B",X"7D",X"C9",X"29",X"84",X"EF",X"06",X"2C",X"26",X"22",
		X"87",X"CD",X"30",X"FC",X"10",X"27",X"D6",X"2B",X"20",X"33",X"16",X"29",X"DD",X"86",X"28",X"DD",
		X"F7",X"28",X"6B",X"7D",X"C9",X"D5",X"4B",X"32",X"96",X"D5",X"D6",X"30",X"5D",X"7F",X"8B",X"0F",
		X"30",X"2B",X"DD",X"35",X"3A",X"DD",X"CB",X"32",X"5E",X"20",X"10",X"21",X"74",X"EF",X"0E",X"2F",
		X"26",X"2A",X"8F",X"C5",X"38",X"FC",X"6B",X"0A",X"C9",X"D5",X"4B",X"3C",X"FE",X"A8",X"8B",X"D5",
		X"36",X"29",X"6A",X"DD",X"36",X"2A",X"40",X"EB",X"AA",X"61",X"DD",X"36",X"29",X"63",X"DD",X"36",
		X"0A",X"E0",X"5D",X"C3",X"1A",X"F6",X"80",X"2F",X"5D",X"C3",X"08",X"4E",X"6B",X"1B",X"C9",X"D5",
		X"CB",X"28",X"AE",X"DD",X"34",X"33",X"CC",X"8A",X"4C",X"CD",X"DC",X"FA",X"DD",X"56",X"08",X"E6",
		X"09",X"D5",X"F7",X"20",X"6B",X"52",X"DE",X"D5",X"B6",X"32",X"58",X"AA",X"16",X"EF",X"5D",X"7D",
		X"29",X"DD",X"74",X"2A",X"DD",X"36",X"38",X"28",X"DD",X"36",X"39",X"28",X"DD",X"36",X"3E",X"29",
		X"5D",X"C3",X"9A",X"FE",X"80",X"ED",X"A1",X"1E",X"6F",X"0E",X"0A",X"8E",X"88",X"D5",X"D6",X"38",
		X"08",X"DD",X"56",X"3A",X"B7",X"D2",X"D9",X"61",X"87",X"CD",X"30",X"FC",X"08",X"DD",X"96",X"38",
		X"80",X"A9",X"5D",X"FE",X"19",X"DF",X"94",X"D5",X"4B",X"3A",X"FE",X"A8",X"0A",X"BD",X"95",X"66",
		X"2F",X"DD",X"77",X"39",X"21",X"EC",X"67",X"3E",X"28",X"19",X"DD",X"56",X"28",X"E6",X"D4",X"B6",
		X"5D",X"7F",X"88",X"C5",X"5F",X"64",X"5D",X"C3",X"BA",X"7E",X"6A",X"1B",X"E9",X"C5",X"B7",X"FB",
		X"5A",X"1B",X"49",X"DD",X"6B",X"BA",X"B6",X"DD",X"96",X"98",X"28",X"DD",X"96",X"9E",X"29",X"DD",
		X"D6",X"28",X"EE",X"D4",X"5D",X"7F",X"88",X"D5",X"B6",X"3C",X"74",X"29",X"06",X"EF",X"06",X"2B",
		X"8E",X"AA",X"27",X"CD",X"30",X"D4",X"5A",X"1B",X"49",X"DD",X"6B",X"88",X"86",X"CD",X"02",X"CC",
		X"5D",X"FE",X"8F",X"C3",X"47",X"40",X"5D",X"C3",X"A8",X"6E",X"80",X"2E",X"DE",X"78",X"58",X"43",
		X"10",X"EF",X"76",X"10",X"58",X"EB",X"10",X"EF",X"81",X"0A",X"67",X"2E",X"2D",X"0E",X"2C",X"87",
		X"4D",X"B8",X"D4",X"52",X"3C",X"61",X"5D",X"FE",X"B8",X"D5",X"F7",X"3A",X"5D",X"FE",X"B9",X"D5",
		X"D7",X"9C",X"7D",X"CB",X"1A",X"2E",X"4B",X"3C",X"49",X"DD",X"F6",X"98",X"17",X"20",X"24",X"DD",
		X"B5",X"3E",X"6A",X"14",X"E9",X"D5",X"D6",X"39",X"DE",X"2C",X"80",X"3B",X"94",X"D5",X"F7",X"39",
		X"7D",X"36",X"3E",X"8C",X"B6",X"89",X"7D",X"86",X"28",X"DD",X"D7",X"88",X"4B",X"3C",X"49",X"DD",
		X"B6",X"3E",X"89",X"29",X"24",X"EF",X"26",X"2E",X"06",X"2C",X"8F",X"C5",X"90",X"FC",X"7A",X"14",
		X"49",X"DD",X"96",X"8E",X"28",X"DD",X"96",X"98",X"2A",X"DD",X"96",X"9E",X"29",X"DD",X"96",X"BA",
		X"E8",X"29",X"2C",X"EF",X"26",X"3C",X"06",X"2C",X"8F",X"C5",X"90",X"FC",X"6B",X"14",X"E9",X"88",
		X"46",X"C0",X"8F",X"2F",X"8F",X"DD",X"6B",X"9A",X"56",X"00",X"09",X"D6",X"29",X"E8",X"81",X"94",
		X"EE",X"43",X"A8",X"64",X"DE",X"2A",X"68",X"29",X"64",X"65",X"6B",X"20",X"EC",X"BA",X"A9",X"4C",
		X"4E",X"A8",X"7D",X"4E",X"09",X"91",X"7A",X"0A",X"4B",X"FE",X"38",X"91",X"5A",X"0A",X"4B",X"02",
		X"0F",X"4C",X"5D",X"DE",X"0F",X"D5",X"76",X"20",X"BF",X"E5",X"72",X"D5",X"D6",X"3A",X"90",X"39",
		X"B7",X"F2",X"5A",X"63",X"4F",X"CD",X"E6",X"63",X"51",X"E8",X"DD",X"36",X"0C",X"20",X"EB",X"B2",
		X"CB",X"37",X"DA",X"E0",X"CB",X"CF",X"D4",X"AF",X"E7",X"FD",X"87",X"EF",X"A3",X"E5",X"53",X"2F",
		X"EC",X"CD",X"E6",X"63",X"51",X"E8",X"DD",X"36",X"0C",X"D0",X"C5",X"6C",X"DD",X"77",X"18",X"DD",
		X"4B",X"32",X"D6",X"D5",X"4B",X"32",X"76",X"D5",X"B6",X"38",X"08",X"D5",X"B6",X"23",X"08",X"29",
		X"8C",X"EF",X"2E",X"3C",X"0E",X"2B",X"87",X"EB",X"30",X"FC",X"DD",X"CB",X"1A",X"6E",X"C8",X"CD",
		X"66",X"63",X"A0",X"AB",X"8F",X"43",X"5E",X"64",X"5D",X"C3",X"9A",X"6E",X"48",X"FC",X"87",X"6F",
		X"55",X"07",X"47",X"23",X"C5",X"5B",X"2F",X"4C",X"CD",X"CE",X"4B",X"20",X"0A",X"F6",X"D7",X"EB",
		X"5E",X"64",X"5D",X"C3",X"9A",X"6E",X"48",X"D5",X"B6",X"38",X"08",X"29",X"02",X"EF",X"26",X"3C",
		X"0E",X"2C",X"87",X"CD",X"30",X"FC",X"DD",X"56",X"1A",X"CB",X"77",X"20",X"2E",X"DD",X"4E",X"3A",
		X"5D",X"79",X"8B",X"76",X"4A",X"D5",X"F7",X"32",X"92",X"3C",X"40",X"5F",X"D1",X"37",X"DA",X"95",
		X"4B",X"1E",X"24",X"52",X"D6",X"30",X"10",X"26",X"1E",X"34",X"EB",X"4E",X"4B",X"1E",X"DC",X"52",
		X"DE",X"30",X"90",X"2A",X"16",X"CC",X"5D",X"7B",X"98",X"D5",X"B6",X"31",X"F0",X"D5",X"B6",X"3C",
		X"28",X"DD",X"36",X"3A",X"28",X"91",X"E2",X"52",X"4B",X"17",X"30",X"2D",X"DD",X"36",X"0C",X"29",
		X"49",X"D5",X"B6",X"24",X"F7",X"C1",X"4B",X"BC",X"4B",X"9D",X"4B",X"BC",X"4B",X"9D",X"4B",X"BC",
		X"CB",X"1D",X"CB",X"14",X"CB",X"1D",X"6D",X"12",X"09",X"4C",X"ED",X"CD",X"78",X"FA",X"E9",X"CB",
		X"E6",X"40",X"A3",X"2B",X"30",X"D1",X"8F",X"C1",X"ED",X"29",X"0A",X"EF",X"26",X"3C",X"06",X"2C",
		X"27",X"DD",X"96",X"98",X"28",X"CD",X"30",X"D4",X"41",X"DD",X"F6",X"BA",X"6B",X"77",X"80",X"8E",
		X"5D",X"CE",X"9A",X"D5",X"F1",X"23",X"FE",X"6A",X"5D",X"7F",X"BA",X"BA",X"9C",X"48",X"2F",X"BC",
		X"FF",X"3E",X"28",X"19",X"F6",X"03",X"7D",X"77",X"19",X"56",X"7D",X"77",X"18",X"DD",X"96",X"9C",
		X"88",X"D5",X"B6",X"3A",X"88",X"B1",X"EA",X"62",X"EC",X"BF",X"B0",X"2D",X"5D",X"3E",X"AC",X"29",
		X"69",X"DD",X"96",X"AC",X"D7",X"C9",X"55",X"DD",X"96",X"98",X"28",X"21",X"AA",X"C7",X"8E",X"9C",
		X"06",X"2C",X"8F",X"C5",X"90",X"FC",X"5D",X"FE",X"BA",X"C3",X"F7",X"28",X"8E",X"D5",X"46",X"3A",
		X"7D",X"71",X"0B",X"F6",X"6A",X"DD",X"D7",X"BA",X"51",X"20",X"2D",X"16",X"30",X"EB",X"AA",X"EC",
		X"96",X"58",X"5D",X"7F",X"B8",X"D5",X"B6",X"31",X"50",X"D5",X"B6",X"3C",X"88",X"D5",X"B6",X"3A",
		X"28",X"91",X"42",X"1E",X"4C",X"17",X"90",X"8D",X"7D",X"36",X"0C",X"89",X"69",X"DD",X"96",X"AC",
		X"77",X"C1",X"92",X"2C",X"48",X"DF",X"92",X"20",X"48",X"F6",X"80",X"B8",X"8A",X"BE",X"BF",X"66",
		X"1C",X"EE",X"E8",X"DD",X"D7",X"BB",X"7D",X"56",X"3A",X"B7",X"52",X"6A",X"4C",X"15",X"76",X"10",
		X"78",X"C3",X"F3",X"A8",X"89",X"BD",X"5D",X"7F",X"9A",X"C1",X"94",X"F6",X"D8",X"50",X"4B",X"7B",
		X"A0",X"89",X"B4",X"DD",X"D7",X"9A",X"69",X"DD",X"F6",X"9A",X"6B",X"57",X"80",X"A9",X"17",X"20",
		X"D8",X"D5",X"4B",X"28",X"CE",X"A8",X"EA",X"D5",X"4B",X"3C",X"F6",X"A8",X"9E",X"3F",X"4D",X"FA",
		X"71",X"87",X"A8",X"51",X"17",X"CA",X"94",X"ED",X"46",X"AC",X"6A",X"10",X"4D",X"CD",X"BE",X"ED",
		X"6B",X"94",X"CD",X"C5",X"25",X"F9",X"ED",X"19",X"40",X"D7",X"11",X"FE",X"E9",X"88",X"D1",X"37",
		X"CA",X"94",X"4D",X"CB",X"7F",X"CA",X"65",X"65",X"E6",X"29",X"20",X"2E",X"CD",X"1E",X"4D",X"EB",
		X"B4",X"65",X"4D",X"4D",X"CD",X"C5",X"16",X"65",X"5D",X"FE",X"9A",X"66",X"F2",X"D5",X"F7",X"32",
		X"C9",X"DD",X"CB",X"3C",X"56",X"EA",X"A9",X"65",X"CD",X"58",X"71",X"E5",X"39",X"48",X"D7",X"19",
		X"D6",X"61",X"00",X"F9",X"BF",X"C2",X"B4",X"65",X"4B",X"4F",X"80",X"31",X"EE",X"2C",X"A0",X"2E",
		X"CD",X"1E",X"4D",X"EB",X"94",X"65",X"CD",X"4D",X"4D",X"CD",X"BE",X"65",X"DD",X"56",X"1A",X"E6",
		X"F2",X"D5",X"F7",X"32",X"49",X"D5",X"4B",X"32",X"16",X"D5",X"4B",X"32",X"06",X"66",X"0A",X"42",
		X"ED",X"65",X"DD",X"CB",X"1A",X"FE",X"EA",X"4D",X"4D",X"CD",X"ED",X"65",X"DD",X"CB",X"1A",X"4E",
		X"49",X"3F",X"4D",X"D5",X"79",X"A7",X"00",X"F9",X"BF",X"C2",X"B4",X"65",X"EE",X"2B",X"80",X"A8",
		X"CD",X"1E",X"4D",X"EB",X"94",X"65",X"DD",X"56",X"3A",X"C5",X"6C",X"DD",X"77",X"3A",X"DD",X"56",
		X"8B",X"E5",X"64",X"D5",X"F7",X"23",X"5D",X"FE",X"8C",X"E5",X"64",X"D5",X"F7",X"24",X"BF",X"C1",
		X"DD",X"56",X"3C",X"B7",X"F2",X"94",X"4D",X"C5",X"6C",X"DD",X"77",X"3C",X"CD",X"92",X"73",X"DD",
		X"4B",X"32",X"56",X"37",X"49",X"D5",X"56",X"29",X"5D",X"5E",X"0A",X"9A",X"4B",X"BF",X"67",X"19",
		X"28",X"C8",X"B7",X"C5",X"7A",X"55",X"0F",X"0F",X"0F",X"E6",X"18",X"47",X"54",X"0F",X"0F",X"0F",
		X"EE",X"C8",X"BD",X"10",X"5D",X"7F",X"89",X"D5",X"B6",X"3C",X"08",X"C1",X"38",X"50",X"AD",X"57",
		X"18",X"50",X"18",X"5C",X"20",X"50",X"20",X"54",X"18",X"5E",X"18",X"5C",X"2E",X"52",X"3F",X"52",
		X"9A",X"50",X"BC",X"50",X"B8",X"56",X"B8",X"50",X"90",X"50",X"AC",X"50",X"98",X"5E",X"A8",X"5E",
		X"18",X"7B",X"0C",X"7C",X"00",X"78",X"3C",X"5C",X"3C",X"78",X"1A",X"78",X"3E",X"5C",X"20",X"7C",
		X"B8",X"5A",X"98",X"5A",X"80",X"5C",X"9C",X"5C",X"9E",X"5C",X"AC",X"5C",X"A0",X"48",X"B8",X"5E",
		X"0C",X"5A",X"18",X"5A",X"F8",X"78",X"E0",X"7F",X"C0",X"78",X"C0",X"5C",X"E0",X"78",X"E0",X"7C",
		X"60",X"5E",X"44",X"54",X"72",X"52",X"61",X"52",X"66",X"50",X"40",X"50",X"60",X"56",X"60",X"50",
		X"F8",X"78",X"F4",X"78",X"F0",X"5E",X"D0",X"5E",X"C0",X"78",X"F0",X"7C",X"D8",X"78",X"C4",X"5C",
		X"64",X"50",X"46",X"50",X"62",X"5C",X"40",X"54",X"60",X"5A",X"50",X"5A",X"40",X"5C",X"64",X"5C",
		X"C2",X"5C",X"F4",X"5C",X"D8",X"5C",X"C0",X"5E",X"F4",X"5A",X"C0",X"5A",X"28",X"4B",X"20",X"4B",
		X"C8",X"4B",X"C0",X"4B",X"08",X"4B",X"00",X"4B",X"48",X"4B",X"40",X"4B",X"88",X"4C",X"80",X"4C",
		X"68",X"4C",X"60",X"4C",X"A8",X"4C",X"A0",X"4C",X"E8",X"4C",X"E0",X"4C",X"28",X"4D",X"20",X"4D",
		X"C8",X"4D",X"C0",X"4D",X"08",X"4D",X"00",X"4D",X"48",X"4D",X"40",X"4D",X"88",X"4E",X"80",X"4E",
		X"68",X"4E",X"60",X"4E",X"A8",X"4E",X"A0",X"4E",X"E8",X"4E",X"E0",X"4E",X"B6",X"77",X"92",X"C6",
		X"48",X"C5",X"00",X"F1",X"8F",X"3A",X"C6",X"48",X"49",X"56",X"8D",X"D0",X"FD",X"65",X"6D",X"29",
		X"A0",X"4D",X"99",X"08",X"ED",X"2E",X"28",X"16",X"2B",X"0E",X"0C",X"C5",X"10",X"0E",X"3C",X"09",
		X"CB",X"89",X"CB",X"BD",X"A0",X"DB",X"69",X"61",X"F9",X"E3",X"A1",X"CE",X"4D",X"3E",X"76",X"2B",
		X"D3",X"23",X"D2",X"23",X"D1",X"23",X"4E",X"8D",X"D7",X"23",X"D0",X"FE",X"2D",X"21",X"E0",X"4D",
		X"B6",X"98",X"A3",X"E3",X"2F",X"CF",X"26",X"28",X"A1",X"65",X"58",X"89",X"CD",X"20",X"CD",X"20",
		X"21",X"0D",X"ED",X"39",X"20",X"28",X"2E",X"2B",X"35",X"19",X"38",X"D4",X"C9",X"DD",X"34",X"2E",
		X"A0",X"2E",X"5D",X"FE",X"8A",X"C5",X"85",X"3F",X"5D",X"FE",X"0E",X"D5",X"9E",X"23",X"6A",X"8C",
		X"6B",X"DD",X"36",X"28",X"28",X"EB",X"02",X"6C",X"21",X"E8",X"ED",X"39",X"68",X"4D",X"29",X"A8",
		X"08",X"E5",X"B8",X"29",X"4D",X"4D",X"B5",X"D5",X"ED",X"29",X"68",X"4D",X"B6",X"98",X"A1",X"EF",
		X"ED",X"DD",X"5E",X"2F",X"73",X"DD",X"7E",X"20",X"23",X"72",X"DD",X"56",X"09",X"DD",X"21",X"E8",
		X"45",X"65",X"4D",X"44",X"7B",X"61",X"A3",X"BD",X"F7",X"2B",X"B6",X"28",X"5D",X"61",X"49",X"D5",
		X"CB",X"28",X"46",X"20",X"2F",X"DD",X"36",X"28",X"28",X"EB",X"02",X"6C",X"DD",X"35",X"0A",X"CA",
		X"7D",X"67",X"5D",X"FE",X"0D",X"07",X"2F",X"07",X"C7",X"2E",X"08",X"A9",X"31",X"29",X"47",X"99",
		X"C3",X"DD",X"56",X"38",X"14",X"D6",X"0A",X"10",X"29",X"87",X"DD",X"77",X"38",X"AF",X"EE",X"58",
		X"C7",X"BE",X"CF",X"C6",X"08",X"6F",X"D6",X"2B",X"E6",X"EF",X"21",X"22",X"08",X"E5",X"B8",X"43",
		X"A4",X"6B",X"28",X"9F",X"4F",X"E7",X"4F",X"2D",X"2D",X"3C",X"28",X"48",X"4F",X"29",X"E8",X"24",
		X"08",X"D7",X"77",X"DE",X"E6",X"9F",X"B7",X"87",X"B6",X"C7",X"08",X"28",X"08",X"28",X"08",X"28",
		X"E4",X"67",X"C6",X"67",X"D0",X"67",X"2A",X"78",X"0C",X"78",X"3E",X"78",X"20",X"78",X"02",X"78",
		X"3C",X"78",X"BE",X"78",X"E0",X"C5",X"F6",X"48",X"B6",X"C0",X"F7",X"D7",X"B4",X"95",X"E7",X"57",
		X"C0",X"C5",X"D6",X"48",X"C0",X"C4",X"E4",X"CD",X"D0",X"1F",X"C7",X"57",X"C0",X"C5",X"F7",X"C6",
		X"D7",X"65",X"47",X"6F",X"50",X"17",X"47",X"D7",X"50",X"65",X"50",X"65",X"E7",X"0F",X"47",X"6F",
		X"D0",X"1F",X"C7",X"D7",X"C7",X"C6",X"57",X"2E",X"EF",X"2F",X"C7",X"EF",X"EF",X"D7",X"A7",X"BE",
		X"56",X"17",X"5F",X"0E",X"E7",X"0F",X"5F",X"3E",X"87",X"AF",X"50",X"E5",X"56",X"17",X"5F",X"0E",
		X"57",X"96",X"95",X"C4",X"96",X"C0",X"D0",X"C5",X"D6",X"1F",X"DF",X"96",X"C6",X"86",X"D6",X"48",
		X"16",X"E0",X"50",X"E5",X"47",X"67",X"97",X"37",X"A8",X"69",X"F8",X"9D",X"6F",X"69",X"F8",X"EA",
		X"78",X"FB",X"78",X"F4",X"78",X"0D",X"78",X"06",X"78",X"1F",X"78",X"88",X"78",X"81",X"78",X"9A",
		X"F8",X"89",X"29",X"C8",X"A8",X"B3",X"F8",X"09",X"E8",X"88",X"29",X"8A",X"F8",X"08",X"13",X"58",
		X"29",X"19",X"20",X"21",X"22",X"78",X"28",X"93",X"78",X"29",X"C3",X"20",X"21",X"22",X"78",X"28",
		X"13",X"58",X"A9",X"4D",X"29",X"89",X"2A",X"58",X"A8",X"B3",X"F8",X"09",X"1F",X"89",X"29",X"8A",
		X"78",X"28",X"93",X"78",X"29",X"D1",X"21",X"21",X"23",X"70",X"28",X"93",X"78",X"29",X"7B",X"22",
		X"29",X"8C",X"E0",X"08",X"13",X"58",X"A9",X"36",X"2A",X"89",X"2C",X"68",X"A8",X"B3",X"F8",X"09",
		X"AA",X"23",X"21",X"24",X"E8",X"28",X"93",X"78",X"29",X"06",X"23",X"28",X"28",X"28",X"B7",X"28",
		X"A8",X"08",X"A8",X"08",X"A8",X"08",X"37",X"08",X"50",X"F0",X"A8",X"36",X"9B",X"4D",X"B5",X"4D",
		X"DD",X"B6",X"28",X"98",X"DD",X"B6",X"25",X"28",X"DD",X"B6",X"3E",X"28",X"DD",X"B6",X"2E",X"28",
		X"5D",X"B6",X"B8",X"08",X"5D",X"F5",X"AF",X"74",X"EE",X"09",X"E7",X"5D",X"F4",X"88",X"5D",X"F1",
		X"21",X"45",X"5B",X"2F",X"4C",X"43",X"B7",X"45",X"7A",X"5A",X"6D",X"79",X"CB",X"34",X"CB",X"3D",
		X"92",X"89",X"44",X"99",X"5A",X"2C",X"59",X"15",X"B0",X"8D",X"4D",X"A0",X"59",X"5D",X"F7",X"1C",
		X"DD",X"B6",X"3A",X"68",X"EB",X"13",X"1A",X"4D",X"98",X"79",X"DD",X"F7",X"3A",X"5D",X"36",X"3C",
		X"28",X"CB",X"93",X"9A",X"CD",X"EC",X"9D",X"B0",X"8F",X"4D",X"A0",X"59",X"CD",X"EC",X"5D",X"F7",
		X"3C",X"5D",X"36",X"3A",X"68",X"6B",X"9B",X"32",X"CD",X"10",X"79",X"5D",X"77",X"3A",X"DD",X"B6",
		X"1C",X"60",X"6B",X"93",X"9A",X"74",X"87",X"E7",X"D5",X"27",X"C7",X"A3",X"4B",X"34",X"4B",X"3D",
		X"12",X"21",X"EC",X"39",X"10",X"37",X"95",X"B0",X"0D",X"4D",X"80",X"79",X"DD",X"F7",X"3C",X"5D",
		X"B6",X"1A",X"40",X"CB",X"93",X"9A",X"4D",X"90",X"59",X"45",X"64",X"5D",X"F7",X"1A",X"5D",X"B6",
		X"3C",X"A8",X"EB",X"13",X"1A",X"CD",X"6C",X"9D",X"30",X"27",X"CD",X"80",X"79",X"CD",X"6C",X"5D",
		X"F7",X"1C",X"5D",X"B6",X"1A",X"40",X"6B",X"93",X"9A",X"4D",X"90",X"59",X"CD",X"EC",X"5D",X"F7",
		X"3A",X"5D",X"36",X"3C",X"E0",X"6B",X"9B",X"32",X"5F",X"D5",X"E6",X"D4",X"0F",X"07",X"67",X"D5",
		X"EE",X"0B",X"07",X"2F",X"C7",X"CB",X"88",X"4D",X"55",X"67",X"EE",X"F0",X"07",X"2F",X"07",X"E7",
		X"55",X"EE",X"2F",X"07",X"0F",X"07",X"47",X"6B",X"08",X"6D",X"12",X"A1",X"E8",X"47",X"DD",X"4B",
		X"9A",X"6E",X"6A",X"5D",X"5A",X"5D",X"D6",X"1E",X"94",X"C6",X"0F",X"5D",X"F7",X"1E",X"67",X"A0",
		X"20",X"05",X"0C",X"A0",X"1C",X"5D",X"56",X"2E",X"D6",X"2A",X"30",X"2C",X"14",X"5D",X"77",X"2E",
		X"A1",X"6D",X"5A",X"BE",X"08",X"8F",X"57",X"39",X"D6",X"5D",X"F7",X"09",X"A3",X"76",X"5D",X"F7",
		X"2A",X"5D",X"56",X"28",X"E6",X"D4",X"5F",X"D0",X"E6",X"2A",X"7F",X"07",X"B2",X"BB",X"DD",X"F7",
		X"A8",X"5D",X"D6",X"0E",X"BF",X"20",X"AE",X"70",X"EE",X"09",X"5D",X"F7",X"2D",X"2C",X"05",X"A0",
		X"AA",X"4D",X"54",X"FA",X"DD",X"76",X"21",X"56",X"30",X"30",X"AB",X"56",X"40",X"B0",X"37",X"5D",
		X"D6",X"0F",X"5D",X"4B",X"28",X"4E",X"80",X"0F",X"DE",X"F0",X"B0",X"1A",X"6B",X"3B",X"FA",X"56",
		X"38",X"30",X"23",X"5D",X"56",X"20",X"E6",X"29",X"DD",X"F7",X"20",X"CB",X"8C",X"6B",X"DD",X"4B",
		X"3A",X"66",X"5D",X"B6",X"BA",X"08",X"5D",X"B6",X"BC",X"08",X"5D",X"B6",X"B8",X"0D",X"5D",X"B6",
		X"3E",X"2C",X"EB",X"BB",X"7A",X"5D",X"CB",X"32",X"8E",X"5D",X"36",X"28",X"28",X"CB",X"A2",X"6C",
		X"A8",X"EB",X"FA",X"B2",X"F9",X"EB",X"FA",X"7C",X"FA",X"FF",X"FA",X"28",X"B8",X"70",X"A9",X"82",
		X"7A",X"29",X"A5",X"BE",X"3A",X"21",X"11",X"28",X"02",X"7A",X"2A",X"A5",X"B0",X"47",X"B0",X"30",
		X"2C",X"1C",X"A9",X"82",X"FA",X"0A",X"F1",X"B9",X"99",X"BA",X"A8",X"F7",X"C7",X"57",X"AF",X"0D",
		X"0C",X"CD",X"AF",X"BF",X"3F",X"2D",X"97",X"F7",X"B7",X"28",X"DD",X"76",X"2D",X"56",X"2A",X"20",
		X"B9",X"22",X"AF",X"43",X"31",X"A8",X"A8",X"39",X"92",X"89",X"CB",X"5D",X"4B",X"08",X"CE",X"CB",
		X"94",X"7A",X"02",X"AF",X"4B",X"B9",X"50",X"D7",X"19",X"32",X"A1",X"4B",X"DD",X"F5",X"2F",X"5D",
		X"F4",X"88",X"CB",X"4D",X"4C",X"7B",X"5D",X"F7",X"29",X"CB",X"1B",X"9A",X"92",X"43",X"C8",X"56",
		X"2A",X"A0",X"2E",X"32",X"3F",X"4B",X"EB",X"54",X"7A",X"32",X"BF",X"4B",X"4F",X"8F",X"5F",X"BE",
		X"A8",X"A1",X"52",X"5A",X"11",X"76",X"5D",X"F7",X"A9",X"A3",X"D6",X"5D",X"F7",X"0A",X"A1",X"0C",
		X"7B",X"79",X"19",X"76",X"DD",X"F7",X"21",X"CB",X"8C",X"6B",X"4C",X"EF",X"93",X"EF",X"93",X"EF",
		X"5C",X"E8",X"5C",X"E8",X"46",X"45",X"43",X"42",X"40",X"30",X"44",X"6F",X"C4",X"5A",X"5D",X"4B",
		X"28",X"E6",X"20",X"2D",X"DD",X"4B",X"28",X"96",X"C9",X"92",X"01",X"48",X"B7",X"6A",X"38",X"71",
		X"5D",X"76",X"9A",X"4B",X"E7",X"CA",X"9C",X"D8",X"4B",X"77",X"6A",X"8C",X"D8",X"4B",X"57",X"CA",
		X"41",X"70",X"CB",X"67",X"EA",X"51",X"58",X"5D",X"56",X"2E",X"CB",X"D7",X"CA",X"57",X"7B",X"4B",
		X"F7",X"20",X"58",X"4B",X"C7",X"A0",X"2E",X"97",X"4D",X"7A",X"79",X"C5",X"31",X"48",X"08",X"39",
		X"CD",X"01",X"72",X"D6",X"E1",X"00",X"51",X"EE",X"0C",X"6A",X"50",X"7D",X"51",X"EE",X"2A",X"4A",
		X"8E",X"5E",X"00",X"AF",X"5A",X"D4",X"5C",X"4D",X"2B",X"D9",X"6B",X"8D",X"D9",X"97",X"4D",X"F5",
		X"71",X"ED",X"39",X"68",X"28",X"11",X"CD",X"F5",X"72",X"D6",X"E1",X"00",X"51",X"EE",X"2B",X"6A",
		X"42",X"5D",X"D1",X"C6",X"0C",X"4A",X"D8",X"5E",X"00",X"AF",X"5A",X"1C",X"5D",X"4D",X"2B",X"D9",
		X"EB",X"25",X"59",X"4B",X"47",X"A0",X"24",X"4D",X"A5",X"F9",X"E5",X"31",X"E8",X"D7",X"19",X"4D",
		X"81",X"7A",X"D6",X"C1",X"00",X"4B",X"71",X"CA",X"E0",X"5D",X"D1",X"C6",X"0A",X"4A",X"FE",X"5E",
		X"08",X"27",X"DA",X"DF",X"7C",X"4D",X"23",X"71",X"EB",X"25",X"59",X"4D",X"F8",X"F9",X"E5",X"31",
		X"40",X"F7",X"11",X"4D",X"FD",X"7A",X"D6",X"C1",X"00",X"4B",X"61",X"CA",X"94",X"5D",X"D1",X"C6",
		X"2A",X"4A",X"34",X"7E",X"08",X"27",X"DA",X"B9",X"7D",X"4D",X"23",X"71",X"EB",X"25",X"59",X"4B",
		X"F7",X"20",X"FD",X"4B",X"C7",X"A0",X"BB",X"97",X"4D",X"7A",X"79",X"5D",X"4B",X"9A",X"CE",X"A0",
		X"39",X"4B",X"69",X"6A",X"A4",X"7E",X"51",X"EE",X"2A",X"4A",X"1A",X"7F",X"CD",X"AB",X"59",X"6B",
		X"2D",X"D9",X"96",X"09",X"5D",X"06",X"A8",X"5D",X"F7",X"08",X"4B",X"E9",X"4A",X"8D",X"79",X"4D",
		X"66",X"7D",X"CD",X"C6",X"71",X"DE",X"2A",X"5D",X"77",X"21",X"DD",X"76",X"2E",X"D6",X"C8",X"CB",
		X"DE",X"5F",X"BF",X"4D",X"55",X"79",X"5D",X"4B",X"3A",X"CE",X"6A",X"BE",X"FC",X"4B",X"51",X"CA",
		X"56",X"7E",X"51",X"C6",X"2C",X"4A",X"74",X"7F",X"CD",X"AB",X"71",X"CB",X"25",X"71",X"16",X"29",
		X"5D",X"06",X"A8",X"5D",X"F7",X"08",X"4B",X"79",X"4A",X"8D",X"79",X"4D",X"6E",X"5D",X"4D",X"E6",
		X"71",X"DE",X"2A",X"5D",X"77",X"21",X"DD",X"76",X"2E",X"D6",X"48",X"C6",X"57",X"CB",X"DA",X"7F",
		X"4B",X"67",X"A0",X"BC",X"4D",X"25",X"F1",X"5D",X"4B",X"9A",X"6E",X"CA",X"77",X"5C",X"4B",X"E9",
		X"EA",X"D4",X"7E",X"71",X"E6",X"2A",X"CA",X"F6",X"7F",X"4D",X"AB",X"71",X"EB",X"25",X"71",X"36",
		X"A9",X"5D",X"8E",X"08",X"5D",X"F7",X"A8",X"4B",X"61",X"4A",X"2D",X"D9",X"4D",X"CE",X"FD",X"4D",
		X"56",X"71",X"14",X"5D",X"77",X"21",X"DD",X"76",X"2E",X"D6",X"88",X"C6",X"97",X"CB",X"DA",X"7F",
		X"4D",X"50",X"F1",X"5D",X"4B",X"9A",X"6E",X"CA",X"13",X"5C",X"4B",X"F9",X"6A",X"40",X"FE",X"71",
		X"E6",X"2A",X"CA",X"B4",X"7F",X"4D",X"AB",X"71",X"EB",X"25",X"71",X"36",X"29",X"5D",X"86",X"28",
		X"5D",X"F7",X"A8",X"4B",X"71",X"4A",X"2D",X"D9",X"4D",X"CE",X"FD",X"4D",X"5E",X"D9",X"94",X"5D",
		X"77",X"21",X"DD",X"76",X"2E",X"D6",X"08",X"C6",X"17",X"CB",X"5E",X"7F",X"CD",X"66",X"7D",X"4D",
		X"AD",X"DA",X"31",X"F2",X"57",X"39",X"5D",X"F5",X"AF",X"74",X"EE",X"09",X"5D",X"F7",X"28",X"5D",
		X"56",X"2E",X"E6",X"37",X"EB",X"88",X"7F",X"4D",X"66",X"7D",X"CD",X"2D",X"72",X"B9",X"D2",X"D7",
		X"11",X"5D",X"F5",X"0F",X"D4",X"C6",X"09",X"5D",X"F7",X"88",X"5D",X"76",X"0E",X"C6",X"DF",X"D6",
		X"68",X"6B",X"94",X"7F",X"CD",X"66",X"7D",X"4D",X"1B",X"72",X"39",X"2E",X"28",X"11",X"DD",X"F5",
		X"0F",X"74",X"EE",X"09",X"5D",X"F7",X"88",X"5D",X"D6",X"0E",X"EE",X"BF",X"FE",X"28",X"6B",X"B4",
		X"7F",X"4D",X"4E",X"7D",X"CD",X"33",X"5A",X"31",X"2E",X"28",X"19",X"5D",X"75",X"2F",X"54",X"EE",
		X"09",X"5D",X"F7",X"88",X"5D",X"76",X"0E",X"C6",X"FF",X"D6",X"68",X"CB",X"20",X"5F",X"ED",X"5D",
		X"CB",X"32",X"DE",X"5D",X"36",X"38",X"28",X"5D",X"36",X"25",X"28",X"5D",X"36",X"3E",X"29",X"26",
		X"0B",X"2E",X"0C",X"5D",X"4B",X"9A",X"CE",X"20",X"0E",X"A1",X"02",X"E8",X"6B",X"7A",X"5D",X"A1",
		X"54",X"E0",X"87",X"4D",X"30",X"FC",X"E1",X"49",X"CD",X"2D",X"5A",X"31",X"D2",X"D7",X"19",X"5D",
		X"F5",X"0F",X"D4",X"C6",X"09",X"5D",X"F7",X"88",X"5D",X"4B",X"9A",X"46",X"5D",X"B6",X"09",X"8B",
		X"DD",X"B6",X"2A",X"E1",X"DD",X"D6",X"2E",X"EE",X"1F",X"6B",X"A0",X"7F",X"CD",X"33",X"5A",X"31",
		X"0E",X"08",X"11",X"5D",X"F5",X"0F",X"D4",X"C6",X"09",X"5D",X"F7",X"88",X"5D",X"4B",X"9A",X"46",
		X"DD",X"B6",X"29",X"23",X"DD",X"B6",X"2A",X"E1",X"DD",X"D6",X"2E",X"EE",X"57",X"FE",X"60",X"6B",
		X"20",X"5F",X"4D",X"9B",X"DA",X"B9",X"0E",X"08",X"11",X"5D",X"F5",X"0F",X"D4",X"C6",X"09",X"5D",
		X"77",X"20",X"DD",X"4B",X"1A",X"4E",X"DD",X"B6",X"29",X"23",X"DD",X"B6",X"2A",X"E1",X"DD",X"D6",
		X"0E",X"C6",X"BF",X"D6",X"28",X"CB",X"B4",X"5F",X"4D",X"0D",X"DA",X"B9",X"F2",X"F7",X"11",X"5D",
		X"75",X"2F",X"54",X"EE",X"29",X"5D",X"77",X"20",X"DD",X"4B",X"1A",X"4E",X"DD",X"B6",X"29",X"23",
		X"5D",X"B6",X"AA",X"E9",X"5D",X"76",X"AE",X"C6",X"7F",X"D6",X"E8",X"CB",X"14",X"5F",X"4D",X"9B",
		X"72",X"B9",X"D4",X"D7",X"19",X"5D",X"75",X"2F",X"54",X"C6",X"29",X"5D",X"77",X"20",X"DD",X"4B",
		X"3A",X"46",X"5D",X"B6",X"A9",X"51",X"5D",X"B6",X"AA",X"E8",X"5D",X"76",X"AE",X"C6",X"77",X"D6",
		X"E8",X"CB",X"94",X"7F",X"CD",X"2D",X"72",X"B9",X"2C",X"28",X"19",X"5D",X"75",X"2F",X"54",X"C6",
		X"A9",X"5D",X"F7",X"88",X"5D",X"4B",X"3A",X"46",X"5D",X"B6",X"A9",X"51",X"5D",X"B6",X"AA",X"E8",
		X"DD",X"76",X"2E",X"C6",X"37",X"CB",X"94",X"7F",X"CD",X"2D",X"72",X"B9",X"2C",X"28",X"19",X"5D",
		X"F5",X"0F",X"D4",X"C6",X"A9",X"5D",X"F7",X"88",X"5D",X"4B",X"3A",X"46",X"5D",X"B6",X"A9",X"51",
		X"DD",X"B6",X"2A",X"E0",X"DD",X"76",X"2E",X"C6",X"77",X"D6",X"68",X"CB",X"88",X"7F",X"CD",X"33",
		X"7A",X"B9",X"54",X"F7",X"11",X"5D",X"F5",X"0F",X"D4",X"C6",X"A9",X"5D",X"F7",X"88",X"5D",X"4B",
		X"32",X"4E",X"DD",X"B6",X"29",X"59",X"DD",X"B6",X"2A",X"E0",X"DD",X"76",X"2E",X"C6",X"B7",X"D6",
		X"A0",X"CB",X"80",X"5F",X"4D",X"E6",X"79",X"DE",X"AB",X"5D",X"F7",X"89",X"5D",X"4B",X"3A",X"46",
		X"DD",X"B6",X"29",X"3C",X"DD",X"B6",X"2A",X"E1",X"DD",X"76",X"2E",X"D6",X"C8",X"CB",X"5E",X"7F",
		X"4D",X"D6",X"79",X"CE",X"AB",X"5D",X"F7",X"89",X"5D",X"4B",X"3A",X"46",X"5D",X"B6",X"A9",X"1C",
		X"DD",X"B6",X"2A",X"E1",X"DD",X"76",X"2E",X"D6",X"08",X"C6",X"17",X"CB",X"5E",X"7F",X"CD",X"C6",
		X"79",X"DE",X"AB",X"5D",X"F7",X"89",X"5D",X"4B",X"3A",X"46",X"5D",X"B6",X"A9",X"1C",X"5D",X"B6",
		X"2A",X"E1",X"DD",X"76",X"2E",X"D6",X"48",X"C6",X"57",X"CB",X"DA",X"7F",X"CD",X"56",X"71",X"CE",
		X"0B",X"5D",X"F7",X"89",X"5D",X"4B",X"9A",X"46",X"5D",X"B6",X"09",X"1C",X"5D",X"B6",X"0A",X"E9",
		X"DD",X"D6",X"2E",X"FE",X"A0",X"EE",X"97",X"6B",X"F2",X"7F",X"39",X"08",X"28",X"11",X"CD",X"56",
		X"D9",X"DE",X"0D",X"5D",X"F7",X"89",X"5D",X"4B",X"9A",X"46",X"5D",X"B6",X"09",X"C0",X"5D",X"B6",
		X"2A",X"E0",X"DD",X"D6",X"2E",X"FE",X"A8",X"EE",X"9F",X"6B",X"F2",X"7F",X"39",X"08",X"D7",X"11",
		X"4D",X"E6",X"D9",X"CE",X"0D",X"5D",X"F7",X"89",X"5D",X"4B",X"9A",X"46",X"5D",X"B6",X"09",X"C0",
		X"DD",X"B6",X"2A",X"E0",X"DD",X"D6",X"2E",X"FE",X"E0",X"6B",X"F2",X"7F",X"39",X"08",X"28",X"11",
		X"4D",X"D6",X"D9",X"DE",X"0D",X"5D",X"F7",X"89",X"5D",X"4B",X"9A",X"46",X"5D",X"B6",X"09",X"C0",
		X"DD",X"B6",X"2A",X"E0",X"DD",X"D6",X"2E",X"FE",X"A0",X"EE",X"97",X"6B",X"FE",X"7F",X"39",X"08",
		X"F7",X"39",X"4D",X"E6",X"D9",X"CE",X"0D",X"5D",X"F7",X"89",X"5D",X"4B",X"9A",X"46",X"5D",X"B6",
		X"29",X"40",X"DD",X"B6",X"2A",X"E0",X"DD",X"D6",X"2E",X"FE",X"E8",X"EE",X"DF",X"6B",X"FE",X"7F",
		X"5D",X"F7",X"0E",X"5D",X"B6",X"1E",X"0B",X"5D",X"B6",X"8D",X"08",X"5D",X"D6",X"1A",X"CD",X"EC",
		X"CB",X"87",X"DD",X"F7",X"3C",X"5D",X"36",X"3A",X"28",X"6B",X"38",X"71",X"DD",X"F7",X"2E",X"5D",
		X"B6",X"1E",X"0B",X"5D",X"B6",X"8D",X"08",X"5D",X"D6",X"1A",X"4B",X"27",X"5D",X"F7",X"1C",X"5D",
		X"36",X"3A",X"28",X"6B",X"38",X"71",X"DD",X"F7",X"2E",X"5D",X"36",X"3E",X"2B",X"5D",X"36",X"25",
		X"08",X"5D",X"D6",X"1C",X"CD",X"EC",X"4B",X"A7",X"5D",X"F7",X"1A",X"5D",X"B6",X"1C",X"08",X"CB",
		X"38",X"71",X"DD",X"F7",X"2E",X"5D",X"36",X"3E",X"2B",X"5D",X"36",X"25",X"28",X"5D",X"56",X"3C",
		X"4B",X"A7",X"5D",X"F7",X"BA",X"5D",X"B6",X"1C",X"A8",X"CB",X"B8",X"D9",X"5D",X"B6",X"3A",X"58",
		X"DD",X"B6",X"38",X"28",X"DD",X"B6",X"25",X"28",X"DD",X"B6",X"3E",X"29",X"DD",X"76",X"38",X"28",
		X"26",X"0A",X"06",X"88",X"A1",X"80",X"60",X"5D",X"D6",X"1A",X"BF",X"52",X"27",X"D8",X"8F",X"4D",
		X"B8",X"FC",X"08",X"5D",X"96",X"38",X"00",X"A9",X"DD",X"76",X"39",X"7F",X"14",X"5D",X"CB",X"3A",
		X"76",X"20",X"AA",X"DE",X"AA",X"C6",X"AF",X"5D",X"F7",X"19",X"A1",X"90",X"60",X"BE",X"A8",X"39",
		X"DD",X"76",X"28",X"C6",X"D4",X"96",X"DD",X"F7",X"28",X"4D",X"B1",X"71",X"CD",X"B7",X"FB",X"DA",
		X"2D",X"D9",X"5D",X"4B",X"A8",X"A6",X"6B",X"AA",X"EC",X"AE",X"AB",X"2E",X"AC",X"5D",X"4B",X"9A",
		X"66",X"A0",X"AB",X"A1",X"F4",X"E0",X"87",X"4D",X"B8",X"FC",X"FA",X"38",X"71",X"5D",X"56",X"32",
		X"FE",X"0A",X"EE",X"77",X"5D",X"F7",X"3A",X"5D",X"B6",X"09",X"AA",X"5D",X"B6",X"0A",X"61",X"5D",
		X"CB",X"32",X"E6",X"CB",X"25",X"71",X"21",X"0A",X"E0",X"07",X"CD",X"B8",X"FC",X"DA",X"38",X"71",
		X"5D",X"76",X"3A",X"C6",X"D5",X"5D",X"F7",X"9A",X"5D",X"B6",X"A9",X"20",X"5D",X"B6",X"AA",X"E8",
		X"DD",X"76",X"2E",X"C6",X"E8",X"AF",X"2F",X"AF",X"C6",X"29",X"4F",X"5D",X"56",X"28",X"E6",X"D4",
		X"B9",X"5D",X"F7",X"08",X"4B",X"6F",X"80",X"8B",X"5D",X"76",X"29",X"DE",X"AA",X"5D",X"F7",X"89",
		X"EB",X"25",X"71",X"5D",X"34",X"21",X"EB",X"25",X"71",X"5D",X"35",X"3E",X"20",X"BA",X"DD",X"76",
		X"AE",X"4B",X"D7",X"20",X"AE",X"A1",X"80",X"E8",X"6B",X"E6",X"78",X"A1",X"5A",X"E8",X"5D",X"F5",
		X"29",X"5D",X"74",X"2A",X"E6",X"C8",X"2F",X"AF",X"2F",X"7F",X"3E",X"28",X"21",X"33",X"71",X"39",
		X"5D",X"76",X"08",X"C6",X"F4",X"96",X"5D",X"F7",X"08",X"5D",X"4B",X"9A",X"06",X"4D",X"D4",X"7A",
		X"DD",X"D6",X"08",X"EE",X"29",X"5D",X"77",X"20",X"EB",X"8C",X"6B",X"28",X"29",X"2A",X"2B",X"29",
		X"08",X"0B",X"0A",X"5D",X"D6",X"8D",X"5D",X"66",X"09",X"5D",X"E6",X"0A",X"31",X"0E",X"08",X"39",
		X"14",X"9E",X"10",X"29",X"87",X"5D",X"77",X"25",X"C9",X"5D",X"CB",X"32",X"BE",X"5D",X"56",X"3A",
		X"BF",X"52",X"CC",X"D9",X"A0",X"3C",X"5D",X"4B",X"08",X"4E",X"80",X"AE",X"5D",X"4B",X"1C",X"FE",
		X"00",X"3A",X"B7",X"4D",X"72",X"F9",X"08",X"D1",X"B7",X"4A",X"CA",X"71",X"E6",X"24",X"EA",X"8C",
		X"D9",X"CB",X"B6",X"D9",X"4D",X"25",X"79",X"28",X"D1",X"97",X"4A",X"C2",X"D9",X"4B",X"77",X"4A",
		X"FB",X"71",X"E6",X"2B",X"EC",X"5B",X"59",X"6B",X"A4",X"71",X"DD",X"4B",X"3C",X"F6",X"EA",X"1E",
		X"D9",X"4D",X"50",X"79",X"00",X"71",X"BF",X"4A",X"C2",X"D9",X"4B",X"EF",X"80",X"4D",X"EE",X"0E",
		X"EC",X"5B",X"59",X"6B",X"A4",X"71",X"B7",X"4D",X"D5",X"F9",X"08",X"D1",X"B7",X"4A",X"CA",X"71",
		X"EE",X"0B",X"80",X"9A",X"5D",X"76",X"1A",X"45",X"64",X"5D",X"F7",X"1A",X"5D",X"76",X"8B",X"45",
		X"6C",X"5D",X"77",X"23",X"DD",X"D6",X"0C",X"CD",X"6C",X"5D",X"77",X"24",X"B7",X"49",X"DD",X"D6",
		X"1C",X"97",X"F8",X"45",X"64",X"5D",X"F7",X"1C",X"BF",X"49",X"4D",X"B2",X"7B",X"5D",X"4B",X"9A",
		X"FE",X"BF",X"C9",X"4D",X"DE",X"71",X"DD",X"F7",X"09",X"5D",X"36",X"3C",X"28",X"49",X"CD",X"7C",
		X"DA",X"4D",X"A8",X"DA",X"38",X"35",X"49",X"4D",X"E6",X"D9",X"5D",X"F7",X"89",X"49",X"4D",X"5C",
		X"5A",X"4D",X"00",X"72",X"A8",X"6E",X"2F",X"49",X"CD",X"2D",X"5A",X"5D",X"75",X"2F",X"54",X"EE",
		X"A9",X"5D",X"F7",X"88",X"49",X"4D",X"7F",X"DA",X"4D",X"BD",X"7A",X"29",X"83",X"49",X"4D",X"9B",
		X"72",X"5D",X"75",X"2F",X"54",X"C6",X"29",X"5D",X"77",X"20",X"C9",X"4D",X"77",X"72",X"CD",X"B5",
		X"7A",X"97",X"CD",X"EA",X"06",X"18",X"01",X"49",X"31",X"08",X"C0",X"97",X"CD",X"FA",X"D5",X"2F",
		X"0F",X"2F",X"E6",X"30",X"47",X"74",X"0F",X"2F",X"0F",X"C6",X"C8",X"95",X"C9",X"B9",X"28",X"C8",
		X"BF",X"45",X"72",X"75",X"EE",X"BE",X"37",X"BF",X"37",X"A6",X"A8",X"4B",X"34",X"67",X"CD",X"7B",
		X"32",X"48",X"19",X"49",X"DD",X"7E",X"29",X"5D",X"7E",X"2A",X"1A",X"4B",X"17",X"EF",X"C9",X"5D",
		X"56",X"09",X"5D",X"FE",X"AA",X"BB",X"12",X"35",X"2F",X"6F",X"26",X"08",X"49",X"5D",X"B6",X"0F",
		X"E8",X"5D",X"36",X"21",X"A8",X"5D",X"36",X"3A",X"2B",X"49",X"DD",X"B6",X"2F",X"08",X"DD",X"B6",
		X"28",X"09",X"5D",X"B6",X"29",X"A8",X"5D",X"B6",X"BA",X"0D",X"49",X"5D",X"B6",X"0F",X"B8",X"5D",
		X"36",X"20",X"2A",X"5D",X"36",X"3C",X"D3",X"5D",X"36",X"26",X"29",X"5D",X"36",X"27",X"2D",X"CB",
		X"BA",X"DB",X"5D",X"B6",X"AF",X"30",X"5D",X"B6",X"28",X"0A",X"5D",X"B6",X"BC",X"F5",X"5D",X"B6",
		X"26",X"29",X"DD",X"B6",X"27",X"2D",X"EB",X"3A",X"73",X"5D",X"36",X"2F",X"78",X"5D",X"36",X"20",
		X"AB",X"5D",X"B6",X"1C",X"57",X"5D",X"B6",X"8E",X"A9",X"5D",X"B6",X"8F",X"AD",X"CB",X"BA",X"DB",
		X"DD",X"B6",X"2F",X"D8",X"DD",X"B6",X"20",X"2B",X"DD",X"B6",X"3C",X"29",X"DD",X"B6",X"26",X"D7",
		X"5D",X"B6",X"2F",X"F3",X"6B",X"1A",X"7B",X"5D",X"B6",X"0F",X"98",X"5D",X"B6",X"88",X"AC",X"5D",
		X"36",X"3C",X"2B",X"5D",X"36",X"26",X"D7",X"5D",X"36",X"27",X"D3",X"CB",X"3A",X"73",X"DD",X"B6",
		X"0F",X"38",X"5D",X"B6",X"88",X"0D",X"5D",X"B6",X"1C",X"0D",X"5D",X"B6",X"8E",X"F7",X"5D",X"B6",
		X"0F",X"D3",X"DD",X"B6",X"09",X"E8",X"DD",X"B6",X"3A",X"D8",X"EB",X"85",X"5C",X"5D",X"36",X"2F",
		X"48",X"5D",X"B6",X"88",X"0A",X"5D",X"B6",X"89",X"1C",X"5D",X"B6",X"1A",X"60",X"49",X"5D",X"B6",
		X"2F",X"68",X"DD",X"B6",X"08",X"2A",X"DD",X"B6",X"09",X"30",X"DD",X"B6",X"3A",X"C8",X"C9",X"49",
		X"4D",X"D4",X"7A",X"5D",X"D6",X"88",X"DE",X"0A",X"6A",X"D2",X"DE",X"5D",X"D6",X"0F",X"DE",X"28",
		X"DA",X"52",X"5E",X"5D",X"36",X"20",X"D7",X"5D",X"36",X"2F",X"E0",X"6B",X"DA",X"76",X"DD",X"D6",
		X"0E",X"8F",X"6E",X"EB",X"C7",X"36",X"DB",X"4E",X"08",X"E7",X"C9",X"38",X"0D",X"38",X"C8",X"CB",
		X"E3",X"73",X"CD",X"85",X"5C",X"80",X"3E",X"5D",X"34",X"2E",X"DD",X"B4",X"0D",X"5D",X"36",X"3A",
		X"08",X"5D",X"B6",X"1E",X"0E",X"36",X"00",X"B2",X"48",X"45",X"6B",X"24",X"4B",X"5D",X"D6",X"1E",
		X"14",X"5D",X"77",X"3E",X"D6",X"22",X"20",X"31",X"DD",X"B6",X"3E",X"28",X"CD",X"7C",X"73",X"B0",
		X"18",X"5D",X"D6",X"8E",X"CD",X"EC",X"5D",X"F7",X"8E",X"5D",X"D6",X"8F",X"CD",X"EC",X"5D",X"F7",
		X"0F",X"4D",X"DC",X"FA",X"EB",X"52",X"5E",X"5D",X"35",X"3E",X"E8",X"5D",X"34",X"2E",X"DD",X"B6",
		X"8D",X"08",X"5D",X"B6",X"08",X"30",X"92",X"43",X"40",X"DE",X"8A",X"8F",X"6E",X"B1",X"C7",X"36",
		X"5C",X"4E",X"28",X"E7",X"56",X"5D",X"77",X"29",X"23",X"D6",X"DD",X"F7",X"2A",X"4D",X"9B",X"32",
		X"6B",X"24",X"4B",X"5D",X"4B",X"08",X"EE",X"48",X"92",X"66",X"44",X"56",X"0A",X"CA",X"85",X"DB",
		X"DD",X"D6",X"2D",X"7E",X"0A",X"C7",X"AF",X"2D",X"EE",X"B3",X"47",X"96",X"5D",X"4E",X"28",X"E7",
		X"56",X"A3",X"76",X"5D",X"46",X"0F",X"5D",X"EE",X"28",X"43",X"CD",X"EA",X"90",X"0E",X"80",X"0D",
		X"2B",X"CB",X"3D",X"74",X"0B",X"28",X"DD",X"F1",X"2F",X"5D",X"70",X"20",X"C3",X"A3",X"DD",X"76",
		X"29",X"16",X"90",X"0E",X"80",X"8B",X"95",X"CB",X"23",X"DC",X"94",X"5D",X"F7",X"89",X"6B",X"24",
		X"6B",X"28",X"EA",X"8C",X"6B",X"5D",X"36",X"28",X"08",X"A1",X"68",X"4C",X"39",X"A8",X"28",X"AE",
		X"AE",X"4B",X"C6",X"CA",X"84",X"4B",X"11",X"B8",X"50",X"A1",X"E4",X"DC",X"A2",X"4B",X"CC",X"36",
		X"48",X"B2",X"7E",X"4C",X"87",X"B2",X"78",X"4C",X"2E",X"2D",X"21",X"E8",X"4C",X"F7",X"19",X"B8",
		X"54",X"CB",X"84",X"4B",X"5D",X"76",X"BE",X"35",X"5D",X"F7",X"BE",X"A0",X"2F",X"07",X"B2",X"48",
		X"4C",X"34",X"32",X"6C",X"48",X"07",X"CD",X"00",X"74",X"CB",X"A3",X"20",X"E6",X"2B",X"E8",X"5D",
		X"D6",X"18",X"94",X"56",X"AE",X"30",X"A9",X"07",X"5D",X"F7",X"B8",X"8F",X"6E",X"8B",X"C7",X"36",
		X"75",X"4E",X"28",X"E7",X"56",X"A3",X"66",X"67",X"16",X"2E",X"39",X"89",X"4F",X"C5",X"29",X"2E",
		X"A8",X"45",X"B8",X"A1",X"2A",X"08",X"11",X"43",X"E9",X"35",X"A0",X"71",X"49",X"A6",X"52",X"5D",
		X"56",X"2D",X"F6",X"68",X"47",X"4B",X"6E",X"F7",X"C9",X"5F",X"74",X"C8",X"74",X"DA",X"74",X"4D",
		X"7C",X"C6",X"7C",X"E1",X"7C",X"2C",X"2C",X"24",X"A9",X"F3",X"7C",X"09",X"9B",X"5D",X"3E",X"8B",
		X"B7",X"29",X"D3",X"74",X"29",X"6B",X"7F",X"36",X"2F",X"43",X"28",X"D3",X"74",X"29",X"05",X"70",
		X"3E",X"8D",X"71",X"09",X"53",X"DC",X"A9",X"DF",X"79",X"9E",X"2C",X"DC",X"A9",X"F3",X"7C",X"09",
		X"CD",X"72",X"AC",X"25",X"4F",X"29",X"D3",X"74",X"29",X"65",X"74",X"C0",X"D7",X"DF",X"C7",X"CF",
		X"17",X"E6",X"08",X"E6",X"D7",X"E7",X"08",X"08",X"08",X"67",X"08",X"1F",X"DD",X"9D",X"DD",X"2B",
		X"5D",X"A1",X"5D",X"A7",X"5D",X"BD",X"5D",X"D7",X"F7",X"C7",X"E7",X"1F",X"E7",X"DF",X"C7",X"CF",
		X"17",X"67",X"77",X"E7",X"67",X"17",X"67",X"F7",X"77",X"67",X"17",X"67",X"F7",X"77",X"E7",X"17",
		X"E7",X"D7",X"F7",X"C7",X"E7",X"CF",X"D7",X"DF",X"C7",X"CF",X"BF",X"56",X"28",X"A4",X"2D",X"29",
		X"AC",X"6B",X"09",X"AA",X"14",X"08",X"AA",X"B6",X"08",X"AC",X"3B",X"09",X"AC",X"5D",X"D6",X"1E",
		X"14",X"EE",X"1F",X"5D",X"77",X"3E",X"DD",X"D6",X"28",X"A0",X"2D",X"CE",X"29",X"5D",X"77",X"28",
		X"EE",X"09",X"82",X"0F",X"45",X"A0",X"0C",X"23",X"6B",X"EC",X"DD",X"A3",X"92",X"08",X"45",X"2F",
		X"30",X"2D",X"03",X"83",X"EB",X"F1",X"5D",X"A3",X"23",X"5D",X"75",X"2F",X"DD",X"F4",X"08",X"5D",
		X"D6",X"0E",X"BF",X"A0",X"3B",X"32",X"89",X"45",X"7E",X"88",X"5D",X"F7",X"89",X"32",X"0E",X"45",
		X"B7",X"4A",X"DA",X"76",X"CB",X"D4",X"EA",X"52",X"5E",X"4B",X"6C",X"D5",X"21",X"3F",X"5E",X"80",
		X"0B",X"A1",X"9A",X"DE",X"21",X"0B",X"08",X"45",X"B9",X"B9",X"9E",X"E8",X"4C",X"9D",X"DE",X"5D",
		X"73",X"29",X"DD",X"F2",X"2A",X"6B",X"DA",X"76",X"DD",X"B5",X"38",X"6A",X"DA",X"76",X"DD",X"B6",
		X"0E",X"08",X"6B",X"D2",X"DE",X"5D",X"D6",X"1E",X"94",X"5D",X"F7",X"1E",X"07",X"B0",X"88",X"5D",
		X"56",X"25",X"C6",X"29",X"DD",X"F7",X"0D",X"5D",X"56",X"2E",X"B7",X"6A",X"D4",X"75",X"CD",X"54",
		X"7A",X"5D",X"D6",X"88",X"BF",X"D2",X"D2",X"DE",X"5D",X"76",X"0F",X"56",X"50",X"DA",X"D2",X"DE",
		X"DD",X"B4",X"2E",X"5D",X"36",X"3A",X"38",X"5D",X"36",X"28",X"B0",X"49",X"CD",X"54",X"72",X"5D",
		X"D6",X"88",X"DE",X"0A",X"6A",X"D2",X"7E",X"5D",X"D6",X"0F",X"DE",X"28",X"5A",X"D2",X"7E",X"07",
		X"32",X"A8",X"4D",X"B2",X"28",X"4D",X"C9",X"68",X"18",X"C8",X"B8",X"08",X"58",X"32",X"68",X"4D",
		X"4B",X"67",X"68",X"36",X"90",X"B2",X"E8",X"45",X"A1",X"4F",X"CD",X"5D",X"D6",X"0F",X"F7",X"A3",
		X"DD",X"76",X"20",X"F7",X"23",X"5D",X"56",X"21",X"EE",X"22",X"77",X"DE",X"2F",X"5D",X"77",X"21",
		X"31",X"DD",X"60",X"07",X"B2",X"5C",X"CD",X"5D",X"B6",X"0E",X"A9",X"5D",X"B6",X"18",X"B8",X"49",
		X"CD",X"92",X"FB",X"4D",X"54",X"FA",X"DD",X"4B",X"28",X"E6",X"EA",X"8C",X"6B",X"5D",X"36",X"28",
		X"A8",X"CB",X"22",X"4C",X"90",X"02",X"7E",X"48",X"7B",X"33",X"0B",X"DE",X"E8",X"DB",X"90",X"24",
		X"76",X"76",X"73",X"98",X"36",X"E0",X"65",X"75",X"99",X"97",X"76",X"4D",X"75",X"28",X"B2",X"E1",
		X"F8",X"DE",X"BC",X"1E",X"82",X"09",X"9C",X"DE",X"A9",X"DE",X"3C",X"1A",X"B9",X"29",X"A9",X"14",
		X"76",X"29",X"3E",X"36",X"28",X"1E",X"4F",X"5F",X"57",X"CF",X"C7",X"DF",X"D7",X"DE",X"D8",X"85",
		X"37",X"38",X"AF",X"08",X"20",X"8D",X"53",X"09",X"07",X"DE",X"AA",X"03",X"F9",X"83",X"FB",X"08",
		X"1E",X"4F",X"5F",X"57",X"CF",X"C7",X"DF",X"D7",X"8E",X"D8",X"85",X"B7",X"B8",X"2F",X"28",X"3C",
		X"2F",X"9D",X"A9",X"C2",X"7E",X"0A",X"E9",X"1E",X"82",X"AD",X"A8",X"F7",X"D6",X"E5",X"9A",X"93",
		X"CC",X"8C",X"2D",X"0F",X"D0",X"B0",X"A0",X"28",X"C6",X"2C",X"DD",X"66",X"29",X"5D",X"66",X"2A",
		X"ED",X"55",X"E9",X"59",X"DD",X"7E",X"A8",X"FB",X"4B",X"33",X"92",X"6D",X"C8",X"C6",X"88",X"5D",
		X"56",X"21",X"00",X"2A",X"EE",X"2A",X"BB",X"B2",X"A8",X"4A",X"AA",X"B2",X"A9",X"4A",X"3E",X"28",
		X"DD",X"7E",X"09",X"3D",X"4B",X"A3",X"5D",X"66",X"0F",X"5D",X"E6",X"88",X"CD",X"FA",X"96",X"08",
		X"D2",X"A9",X"5F",X"ED",X"39",X"28",X"2A",X"BF",X"C5",X"72",X"E1",X"7A",X"A0",X"77",X"EB",X"69",
		X"DF",X"55",X"D6",X"09",X"95",X"8F",X"2F",X"8D",X"7A",X"20",X"DF",X"75",X"CD",X"EC",X"C7",X"4B",
		X"15",X"4B",X"15",X"EE",X"2B",X"80",X"29",X"84",X"4D",X"CD",X"6C",X"EE",X"2B",X"A6",X"28",X"C7",
		X"D1",X"A2",X"2A",X"42",X"59",X"6F",X"26",X"08",X"5D",X"76",X"8D",X"8F",X"6E",X"0F",X"57",X"BE",
		X"28",X"11",X"56",X"A3",X"66",X"C7",X"12",X"ED",X"E8",X"EE",X"A8",X"5D",X"56",X"28",X"00",X"2A",
		X"CE",X"0A",X"17",X"B0",X"8E",X"55",X"56",X"09",X"15",X"3D",X"11",X"4B",X"DC",X"97",X"CD",X"EA",
		X"EB",X"FC",X"5F",X"01",X"E6",X"29",X"00",X"2F",X"D5",X"56",X"2A",X"DD",X"7E",X"2B",X"19",X"A2",
		X"2E",X"42",X"DD",X"66",X"09",X"A6",X"08",X"97",X"80",X"0E",X"31",X"08",X"08",X"43",X"CD",X"FA",
		X"22",X"AC",X"EA",X"CB",X"02",X"AE",X"EA",X"BF",X"C5",X"72",X"22",X"AE",X"EA",X"6B",X"32",X"6C",
		X"5D",X"4B",X"08",X"A6",X"6B",X"AA",X"4C",X"6A",X"6C",X"6E",X"6B",X"6D",X"6F",X"EC",X"EE",X"78",
		X"45",X"E7",X"71",X"FE",X"50",X"F2",X"A8",X"CC",X"AE",X"CC",X"8C",X"CC",X"BA",X"CC",X"98",X"CC",
		X"34",X"64",X"B2",X"64",X"00",X"80",X"10",X"90",X"01",X"81",X"11",X"91",X"02",X"82",X"12",X"92",
		X"AB",X"03",X"BB",X"13",X"AC",X"04",X"BC",X"14",X"AD",X"05",X"BD",X"15",X"E8",X"CD",X"C8",X"CD",
		X"50",X"65",X"D0",X"65",X"60",X"65",X"E0",X"65",X"70",X"65",X"F0",X"65",X"E8",X"20",X"20",X"20",
		X"A0",X"88",X"A0",X"88",X"A0",X"88",X"60",X"E1",X"A0",X"88",X"A0",X"88",X"84",X"98",X"B4",X"90",
		X"00",X"E9",X"D2",X"88",X"00",X"88",X"21",X"85",X"11",X"9D",X"31",X"95",X"E2",X"FB",X"02",X"8E",
		X"82",X"26",X"86",X"26",X"86",X"26",X"86",X"E3",X"54",X"03",X"A3",X"03",X"A3",X"03",X"A3",X"03",
		X"03",X"8B",X"D4",X"99",X"12",X"EF",X"E4",X"E8",X"11",X"88",X"E0",X"F2",X"C0",X"E8",X"88",X"F4",
		X"20",X"89",X"54",X"21",X"23",X"C0",X"99",X"80",X"ED",X"29",X"2D",X"88",X"65",X"B0",X"81",X"A5",
		X"C0",X"19",X"87",X"4D",X"6B",X"70",X"C0",X"29",X"A0",X"E8",X"31",X"28",X"4D",X"09",X"8D",X"28",
		X"65",X"B0",X"81",X"90",X"60",X"39",X"2F",X"4D",X"89",X"8B",X"28",X"C5",X"10",X"DD",X"96",X"9E",
		X"8A",X"D5",X"B6",X"38",X"88",X"D5",X"B6",X"25",X"88",X"43",X"3B",X"32",X"26",X"2A",X"06",X"2F",
		X"27",X"21",X"74",X"C7",X"6D",X"90",X"74",X"EB",X"A4",X"CB",X"7D",X"35",X"3E",X"E8",X"7D",X"36",
		X"9E",X"2A",X"5D",X"FE",X"AD",X"BC",X"DE",X"2B",X"90",X"29",X"8F",X"D5",X"F7",X"25",X"6B",X"8C",
		X"6B",X"21",X"DE",X"C0",X"F6",X"32",X"37",X"48",X"99",X"D9",X"DA",X"2E",X"2C",X"76",X"65",X"A0",
		X"ED",X"29",X"B7",X"28",X"11",X"E3",X"E9",X"18",X"55",X"29",X"42",X"E8",X"96",X"20",X"31",X"14",
		X"C2",X"29",X"D7",X"8C",X"6D",X"C0",X"51",X"39",X"38",X"63",X"8E",X"8E",X"B4",X"CD",X"60",X"F1",
		X"31",X"A0",X"63",X"0E",X"8E",X"BC",X"4D",X"E8",X"F1",X"19",X"58",X"C3",X"26",X"20",X"94",X"C5",
		X"60",X"F1",X"99",X"60",X"C3",X"2E",X"2D",X"14",X"6D",X"C0",X"51",X"EB",X"D7",X"C0",X"07",X"67",
		X"70",X"B7",X"CB",X"69",X"DB",X"7C",X"CE",X"64",X"E9",X"6B",X"EB",X"71",X"D8",X"61",X"EF",X"78",
		X"49",X"EF",X"4E",X"F9",X"69",X"EE",X"4E",X"F9",X"69",X"EE",X"6B",X"E8",X"4F",X"DA",X"4F",X"21",
		X"9D",X"E9",X"31",X"7E",X"E5",X"8E",X"F7",X"BE",X"0C",X"0E",X"8A",X"88",X"96",X"20",X"4D",X"E8",
		X"51",X"E5",X"21",X"A4",X"28",X"19",X"C3",X"E1",X"08",X"15",X"20",X"C5",X"C9",X"08",X"AC",X"00",
		X"04",X"05",X"04",X"1B",X"16",X"11",X"95",X"09",X"05",X"01",X"84",X"06",X"11",X"1C",X"17",X"12",
		X"9E",X"0A",X"AE",X"02",X"8C",X"07",X"BA",X"1D",X"98",X"13",X"9F",X"0B",X"AF",X"03",X"AB",X"18",
		X"03",X"0B",X"03",X"14",X"97",X"CF",X"92",X"A4",X"40",X"37",X"68",X"F9",X"DE",X"20",X"80",X"2E",
		X"16",X"D7",X"32",X"34",X"E8",X"C9",X"12",X"30",X"E8",X"21",X"A3",X"EA",X"2E",X"2E",X"96",X"00",
		X"0E",X"2B",X"30",X"D2",X"6B",X"E3",X"69",X"A7",X"B2",X"34",X"40",X"BA",X"9C",X"48",X"BF",X"40",
		X"02",X"39",X"E8",X"54",X"B5",X"00",X"2E",X"16",X"D7",X"32",X"1C",X"48",X"C9",X"12",X"18",X"48",
		X"A1",X"81",X"6A",X"0E",X"0E",X"B6",X"90",X"2E",X"80",X"27",X"A3",X"18",X"F0",X"C1",X"4D",X"1E",
		X"62",X"93",X"D8",X"16",X"D7",X"32",X"1C",X"48",X"C9",X"CD",X"BE",X"EA",X"93",X"F8",X"DD",X"E5",
		X"6D",X"29",X"35",X"EA",X"50",X"1E",X"08",X"99",X"11",X"FE",X"A3",X"6E",X"C7",X"DE",X"A3",X"5E",
		X"23",X"56",X"76",X"32",X"F7",X"55",X"23",X"56",X"23",X"E5",X"B7",X"00",X"0F",X"21",X"2B",X"EB",
		X"4D",X"3F",X"6A",X"C5",X"38",X"EA",X"A1",X"21",X"6B",X"43",X"D0",X"E9",X"A1",X"DF",X"6A",X"C5",
		X"3F",X"EA",X"CD",X"B8",X"62",X"21",X"D5",X"EA",X"CD",X"3F",X"62",X"E1",X"DD",X"21",X"A8",X"4D",
		X"56",X"2B",X"76",X"E5",X"73",X"09",X"45",X"55",X"5D",X"3E",X"08",X"28",X"5D",X"3E",X"8D",X"28",
		X"23",X"5E",X"23",X"7E",X"E5",X"02",X"1A",X"48",X"19",X"54",X"E6",X"29",X"67",X"C3",X"E1",X"C5",
		X"73",X"0F",X"4D",X"2B",X"D6",X"D5",X"F7",X"21",X"4D",X"13",X"BA",X"F5",X"E9",X"41",X"A1",X"BE",
		X"62",X"58",X"9E",X"88",X"B9",X"19",X"61",X"16",X"2B",X"FD",X"A8",X"16",X"2F",X"29",X"D7",X"8A",
		X"4D",X"E8",X"F1",X"65",X"A1",X"B4",X"88",X"99",X"CB",X"61",X"00",X"BD",X"A0",X"C4",X"79",X"C1",
		X"8E",X"8B",X"D6",X"38",X"D5",X"C9",X"B8",X"AA",X"B8",X"A8",X"B8",X"AE",X"B8",X"9C",X"B8",X"BA",
		X"10",X"A8",X"21",X"28",X"D8",X"BE",X"9C",X"43",X"C7",X"EA",X"21",X"28",X"D8",X"BE",X"AA",X"43",
		X"67",X"C2",X"89",X"88",X"38",X"16",X"0A",X"EB",X"67",X"C2",X"89",X"88",X"2D",X"16",X"0A",X"EB",
		X"C7",X"EA",X"21",X"28",X"89",X"BE",X"AA",X"45",X"FD",X"F5",X"ED",X"C5",X"02",X"3F",X"26",X"20",
		X"D6",X"38",X"D5",X"D5",X"41",X"DD",X"F6",X"AD",X"B4",X"D5",X"36",X"8E",X"B0",X"89",X"27",X"DD",
		X"F7",X"25",X"DD",X"65",X"4D",X"8C",X"CB",X"F5",X"E9",X"BE",X"19",X"C5",X"95",X"6D",X"F9",X"41",
		X"B5",X"20",X"FC",X"DD",X"41",X"C9",X"81",X"27",X"62",X"2D",X"F8",X"3E",X"28",X"19",X"FE",X"12",
		X"98",X"48",X"49",X"2B",X"AB",X"3B",X"BB",X"AB",X"A3",X"21",X"99",X"31",X"81",X"A1",X"91",X"E8",
		X"60",X"D8",X"68",X"95",X"30",X"66",X"62",X"45",X"62",X"7C",X"62",X"5B",X"62",X"6A",X"62",X"49",
		X"C2",X"56",X"43",X"8D",X"88",X"27",X"C3",X"D5",X"88",X"0E",X"14",X"C9",X"8A",X"29",X"BA",X"EB",
		X"86",X"89",X"15",X"C6",X"E1",X"25",X"28",X"A1",X"63",X"B6",X"29",X"94",X"76",X"42",X"1C",X"88",
		X"94",X"EB",X"36",X"29",X"DE",X"C8",X"41",X"28",X"88",X"B7",X"C3",X"26",X"89",X"6D",X"1A",X"CA",
		X"03",X"89",X"0F",X"C3",X"9E",X"88",X"5E",X"48",X"EB",X"49",X"EC",X"4A",X"ED",X"4E",X"C9",X"4F",
		X"C2",X"40",X"C3",X"58",X"53",X"59",X"54",X"5A",X"55",X"5E",X"D1",X"5F",X"D2",X"50",X"D3",X"38",
		X"08",X"F0",X"28",X"62",X"63",X"2A",X"21",X"76",X"A1",X"76",X"39",X"20",X"A8",X"28",X"5A",X"EB",
		X"0C",X"A9",X"DF",X"81",X"DF",X"B9",X"68",X"91",X"68",X"3B",X"0E",X"E4",X"08",X"E2",X"6B",X"2A",
		X"69",X"E9",X"B3",X"E9",X"38",X"20",X"50",X"28",X"52",X"EB",X"2A",X"AD",X"62",X"8D",X"62",X"3A",
		X"88",X"00",X"08",X"02",X"6B",X"2A",X"2D",X"EB",X"35",X"EB",X"08",X"D7",X"F0",X"BF",X"AF",X"A6",
		X"26",X"85",X"B6",X"97",X"28",X"DE",X"EF",X"8C",X"17",X"28",X"28",X"68",X"2D",X"2F",X"00",X"A7",
		X"F7",X"B7",X"38",X"B0",X"07",X"4F",X"D7",X"C7",X"76",X"28",X"08",X"A7",X"2F",X"37",X"BF",X"D4",
		X"C3",X"C7",X"3D",X"DF",X"D7",X"97",X"84",X"33",X"EF",X"28",X"28",X"D7",X"2F",X"C7",X"D0",X"88",
		X"A5",X"08",X"BF",X"DE",X"B8",X"A6",X"08",X"4F",X"F0",X"28",X"08",X"B7",X"3F",X"9F",X"A7",X"86",
		X"85",X"28",X"D7",X"97",X"34",X"A3",X"22",X"2F",X"C5",X"28",X"DD",X"56",X"2D",X"D6",X"0C",X"DA",
		X"93",X"32",X"DE",X"3A",X"7A",X"13",X"9A",X"F6",X"8D",X"A8",X"8C",X"BA",X"EF",X"48",X"4B",X"4F",
		X"00",X"2D",X"DD",X"36",X"28",X"28",X"C9",X"DD",X"56",X"28",X"E6",X"DC",X"F6",X"A8",X"DD",X"77",
		X"08",X"A7",X"5D",X"7F",X"0E",X"D5",X"F7",X"25",X"5D",X"7F",X"8A",X"D5",X"F7",X"3C",X"5D",X"7F",
		X"1A",X"DD",X"77",X"23",X"DD",X"77",X"0C",X"12",X"18",X"48",X"26",X"28",X"47",X"1E",X"0F",X"CD",
		X"88",X"6D",X"D4",X"07",X"57",X"1E",X"08",X"29",X"4E",X"EF",X"11",X"DE",X"A3",X"5E",X"5D",X"7B",
		X"29",X"DD",X"72",X"2A",X"DD",X"36",X"3E",X"2A",X"3E",X"28",X"12",X"3C",X"E8",X"AF",X"5F",X"21",
		X"EE",X"ED",X"11",X"FE",X"A3",X"6E",X"C7",X"D5",X"D6",X"2D",X"7E",X"24",X"2F",X"DF",X"11",X"FE",
		X"0F",X"5F",X"9E",X"88",X"6B",X"3A",X"63",X"C5",X"EB",X"BA",X"E8",X"09",X"63",X"52",X"46",X"89",
		X"5D",X"7B",X"8F",X"D5",X"F7",X"20",X"A3",X"FE",X"4D",X"44",X"D3",X"D5",X"F7",X"21",X"5D",X"3E",
		X"3A",X"88",X"4B",X"3B",X"1A",X"D9",X"A8",X"21",X"B7",X"C4",X"7D",X"E5",X"59",X"29",X"2B",X"88",
		X"CD",X"30",X"A1",X"20",X"88",X"99",X"55",X"5C",X"33",X"3E",X"88",X"09",X"98",X"28",X"CD",X"30",
		X"79",X"DD",X"D5",X"8F",X"F4",X"E6",X"29",X"DD",X"D7",X"A8",X"C7",X"C3",X"A8",X"CD",X"CC",X"D3",
		X"7E",X"2C",X"5D",X"7F",X"A9",X"D5",X"B6",X"2E",X"89",X"D5",X"B6",X"3E",X"A8",X"C5",X"96",X"ED",
		X"B2",X"8C",X"E8",X"5F",X"B2",X"87",X"E8",X"4F",X"B2",X"B8",X"E8",X"CB",X"D3",X"20",X"0E",X"CB",
		X"97",X"46",X"80",X"01",X"DE",X"B8",X"90",X"26",X"96",X"B8",X"6B",X"1E",X"C4",X"46",X"80",X"01",
		X"76",X"C8",X"B0",X"8A",X"B6",X"C8",X"7D",X"CB",X"2D",X"CE",X"A0",X"AB",X"7D",X"CB",X"28",X"4E",
		X"5D",X"3E",X"AC",X"20",X"6B",X"99",X"C4",X"E5",X"64",X"D5",X"4B",X"28",X"0E",X"D5",X"B6",X"24",
		X"D0",X"DD",X"D7",X"B8",X"4B",X"3B",X"1A",X"10",X"1E",X"E0",X"79",X"08",X"81",X"93",X"65",X"DD",
		X"ED",X"51",X"21",X"2B",X"88",X"E5",X"B8",X"29",X"A8",X"28",X"11",X"DD",X"74",X"1B",X"B6",X"28",
		X"89",X"98",X"28",X"C5",X"10",X"DD",X"96",X"9E",X"29",X"CD",X"36",X"C5",X"79",X"DD",X"D5",X"8F",
		X"D4",X"66",X"89",X"D5",X"F7",X"20",X"77",X"DD",X"00",X"C5",X"6C",X"FB",X"5D",X"7F",X"A9",X"BA",
		X"2C",X"48",X"FF",X"12",X"27",X"48",X"EF",X"12",X"18",X"48",X"6B",X"73",X"80",X"A8",X"6B",X"17",
		X"6E",X"A8",X"29",X"43",X"89",X"ED",X"6E",X"A0",X"29",X"F6",X"78",X"B8",X"0A",X"BE",X"78",X"D5",
		X"CB",X"2D",X"6E",X"00",X"0E",X"DD",X"77",X"3A",X"DD",X"36",X"2E",X"88",X"DD",X"CB",X"28",X"0E",
		X"6B",X"13",X"9A",X"E5",X"64",X"D5",X"F7",X"3A",X"5D",X"3E",X"0E",X"08",X"5D",X"C3",X"08",X"4E",
		X"EB",X"13",X"1A",X"98",X"A0",X"E0",X"DD",X"56",X"2D",X"0F",X"0F",X"0F",X"4F",X"E6",X"2B",X"F6",
		X"F0",X"5F",X"D1",X"66",X"60",X"76",X"08",X"DF",X"21",X"20",X"08",X"E5",X"B8",X"C1",X"16",X"ED",
		X"A2",X"ED",X"86",X"ED",X"92",X"ED",X"EE",X"ED",X"FA",X"ED",X"DE",X"ED",X"C2",X"ED",X"F6",X"ED",
		X"0A",X"EE",X"8E",X"EE",X"9A",X"EE",X"2E",X"EE",X"3A",X"EE",X"BE",X"EE",X"CA",X"EE",X"5E",X"EE",
		X"62",X"EE",X"46",X"EE",X"52",X"EE",X"AE",X"EE",X"BA",X"EE",X"9E",X"EE",X"82",X"EE",X"B6",X"EE",
		X"42",X"EE",X"C6",X"EE",X"D2",X"EE",X"66",X"EE",X"72",X"EE",X"F6",X"EE",X"8A",X"EF",X"1E",X"EF",
		X"22",X"EF",X"06",X"EF",X"12",X"EF",X"F8",X"B0",X"30",X"B0",X"F8",X"E0",X"30",X"E0",X"F8",X"10",
		X"38",X"10",X"20",X"B8",X"68",X"B8",X"20",X"E8",X"68",X"E8",X"20",X"18",X"68",X"18",X"40",X"A0",
		X"30",X"A0",X"E8",X"70",X"20",X"F0",X"E8",X"00",X"30",X"80",X"E0",X"B0",X"20",X"B0",X"C8",X"E0",
		X"38",X"E0",X"50",X"10",X"38",X"10",X"E8",X"B0",X"E8",X"70",X"E8",X"10",X"C0",X"10",X"E8",X"40",
		X"C8",X"40",X"78",X"60",X"B0",X"60",X"28",X"E0",X"78",X"00",X"B0",X"00",X"A8",X"80",X"78",X"B0",
		X"40",X"B0",X"40",X"E0",X"58",X"E0",X"40",X"10",X"58",X"10",X"00",X"E0",X"00",X"10",X"70",X"30",
		X"F0",X"60",X"F0",X"F0",X"F0",X"80",X"30",X"30",X"78",X"30",X"70",X"30",X"B8",X"30",X"B0",X"30",
		X"58",X"30",X"C0",X"A8",X"00",X"68",X"C0",X"08",X"00",X"08",X"C0",X"80",X"00",X"80",X"98",X"80",
		X"10",X"F0",X"60",X"E8",X"A0",X"E8",X"C8",X"F0",X"F0",X"20",X"58",X"80",X"F8",X"80",X"40",X"D8",
		X"10",X"08",X"F0",X"88",X"B0",X"80",X"E0",X"60",X"38",X"60",X"F8",X"00",X"20",X"00",X"A8",X"80",
		X"D0",X"20",X"68",X"B8",X"78",X"B8",X"60",X"B8",X"A0",X"B8",X"B0",X"B8",X"E8",X"B8",X"78",X"A0",
		X"10",X"A0",X"D8",X"78",X"10",X"78",X"D8",X"88",X"10",X"88",X"08",X"B0",X"08",X"70",X"D0",X"F0",
		X"B8",X"F0",X"60",X"00",X"A0",X"00",X"78",X"B8",X"B0",X"B8",X"D7",X"80",X"78",X"F0",X"B0",X"F0",
		X"77",X"08",X"E0",X"A8",X"38",X"A8",X"D8",X"60",X"10",X"60",X"B0",X"F8",X"68",X"F8",X"10",X"E8",
		X"90",X"C0",X"E8",X"C0",X"20",X"00",X"00",X"00",X"30",X"00",X"38",X"80",X"98",X"08",X"A0",X"08",
		X"20",X"08",X"F8",X"88",X"C0",X"88",X"D8",X"68",X"20",X"68",X"08",X"E8",X"D8",X"08",X"10",X"08",
		X"A8",X"00",X"40",X"E8",X"E8",X"E8",X"40",X"D0",X"E8",X"D0",X"40",X"00",X"E8",X"00",X"00",X"C8",
		X"20",X"68",X"77",X"F8",X"F0",X"F8",X"90",X"40",X"10",X"40",X"D8",X"60",X"20",X"60",X"D8",X"F0",
		X"80",X"F0",X"78",X"00",X"80",X"00",X"18",X"80",X"F0",X"80",X"18",X"18",X"F0",X"18",X"18",X"68",
		X"50",X"40",X"C0",X"30",X"38",X"30",X"C0",X"60",X"38",X"60",X"C0",X"F0",X"38",X"F0",X"E0",X"A8",
		X"A0",X"80",X"40",X"F8",X"A0",X"F8",X"40",X"18",X"A0",X"18",X"68",X"B0",X"48",X"18",X"00",X"18",
		X"38",X"30",X"30",X"18",X"40",X"70",X"D8",X"10",X"10",X"10",X"88",X"10",X"A0",X"40",X"08",X"40",
		X"D8",X"68",X"D8",X"B8",X"D8",X"B0",X"D8",X"C0",X"D8",X"08",X"D8",X"20",X"D8",X"68",X"60",X"B0",
		X"A0",X"B0",X"48",X"70",X"00",X"70",X"40",X"70",X"00",X"10",X"A8",X"A8",X"E8",X"A8",X"A0",X"A8",
		X"C0",X"A8",X"68",X"40",X"C8",X"40",X"74",X"A8",X"74",X"A8",X"74",X"A8",X"74",X"A8",X"74",X"A8",
		X"7C",X"A8",X"0C",X"A8",X"BC",X"78",X"44",X"78",X"F8",X"F0",X"10",X"F0",X"0C",X"08",X"DC",X"40",
		X"8C",X"F8",X"BC",X"80",X"A4",X"80",X"74",X"F8",X"A8",X"60",X"38",X"70",X"60",X"70",X"80",X"70",
		X"F0",X"70",X"98",X"18",X"70",X"18",X"BA",X"E1",X"AD",X"E1",X"4F",X"E1",X"6C",X"E1",X"79",X"E1",
		X"56",X"E1",X"8B",X"E1",X"98",X"E1",X"A5",X"E1",X"B2",X"E1",X"97",X"E1",X"CC",X"E1",X"D9",X"E1",
		X"66",X"E1",X"73",X"E1",X"08",X"28",X"08",X"2A",X"0B",X"2B",X"09",X"29",X"08",X"29",X"0A",X"29",
		X"28",X"29",X"2A",X"29",X"B2",X"EF",X"93",X"EF",X"EC",X"EF",X"CD",X"EF",X"FE",X"EF",X"EC",X"EF",
		X"B3",X"EF",X"32",X"EF",X"B3",X"EF",X"B9",X"E0",X"4A",X"E0",X"CB",X"E0",X"32",X"EF",X"E0",X"EF",
		X"DF",X"EF",X"C0",X"EF",X"B2",X"EF",X"DF",X"EF",X"F1",X"EF",X"D2",X"EF",X"F1",X"EF",X"DF",X"EF",
		X"71",X"EF",X"F2",X"EF",X"71",X"EF",X"0B",X"E0",X"8C",X"E0",X"1D",X"E0",X"9E",X"E0",X"2F",X"E0",
		X"30",X"E0",X"3C",X"21",X"83",X"28",X"66",X"E0",X"29",X"D0",X"21",X"3C",X"0A",X"96",X"28",X"EE",
		X"E8",X"29",X"A4",X"AA",X"1C",X"22",X"B6",X"28",X"6E",X"E0",X"09",X"FC",X"2B",X"3C",X"8B",X"59",
		X"28",X"EE",X"40",X"29",X"14",X"AC",X"3C",X"23",X"F9",X"28",X"66",X"E0",X"29",X"30",X"25",X"3C",
		X"0F",X"0D",X"08",X"EE",X"E8",X"29",X"14",X"AE",X"1C",X"2F",X"05",X"28",X"6E",X"E0",X"09",X"A8",
		X"27",X"3C",X"0B",X"59",X"28",X"EE",X"40",X"29",X"84",X"AF",X"3C",X"22",X"96",X"28",X"66",X"E0",
		X"89",X"00",X"A0",X"20",X"8D",X"AB",X"88",X"EE",X"E0",X"29",X"D8",X"A1",X"8D",X"2C",X"98",X"28",
		X"66",X"E0",X"29",X"F0",X"01",X"8B",X"2C",X"A8",X"28",X"C6",X"40",X"89",X"8C",X"A1",X"09",X"8F",
		X"B0",X"28",X"C6",X"E0",X"89",X"10",X"A1",X"23",X"8F",X"6E",X"88",X"EE",X"E0",X"29",X"38",X"A1",
		X"0E",X"8F",X"5B",X"88",X"66",X"E0",X"29",X"45",X"01",X"9D",X"0A",X"68",X"28",X"C6",X"40",X"89",
		X"CF",X"A2",X"9A",X"22",X"22",X"28",X"C6",X"E0",X"89",X"31",X"A3",X"3A",X"AB",X"93",X"88",X"EE",
		X"40",X"89",X"CD",X"A3",X"3C",X"A9",X"83",X"88",X"66",X"E0",X"29",X"1B",X"04",X"AD",X"2F",X"DC",
		X"88",X"EE",X"E0",X"29",X"CF",X"A5",X"88",X"D7",X"37",X"9F",X"97",X"A7",X"86",X"35",X"9C",X"7A",
		X"9B",X"8E",X"B6",X"57",X"A4",X"88",X"85",X"E0",X"B6",X"E0",X"97",X"E0",X"E7",X"E0",X"F0",X"E0",
		X"71",X"E0",X"71",X"E0",X"50",X"E0",X"47",X"E0",X"00",X"E0",X"59",X"E0",X"7A",X"E0",X"68",X"E0",
		X"A0",X"E0",X"F9",X"E0",X"DA",X"E0",X"C8",X"E0",X"28",X"88",X"28",X"88",X"2B",X"8B",X"2B",X"8B",
		X"A9",X"20",X"C8",X"28",X"BD",X"E1",X"8B",X"73",X"91",X"8B",X"91",X"C3",X"91",X"21",X"A8",X"68",
		X"28",X"BD",X"41",X"89",X"33",X"92",X"09",X"8F",X"10",X"88",X"1D",X"E1",X"29",X"F3",X"32",X"A9",
		X"8E",X"B8",X"88",X"35",X"E1",X"29",X"32",X"BA",X"AD",X"2F",X"DC",X"28",X"BD",X"E1",X"89",X"D8",
		X"32",X"AB",X"08",X"D8",X"28",X"BD",X"41",X"89",X"4B",X"93",X"0F",X"8D",X"6E",X"88",X"1D",X"E1",
		X"8B",X"8B",X"93",X"C6",X"93",X"B1",X"94",X"21",X"8F",X"B0",X"88",X"35",X"E1",X"29",X"0C",X"BC",
		X"09",X"8E",X"30",X"88",X"1D",X"E1",X"29",X"4B",X"34",X"AC",X"2D",X"97",X"28",X"BD",X"41",X"89",
		X"F1",X"BC",X"8F",X"2E",X"5C",X"28",X"9D",X"E1",X"09",X"BD",X"3D",X"22",X"88",X"60",X"08",X"35",
		X"41",X"29",X"8F",X"BD",X"0D",X"2E",X"48",X"28",X"1D",X"E1",X"29",X"57",X"35",X"28",X"38",X"30",
		X"28",X"A0",X"3C",X"B5",X"B7",X"3C",X"1D",X"AF",X"A5",X"D7",X"47",X"28",X"A3",X"20",X"0D",X"AB",
		X"28",X"7C",X"41",X"29",X"6D",X"EC",X"45",X"EC",X"BD",X"EC",X"08",X"2D",X"23",X"28",X"7C",X"E1",
		X"09",X"95",X"6C",X"CD",X"6C",X"25",X"6D",X"22",X"0E",X"BE",X"08",X"7C",X"E9",X"29",X"25",X"E5",
		X"E1",X"E5",X"1D",X"E6",X"28",X"2F",X"2D",X"2B",X"27",X"A7",X"28",X"2C",X"D7",X"2F",X"10",X"B7",
		X"F6",X"D5",X"F0",X"EF",X"89",X"2E",X"38",X"28",X"08",X"E2",X"09",X"55",X"6D",X"3B",X"6E",X"61",
		X"66",X"21",X"2E",X"B8",X"28",X"28",X"42",X"29",X"57",X"EE",X"B5",X"EE",X"C3",X"EE",X"0A",X"2D",
		X"AD",X"28",X"08",X"E2",X"09",X"A9",X"6F",X"7B",X"6F",X"0D",X"6F",X"21",X"0E",X"B8",X"08",X"38",
		X"42",X"29",X"B7",X"EF",X"C5",X"EF",X"23",X"E0",X"08",X"2D",X"23",X"28",X"20",X"E2",X"29",X"71",
		X"E8",X"09",X"E8",X"81",X"E8",X"20",X"0E",X"A2",X"08",X"38",X"EA",X"29",X"51",X"E0",X"09",X"E1",
		X"31",X"E1",X"0A",X"2E",X"36",X"28",X"30",X"E2",X"29",X"E9",X"41",X"15",X"41",X"51",X"41",X"20",
		X"0D",X"AB",X"08",X"68",X"EA",X"29",X"1D",X"E2",X"BD",X"E2",X"6D",X"E2",X"8A",X"2E",X"3E",X"28",
		X"68",X"E2",X"29",X"05",X"42",X"41",X"42",X"2D",X"43",X"22",X"2E",X"BE",X"28",X"68",X"42",X"29",
		X"49",X"E3",X"FD",X"E3",X"B1",X"E3",X"8C",X"2F",X"CD",X"28",X"48",X"E2",X"09",X"DD",X"EB",X"61",
		X"44",X"15",X"44",X"22",X"2E",X"A2",X"28",X"68",X"42",X"29",X"F1",X"E4",X"05",X"E5",X"41",X"E5",
		X"88",X"D7",X"36",X"8C",X"23",X"85",X"34",X"D0",X"8F",X"2C",X"BC",X"AD",X"F7",X"A5",X"88",X"A8",
		X"28",X"77",X"F7",X"47",X"83",X"87",X"20",X"25",X"2F",X"8C",X"30",X"A5",X"E8",X"08",X"28",X"98",
		X"88",X"D7",X"57",X"CF",X"23",X"A7",X"80",X"94",X"8F",X"2C",X"90",X"D5",X"48",X"08",X"88",X"A8",
		X"28",X"77",X"C5",X"47",X"AD",X"8C",X"20",X"44",X"2F",X"84",X"30",X"A5",X"57",X"A7",X"28",X"80",
		X"88",X"28",X"8C",X"AC",X"80",X"B8",X"37",X"B7",X"47",X"2F",X"08",X"C6",X"9D",X"D5",X"77",X"28",
		X"E0",X"E2",X"F2",X"E2",X"38",X"E3",X"06",X"E3",X"68",X"E3",X"7E",X"E3",X"44",X"E3",X"52",X"E3",
		X"02",X"E3",X"30",X"E3",X"64",X"E3",X"76",X"E3",X"BC",X"E4",X"CE",X"E4",X"F8",X"E4",X"E2",X"E4",
		X"A8",X"E4",X"A2",X"E4",X"90",X"E4",X"CE",X"E4",X"E0",X"E4",X"F6",X"E4",X"2C",X"E5",X"3C",X"E5",
		X"86",X"E5",X"B0",X"E5",X"DE",X"E5",X"F4",X"E5",X"3A",X"E5",X"10",X"E5",X"4A",X"E5",X"9C",X"E6",
		X"06",X"E6",X"14",X"E6",X"5A",X"E6",X"74",X"E6",X"C1",X"E2",X"29",X"E3",X"1F",X"E3",X"31",X"E3",
		X"ED",X"E3",X"C1",X"E3",X"D3",X"E3",X"19",X"E3",X"25",X"E3",X"5B",X"E3",X"55",X"E3",X"AD",X"E4",
		X"31",X"E4",X"4F",X"E4",X"61",X"E4",X"75",X"E4",X"B9",X"E4",X"85",X"E4",X"E9",X"E4",X"FB",X"E4",
		X"63",X"E4",X"73",X"E4",X"8D",X"E5",X"BD",X"E5",X"A7",X"E5",X"CF",X"E5",X"E1",X"E5",X"2D",X"E5",
		X"A5",X"E5",X"B5",X"E5",X"C3",X"E5",X"05",X"E6",X"35",X"E6",X"4B",X"E6",X"67",X"E6",X"A9",X"E6",
		X"8C",X"CE",X"41",X"EE",X"43",X"CE",X"44",X"EE",X"46",X"2C",X"78",X"C9",X"F8",X"CB",X"78",X"CC",
		X"58",X"46",X"2F",X"1C",X"E1",X"D4",X"E2",X"9C",X"E3",X"54",X"E3",X"1C",X"E4",X"D4",X"E5",X"DC",
		X"66",X"2F",X"A2",X"C9",X"CA",X"CA",X"AA",X"CB",X"C2",X"CB",X"A2",X"CC",X"CA",X"CD",X"EA",X"CE",
		X"2F",X"EE",X"E1",X"F6",X"E1",X"D6",X"E2",X"F6",X"E4",X"7C",X"E5",X"CC",X"E2",X"F4",X"E5",X"2F",
		X"D8",X"C9",X"D2",X"CA",X"7A",X"C9",X"72",X"CA",X"7A",X"CC",X"DC",X"CE",X"7A",X"CE",X"09",X"D0",
		X"E1",X"2F",X"6A",X"CE",X"4E",X"CB",X"D8",X"CC",X"62",X"CE",X"C6",X"C9",X"46",X"CB",X"D0",X"CC",
		X"0E",X"4E",X"62",X"7E",X"63",X"DE",X"63",X"DC",X"64",X"7E",X"66",X"E4",X"66",X"2C",X"66",X"C9",
		X"C8",X"CA",X"C6",X"CC",X"62",X"CE",X"2D",X"E6",X"E2",X"F6",X"E3",X"66",X"E4",X"76",X"E5",X"E6",
		X"66",X"2D",X"58",X"CA",X"48",X"CB",X"78",X"CC",X"68",X"CD",X"58",X"CE",X"0B",X"6A",X"63",X"CA",
		X"E4",X"6A",X"E6",X"2B",X"54",X"CB",X"DC",X"CC",X"54",X"CE",X"0B",X"64",X"E1",X"10",X"E1",X"DC",
		X"61",X"44",X"62",X"30",X"63",X"D4",X"63",X"64",X"64",X"10",X"64",X"D8",X"64",X"FA",X"63",X"66",
		X"E6",X"20",X"A6",X"C9",X"B2",X"C9",X"CE",X"CA",X"26",X"CB",X"4E",X"CC",X"A6",X"CC",X"78",X"CE",
		X"E8",X"CE",X"0D",X"B4",X"62",X"36",X"63",X"AE",X"64",X"E2",X"65",X"E6",X"66",X"2D",X"0A",X"CA",
		X"20",X"CB",X"18",X"CC",X"7C",X"CD",X"78",X"CE",X"0D",X"04",X"E1",X"90",X"E1",X"A0",X"E2",X"B8",
		X"63",X"32",X"64",X"B2",X"64",X"2A",X"65",X"EA",X"65",X"62",X"66",X"F8",X"66",X"24",X"63",X"A0",
		X"E4",X"22",X"E4",X"24",X"AA",X"C9",X"2C",X"CC",X"24",X"CC",X"5C",X"CD",X"14",X"CD",X"4E",X"CE",
		X"7C",X"CE",X"86",X"C9",X"AA",X"CA",X"1E",X"CC",X"3A",X"CB",X"3C",X"CC",X"0C",X"E6",X"62",X"D0",
		X"E3",X"6A",X"E5",X"62",X"E6",X"2C",X"78",X"CA",X"EE",X"CB",X"54",X"CD",X"74",X"CE",X"2F",X"14",
		X"41",X"08",X"42",X"38",X"44",X"BA",X"44",X"AE",X"45",X"68",X"45",X"F8",X"46",X"2F",X"24",X"C9",
		X"AE",X"42",X"3A",X"44",X"30",X"44",X"48",X"45",X"7C",X"46",X"52",X"46",X"0A",X"EA",X"E2",X"E2",
		X"42",X"7A",X"43",X"FA",X"43",X"72",X"44",X"F2",X"44",X"6A",X"45",X"EA",X"45",X"E2",X"46",X"62",
		X"E6",X"AA",X"7C",X"42",X"74",X"42",X"4C",X"43",X"44",X"43",X"6C",X"44",X"64",X"44",X"5C",X"45",
		X"F4",X"CD",X"DC",X"CE",X"D4",X"CE",X"8C",X"4C",X"43",X"F2",X"42",X"70",X"45",X"EC",X"46",X"2C",
		X"6C",X"42",X"D2",X"43",X"66",X"45",X"5A",X"46",X"2C",X"04",X"E2",X"56",X"E3",X"9E",X"E5",X"CC",
		X"46",X"2C",X"3A",X"CA",X"68",X"CB",X"A0",X"CD",X"F2",X"CE",X"8D",X"CE",X"41",X"C4",X"42",X"DA",
		X"E3",X"B0",X"E5",X"F6",X"E6",X"8D",X"D8",X"41",X"FA",X"42",X"CC",X"43",X"2E",X"45",X"68",X"46",
		X"A8",X"64",X"42",X"FE",X"42",X"50",X"43",X"28",X"44",X"66",X"45",X"A8",X"45",X"FE",X"45",X"7C",
		X"E6",X"A8",X"48",X"42",X"72",X"42",X"C0",X"43",X"16",X"44",X"1E",X"45",X"48",X"45",X"70",X"45",
		X"E2",X"CE",X"8D",X"E6",X"42",X"9C",X"43",X"D2",X"44",X"68",X"46",X"F8",X"46",X"2D",X"D8",X"CA",
		X"8A",X"43",X"EC",X"44",X"78",X"46",X"56",X"46",X"2C",X"92",X"E2",X"B4",X"E2",X"BA",X"E3",X"CA",
		X"46",X"2E",X"90",X"CA",X"B6",X"CA",X"8C",X"CC",X"96",X"CC",X"B8",X"CD",X"F6",X"CE",X"8A",X"A4",
		X"E1",X"D4",X"E6",X"8E",X"26",X"42",X"1C",X"43",X"3C",X"44",X"0C",X"45",X"6C",X"46",X"1E",X"45",
		X"8D",X"2A",X"42",X"AC",X"43",X"2A",X"44",X"AC",X"45",X"6A",X"46",X"2D",X"B4",X"CA",X"BA",X"CB",
		X"14",X"44",X"1A",X"45",X"54",X"46",X"2A",X"B0",X"E5",X"F6",X"E6",X"8C",X"56",X"42",X"BA",X"43",
		X"8A",X"CD",X"48",X"CE",X"08",X"2F",X"0C",X"CA",X"2C",X"CA",X"90",X"CB",X"B0",X"CB",X"C4",X"CC",
		X"C4",X"CC",X"68",X"CE",X"2C",X"EC",X"E2",X"CC",X"E3",X"AA",X"E5",X"FE",X"E6",X"2C",X"58",X"CA",
		X"D0",X"CB",X"9A",X"CD",X"4E",X"CE",X"0C",X"CA",X"62",X"82",X"64",X"96",X"64",X"EA",X"66",X"2C",
		X"DC",X"CA",X"A8",X"CC",X"BC",X"CC",X"5C",X"CE",X"2F",X"7C",X"E2",X"5C",X"E3",X"7C",X"E5",X"9C",
		X"61",X"BC",X"63",X"9C",X"64",X"FC",X"66",X"2F",X"84",X"C9",X"8C",X"CB",X"84",X"CC",X"CC",X"CE",
		X"44",X"CA",X"C4",X"CB",X"44",X"CD",X"09",X"AC",X"E1",X"50",X"E2",X"CC",X"E2",X"DE",X"E2",X"10",
		X"64",X"8C",X"64",X"9E",X"64",X"78",X"66",X"EC",X"66",X"21",X"C2",X"CA",X"82",X"CC",X"9C",X"C9",
		X"DC",X"CA",X"5C",X"CE",X"C0",X"CA",X"80",X"CC",X"70",X"CE",X"9C",X"CC",X"08",X"0C",X"E4",X"74",
		X"65",X"CA",X"62",X"C6",X"61",X"D0",X"62",X"86",X"64",X"68",X"66",X"E4",X"66",X"2E",X"46",X"CA",
		X"FA",X"C9",X"54",X"CE",X"62",X"CD",X"D4",X"CA",X"AA",X"CC",X"2D",X"66",X"E6",X"34",X"E3",X"EA",
		X"66",X"C4",X"64",X"F2",X"66",X"2D",X"4C",X"CE",X"52",X"CC",X"DC",X"CE",X"2A",X"CB",X"78",X"CE",
		X"2A",X"30",X"E4",X"7E",X"E6",X"2E",X"FE",X"C9",X"3E",X"CC",X"26",X"CB",X"40",X"CD",X"14",X"CB",
		X"FC",X"CD",X"1C",X"4A",X"62",X"4A",X"64",X"42",X"61",X"42",X"63",X"62",X"66",X"5A",X"62",X"5A",
		X"E4",X"52",X"E1",X"52",X"E3",X"72",X"E6",X"CA",X"E2",X"CA",X"E4",X"C2",X"E1",X"C2",X"E3",X"E2",
		X"66",X"DA",X"62",X"DA",X"64",X"D2",X"61",X"D2",X"63",X"F2",X"66",X"3C",X"46",X"C9",X"46",X"CB",
		X"6E",X"CE",X"CE",X"CA",X"CA",X"CC",X"FE",X"C9",X"FE",X"CB",X"7E",X"CE",X"DE",X"CA",X"DE",X"CC",
		X"46",X"C9",X"46",X"CB",X"C6",X"CE",X"66",X"CA",X"66",X"CC",X"56",X"C9",X"56",X"CB",X"D6",X"CE",
		X"D6",X"42",X"D6",X"44",X"0C",X"4A",X"E2",X"28",X"E4",X"EE",X"E6",X"5A",X"E2",X"38",X"E4",X"FE",
		X"46",X"CA",X"42",X"80",X"44",X"E6",X"46",X"DA",X"42",X"90",X"44",X"F6",X"46",X"28",X"8B",X"0C",
		X"E4",X"C0",X"E6",X"52",X"E2",X"8B",X"AA",X"44",X"7C",X"46",X"F0",X"42",X"2F",X"2E",X"E2",X"7C",
		X"43",X"E4",X"45",X"86",X"42",X"B6",X"44",X"F2",X"46",X"EC",X"46",X"2F",X"8A",X"CC",X"CE",X"CE",
		X"BA",X"42",X"7C",X"45",X"E4",X"43",X"B2",X"42",X"5C",X"46",X"2E",X"C8",X"E6",X"06",X"E3",X"E4",
		X"45",X"FC",X"46",X"DC",X"42",X"92",X"44",X"2E",X"0C",X"CC",X"6A",X"CA",X"EC",X"CE",X"DA",X"CD",
		X"98",X"43",X"5A",X"46",X"2E",X"4A",X"E2",X"18",X"E4",X"FA",X"E6",X"42",X"E2",X"14",X"E4",X"E2",
		X"46",X"2E",X"2C",X"CC",X"7E",X"CA",X"DE",X"CE",X"C6",X"CE",X"10",X"CC",X"76",X"CA",X"5E",X"E6",
		X"E3",X"E6",X"28",X"E7",X"39",X"E7",X"3E",X"E7",X"1F",X"E7",X"14",X"E7",X"49",X"E7",X"5E",X"E7",
		X"D3",X"E7",X"1C",X"E7",X"25",X"E7",X"36",X"E7",X"57",X"E7",X"AC",X"F8",X"BD",X"F8",X"92",X"F8",
		X"4F",X"D0",X"58",X"D0",X"65",X"D0",X"46",X"D0",X"AB",X"D0",X"B8",X"D0",X"B9",X"D0",X"9E",X"D0",
		X"23",X"F8",X"34",X"F8",X"49",X"F8",X"6A",X"F8",X"7B",X"F8",X"44",X"F8",X"95",X"F9",X"96",X"F9",
		X"6B",X"D1",X"5C",X"D1",X"5D",X"D1",X"2E",X"F4",X"E2",X"F4",X"E3",X"74",X"E3",X"74",X"E4",X"F4",
		X"45",X"F4",X"46",X"26",X"BA",X"CA",X"BA",X"CB",X"3A",X"CB",X"FA",X"CC",X"BA",X"CD",X"FA",X"CE",
		X"54",X"41",X"54",X"42",X"D4",X"42",X"D4",X"43",X"54",X"44",X"54",X"45",X"D4",X"45",X"54",X"46",
		X"88",X"42",X"61",X"42",X"62",X"4C",X"64",X"6C",X"65",X"C4",X"61",X"C4",X"62",X"CE",X"64",X"CE",
		X"E5",X"2A",X"FC",X"CB",X"FC",X"CC",X"2C",X"E8",X"E2",X"E8",X"E3",X"E8",X"E5",X"E8",X"E6",X"26",
		X"C6",X"CA",X"CE",X"CC",X"C6",X"CC",X"CE",X"CE",X"D6",X"C9",X"DE",X"CD",X"D6",X"CD",X"DE",X"CE",
		X"C6",X"CA",X"46",X"CC",X"C6",X"CC",X"46",X"CE",X"D4",X"CB",X"54",X"CE",X"2E",X"76",X"E2",X"56",
		X"64",X"76",X"65",X"76",X"66",X"DA",X"63",X"DA",X"64",X"22",X"9E",X"CA",X"9E",X"CB",X"96",X"CB",
		X"9E",X"CC",X"1E",X"CD",X"5E",X"CE",X"D4",X"CA",X"D4",X"CB",X"D4",X"CD",X"54",X"CE",X"0A",X"76",
		X"61",X"36",X"63",X"EE",X"61",X"AE",X"62",X"16",X"63",X"36",X"64",X"14",X"64",X"74",X"65",X"56",
		X"E5",X"76",X"E6",X"38",X"AE",X"CC",X"6E",X"CE",X"38",X"CA",X"38",X"CB",X"98",X"CC",X"58",X"CD",
		X"D6",X"CD",X"DE",X"CE",X"26",X"CC",X"6E",X"CD",X"36",X"CC",X"7E",X"CE",X"BE",X"CA",X"BE",X"CD",
		X"96",X"CD",X"56",X"CE",X"0C",X"60",X"E4",X"60",X"E6",X"5A",X"E2",X"7A",X"E6",X"16",X"E1",X"76",
		X"66",X"C2",X"62",X"E2",X"66",X"FC",X"64",X"FC",X"66",X"D6",X"65",X"F6",X"66",X"20",X"2A",X"CA",
		X"A2",X"CA",X"2A",X"CB",X"6A",X"CD",X"CE",X"CD",X"4E",X"CE",X"A2",X"CD",X"62",X"CE",X"1C",X"4E",
		X"62",X"6E",X"64",X"4E",X"64",X"6E",X"66",X"46",X"63",X"66",X"66",X"5E",X"62",X"7E",X"64",X"5E",
		X"E4",X"7E",X"E6",X"56",X"E1",X"76",X"E5",X"56",X"E5",X"76",X"E6",X"CE",X"E2",X"EE",X"E4",X"CE",
		X"64",X"EE",X"66",X"C6",X"63",X"E6",X"66",X"DE",X"62",X"FE",X"64",X"DE",X"64",X"FE",X"66",X"D6",
		X"E1",X"F6",X"E5",X"D6",X"E5",X"F6",X"E6",X"22",X"CA",X"CA",X"CA",X"CB",X"FA",X"CD",X"7A",X"CE",
		X"7E",X"62",X"7E",X"66",X"42",X"65",X"62",X"66",X"D4",X"62",X"D4",X"63",X"28",X"CC",X"C4",X"8C",
		X"CD",X"06",X"CD",X"66",X"CE",X"FA",X"CC",X"BA",X"CD",X"98",X"CD",X"F8",X"CE",X"22",X"E8",X"C9",
		X"C0",X"61",X"7C",X"62",X"5C",X"62",X"E6",X"63",X"C6",X"63",X"FC",X"64",X"BC",X"65",X"02",X"65",
		X"E2",X"CE",X"26",X"7C",X"C9",X"5C",X"CB",X"DC",X"CA",X"FC",X"CD",X"44",X"CD",X"64",X"CE",X"12",
		X"C5",X"DA",X"C6",X"C2",X"C2",X"CA",X"C5",X"EA",X"C1",X"E2",X"C3",X"B6",X"C1",X"BE",X"C4",X"0C",
		X"5E",X"CD",X"7E",X"CE",X"C0",X"CD",X"70",X"CE",X"2E",X"18",X"CA",X"38",X"CB",X"8A",X"CC",X"AA",
		X"C5",X"B0",X"C5",X"F8",X"C6",X"0C",X"F2",X"60",X"B2",X"61",X"02",X"65",X"62",X"66",X"2A",X"34",
		X"C9",X"BC",X"CA",X"1E",X"CA",X"3E",X"CB",X"9C",X"CB",X"BC",X"CC",X"1E",X"CC",X"3E",X"CD",X"84",
		X"C5",X"EC",X"C6",X"0E",X"5A",X"62",X"1A",X"63",X"26",X"64",X"26",X"65",X"96",X"65",X"F6",X"66",
		X"28",X"2E",X"7E",X"CC",X"3E",X"CD",X"EE",X"CC",X"AE",X"CD",X"82",X"CD",X"E2",X"CE",X"2E",X"1E",
		X"C1",X"16",X"C4",X"DE",X"C3",X"DE",X"C6",X"3C",X"C5",X"7C",X"C6",X"88",X"2A",X"65",X"6A",X"66",
		X"5E",X"CD",X"7E",X"CE",X"C2",X"CD",X"E2",X"CE",X"BE",X"CD",X"FE",X"CE",X"2A",X"B0",X"CD",X"90",
		X"C5",X"0C",X"E4",X"61",X"C4",X"62",X"C4",X"65",X"E4",X"66",X"28",X"5A",X"C5",X"5A",X"C6",X"96",
		X"CB",X"76",X"CE",X"E4",X"CD",X"E4",X"CE",X"F6",X"CD",X"F6",X"CE",X"2C",X"64",X"C9",X"44",X"C9",
		X"54",X"65",X"74",X"66",X"20",X"48",X"C1",X"40",X"C2",X"48",X"C3",X"40",X"C4",X"48",X"C5",X"48",
		X"CE",X"60",X"CA",X"40",X"CB",X"60",X"CC",X"60",X"CE",X"78",X"C9",X"58",X"CA",X"78",X"CB",X"58",
		X"64",X"58",X"65",X"58",X"66",X"D8",X"62",X"D0",X"63",X"D8",X"64",X"D8",X"66",X"68",X"61",X"60",
		X"E2",X"E8",X"E3",X"C8",X"E4",X"E8",X"E5",X"E8",X"E6",X"E0",X"E2",X"C0",X"E3",X"E0",X"E4",X"E0",
		X"66",X"78",X"61",X"70",X"62",X"78",X"63",X"70",X"64",X"78",X"65",X"78",X"66",X"F8",X"62",X"F0",
		X"E3",X"F0",X"E4",X"F0",X"E6",X"28",X"2E",X"2E",X"E5",X"6E",X"E6",X"16",X"E1",X"76",X"E6",X"F8",
		X"63",X"78",X"66",X"8C",X"48",X"62",X"08",X"64",X"48",X"65",X"48",X"66",X"50",X"63",X"58",X"66",
		X"60",X"CA",X"E0",X"CB",X"60",X"CC",X"60",X"CE",X"F0",X"CB",X"70",X"CE",X"28",X"22",X"2E",X"CC",
		X"06",X"64",X"D8",X"62",X"D0",X"62",X"28",X"64",X"20",X"64",X"EA",X"62",X"E2",X"62",X"20",X"65",
		X"60",X"CE",X"08",X"4D",X"69",X"FA",X"08",X"5D",X"56",X"21",X"30",X"2C",X"A8",X"6B",X"AB",X"F9",
		X"38",X"CE",X"18",X"AE",X"08",X"5D",X"C6",X"0F",X"5D",X"E6",X"88",X"45",X"62",X"43",X"4D",X"58",
		X"72",X"31",X"E8",X"D7",X"29",X"28",X"2B",X"4D",X"33",X"FA",X"CD",X"F5",X"72",X"ED",X"2E",X"29",
		X"4D",X"3B",X"7A",X"C1",X"49",X"4D",X"49",X"7A",X"5D",X"76",X"89",X"DE",X"0F",X"88",X"26",X"08",
		X"DD",X"C6",X"2F",X"5D",X"66",X"20",X"C5",X"62",X"C3",X"4D",X"78",X"FA",X"39",X"68",X"28",X"21",
		X"08",X"0A",X"4D",X"3B",X"7A",X"4D",X"FD",X"7A",X"ED",X"AE",X"09",X"4D",X"3B",X"7A",X"E9",X"49",
		X"CD",X"69",X"72",X"5D",X"56",X"21",X"A8",X"94",X"DD",X"C6",X"2F",X"5D",X"66",X"20",X"2E",X"28",
		X"01",X"2E",X"18",X"45",X"62",X"43",X"4D",X"58",X"7A",X"C5",X"21",X"08",X"09",X"4D",X"3B",X"7A",
		X"CD",X"F5",X"72",X"31",X"E8",X"D7",X"2E",X"2A",X"CD",X"BB",X"72",X"E9",X"C9",X"00",X"CD",X"69",
		X"F2",X"28",X"5D",X"76",X"29",X"B0",X"AE",X"88",X"7E",X"18",X"6B",X"8E",X"F2",X"98",X"5D",X"66",
		X"2F",X"5D",X"66",X"20",X"2E",X"28",X"09",X"2E",X"38",X"45",X"6A",X"43",X"CD",X"78",X"FA",X"C5",
		X"21",X"08",X"A9",X"4D",X"B3",X"7A",X"4D",X"FD",X"F2",X"B9",X"E8",X"08",X"26",X"0B",X"4D",X"3B",
		X"FA",X"C1",X"C9",X"4B",X"29",X"4B",X"66",X"20",X"29",X"2C",X"38",X"29",X"C9",X"39",X"EB",X"BB",
		X"F2",X"5D",X"C6",X"09",X"5D",X"E6",X"AA",X"EE",X"4B",X"30",X"A3",X"6E",X"05",X"4B",X"A1",X"49",
		X"6F",X"C6",X"30",X"AF",X"2F",X"AF",X"4F",X"70",X"E6",X"C8",X"2F",X"AF",X"2F",X"D6",X"C8",X"EF",
		X"CB",X"A4",X"A4",X"45",X"53",X"9A",X"C8",X"72",X"EE",X"09",X"77",X"45",X"72",X"74",X"EE",X"09",
		X"1F",X"75",X"1F",X"3F",X"1F",X"C6",X"B6",X"34",X"47",X"A6",X"28",X"29",X"C9",X"75",X"E6",X"48",
		X"57",X"75",X"6E",X"0A",X"EE",X"BF",X"BB",X"67",X"49",X"75",X"EE",X"40",X"57",X"75",X"7E",X"0A",
		X"E6",X"B7",X"B3",X"67",X"C9",X"32",X"4B",X"48",X"0F",X"2F",X"0F",X"67",X"E6",X"2B",X"F6",X"D0",
		X"E7",X"75",X"EE",X"60",X"FE",X"89",X"C7",X"B9",X"B0",X"42",X"96",X"89",X"26",X"08",X"4B",X"EE",
		X"00",X"2C",X"77",X"BA",X"3B",X"AC",X"23",X"34",X"D6",X"24",X"20",X"DA",X"16",X"D7",X"3A",X"AD",
		X"24",X"49",X"92",X"43",X"C8",X"2F",X"07",X"2F",X"C7",X"C6",X"AB",X"D6",X"50",X"E7",X"D5",X"C6",
		X"C8",X"D6",X"21",X"67",X"29",X"2B",X"28",X"7D",X"7C",X"45",X"B0",X"49",X"DD",X"76",X"3A",X"5D",
		X"56",X"1B",X"4D",X"2A",X"F3",X"5D",X"F3",X"1B",X"80",X"1C",X"5D",X"66",X"AF",X"5D",X"E6",X"88",
		X"3E",X"28",X"F2",X"DE",X"FA",X"BD",X"5F",X"39",X"DD",X"F5",X"2F",X"5D",X"74",X"20",X"DD",X"76",
		X"1C",X"97",X"48",X"5D",X"56",X"1D",X"4D",X"2A",X"7B",X"5D",X"F3",X"1D",X"5D",X"66",X"89",X"5D",
		X"66",X"22",X"3E",X"28",X"B7",X"FA",X"19",X"FB",X"3D",X"57",X"19",X"5D",X"75",X"21",X"DD",X"F4",
		X"8A",X"49",X"2B",X"FF",X"CA",X"3C",X"7B",X"C6",X"8F",X"7F",X"D2",X"4B",X"87",X"4B",X"87",X"4B",
		X"07",X"4B",X"07",X"49",X"E6",X"27",X"5F",X"D2",X"E6",X"D8",X"2F",X"27",X"2F",X"27",X"C9",X"5D",
		X"46",X"8C",X"5D",X"EE",X"1A",X"5D",X"56",X"8B",X"4D",X"E9",X"7B",X"5D",X"F7",X"1A",X"78",X"5D",
		X"CB",X"28",X"DE",X"49",X"DD",X"46",X"0E",X"5D",X"6E",X"3C",X"DD",X"56",X"0F",X"4D",X"41",X"FB",
		X"5D",X"F7",X"1C",X"D8",X"5D",X"4B",X"08",X"D6",X"49",X"71",X"BF",X"70",X"DA",X"13",X"7B",X"97",
		X"D2",X"F5",X"73",X"29",X"4F",X"D3",X"91",X"DA",X"B4",X"FB",X"EB",X"9F",X"73",X"D3",X"B7",X"D0",
		X"DA",X"83",X"7B",X"89",X"47",X"D2",X"7D",X"7B",X"6B",X"37",X"7B",X"89",X"47",X"52",X"7D",X"7B",
		X"EB",X"9C",X"73",X"BF",X"F2",X"89",X"73",X"29",X"4F",X"D1",X"93",X"FA",X"B7",X"FB",X"EB",X"9C",
		X"7B",X"73",X"BF",X"70",X"FA",X"A7",X"7B",X"89",X"47",X"52",X"91",X"7B",X"6B",X"37",X"7B",X"89",
		X"4F",X"FA",X"99",X"FB",X"53",X"B7",X"C9",X"D1",X"B7",X"49",X"DD",X"D6",X"3C",X"94",X"D2",X"40",
		X"7B",X"56",X"39",X"5D",X"F7",X"1C",X"58",X"35",X"5D",X"F7",X"1C",X"49",X"4D",X"64",X"7B",X"C5",
		X"CD",X"D6",X"73",X"11",X"0C",X"4B",X"66",X"80",X"D2",X"E9",X"51",X"2F",X"AF",X"2F",X"4E",X"4B",
		X"91",X"99",X"95",X"49",X"5D",X"66",X"09",X"5D",X"E6",X"0A",X"46",X"2D",X"4B",X"31",X"39",X"4B",
		X"11",X"4B",X"11",X"61",X"2C",X"FD",X"E6",X"D0",X"0F",X"07",X"0F",X"47",X"F1",X"49",X"ED",X"4D",
		X"F8",X"7A",X"69",X"B9",X"E8",X"08",X"D0",X"4B",X"E6",X"20",X"AE",X"EF",X"11",X"2C",X"6B",X"0F",
		X"FC",X"B8",X"29",X"49",X"19",X"2C",X"CB",X"E6",X"20",X"D9",X"38",X"D0",X"C9",X"BE",X"4F",X"8F",
		X"2F",X"8F",X"B0",X"09",X"34",X"8F",X"2E",X"A3",X"57",X"6E",X"A3",X"AE",X"A8",X"45",X"B8",X"49",
		X"B7",X"5D",X"35",X"3E",X"E8",X"5D",X"70",X"3E",X"F5",X"5D",X"56",X"38",X"6F",X"8F",X"5F",X"BE",
		X"A8",X"39",X"D6",X"A3",X"5D",X"F7",X"A9",X"76",X"5D",X"F7",X"AA",X"D1",X"BF",X"70",X"A0",X"88",
		X"14",X"11",X"10",X"23",X"87",X"CB",X"77",X"FC",X"FE",X"29",X"17",X"30",X"2A",X"71",X"15",X"5D",
		X"F7",X"18",X"97",X"49",X"A1",X"FB",X"F4",X"B9",X"A8",X"67",X"21",X"39",X"A8",X"45",X"B8",X"A1",
		X"F3",X"FC",X"39",X"5D",X"48",X"A9",X"2B",X"28",X"C5",X"90",X"C9",X"28",X"38",X"28",X"28",X"21",
		X"A8",X"08",X"28",X"08",X"A8",X"0F",X"A8",X"08",X"AE",X"08",X"A8",X"0D",X"A8",X"08",X"AC",X"08",
		X"2B",X"2B",X"2B",X"2A",X"2A",X"2A",X"29",X"60",X"74",X"61",X"61",X"6B",X"61",X"71",X"74",X"63",
		X"6B",X"5C",X"EF",X"CD",X"7C",X"5C",X"FB",X"4D",X"A0",X"28",X"EF",X"49",X"92",X"08",X"C8",X"4B",
		X"6F",X"CA",X"66",X"FE",X"CD",X"4C",X"FE",X"56",X"2F",X"D8",X"32",X"B9",X"CF",X"4D",X"E8",X"FF",
		X"A1",X"08",X"C7",X"B9",X"DD",X"40",X"21",X"0B",X"A8",X"45",X"B8",X"36",X"8B",X"4D",X"B5",X"4D",
		X"12",X"B9",X"CF",X"34",X"F6",X"20",X"08",X"32",X"B9",X"CF",X"CD",X"34",X"F0",X"A2",X"BA",X"CF",
		X"F6",X"76",X"FD",X"B9",X"28",X"08",X"11",X"76",X"FD",X"4D",X"52",X"7C",X"F9",X"6F",X"F9",X"22",
		X"BA",X"CF",X"76",X"F7",X"39",X"20",X"28",X"39",X"71",X"49",X"12",X"B9",X"CF",X"6F",X"AF",X"D5",
		X"29",X"6F",X"26",X"08",X"A1",X"9C",X"67",X"29",X"B6",X"DE",X"59",X"B9",X"8B",X"1E",X"F9",X"8B",
		X"5F",X"21",X"28",X"28",X"C5",X"63",X"35",X"CF",X"2C",X"59",X"12",X"BD",X"E7",X"EE",X"20",X"D6",
		X"80",X"0A",X"96",X"DD",X"59",X"4D",X"04",X"F8",X"59",X"32",X"09",X"40",X"06",X"08",X"26",X"08",
		X"CB",X"67",X"00",X"2E",X"CB",X"D7",X"20",X"2A",X"0E",X"2C",X"C5",X"D0",X"5F",X"92",X"34",X"CF",
		X"94",X"B2",X"3C",X"67",X"4D",X"09",X"F8",X"32",X"3C",X"67",X"94",X"B2",X"3C",X"67",X"4D",X"09",
		X"50",X"CD",X"50",X"9B",X"20",X"2B",X"14",X"A0",X"12",X"92",X"36",X"CF",X"D6",X"2F",X"30",X"A0",
		X"59",X"2E",X"08",X"59",X"8F",X"5B",X"88",X"27",X"47",X"4B",X"71",X"B2",X"0E",X"40",X"A0",X"98",
		X"E6",X"B8",X"CA",X"32",X"75",X"B2",X"2E",X"48",X"12",X"78",X"E8",X"BF",X"CA",X"32",X"75",X"DE",
		X"0A",X"B0",X"0D",X"4B",X"E1",X"4A",X"9A",X"7D",X"D6",X"56",X"DE",X"20",X"0B",X"56",X"DF",X"C8",
		X"36",X"75",X"C9",X"95",X"07",X"57",X"E6",X"2A",X"2F",X"BB",X"5F",X"4B",X"7B",X"6A",X"EF",X"FD",
		X"59",X"4B",X"39",X"59",X"4B",X"73",X"6A",X"1A",X"7E",X"59",X"4B",X"11",X"59",X"4B",X"F3",X"CA",
		X"30",X"FE",X"D9",X"4B",X"B1",X"59",X"EB",X"71",X"75",X"8F",X"32",X"BE",X"E7",X"6B",X"1A",X"FD",
		X"8F",X"B2",X"3D",X"67",X"6B",X"B1",X"7D",X"59",X"4B",X"F9",X"59",X"CA",X"40",X"7D",X"59",X"4B",
		X"F9",X"59",X"16",X"03",X"CD",X"BD",X"6D",X"D6",X"D6",X"77",X"20",X"30",X"16",X"75",X"77",X"59",
		X"4D",X"04",X"F8",X"BD",X"25",X"59",X"83",X"CA",X"B1",X"7D",X"59",X"BC",X"24",X"59",X"A3",X"B6",
		X"5F",X"6B",X"91",X"FD",X"D6",X"76",X"20",X"20",X"16",X"75",X"77",X"59",X"CD",X"0C",X"50",X"49",
		X"D6",X"A3",X"59",X"4D",X"8C",X"F8",X"34",X"AC",X"D0",X"59",X"DE",X"0C",X"78",X"B6",X"7E",X"CB",
		X"91",X"FD",X"D9",X"4B",X"51",X"59",X"00",X"20",X"12",X"BD",X"CF",X"56",X"27",X"5A",X"91",X"FD",
		X"59",X"4B",X"D9",X"59",X"D6",X"35",X"DE",X"49",X"B0",X"0A",X"96",X"DF",X"F7",X"CB",X"C8",X"7D",
		X"D9",X"4B",X"71",X"59",X"00",X"20",X"12",X"BD",X"CF",X"56",X"27",X"5A",X"91",X"FD",X"D9",X"4B",
		X"F9",X"59",X"D6",X"34",X"DE",X"68",X"A0",X"0A",X"96",X"49",X"F7",X"CB",X"C8",X"7D",X"4D",X"68",
		X"FF",X"2E",X"2C",X"07",X"32",X"B9",X"CF",X"4D",X"34",X"F0",X"22",X"BA",X"CF",X"F6",X"56",X"D5",
		X"31",X"88",X"A8",X"39",X"D6",X"D5",X"26",X"0E",X"50",X"3D",X"36",X"08",X"A1",X"B6",X"70",X"39",
		X"56",X"22",X"BA",X"CF",X"E5",X"B9",X"20",X"28",X"19",X"F6",X"5F",X"07",X"DB",X"20",X"07",X"C6",
		X"B0",X"B2",X"AE",X"40",X"D3",X"20",X"3A",X"32",X"F8",X"40",X"BF",X"73",X"80",X"1B",X"92",X"58",
		X"48",X"56",X"2A",X"B0",X"20",X"32",X"2E",X"48",X"CB",X"E7",X"53",X"20",X"2C",X"C1",X"F1",X"D1",
		X"49",X"F6",X"F7",X"C1",X"F7",X"B8",X"C9",X"CD",X"ED",X"4D",X"91",X"8B",X"E9",X"C9",X"F9",X"28",
		X"F1",X"F7",X"39",X"20",X"28",X"39",X"08",X"F7",X"12",X"B9",X"CF",X"34",X"D6",X"2F",X"20",X"1C",
		X"05",X"A0",X"98",X"49",X"ED",X"55",X"E9",X"A1",X"A8",X"67",X"31",X"0B",X"A8",X"AE",X"AF",X"6A",
		X"D5",X"76",X"28",X"16",X"30",X"2F",X"19",X"2C",X"38",X"D1",X"16",X"D7",X"C9",X"CA",X"D2",X"FE",
		X"ED",X"A3",X"DD",X"76",X"A9",X"16",X"B0",X"0F",X"E9",X"55",X"D6",X"08",X"6B",X"56",X"F6",X"CA",
		X"D1",X"FE",X"23",X"55",X"56",X"2A",X"96",X"30",X"C7",X"C1",X"51",X"43",X"21",X"3C",X"CF",X"97",
		X"CD",X"FA",X"64",X"6D",X"31",X"1C",X"67",X"20",X"9F",X"CD",X"A1",X"19",X"67",X"45",X"98",X"C9",
		X"39",X"B8",X"E7",X"A1",X"05",X"CF",X"C5",X"98",X"39",X"33",X"E7",X"A1",X"1A",X"CF",X"6F",X"96",
		X"0F",X"98",X"47",X"70",X"26",X"08",X"CD",X"10",X"47",X"8F",X"29",X"7F",X"36",X"08",X"A1",X"9C",
		X"E7",X"11",X"51",X"06",X"2A",X"B6",X"5D",X"55",X"7C",X"33",X"C5",X"B8",X"4F",X"A1",X"3D",X"CF",
		X"36",X"08",X"57",X"39",X"92",X"88",X"40",X"CE",X"09",X"A7",X"F7",X"71",X"A1",X"08",X"67",X"8F",
		X"A9",X"57",X"51",X"36",X"28",X"11",X"C3",X"DD",X"E5",X"E9",X"29",X"2B",X"28",X"CD",X"B0",X"49",
		X"A1",X"AA",X"F8",X"AE",X"0B",X"36",X"88",X"CD",X"4D",X"11",X"F8",X"A3",X"69",X"B8",X"F0",X"34",
		X"CD",X"19",X"50",X"A3",X"D6",X"27",X"20",X"DF",X"21",X"28",X"E7",X"16",X"0B",X"96",X"09",X"36",
		X"8B",X"28",X"26",X"0B",X"D6",X"97",X"A0",X"0D",X"34",X"BC",X"A3",X"B8",X"77",X"56",X"18",X"30",
		X"0D",X"47",X"2F",X"27",X"2F",X"27",X"E6",X"27",X"F6",X"B8",X"CD",X"0C",X"50",X"D1",X"3C",X"EE",
		X"8F",X"D6",X"38",X"4D",X"04",X"F8",X"34",X"A3",X"D6",X"B8",X"66",X"36",X"38",X"4D",X"04",X"F8",
		X"1C",X"14",X"08",X"94",X"D6",X"38",X"EA",X"F7",X"77",X"A1",X"3D",X"CF",X"39",X"23",X"3B",X"96",
		X"89",X"28",X"D6",X"EF",X"27",X"AF",X"27",X"AF",X"EE",X"8F",X"FE",X"38",X"4D",X"04",X"F8",X"BC",
		X"50",X"EE",X"0F",X"FE",X"30",X"4D",X"AC",X"F0",X"3D",X"14",X"1C",X"A3",X"08",X"94",X"D6",X"38",
		X"A0",X"D7",X"A1",X"9C",X"67",X"3E",X"8B",X"36",X"89",X"BE",X"1E",X"28",X"26",X"0B",X"D6",X"4D",
		X"AC",X"F0",X"23",X"34",X"38",X"D0",X"1C",X"14",X"08",X"94",X"D6",X"38",X"20",X"C3",X"EB",X"D3",
		X"29",X"C5",X"7D",X"22",X"B2",X"67",X"ED",X"B9",X"28",X"08",X"11",X"32",X"B4",X"67",X"F6",X"F7",
		X"E1",X"F7",X"02",X"BD",X"CF",X"A3",X"22",X"BD",X"CF",X"D9",X"E1",X"49",X"AF",X"8F",X"AF",X"8F",
		X"C7",X"A6",X"A8",X"21",X"81",X"B9",X"69",X"D2",X"11",X"49",X"AB",X"8D",X"EE",X"CC",X"69",X"4B",
		X"63",X"71",X"28",X"2E",X"21",X"7B",X"7D",X"78",X"6D",X"7A",X"A8",X"78",X"64",X"69",X"71",X"6D",
		X"FA",X"5B",X"A8",X"89",X"AE",X"5A",X"E9",X"CE",X"6B",X"28",X"A0",X"28",X"FB",X"4B",X"6F",X"5A",
		X"6D",X"A8",X"7A",X"6C",X"74",X"66",X"69",X"65",X"6D",X"28",X"23",X"2F",X"B9",X"7B",X"7C",X"28",
		X"2D",X"0F",X"B2",X"CE",X"EC",X"08",X"2F",X"0F",X"B3",X"5A",X"EC",X"08",X"B9",X"0F",X"B4",X"5C",
		X"60",X"28",X"3B",X"2F",X"BD",X"7C",X"60",X"28",X"3D",X"2F",X"BE",X"7C",X"60",X"28",X"3F",X"2F",
		X"B7",X"5C",X"68",X"08",X"ED",X"CD",X"4D",X"A0",X"70",X"F7",X"A3",X"28",X"F7",X"28",X"69",X"C1",
		X"C9",X"28",X"87",X"7E",X"23",X"FE",X"23",X"C5",X"CD",X"80",X"F0",X"43",X"E1",X"28",X"C5",X"80",
		X"32",X"BB",X"00",X"16",X"A0",X"77",X"00",X"49",X"FD",X"DD",X"C3",X"A6",X"A8",X"21",X"81",X"21",
		X"01",X"21",X"01",X"72",X"2F",X"8D",X"47",X"B9",X"28",X"C0",X"19",X"D9",X"F1",X"49",X"28",X"2F",
		X"57",X"BF",X"57",X"0F",X"ED",X"32",X"1C",X"F9",X"B2",X"3F",X"C8",X"B2",X"65",X"40",X"31",X"C9",
		X"52",X"A1",X"14",X"F1",X"2E",X"2C",X"56",X"F6",X"3A",X"C5",X"21",X"20",X"28",X"39",X"C3",X"C1",
		X"32",X"A3",X"ED",X"A1",X"30",X"08",X"11",X"43",X"E9",X"B8",X"43",X"C1",X"CB",X"A1",X"E7",X"F9",
		X"29",X"D7",X"24",X"36",X"21",X"4D",X"E8",X"F1",X"21",X"EE",X"28",X"39",X"C3",X"32",X"2C",X"48",
		X"EE",X"38",X"07",X"2F",X"07",X"A1",X"7B",X"F9",X"47",X"AE",X"08",X"29",X"D6",X"A3",X"E6",X"67",
		X"16",X"22",X"E5",X"A1",X"5C",X"F0",X"CD",X"6F",X"51",X"E9",X"2E",X"2A",X"CD",X"E8",X"51",X"4D",
		X"58",X"F9",X"94",X"C5",X"A1",X"6A",X"F8",X"4D",X"4F",X"F9",X"E9",X"AE",X"0A",X"4D",X"68",X"F9",
		X"CD",X"78",X"51",X"94",X"E5",X"A1",X"40",X"F0",X"CD",X"6F",X"51",X"E9",X"2E",X"2A",X"CD",X"E8",
		X"F9",X"4D",X"58",X"F9",X"6B",X"F7",X"68",X"A9",X"F7",X"0B",X"4D",X"68",X"F9",X"BB",X"33",X"49",
		X"E5",X"A1",X"BB",X"F1",X"2E",X"21",X"CD",X"E8",X"51",X"A1",X"22",X"28",X"19",X"CB",X"E1",X"49",
		X"CD",X"80",X"32",X"BB",X"30",X"F2",X"49",X"4D",X"D8",X"5C",X"5A",X"49",X"28",X"58",X"CC",X"49",
		X"59",X"6D",X"7A",X"F3",X"51",X"09",X"51",X"0F",X"51",X"05",X"51",X"A8",X"33",X"A8",X"10",X"B9",
		X"3E",X"28",X"3B",X"39",X"38",X"3A",X"38",X"28",X"3C",X"39",X"3A",X"3A",X"3C",X"28",X"3C",X"39",
		X"34",X"BA",X"10",X"B8",X"30",X"B8",X"30",X"A8",X"78",X"7C",X"7B",X"74",X"C7",X"B0",X"17",X"D0",
		X"8F",X"DB",X"98",X"4D",X"A7",X"F9",X"4D",X"76",X"FA",X"4D",X"D2",X"FB",X"6B",X"D9",X"FC",X"4D",
		X"AD",X"F2",X"21",X"28",X"E0",X"21",X"28",X"38",X"CD",X"B8",X"52",X"B0",X"0A",X"96",X"28",X"4D",
		X"E1",X"FA",X"96",X"09",X"4D",X"E1",X"FA",X"A1",X"08",X"D0",X"21",X"08",X"88",X"4D",X"38",X"FA",
		X"16",X"2A",X"DC",X"C1",X"52",X"A1",X"28",X"48",X"29",X"28",X"38",X"4D",X"30",X"F2",X"16",X"2B",
		X"5C",X"E1",X"FA",X"A1",X"08",X"50",X"21",X"08",X"88",X"4D",X"38",X"FA",X"B0",X"1C",X"96",X"0C",
		X"CD",X"C1",X"52",X"96",X"2D",X"4D",X"C1",X"F2",X"16",X"2E",X"CD",X"C1",X"52",X"96",X"2F",X"4D",
		X"41",X"FA",X"4D",X"D4",X"74",X"4D",X"C7",X"FC",X"90",X"F3",X"4D",X"37",X"72",X"A1",X"A0",X"08",
		X"D9",X"A1",X"28",X"28",X"CD",X"6A",X"F2",X"36",X"28",X"5C",X"C1",X"F2",X"21",X"28",X"68",X"4D",
		X"EA",X"FA",X"96",X"09",X"5C",X"E1",X"72",X"4D",X"5C",X"FC",X"4D",X"67",X"74",X"30",X"53",X"49",
		X"56",X"FF",X"07",X"F7",X"07",X"8E",X"D6",X"D7",X"37",X"C8",X"72",X"A3",X"0B",X"70",X"B1",X"A0",
		X"47",X"49",X"21",X"08",X"A0",X"4D",X"FF",X"FA",X"D3",X"59",X"9E",X"A3",X"A0",X"0C",X"59",X"72",
		X"D9",X"16",X"23",X"59",X"C8",X"B7",X"C9",X"B9",X"28",X"28",X"E5",X"DD",X"39",X"A8",X"28",X"87",
		X"CD",X"FA",X"79",X"C1",X"A0",X"0B",X"A3",X"A3",X"03",X"73",X"8E",X"7F",X"A3",X"72",X"8E",X"FF",
		X"23",X"4B",X"12",X"4B",X"1B",X"B0",X"20",X"72",X"C6",X"00",X"7F",X"73",X"C6",X"38",X"5F",X"2B",
		X"D0",X"91",X"A0",X"56",X"49",X"4D",X"2B",X"FD",X"4D",X"61",X"74",X"A1",X"1D",X"FD",X"4D",X"39",
		X"F5",X"A1",X"8B",X"F5",X"CD",X"B9",X"F5",X"45",X"5B",X"82",X"F5",X"A1",X"84",X"F5",X"2E",X"20",
		X"4D",X"DA",X"75",X"A1",X"07",X"FD",X"26",X"88",X"4D",X"E8",X"75",X"45",X"53",X"D3",X"75",X"A1",
		X"55",X"F5",X"2E",X"20",X"EB",X"72",X"F5",X"4D",X"23",X"F5",X"CD",X"C9",X"F4",X"A1",X"CA",X"F5",
		X"4D",X"39",X"75",X"A1",X"83",X"FD",X"4D",X"39",X"75",X"45",X"53",X"A2",X"75",X"A1",X"04",X"FD",
		X"2E",X"2A",X"CD",X"72",X"F5",X"A1",X"C0",X"F5",X"2E",X"2A",X"CD",X"E0",X"F5",X"45",X"5B",X"53",
		X"75",X"A1",X"5D",X"FD",X"26",X"0A",X"6B",X"DA",X"75",X"45",X"53",X"D3",X"75",X"8F",X"2B",X"7F",
		X"21",X"DC",X"F5",X"CB",X"BD",X"F5",X"CD",X"D7",X"F4",X"4D",X"23",X"F5",X"87",X"5B",X"38",X"4B",
		X"D7",X"20",X"0B",X"07",X"5B",X"8D",X"59",X"6F",X"59",X"4D",X"9A",X"FB",X"4D",X"69",X"FB",X"58",
		X"D9",X"4B",X"69",X"59",X"EC",X"88",X"53",X"B0",X"F0",X"49",X"87",X"5B",X"38",X"4B",X"57",X"80",
		X"0B",X"07",X"5B",X"8D",X"59",X"11",X"47",X"59",X"6C",X"8B",X"FD",X"A1",X"F1",X"FD",X"26",X"0F",
		X"CD",X"E0",X"55",X"4D",X"7D",X"F3",X"21",X"B2",X"56",X"26",X"2D",X"4D",X"71",X"F5",X"D9",X"4B",
		X"61",X"59",X"48",X"A1",X"DD",X"FE",X"4D",X"39",X"FD",X"A1",X"BE",X"FE",X"31",X"08",X"8A",X"AE",
		X"2C",X"4D",X"71",X"F5",X"C9",X"59",X"CB",X"61",X"D9",X"31",X"28",X"28",X"E8",X"31",X"28",X"2D",
		X"49",X"07",X"5B",X"88",X"31",X"0D",X"1B",X"AE",X"0E",X"A1",X"69",X"FE",X"07",X"B0",X"0C",X"A1",
		X"64",X"F6",X"B7",X"00",X"ED",X"7D",X"CD",X"BD",X"55",X"79",X"E9",X"D0",X"D6",X"2D",X"20",X"2D",
		X"00",X"2F",X"97",X"28",X"25",X"28",X"58",X"28",X"D3",X"CE",X"0A",X"7F",X"00",X"B8",X"D2",X"4D",
		X"7D",X"F3",X"C3",X"8F",X"DB",X"28",X"39",X"39",X"0E",X"11",X"C3",X"4D",X"83",X"F3",X"B7",X"49",
		X"8F",X"5B",X"0C",X"B9",X"19",X"98",X"4D",X"A3",X"FB",X"97",X"49",X"27",X"47",X"AF",X"27",X"AF",
		X"E6",X"2E",X"6F",X"D1",X"0F",X"EE",X"29",X"B8",X"6F",X"D1",X"0F",X"07",X"E6",X"29",X"B0",X"47",
		X"26",X"0B",X"A1",X"69",X"FE",X"4B",X"91",X"30",X"0B",X"A1",X"6C",X"FE",X"6D",X"DD",X"4D",X"3D",
		X"55",X"79",X"E9",X"D3",X"EE",X"2A",X"5F",X"30",X"C1",X"49",X"CD",X"D7",X"54",X"4D",X"0B",X"F5",
		X"8F",X"DB",X"98",X"A1",X"6F",X"FE",X"26",X"0B",X"4D",X"E8",X"FD",X"A1",X"00",X"FE",X"8F",X"28",
		X"16",X"38",X"18",X"2D",X"76",X"F6",X"87",X"5B",X"08",X"4B",X"67",X"4C",X"0C",X"F4",X"CB",X"C7",
		X"4C",X"8C",X"74",X"4B",X"77",X"A0",X"45",X"F6",X"8F",X"DB",X"38",X"49",X"8F",X"DB",X"39",X"DB",
		X"30",X"F6",X"CD",X"A7",X"F4",X"32",X"F7",X"F6",X"4F",X"43",X"56",X"DB",X"30",X"A3",X"08",X"CE",
		X"A9",X"A7",X"99",X"30",X"AC",X"07",X"A1",X"00",X"76",X"28",X"4D",X"CE",X"74",X"35",X"49",X"B9",
		X"8C",X"C4",X"C3",X"28",X"4F",X"28",X"51",X"C6",X"D8",X"AF",X"2F",X"AF",X"2F",X"D6",X"B8",X"F7",
		X"A3",X"B6",X"A8",X"A3",X"D1",X"C6",X"2F",X"D6",X"B0",X"F7",X"A3",X"B6",X"A8",X"49",X"F6",X"F6",
		X"87",X"5B",X"20",X"27",X"E6",X"B8",X"20",X"DE",X"C9",X"4D",X"D7",X"F4",X"CD",X"23",X"F5",X"A1",
		X"AA",X"E0",X"96",X"29",X"31",X"09",X"A8",X"EB",X"4D",X"54",X"74",X"AE",X"3C",X"36",X"A2",X"4D",
		X"5C",X"F4",X"16",X"AB",X"6B",X"B9",X"B7",X"28",X"CD",X"5C",X"F4",X"36",X"A0",X"AE",X"32",X"4D",
		X"DC",X"FC",X"96",X"2E",X"26",X"09",X"31",X"F5",X"57",X"4D",X"DC",X"FC",X"96",X"2D",X"26",X"9C",
		X"CD",X"5C",X"F4",X"36",X"AC",X"AE",X"29",X"B9",X"97",X"D7",X"CD",X"5C",X"F4",X"36",X"AF",X"AE",
		X"3A",X"4D",X"DC",X"FC",X"A1",X"10",X"76",X"B9",X"A9",X"D0",X"96",X"0C",X"21",X"0F",X"A8",X"45",
		X"B0",X"43",X"29",X"21",X"28",X"29",X"C3",X"35",X"EA",X"84",X"F4",X"A1",X"84",X"F6",X"39",X"28",
		X"D8",X"36",X"AC",X"A9",X"28",X"08",X"CD",X"90",X"CB",X"A9",X"28",X"08",X"01",X"43",X"95",X"A0",
		X"DD",X"CB",X"CF",X"F4",X"77",X"A3",X"36",X"28",X"19",X"B8",X"D1",X"49",X"87",X"DB",X"31",X"53",
		X"49",X"D3",X"96",X"18",X"7B",X"99",X"49",X"07",X"5B",X"88",X"4B",X"FF",X"B7",X"48",X"F6",X"07",
		X"DB",X"20",X"CB",X"FF",X"20",X"D0",X"76",X"07",X"DB",X"20",X"CB",X"FF",X"20",X"C1",X"C9",X"F6",
		X"F6",X"F6",X"8F",X"5B",X"88",X"27",X"EE",X"0C",X"A0",X"75",X"49",X"4D",X"61",X"FC",X"A1",X"08",
		X"F8",X"31",X"29",X"58",X"29",X"D7",X"3E",X"B6",X"28",X"CD",X"B0",X"A1",X"28",X"58",X"39",X"28",
		X"E0",X"A9",X"08",X"88",X"CD",X"90",X"96",X"F7",X"B2",X"89",X"D2",X"B2",X"19",X"D2",X"6B",X"D4",
		X"54",X"56",X"23",X"76",X"23",X"ED",X"CD",X"6C",X"55",X"CB",X"E1",X"8F",X"C5",X"A8",X"3A",X"33",
		X"9E",X"A0",X"F1",X"49",X"FD",X"DD",X"C3",X"A6",X"08",X"21",X"81",X"21",X"81",X"21",X"81",X"72",
		X"2F",X"BD",X"47",X"31",X"28",X"C0",X"19",X"79",X"F1",X"49",X"ED",X"7D",X"E5",X"4D",X"35",X"F5",
		X"E9",X"D9",X"69",X"3C",X"14",X"B8",X"73",X"49",X"6D",X"4D",X"39",X"FD",X"A3",X"C9",X"30",X"F0",
		X"C9",X"6D",X"FD",X"46",X"23",X"66",X"23",X"CB",X"09",X"CB",X"CD",X"BD",X"55",X"A3",X"F9",X"69",
		X"30",X"E7",X"49",X"DD",X"6D",X"BE",X"08",X"A9",X"48",X"08",X"4D",X"10",X"FD",X"C9",X"79",X"49",
		X"E5",X"4D",X"6C",X"F5",X"7C",X"55",X"3B",X"B6",X"28",X"CD",X"B0",X"E9",X"C9",X"2B",X"0C",X"7A",
		X"49",X"CD",X"08",X"0B",X"18",X"5C",X"4D",X"5B",X"5C",X"08",X"0F",X"89",X"C9",X"4B",X"08",X"0F",
		X"0C",X"BF",X"33",X"28",X"09",X"24",X"10",X"BC",X"28",X"23",X"0C",X"B0",X"35",X"28",X"0D",X"24",
		X"B8",X"B9",X"08",X"8F",X"8C",X"39",X"38",X"38",X"08",X"19",X"8C",X"39",X"38",X"39",X"08",X"1B",
		X"0C",X"B9",X"30",X"BA",X"28",X"3D",X"0C",X"B9",X"30",X"BB",X"28",X"2F",X"3A",X"6F",X"4F",X"67",
		X"4C",X"08",X"0B",X"8C",X"5A",X"CF",X"CD",X"08",X"0F",X"8C",X"39",X"39",X"B9",X"08",X"89",X"8C",
		X"31",X"B8",X"36",X"28",X"6A",X"69",X"6C",X"A8",X"28",X"2A",X"0B",X"61",X"4E",X"78",X"7D",X"7C",
		X"A8",X"0A",X"B9",X"5C",X"ED",X"5B",X"FC",X"08",X"AD",X"8C",X"EB",X"CF",X"69",X"CE",X"A0",X"39",
		X"28",X"2F",X"24",X"6B",X"67",X"61",X"66",X"A8",X"BA",X"28",X"21",X"23",X"7B",X"6D",X"7A",X"7E",
		X"69",X"4B",X"ED",X"08",X"2B",X"8A",X"B1",X"58",X"A0",X"5B",X"FC",X"49",X"FA",X"5C",X"A8",X"8D",
		X"22",X"BA",X"78",X"A8",X"7B",X"7C",X"69",X"7A",X"7C",X"28",X"27",X"2F",X"B9",X"28",X"27",X"21",
		X"F8",X"CC",X"E9",X"D9",X"ED",X"5A",X"A8",X"19",X"28",X"CA",X"FD",X"CD",X"F8",X"08",X"BB",X"0F",
		X"7A",X"61",X"6F",X"60",X"7C",X"28",X"3D",X"20",X"64",X"6D",X"6E",X"7C",X"28",X"27",X"39",X"BA",
		X"A8",X"CF",X"6E",X"08",X"A0",X"28",X"A8",X"89",X"2B",X"5B",X"6F",X"5D",X"6E",X"4C",X"A8",X"89",
		X"39",X"7C",X"6D",X"7B",X"7C",X"28",X"3A",X"24",X"7B",X"67",X"7D",X"66",X"6C",X"A8",X"28",X"3E",
		X"89",X"02",X"8B",X"04",X"8D",X"06",X"8F",X"80",X"09",X"82",X"0B",X"86",X"0F",X"10",X"99",X"13",
		X"2F",X"B0",X"B7",X"48",X"4F",X"D0",X"D7",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"20",X"38",
		X"38",X"28",X"20",X"38",X"30",X"48",X"E8",X"48",X"88",X"00",X"C8",X"40",X"B8",X"BF",X"B0",X"08",
		X"28",X"28",X"1E",X"F7",X"68",X"E7",X"B8",X"28",X"28",X"28",X"1E",X"F7",X"F8",X"17",X"B8",X"28",
		X"A8",X"08",X"9E",X"FF",X"80",X"C7",X"B0",X"08",X"A8",X"08",X"9E",X"FF",X"A8",X"08",X"57",X"F7",
		X"28",X"28",X"D7",X"D7",X"28",X"28",X"D7",X"D7",X"28",X"28",X"D7",X"D7",X"31",X"39",X"38",X"34",
		X"2F",X"30",X"35",X"2F",X"32",X"34",X"20",X"53",X"45",X"47",X"41",X"20",X"52",X"2F",X"44",X"20",
		X"5B",X"5B",X"20",X"46",X"4C",X"49",X"43",X"4B",X"59",X"20",X"21",X"21",X"5D",X"5D",X"20",X"20",
		X"4F",X"4C",X"44",X"20",X"4E",X"41",X"4D",X"45",X"20",X"31",X"29",X"20",X"42",X"55",X"53",X"54",
		X"59",X"20",X"32",X"29",X"20",X"46",X"4C",X"49",X"50",X"50",X"20",X"50",X"52",X"4F",X"47",X"52",
		X"41",X"4D",X"45",X"44",X"20",X"42",X"59",X"20",X"48",X"49",X"44",X"45",X"4B",X"49",X"2E",X"49",
		X"53",X"48",X"49",X"4B",X"41",X"57",X"41",X"20",X"53",X"48",X"55",X"49",X"43",X"48",X"49",X"2E",
		X"4B",X"41",X"54",X"41",X"47",X"49",X"20",X"47",X"41",X"4D",X"45",X"20",X"44",X"45",X"53",X"49",
		X"47",X"4E",X"45",X"44",X"20",X"42",X"59",X"20",X"59",X"4F",X"4A",X"49",X"2E",X"49",X"53",X"48",
		X"49",X"49",X"20",X"43",X"48",X"41",X"52",X"41",X"43",X"54",X"4F",X"52",X"20",X"44",X"45",X"53",
		X"49",X"47",X"4E",X"45",X"44",X"20",X"42",X"59",X"20",X"59",X"4F",X"53",X"48",X"49",X"4B",X"49",
		X"2E",X"4B",X"41",X"57",X"41",X"53",X"41",X"4B",X"49",X"20",X"53",X"45",X"43",X"55",X"52",X"49",
		X"54",X"59",X"20",X"42",X"59",X"20",X"53",X"2E",X"4B",X"41",X"54",X"41",X"47",X"49",X"20",X"41",
		X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",
		X"44",X"20",X"5B",X"5B",X"20",X"44",X"4F",X"4E",X"27",X"54",X"20",X"43",X"4F",X"50",X"59",X"20",
		X"21",X"21",X"20",X"5D",X"5D",X"20",X"5B",X"5B",X"20",X"44",X"4F",X"4E",X"27",X"54",X"20",X"43",
		X"4F",X"50",X"59",X"20",X"21",X"21",X"20",X"5D",X"5D",X"20",X"5B",X"5B",X"20",X"44",X"4F",X"4E",
		X"27",X"54",X"20",X"43",X"4F",X"50",X"59",X"20",X"21",X"21",X"20",X"5D",X"5D",X"20",X"5B",X"5B",
		X"20",X"44",X"4F",X"4E",X"27",X"54",X"20",X"43",X"4F",X"50",X"59",X"20",X"21",X"21",X"20",X"5D");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
