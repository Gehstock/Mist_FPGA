library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpa_23l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpa_23l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"0E",X"12",X"F0",X"10",X"00",X"01",X"00",X"01",X"0F",X"12",X"F0",X"10",X"00",X"01",X"00",
		X"02",X"10",X"12",X"F0",X"10",X"00",X"01",X"00",X"03",X"11",X"12",X"F0",X"10",X"00",X"01",X"00",
		X"0D",X"25",X"12",X"FD",X"06",X"10",X"00",X"00",X"0A",X"21",X"1D",X"F0",X"05",X"10",X"00",X"00",
		X"04",X"12",X"16",X"F4",X"18",X"10",X"01",X"00",X"05",X"16",X"16",X"F2",X"18",X"10",X"01",X"00",
		X"06",X"1B",X"16",X"F0",X"18",X"10",X"01",X"00",X"0B",X"23",X"17",X"F0",X"01",X"20",X"00",X"00",
		X"13",X"00",X"10",X"00",X"00",X"00",X"4A",X"14",X"00",X"03",X"40",X"00",X"00",X"EB",X"DD",X"21",
		X"00",X"00",X"DD",X"19",X"DD",X"71",X"0D",X"DD",X"36",X"09",X"00",X"DD",X"36",X"08",X"00",X"FD",
		X"56",X"07",X"DD",X"72",X"07",X"FD",X"7E",X"00",X"D6",X"1E",X"FE",X"0A",X"D0",X"CB",X"4F",X"C0",
		X"FD",X"7E",X"03",X"D6",X"10",X"FE",X"E0",X"D0",X"79",X"FE",X"3A",X"28",X"36",X"CD",X"92",X"20",
		X"ED",X"5F",X"E6",X"7F",X"47",X"3A",X"03",X"E3",X"80",X"D6",X"2F",X"4F",X"DD",X"96",X"03",X"C6",
		X"08",X"FE",X"11",X"79",X"30",X"03",X"EE",X"10",X"4F",X"FD",X"BE",X"03",X"17",X"DD",X"77",X"0C",
		X"79",X"CD",X"38",X"15",X"92",X"1F",X"1F",X"1F",X"E6",X"1F",X"C6",X"02",X"41",X"CB",X"38",X"0E",
		X"2E",X"18",X"0F",X"01",X"2A",X"8F",X"CB",X"3A",X"CB",X"3A",X"CB",X"3A",X"3A",X"14",X"E5",X"EE",
		X"1F",X"92",X"21",X"00",X"31",X"85",X"6F",X"56",X"FD",X"7E",X"03",X"DD",X"77",X"03",X"CB",X"3F",
		X"90",X"30",X"02",X"ED",X"44",X"1E",X"FF",X"1C",X"92",X"30",X"FC",X"82",X"DD",X"73",X"05",X"06",
		X"08",X"CB",X"27",X"BA",X"CB",X"13",X"CB",X"43",X"20",X"01",X"92",X"10",X"F4",X"7B",X"2F",X"DD",
		X"77",X"04",X"DD",X"71",X"00",X"C9",X"21",X"D9",X"E1",X"7E",X"A7",X"C2",X"9A",X"11",X"3A",X"08",
		X"E5",X"FE",X"03",X"30",X"79",X"47",X"05",X"21",X"B4",X"2C",X"3A",X"E2",X"E1",X"1F",X"1F",X"1F",
		X"E6",X"1F",X"85",X"10",X"02",X"C6",X"20",X"6F",X"4E",X"3A",X"E2",X"E1",X"1F",X"1F",X"1F",X"E6",
		X"1F",X"5F",X"16",X"83",X"FD",X"21",X"00",X"04",X"FD",X"19",X"EB",X"11",X"20",X"00",X"06",X"07",
		X"3A",X"14",X"E5",X"B8",X"28",X"07",X"36",X"00",X"19",X"FD",X"19",X"10",X"F6",X"22",X"E4",X"E0",
		X"71",X"FD",X"36",X"00",X"04",X"19",X"FD",X"19",X"36",X"F3",X"FD",X"36",X"00",X"04",X"10",X"F5",
		X"3A",X"E2",X"E1",X"1F",X"1F",X"E6",X"3E",X"C6",X"00",X"6F",X"26",X"E2",X"3A",X"14",X"E5",X"EE",
		X"1F",X"57",X"FD",X"21",X"24",X"2C",X"FD",X"09",X"FD",X"7E",X"00",X"5F",X"E6",X"70",X"07",X"B2",
		X"07",X"07",X"07",X"77",X"E6",X"F8",X"57",X"7B",X"E6",X"07",X"B2",X"23",X"77",X"C9",X"87",X"C6",
		X"7A",X"77",X"87",X"28",X"02",X"3E",X"0A",X"32",X"D8",X"E1",X"4E",X"CB",X"19",X"D8",X"CB",X"19",
		X"21",X"D8",X"E1",X"35",X"F2",X"B6",X"11",X"36",X"0B",X"3A",X"14",X"E5",X"38",X"3C",X"FE",X"07",
		X"28",X"3E",X"3E",X"0B",X"18",X"27",X"7E",X"21",X"14",X"E5",X"30",X"1C",X"A7",X"20",X"01",X"35",
		X"C6",X"F3",X"FE",X"FC",X"38",X"02",X"D6",X"0C",X"4F",X"C6",X"03",X"FA",X"C9",X"11",X"C2",X"29",
		X"11",X"79",X"D6",X"10",X"4F",X"C3",X"29",X"11",X"FE",X"09",X"20",X"01",X"34",X"2F",X"C6",X"F2",
		X"FE",X"F0",X"30",X"02",X"C6",X"0C",X"4F",X"C3",X"29",X"11",X"FE",X"04",X"3E",X"0B",X"20",X"D0",
		X"21",X"D9",X"E1",X"34",X"2A",X"E1",X"E1",X"22",X"F1",X"E0",X"21",X"00",X"00",X"22",X"EF",X"E0",
		X"C9",X"21",X"44",X"2D",X"ED",X"53",X"EB",X"E0",X"22",X"E9",X"E0",X"3A",X"4E",X"E0",X"C6",X"03",
		X"DD",X"77",X"01",X"DD",X"36",X"00",X"0B",X"C9",X"3A",X"4E",X"E0",X"DD",X"BE",X"01",X"20",X"F3",
		X"2A",X"EB",X"E0",X"23",X"22",X"EB",X"E0",X"2B",X"EB",X"FD",X"21",X"00",X"04",X"FD",X"19",X"2A",
		X"E9",X"E0",X"01",X"20",X"00",X"7E",X"23",X"3D",X"FE",X"03",X"38",X"0D",X"3C",X"12",X"FD",X"36",
		X"00",X"80",X"EB",X"09",X"EB",X"FD",X"09",X"18",X"EC",X"3D",X"FA",X"55",X"12",X"28",X"B9",X"5E",
		X"23",X"56",X"23",X"18",X"AF",X"21",X"97",X"2C",X"C3",X"00",X"03",X"3A",X"0D",X"E5",X"3D",X"F8",
		X"21",X"AB",X"2C",X"3A",X"4E",X"E0",X"E6",X"3F",X"28",X"1B",X"E6",X"1F",X"C0",X"CD",X"7B",X"03",
		X"CD",X"88",X"12",X"36",X"02",X"EB",X"36",X"12",X"21",X"0B",X"E5",X"7E",X"23",X"96",X"FE",X"40",
		X"D8",X"23",X"36",X"00",X"C9",X"CD",X"00",X"03",X"3A",X"0D",X"E5",X"21",X"55",X"80",X"01",X"02",
		X"13",X"11",X"20",X"00",X"3D",X"28",X"08",X"19",X"0C",X"05",X"3D",X"28",X"02",X"04",X"19",X"70",
		X"11",X"00",X"04",X"EB",X"19",X"71",X"C9",X"21",X"70",X"E3",X"11",X"10",X"00",X"01",X"02",X"19",
		X"7E",X"FE",X"14",X"28",X"2A",X"FE",X"1E",X"38",X"1B",X"FE",X"20",X"38",X"08",X"FE",X"22",X"38",
		X"13",X"FE",X"2A",X"30",X"0F",X"3A",X"DF",X"E1",X"1F",X"1F",X"D8",X"79",X"32",X"DF",X"E1",X"C6",
		X"15",X"C3",X"6F",X"0D",X"19",X"10",X"D9",X"3A",X"DF",X"E1",X"A7",X"C8",X"AF",X"18",X"ED",X"3A",
		X"DF",X"E1",X"1F",X"0D",X"30",X"E5",X"C9",X"3A",X"DC",X"E1",X"A7",X"C8",X"3A",X"4E",X"E0",X"E6",
		X"0F",X"28",X"04",X"E6",X"07",X"C0",X"3C",X"3C",X"4F",X"2A",X"DA",X"E1",X"7E",X"D6",X"5A",X"28",
		X"0A",X"3C",X"06",X"04",X"C6",X"05",X"28",X"03",X"10",X"FA",X"C9",X"11",X"00",X"04",X"19",X"71",
		X"C9",X"21",X"00",X"40",X"22",X"02",X"E3",X"3A",X"4E",X"E0",X"E6",X"03",X"20",X"48",X"DD",X"35",
		X"0A",X"F2",X"66",X"13",X"21",X"5F",X"2A",X"CD",X"7B",X"03",X"3E",X"18",X"CD",X"75",X"0D",X"18",
		X"29",X"CD",X"48",X"15",X"07",X"07",X"30",X"2B",X"2A",X"1A",X"E3",X"11",X"79",X"FF",X"19",X"7C",
		X"A7",X"20",X"05",X"7D",X"FE",X"D1",X"38",X"02",X"3E",X"D1",X"5F",X"CB",X"3B",X"83",X"2F",X"6F",
		X"3E",X"FF",X"DE",X"00",X"67",X"2B",X"67",X"22",X"08",X"E3",X"DD",X"34",X"00",X"CD",X"76",X"15",
		X"C3",X"B8",X"08",X"CD",X"8A",X"14",X"CD",X"33",X"15",X"D6",X"1C",X"32",X"07",X"E3",X"18",X"ED",
		X"DD",X"34",X"00",X"3E",X"14",X"CD",X"75",X"0D",X"CD",X"48",X"15",X"2A",X"0E",X"E3",X"CD",X"A4",
		X"14",X"CD",X"33",X"15",X"D6",X"1E",X"18",X"E3",X"CD",X"48",X"15",X"2A",X"0E",X"E3",X"CD",X"A4",
		X"14",X"2A",X"06",X"E3",X"ED",X"5B",X"08",X"E3",X"19",X"22",X"06",X"E3",X"21",X"0C",X"00",X"19",
		X"22",X"08",X"E3",X"CB",X"14",X"38",X"0F",X"CD",X"33",X"15",X"D6",X"1D",X"47",X"3A",X"07",X"E3",
		X"B8",X"38",X"03",X"DD",X"34",X"00",X"CD",X"AC",X"15",X"C3",X"B8",X"08",X"DD",X"36",X"00",X"02",
		X"18",X"B6",X"2A",X"02",X"E3",X"ED",X"5B",X"04",X"E3",X"19",X"22",X"02",X"E3",X"2A",X"06",X"E3",
		X"ED",X"5B",X"08",X"E3",X"19",X"22",X"06",X"E3",X"CD",X"B8",X"08",X"DD",X"35",X"0A",X"C0",X"DD",
		X"34",X"00",X"DD",X"36",X"0D",X"03",X"3E",X"1F",X"C3",X"75",X"0D",X"AF",X"32",X"A2",X"E1",X"DD",
		X"35",X"0A",X"F0",X"DD",X"7E",X"0D",X"FE",X"09",X"D2",X"18",X"01",X"FE",X"05",X"38",X"0B",X"CD",
		X"B8",X"08",X"DD",X"34",X"0D",X"DD",X"36",X"0A",X"0E",X"C9",X"DD",X"CB",X"0A",X"4E",X"C0",X"EE",
		X"07",X"DD",X"77",X"0D",X"DD",X"7E",X"0A",X"FE",X"C0",X"D2",X"B8",X"08",X"DD",X"36",X"0D",X"05",
		X"C9",X"DD",X"35",X"0A",X"DD",X"7E",X"0A",X"FE",X"50",X"D0",X"21",X"4D",X"E0",X"34",X"DD",X"36",
		X"00",X"04",X"C9",X"CD",X"DB",X"20",X"22",X"D6",X"E0",X"7C",X"D6",X"08",X"FE",X"F0",X"D2",X"52",
		X"08",X"2A",X"D8",X"E0",X"23",X"CB",X"7C",X"20",X"02",X"2B",X"2B",X"22",X"D8",X"E0",X"2A",X"DA",
		X"E0",X"ED",X"5B",X"DC",X"E0",X"19",X"4C",X"22",X"DA",X"E0",X"21",X"24",X"00",X"19",X"22",X"DC",
		X"E0",X"CB",X"14",X"38",X"1F",X"C6",X"0B",X"CD",X"38",X"15",X"D6",X"08",X"B9",X"30",X"15",X"ED",
		X"5B",X"DC",X"E0",X"21",X"00",X"00",X"ED",X"52",X"CB",X"3A",X"CB",X"1B",X"CB",X"3A",X"CB",X"1B",
		X"19",X"22",X"DC",X"E0",X"CD",X"B8",X"08",X"C3",X"EF",X"20",X"3A",X"49",X"E0",X"87",X"21",X"28",
		X"30",X"85",X"6F",X"5E",X"23",X"66",X"2E",X"00",X"22",X"0E",X"E3",X"AF",X"CB",X"13",X"17",X"57",
		X"ED",X"53",X"1C",X"E3",X"ED",X"5B",X"02",X"E3",X"AF",X"ED",X"52",X"4F",X"7C",X"30",X"03",X"ED",
		X"44",X"0C",X"FE",X"18",X"38",X"02",X"3E",X"18",X"21",X"30",X"30",X"85",X"6F",X"5E",X"16",X"00",
		X"2A",X"04",X"E3",X"7C",X"A7",X"F2",X"D4",X"14",X"0D",X"20",X"11",X"2F",X"67",X"7D",X"2F",X"6F",
		X"23",X"EB",X"18",X"03",X"0D",X"28",X"57",X"A7",X"ED",X"52",X"30",X"52",X"11",X"02",X"00",X"3A",
		X"4E",X"E0",X"1F",X"2A",X"04",X"E3",X"ED",X"5A",X"22",X"04",X"E3",X"ED",X"5B",X"02",X"E3",X"19",
		X"22",X"02",X"E3",X"54",X"21",X"DC",X"E1",X"7E",X"3D",X"C0",X"3A",X"0B",X"E5",X"87",X"87",X"87",
		X"C6",X"08",X"82",X"D0",X"36",X"00",X"21",X"0E",X"E5",X"34",X"7E",X"06",X"09",X"FE",X"19",X"28",
		X"0F",X"38",X"01",X"3D",X"D6",X"05",X"CA",X"C0",X"27",X"10",X"F9",X"FE",X"06",X"CA",X"C0",X"27",
		X"3E",X"10",X"CD",X"75",X"0D",X"AF",X"0E",X"01",X"CD",X"C2",X"02",X"C3",X"12",X"0D",X"11",X"FD",
		X"FF",X"18",X"AC",X"3A",X"03",X"E3",X"C6",X"20",X"47",X"3A",X"E2",X"E1",X"80",X"C6",X"06",X"CB",
		X"3F",X"CB",X"3F",X"6F",X"26",X"E2",X"7E",X"C9",X"2A",X"4A",X"E0",X"7C",X"AD",X"A5",X"07",X"D0",
		X"4F",X"3A",X"20",X"E3",X"A7",X"20",X"05",X"3E",X"0A",X"32",X"20",X"E3",X"21",X"30",X"E3",X"06",
		X"04",X"11",X"10",X"00",X"7E",X"A7",X"28",X"05",X"19",X"10",X"F9",X"79",X"C9",X"36",X"0E",X"3E",
		X"12",X"CD",X"75",X"0D",X"79",X"C9",X"3A",X"03",X"E3",X"4F",X"C6",X"04",X"CD",X"38",X"15",X"D6",
		X"09",X"CD",X"C9",X"15",X"7A",X"EE",X"03",X"57",X"3E",X"09",X"CD",X"92",X"15",X"2C",X"14",X"14",
		X"3E",X"0D",X"81",X"4F",X"2C",X"2C",X"7D",X"E6",X"3F",X"6F",X"7E",X"D6",X"09",X"CD",X"ED",X"08",
		X"47",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"C3",X"76",X"09",X"3A",X"03",X"E3",X"4F",
		X"3A",X"07",X"E3",X"C6",X"11",X"CD",X"C9",X"15",X"7A",X"EE",X"03",X"57",X"3E",X"09",X"CD",X"C5",
		X"15",X"14",X"14",X"3E",X"0D",X"81",X"4F",X"18",X"D8",X"0C",X"CD",X"ED",X"08",X"47",X"11",X"00",
		X"05",X"3A",X"E2",X"E1",X"CB",X"67",X"20",X"01",X"14",X"FD",X"21",X"A4",X"E1",X"C3",X"76",X"09",
		X"DD",X"36",X"0A",X"0C",X"3A",X"07",X"E3",X"C6",X"0A",X"32",X"27",X"E3",X"2A",X"02",X"E3",X"11",
		X"00",X"1C",X"19",X"22",X"22",X"E3",X"DD",X"34",X"00",X"C9",X"DD",X"35",X"0A",X"28",X"19",X"2A",
		X"22",X"E3",X"11",X"5D",X"04",X"19",X"22",X"22",X"E3",X"DD",X"7E",X"0A",X"1F",X"3E",X"09",X"38",
		X"01",X"3C",X"DD",X"77",X"0D",X"C3",X"B8",X"08",X"DD",X"34",X"00",X"DD",X"36",X"0A",X"03",X"DD",
		X"36",X"0D",X"0B",X"3A",X"E2",X"E1",X"DD",X"86",X"03",X"DD",X"77",X"0F",X"C9",X"CD",X"31",X"08",
		X"DD",X"35",X"0A",X"F0",X"DD",X"7E",X"0D",X"FE",X"0D",X"CA",X"52",X"08",X"FE",X"29",X"CA",X"52",
		X"08",X"DD",X"34",X"0D",X"DD",X"36",X"0A",X"03",X"C9",X"3A",X"03",X"E3",X"C6",X"0A",X"DD",X"77",
		X"03",X"3A",X"07",X"E3",X"C6",X"02",X"DD",X"77",X"07",X"DD",X"34",X"00",X"C9",X"3A",X"00",X"E3",
		X"FE",X"06",X"30",X"2B",X"DD",X"7E",X"07",X"D6",X"03",X"FE",X"3A",X"38",X"22",X"DD",X"77",X"07",
		X"CD",X"1B",X"08",X"DD",X"7E",X"07",X"1F",X"1F",X"1F",X"7A",X"17",X"E6",X"07",X"F6",X"60",X"77",
		X"11",X"00",X"04",X"19",X"36",X"00",X"1F",X"D0",X"11",X"20",X"FC",X"19",X"36",X"00",X"C9",X"CD",
		X"1B",X"08",X"36",X"00",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"4E",X"03",X"DD",X"7E",X"0C",X"87",
		X"87",X"87",X"21",X"1C",X"31",X"85",X"6F",X"3A",X"20",X"E3",X"11",X"04",X"F8",X"D6",X"0B",X"28",
		X"06",X"3D",X"20",X"17",X"11",X"0A",X"F0",X"3A",X"23",X"E3",X"82",X"91",X"FE",X"E8",X"38",X"0B",
		X"3A",X"27",X"E3",X"DD",X"96",X"07",X"86",X"83",X"F2",X"4E",X"17",X"DD",X"7E",X"0C",X"A7",X"F8",
		X"23",X"3A",X"03",X"E3",X"91",X"86",X"23",X"46",X"23",X"B8",X"38",X"05",X"96",X"30",X"01",X"AF",
		X"80",X"23",X"BE",X"D2",X"C4",X"17",X"23",X"46",X"23",X"86",X"6F",X"24",X"3A",X"07",X"E3",X"86",
		X"DD",X"96",X"07",X"3D",X"80",X"F8",X"3A",X"04",X"D0",X"CB",X"77",X"C8",X"E1",X"3E",X"07",X"32",
		X"00",X"E3",X"3E",X"03",X"32",X"0D",X"E3",X"AF",X"32",X"0A",X"E3",X"32",X"B0",X"E3",X"32",X"72",
		X"E1",X"CD",X"52",X"08",X"06",X"03",X"3A",X"07",X"E3",X"C6",X"14",X"4F",X"3A",X"03",X"E3",X"21",
		X"D3",X"E1",X"34",X"21",X"C0",X"E3",X"FD",X"21",X"DF",X"30",X"36",X"1C",X"23",X"23",X"23",X"77",
		X"C6",X"10",X"CD",X"F8",X"17",X"71",X"CD",X"F8",X"17",X"23",X"23",X"FD",X"5E",X"00",X"73",X"FD",
		X"23",X"23",X"23",X"23",X"10",X"E4",X"CD",X"A1",X"08",X"3E",X"1F",X"C3",X"75",X"0D",X"3A",X"E2",
		X"E1",X"DD",X"86",X"03",X"32",X"2F",X"E3",X"3E",X"0D",X"32",X"20",X"E3",X"3E",X"26",X"32",X"2D",
		X"E3",X"3E",X"03",X"32",X"2A",X"E3",X"3E",X"01",X"CD",X"75",X"0D",X"11",X"07",X"00",X"19",X"7E",
		X"E6",X"0F",X"0E",X"01",X"FE",X"0E",X"30",X"07",X"CD",X"C2",X"02",X"E1",X"C3",X"52",X"08",X"20",
		X"13",X"CD",X"F0",X"17",X"C6",X"05",X"DD",X"77",X"08",X"CD",X"C2",X"02",X"DD",X"34",X"00",X"DD",
		X"36",X"0A",X"00",X"C9",X"CD",X"56",X"08",X"CD",X"F0",X"17",X"21",X"10",X"FB",X"C6",X"06",X"DD",
		X"77",X"08",X"E5",X"CD",X"C2",X"02",X"E1",X"DD",X"7E",X"07",X"84",X"DD",X"77",X"07",X"DD",X"7E",
		X"03",X"85",X"DD",X"77",X"03",X"DD",X"36",X"0D",X"54",X"DD",X"36",X"00",X"21",X"DD",X"36",X"0A",
		X"3B",X"C3",X"56",X"08",X"47",X"DD",X"7E",X"0C",X"C6",X"80",X"4F",X"FE",X"8B",X"28",X"1B",X"FE",
		X"8E",X"28",X"17",X"78",X"96",X"FE",X"04",X"D0",X"DD",X"71",X"0C",X"23",X"23",X"23",X"7E",X"1F",
		X"1F",X"1F",X"1F",X"E6",X"0F",X"0E",X"01",X"C3",X"C2",X"02",X"78",X"FE",X"FC",X"30",X"E9",X"C9",
		X"ED",X"5F",X"E6",X"03",X"C0",X"3E",X"02",X"C9",X"23",X"FD",X"5E",X"00",X"73",X"23",X"FD",X"5E",
		X"01",X"73",X"23",X"23",X"FD",X"23",X"FD",X"23",X"C9",X"3A",X"00",X"E3",X"FE",X"06",X"D0",X"FE",
		X"01",X"26",X"00",X"28",X"76",X"2A",X"1C",X"E3",X"ED",X"5B",X"1A",X"E3",X"7A",X"A7",X"FA",X"23",
		X"18",X"ED",X"52",X"21",X"03",X"00",X"30",X"03",X"21",X"FE",X"FF",X"3A",X"4E",X"E0",X"1F",X"38",
		X"01",X"1D",X"19",X"22",X"1A",X"E3",X"ED",X"5B",X"04",X"E3",X"A7",X"ED",X"52",X"22",X"14",X"E3",
		X"EB",X"2A",X"E1",X"E1",X"19",X"22",X"E1",X"E1",X"3A",X"D9",X"E1",X"1F",X"30",X"3D",X"2A",X"EF",
		X"E0",X"19",X"7C",X"C6",X"06",X"FE",X"0C",X"38",X"17",X"D6",X"12",X"67",X"E5",X"21",X"3F",X"E2",
		X"11",X"42",X"E2",X"01",X"40",X"00",X"ED",X"B8",X"21",X"42",X"E2",X"0E",X"03",X"ED",X"B8",X"E1",
		X"22",X"EF",X"E0",X"ED",X"5B",X"F1",X"E0",X"19",X"3A",X"08",X"E5",X"FE",X"03",X"30",X"0C",X"3A",
		X"E2",X"E1",X"94",X"FE",X"F4",X"38",X"04",X"AF",X"32",X"D9",X"E1",X"7C",X"2F",X"21",X"3D",X"E0",
		X"86",X"32",X"C0",X"E1",X"2A",X"14",X"E3",X"54",X"5D",X"CB",X"3C",X"CB",X"1D",X"19",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"EB",X"2A",X"04",X"E5",X"19",X"22",X"04",X"E5",X"7C",X"2F",
		X"32",X"C1",X"E1",X"CB",X"3A",X"CB",X"1B",X"2A",X"06",X"E5",X"19",X"22",X"06",X"E5",X"7C",X"2F",
		X"32",X"C2",X"E1",X"CD",X"33",X"15",X"FE",X"C4",X"30",X"02",X"3E",X"C4",X"C6",X"28",X"30",X"01",
		X"AF",X"47",X"C6",X"94",X"32",X"C3",X"E1",X"CB",X"28",X"78",X"C6",X"72",X"32",X"C4",X"E1",X"C9",
		X"CD",X"31",X"08",X"CD",X"99",X"16",X"DD",X"35",X"0A",X"F0",X"DD",X"34",X"0A",X"DD",X"7E",X"03",
		X"FE",X"E0",X"D0",X"DD",X"7E",X"0C",X"17",X"D8",X"3A",X"C0",X"E3",X"A7",X"C0",X"FD",X"21",X"70",
		X"E3",X"11",X"10",X"00",X"06",X"05",X"FD",X"7E",X"00",X"FE",X"1D",X"20",X"0D",X"FD",X"7E",X"0C",
		X"17",X"38",X"07",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"D8",X"FD",X"19",X"10",X"E8",X"DD",X"7E",
		X"07",X"FD",X"77",X"07",X"DD",X"7E",X"0F",X"D6",X"04",X"FD",X"77",X"0F",X"FD",X"36",X"00",X"11",
		X"FD",X"36",X"0D",X"22",X"FD",X"36",X"0C",X"0C",X"DD",X"36",X"0A",X"43",X"C9",X"3A",X"00",X"E3",
		X"FE",X"06",X"D0",X"DD",X"7E",X"04",X"C6",X"DD",X"DD",X"77",X"04",X"30",X"03",X"DD",X"35",X"0F",
		X"CD",X"38",X"08",X"CD",X"99",X"16",X"C9",X"CD",X"31",X"08",X"CD",X"99",X"16",X"C9",X"CD",X"31",
		X"08",X"DD",X"7E",X"0C",X"A7",X"C0",X"DD",X"7E",X"0D",X"07",X"07",X"E6",X"1C",X"21",X"00",X"2E",
		X"85",X"6F",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"86",X"23",X"BE",X"30",X"45",X"47",X"3A",X"00",
		X"E3",X"FE",X"04",X"C8",X"3A",X"04",X"D0",X"CB",X"77",X"C8",X"78",X"46",X"0E",X"02",X"CB",X"38",
		X"50",X"CB",X"38",X"BA",X"38",X"04",X"78",X"82",X"47",X"0D",X"DD",X"7E",X"03",X"80",X"D6",X"1C",
		X"32",X"03",X"E3",X"79",X"32",X"0D",X"E3",X"3D",X"3D",X"32",X"05",X"E3",X"3E",X"80",X"32",X"04",
		X"E3",X"23",X"7E",X"32",X"0A",X"E3",X"21",X"00",X"02",X"22",X"08",X"E3",X"3E",X"06",X"32",X"00",
		X"E3",X"C9",X"96",X"FE",X"04",X"D0",X"DD",X"34",X"0C",X"23",X"23",X"7E",X"0E",X"01",X"C3",X"C2",
		X"02",X"DD",X"35",X"0A",X"F2",X"0D",X"1A",X"DD",X"7E",X"0E",X"47",X"3C",X"0E",X"07",X"FE",X"06",
		X"38",X"0B",X"3A",X"4E",X"E0",X"E6",X"30",X"20",X"02",X"3E",X"30",X"4F",X"AF",X"DD",X"77",X"0E",
		X"DD",X"71",X"0A",X"78",X"FE",X"04",X"38",X"04",X"EE",X"07",X"3D",X"47",X"C6",X"06",X"DD",X"46",
		X"0C",X"04",X"FA",X"08",X"1A",X"DD",X"77",X"0C",X"C6",X"45",X"DD",X"77",X"0D",X"3A",X"20",X"E3",
		X"FE",X"0F",X"38",X"0E",X"C0",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"C6",X"10",X"FE",X"30",X"DA",
		X"FD",X"16",X"CD",X"38",X"08",X"DD",X"7E",X"0C",X"FE",X"06",X"C8",X"CD",X"99",X"16",X"C9",X"CD",
		X"31",X"08",X"DD",X"35",X"0A",X"F0",X"DD",X"7E",X"0D",X"FE",X"4A",X"C8",X"DD",X"35",X"0D",X"DD",
		X"36",X"0A",X"07",X"C9",X"3A",X"00",X"E3",X"FE",X"06",X"D0",X"DD",X"35",X"0E",X"F2",X"66",X"1A",
		X"DD",X"36",X"0E",X"06",X"DD",X"7E",X"0D",X"3D",X"01",X"03",X"00",X"21",X"8E",X"1A",X"ED",X"B1",
		X"20",X"01",X"7E",X"DD",X"77",X"0D",X"DD",X"7E",X"04",X"C6",X"C0",X"DD",X"77",X"04",X"30",X"03",
		X"DD",X"35",X"0F",X"CD",X"38",X"08",X"DD",X"7E",X"0C",X"D6",X"04",X"CB",X"27",X"C6",X"0C",X"4F",
		X"DD",X"7E",X"03",X"CD",X"38",X"15",X"91",X"DD",X"77",X"07",X"CD",X"99",X"16",X"C9",X"11",X"15",
		X"1A",X"20",X"DD",X"36",X"0B",X"01",X"3A",X"00",X"E3",X"FE",X"06",X"D0",X"2A",X"72",X"E3",X"7C",
		X"FE",X"08",X"28",X"09",X"11",X"70",X"00",X"19",X"22",X"72",X"E3",X"18",X"2C",X"DD",X"36",X"0A",
		X"00",X"DD",X"34",X"00",X"DD",X"36",X"0E",X"80",X"C9",X"3A",X"4E",X"E0",X"1F",X"D8",X"3A",X"00",
		X"E3",X"FE",X"06",X"D0",X"3A",X"4E",X"E0",X"47",X"E6",X"03",X"20",X"0D",X"DD",X"34",X"03",X"CB",
		X"68",X"28",X"06",X"DD",X"35",X"03",X"DD",X"35",X"03",X"3A",X"4E",X"E0",X"E6",X"07",X"20",X"0D",
		X"DD",X"7E",X"03",X"C6",X"18",X"CD",X"38",X"15",X"D6",X"10",X"DD",X"77",X"07",X"C3",X"B8",X"08",
		X"DD",X"35",X"0E",X"20",X"CF",X"DD",X"36",X"0A",X"58",X"DD",X"34",X"00",X"DD",X"36",X"0D",X"52",
		X"C9",X"DD",X"35",X"0A",X"28",X"15",X"2A",X"72",X"E3",X"11",X"80",X"01",X"19",X"22",X"72",X"E3",
		X"7C",X"FE",X"F0",X"D2",X"52",X"08",X"CD",X"99",X"16",X"18",X"BE",X"DD",X"34",X"00",X"DD",X"36",
		X"0A",X"6E",X"DD",X"36",X"0D",X"23",X"C9",X"CD",X"99",X"16",X"DD",X"35",X"0A",X"20",X"95",X"DD",
		X"35",X"00",X"DD",X"35",X"0B",X"DD",X"36",X"0D",X"52",X"C9",X"21",X"EE",X"E0",X"3A",X"4E",X"E0",
		X"96",X"F8",X"01",X"00",X"10",X"ED",X"5F",X"E6",X"F0",X"26",X"E4",X"51",X"59",X"6F",X"7E",X"D6",
		X"1E",X"FE",X"0A",X"30",X"0A",X"CB",X"4F",X"20",X"06",X"FE",X"04",X"38",X"63",X"0C",X"5D",X"7D",
		X"C6",X"10",X"10",X"E9",X"ED",X"53",X"D4",X"E1",X"0D",X"F8",X"3A",X"10",X"E5",X"E6",X"03",X"FE",
		X"01",X"89",X"4F",X"FE",X"09",X"DA",X"7A",X"1B",X"0E",X"08",X"21",X"FF",X"2F",X"09",X"4E",X"06",
		X"05",X"21",X"70",X"E3",X"11",X"00",X"00",X"7E",X"A7",X"28",X"39",X"D6",X"2F",X"20",X"01",X"14",
		X"7D",X"C6",X"10",X"6F",X"10",X"F1",X"7A",X"B9",X"D0",X"1C",X"1D",X"C8",X"ED",X"5F",X"E6",X"0F",
		X"C6",X"19",X"21",X"4E",X"E0",X"86",X"32",X"EE",X"E0",X"16",X"00",X"DD",X"21",X"00",X"E3",X"DD",
		X"19",X"21",X"D4",X"E1",X"5E",X"FD",X"21",X"00",X"E4",X"FD",X"19",X"0E",X"3B",X"C3",X"64",X"10",
		X"55",X"14",X"18",X"9B",X"5D",X"18",X"C9",X"3A",X"4E",X"E0",X"21",X"52",X"E0",X"AE",X"E6",X"1F",
		X"C0",X"ED",X"5F",X"77",X"21",X"C6",X"E1",X"06",X"03",X"7E",X"A7",X"20",X"04",X"23",X"10",X"F9",
		X"C9",X"DD",X"21",X"00",X"E4",X"04",X"78",X"48",X"06",X"10",X"FE",X"04",X"28",X"0F",X"3A",X"D6",
		X"E1",X"3D",X"FA",X"FD",X"1B",X"0D",X"0D",X"DD",X"21",X"70",X"E3",X"06",X"05",X"11",X"10",X"00",
		X"DD",X"7E",X"00",X"A7",X"28",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"35",X"79",X"FE",X"02",X"30",
		X"43",X"ED",X"5F",X"E6",X"1F",X"C6",X"20",X"DD",X"77",X"0F",X"21",X"D6",X"E1",X"35",X"ED",X"5F",
		X"E6",X"1E",X"5F",X"16",X"00",X"FE",X"0E",X"3E",X"82",X"38",X"04",X"ED",X"5F",X"E6",X"80",X"DD",
		X"77",X"0C",X"21",X"08",X"30",X"19",X"7E",X"DD",X"77",X"07",X"23",X"7E",X"DD",X"77",X"03",X"06",
		X"00",X"21",X"59",X"1C",X"09",X"09",X"7E",X"DD",X"77",X"0D",X"DD",X"36",X"0E",X"00",X"23",X"7E",
		X"DD",X"77",X"00",X"C9",X"CD",X"0A",X"08",X"18",X"C5",X"2B",X"26",X"2A",X"26",X"2B",X"22",X"2A",
		X"22",X"31",X"1E",X"DD",X"7E",X"0D",X"FE",X"2B",X"D8",X"DD",X"CB",X"0E",X"7E",X"20",X"18",X"DD",
		X"35",X"0E",X"F0",X"DD",X"34",X"0D",X"FE",X"2F",X"28",X"1C",X"FE",X"34",X"20",X"04",X"DD",X"36",
		X"0D",X"31",X"DD",X"36",X"0E",X"08",X"C9",X"DD",X"34",X"0E",X"F8",X"DD",X"35",X"0D",X"FE",X"2C",
		X"28",X"F0",X"FE",X"32",X"28",X"EC",X"DD",X"36",X"0E",X"F8",X"C9",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"CB",X"3C",X"CB",X"1D",X"DD",X"CB",X"0C",X"46",X"28",X"07",X"EB",X"21",X"00",X"00",X"A7",
		X"ED",X"52",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"34",X"00",X"C9",X"0E",X"3D",X"DD",X"7E",
		X"09",X"A7",X"20",X"13",X"0E",X"3B",X"DD",X"46",X"05",X"CB",X"10",X"30",X"02",X"0E",X"50",X"DD",
		X"7E",X"08",X"FE",X"60",X"38",X"01",X"0C",X"DD",X"71",X"0D",X"CD",X"FB",X"20",X"7C",X"FE",X"06",
		X"DA",X"52",X"08",X"01",X"05",X"00",X"22",X"D6",X"E0",X"7C",X"2A",X"DC",X"E0",X"09",X"22",X"DC",
		X"E0",X"ED",X"5B",X"DA",X"E0",X"19",X"22",X"DA",X"E0",X"54",X"CD",X"38",X"15",X"D6",X"08",X"BA",
		X"CD",X"EF",X"20",X"30",X"35",X"DD",X"77",X"07",X"DD",X"34",X"00",X"DD",X"36",X"0B",X"00",X"DD",
		X"7E",X"00",X"FE",X"2A",X"3E",X"03",X"20",X"05",X"DD",X"36",X"00",X"30",X"3D",X"CD",X"75",X"0D",
		X"C3",X"56",X"08",X"CD",X"DB",X"20",X"ED",X"5B",X"14",X"E3",X"CB",X"2A",X"CB",X"1B",X"ED",X"52",
		X"11",X"8E",X"00",X"ED",X"52",X"01",X"10",X"00",X"18",X"AC",X"3A",X"00",X"E3",X"FE",X"06",X"D2",
		X"B8",X"08",X"21",X"05",X"06",X"DD",X"7E",X"00",X"FE",X"2A",X"30",X"03",X"21",X"0B",X"02",X"FD",
		X"21",X"30",X"E3",X"11",X"10",X"00",X"06",X"04",X"FD",X"7E",X"00",X"FE",X"0F",X"20",X"14",X"FD",
		X"7E",X"07",X"DD",X"96",X"07",X"FE",X"0A",X"30",X"0A",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"94",
		X"BD",X"38",X"2B",X"FD",X"19",X"10",X"E1",X"3A",X"07",X"E3",X"DD",X"96",X"07",X"FE",X"F0",X"DA",
		X"B8",X"08",X"57",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"D6",X"04",X"FE",X"EA",X"DA",X"B8",X"08",
		X"3A",X"04",X"D0",X"CB",X"77",X"CA",X"B8",X"08",X"CD",X"52",X"08",X"C3",X"FD",X"16",X"FD",X"34",
		X"00",X"DD",X"7E",X"0D",X"FE",X"37",X"38",X"11",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"00",X"2D",
		X"DD",X"36",X"0A",X"0A",X"DD",X"36",X"0D",X"4F",X"C9",X"21",X"C9",X"E1",X"01",X"01",X"05",X"FE",
		X"31",X"30",X"07",X"23",X"05",X"FE",X"2A",X"28",X"01",X"23",X"3E",X"11",X"CD",X"75",X"0D",X"35",
		X"20",X"08",X"23",X"23",X"23",X"7E",X"FE",X"03",X"30",X"11",X"DD",X"36",X"00",X"20",X"DD",X"36",
		X"0A",X"06",X"DD",X"36",X"0D",X"37",X"78",X"CD",X"C2",X"02",X"C9",X"21",X"00",X"FC",X"D6",X"02",
		X"C3",X"9D",X"17",X"DD",X"36",X"0D",X"3E",X"CD",X"23",X"16",X"D6",X"03",X"E6",X"F8",X"C6",X"06",
		X"DD",X"77",X"0F",X"21",X"D1",X"E1",X"7E",X"A7",X"28",X"13",X"23",X"36",X"01",X"23",X"7E",X"A7",
		X"C8",X"C3",X"52",X"08",X"DD",X"36",X"0D",X"43",X"CD",X"23",X"16",X"18",X"E6",X"34",X"DD",X"34",
		X"00",X"DD",X"36",X"0A",X"04",X"CD",X"31",X"08",X"C9",X"21",X"D2",X"E1",X"7E",X"23",X"B6",X"A7",
		X"C2",X"52",X"08",X"DD",X"7E",X"03",X"FE",X"F8",X"D2",X"52",X"08",X"DD",X"35",X"0A",X"20",X"E5",
		X"DD",X"7E",X"0D",X"FE",X"49",X"CA",X"52",X"08",X"DD",X"34",X"0D",X"DD",X"36",X"0A",X"05",X"18",
		X"D4",X"3A",X"D3",X"E1",X"A7",X"C2",X"52",X"08",X"DD",X"35",X"0A",X"20",X"C8",X"DD",X"7E",X"0D",
		X"FE",X"42",X"30",X"1F",X"DD",X"34",X"0D",X"FE",X"3F",X"20",X"12",X"DD",X"7E",X"0F",X"1F",X"1F",
		X"1F",X"E6",X"1F",X"5F",X"16",X"83",X"0E",X"09",X"3E",X"01",X"CD",X"C2",X"02",X"DD",X"36",X"0A",
		X"02",X"18",X"A2",X"DD",X"7E",X"07",X"C6",X"08",X"DD",X"77",X"07",X"CD",X"56",X"08",X"DD",X"36",
		X"0C",X"00",X"DD",X"36",X"0D",X"81",X"DD",X"36",X"00",X"13",X"C9",X"DD",X"35",X"0A",X"CA",X"52",
		X"08",X"C3",X"B8",X"08",X"DD",X"35",X"0F",X"CA",X"4D",X"20",X"DD",X"34",X"00",X"DD",X"7E",X"0C",
		X"CB",X"27",X"28",X"3D",X"3F",X"1F",X"E6",X"80",X"DD",X"77",X"0C",X"4F",X"ED",X"5F",X"E6",X"3F",
		X"5F",X"16",X"00",X"21",X"26",X"01",X"19",X"0C",X"F2",X"D2",X"1E",X"EB",X"A7",X"21",X"00",X"00",
		X"ED",X"52",X"DD",X"74",X"05",X"DD",X"75",X"04",X"EE",X"3F",X"D6",X"20",X"87",X"DD",X"77",X"08",
		X"3E",X"00",X"DE",X"00",X"DD",X"77",X"09",X"ED",X"5F",X"E6",X"7F",X"C6",X"20",X"DD",X"77",X"0A",
		X"C9",X"06",X"01",X"DD",X"7E",X"07",X"FE",X"44",X"38",X"0C",X"06",X"03",X"FE",X"58",X"30",X"06",
		X"ED",X"5F",X"E6",X"02",X"3C",X"47",X"78",X"DD",X"86",X"0C",X"DD",X"77",X"0C",X"ED",X"5F",X"E6",
		X"0F",X"C6",X"24",X"DD",X"77",X"0B",X"21",X"66",X"01",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",
		X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"C9",X"CD",X"63",X"1C",X"CD",X"DB",X"20",X"DD",X"7E",
		X"0C",X"CB",X"27",X"20",X"52",X"DD",X"35",X"0A",X"28",X"49",X"2A",X"D6",X"E0",X"ED",X"5B",X"D8",
		X"E0",X"19",X"7A",X"ED",X"5B",X"04",X"E3",X"ED",X"52",X"22",X"D6",X"E0",X"17",X"38",X"2F",X"DD",
		X"7E",X"0D",X"06",X"A0",X"D6",X"2A",X"28",X"08",X"06",X"80",X"D6",X"07",X"38",X"02",X"06",X"D0",
		X"7C",X"B8",X"30",X"1F",X"2A",X"DA",X"E0",X"ED",X"5B",X"DC",X"E0",X"19",X"22",X"DA",X"E0",X"7C",
		X"FE",X"38",X"38",X"0F",X"FE",X"70",X"30",X"0B",X"CD",X"EF",X"20",X"C3",X"4C",X"1D",X"7C",X"FE",
		X"16",X"30",X"E1",X"DD",X"35",X"00",X"C9",X"2A",X"D8",X"E0",X"DD",X"5E",X"0B",X"16",X"00",X"A7",
		X"ED",X"52",X"22",X"D8",X"E0",X"30",X"16",X"DD",X"7E",X"03",X"D6",X"30",X"FE",X"40",X"3E",X"00",
		X"30",X"04",X"ED",X"5F",X"E6",X"80",X"DD",X"86",X"0C",X"3C",X"DD",X"77",X"0C",X"EB",X"2A",X"D6",
		X"E0",X"ED",X"52",X"DD",X"7E",X"0C",X"07",X"38",X"02",X"19",X"19",X"ED",X"5B",X"04",X"E3",X"ED",
		X"52",X"22",X"D6",X"E0",X"2A",X"DC",X"E0",X"DD",X"5E",X"0B",X"16",X"00",X"0F",X"3D",X"0F",X"30",
		X"1A",X"A7",X"ED",X"52",X"38",X"AD",X"22",X"DC",X"E0",X"EB",X"2A",X"DA",X"E0",X"A7",X"ED",X"52",
		X"0F",X"38",X"02",X"19",X"19",X"22",X"DA",X"E0",X"C3",X"78",X"1F",X"19",X"18",X"E8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
