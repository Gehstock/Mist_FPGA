library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_1R is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_1R is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"60",X"C0",X"7C",X"C0",X"94",X"C0",X"AC",X"C0",X"C4",X"C0",X"DC",X"C0",X"F4",X"C0",X"0C",X"C1",
		X"24",X"C1",X"3C",X"C1",X"54",X"C1",X"6E",X"C1",X"03",X"08",X"46",X"0F",X"41",X"0F",X"4E",X"0F",
		X"54",X"0F",X"41",X"0F",X"53",X"0F",X"54",X"0F",X"49",X"0F",X"43",X"0F",X"00",X"00",X"53",X"0F",
		X"43",X"0F",X"4F",X"0F",X"52",X"0F",X"45",X"0F",X"3F",X"0F",X"FF",X"FF",X"05",X"08",X"52",X"05",
		X"45",X"05",X"43",X"05",X"4F",X"05",X"52",X"05",X"44",X"05",X"00",X"00",X"59",X"05",X"4F",X"05",
		X"55",X"05",X"52",X"05",X"00",X"00",X"4E",X"05",X"41",X"05",X"4D",X"05",X"45",X"05",X"FF",X"FF",
		X"04",X"0A",X"42",X"06",X"45",X"06",X"53",X"06",X"54",X"06",X"00",X"00",X"50",X"06",X"4C",X"06",
		X"41",X"06",X"59",X"06",X"45",X"06",X"52",X"06",X"53",X"06",X"FF",X"FF",X"07",X"04",X"31",X"05",
		X"53",X"05",X"54",X"05",X"0F",X"FF",X"00",X"00",X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",
		X"44",X"05",X"FF",X"FF",X"09",X"04",X"32",X"05",X"4E",X"05",X"44",X"05",X"0F",X"FF",X"00",X"00",
		X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",X"44",X"05",X"FF",X"FF",X"0B",X"04",X"33",X"05",
		X"52",X"05",X"44",X"05",X"0F",X"FF",X"00",X"00",X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",
		X"44",X"05",X"FF",X"FF",X"0D",X"04",X"34",X"05",X"54",X"05",X"48",X"05",X"0F",X"FF",X"00",X"00",
		X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",X"44",X"05",X"FF",X"FF",X"0F",X"04",X"35",X"05",
		X"54",X"05",X"48",X"05",X"0F",X"FF",X"00",X"00",X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",
		X"44",X"05",X"FF",X"FF",X"11",X"04",X"36",X"05",X"54",X"05",X"48",X"05",X"0F",X"FF",X"00",X"00",
		X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",X"44",X"05",X"FF",X"FF",X"13",X"04",X"37",X"05",
		X"54",X"05",X"48",X"05",X"0F",X"FF",X"00",X"00",X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",
		X"44",X"05",X"FF",X"FF",X"15",X"04",X"38",X"05",X"54",X"05",X"48",X"05",X"0F",X"FF",X"00",X"00",
		X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",X"44",X"05",X"FF",X"FF",X"17",X"04",X"39",X"05",
		X"54",X"05",X"48",X"05",X"0F",X"FF",X"00",X"00",X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",
		X"44",X"05",X"FF",X"FF",X"19",X"03",X"31",X"05",X"30",X"05",X"54",X"05",X"48",X"05",X"0F",X"FF",
		X"00",X"00",X"52",X"05",X"4F",X"05",X"55",X"05",X"4E",X"05",X"44",X"05",X"FF",X"FF",X"1C",X"07",
		X"3A",X"05",X"3B",X"05",X"31",X"05",X"39",X"05",X"38",X"05",X"34",X"05",X"00",X"00",X"54",X"0F",
		X"45",X"0F",X"48",X"0F",X"4B",X"0F",X"41",X"0F",X"4E",X"0F",X"00",X"00",X"4C",X"05",X"54",X"05",
		X"44",X"05",X"2E",X"05",X"FF",X"FF",X"AA",X"C1",X"B0",X"C1",X"B6",X"C1",X"BC",X"C1",X"C2",X"C1",
		X"C8",X"C1",X"CE",X"C1",X"D4",X"C1",X"DA",X"C1",X"E0",X"C1",X"07",X"08",X"00",X"81",X"0F",X"08",
		X"09",X"08",X"04",X"81",X"05",X"08",X"0B",X"08",X"08",X"81",X"05",X"08",X"0D",X"08",X"0C",X"81",
		X"05",X"08",X"0F",X"08",X"10",X"81",X"05",X"08",X"11",X"08",X"14",X"81",X"05",X"08",X"13",X"08",
		X"18",X"81",X"05",X"08",X"15",X"08",X"1C",X"81",X"05",X"08",X"17",X"08",X"20",X"81",X"05",X"08",
		X"19",X"08",X"24",X"81",X"05",X"08",X"32",X"81",X"3C",X"81",X"46",X"81",X"50",X"81",X"5A",X"81",
		X"64",X"81",X"6E",X"81",X"78",X"81",X"82",X"81",X"8C",X"81",X"0E",X"C2",X"14",X"C2",X"1A",X"C2",
		X"20",X"C2",X"26",X"C2",X"2C",X"C2",X"32",X"C2",X"38",X"C2",X"3E",X"C2",X"44",X"C2",X"07",X"1B",
		X"28",X"81",X"05",X"02",X"09",X"1B",X"29",X"81",X"05",X"02",X"0B",X"1B",X"2A",X"81",X"05",X"02",
		X"0D",X"1B",X"2B",X"81",X"05",X"02",X"0F",X"1B",X"2C",X"81",X"05",X"02",X"11",X"1B",X"2D",X"81",
		X"05",X"02",X"13",X"1B",X"2E",X"81",X"05",X"02",X"15",X"1B",X"2F",X"81",X"05",X"02",X"17",X"1B",
		X"30",X"81",X"05",X"02",X"19",X"1B",X"31",X"81",X"05",X"02",X"18",X"C0",X"3C",X"C0",X"64",X"C2",
		X"7C",X"C2",X"94",X"C2",X"AC",X"C2",X"C4",X"C2",X"DC",X"C2",X"F4",X"C2",X"0C",X"C3",X"24",X"C3",
		X"3C",X"C3",X"6E",X"C1",X"07",X"04",X"31",X"02",X"53",X"02",X"54",X"02",X"0F",X"FF",X"00",X"00",
		X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",X"44",X"01",X"FF",X"FF",X"09",X"04",X"32",X"00",
		X"4E",X"00",X"44",X"00",X"0F",X"FF",X"00",X"00",X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",
		X"44",X"01",X"FF",X"FF",X"0B",X"04",X"33",X"00",X"52",X"00",X"44",X"00",X"0F",X"FF",X"00",X"00",
		X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",X"44",X"01",X"FF",X"FF",X"0D",X"04",X"34",X"00",
		X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",
		X"44",X"01",X"FF",X"FF",X"0F",X"04",X"35",X"00",X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",
		X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",X"44",X"01",X"FF",X"FF",X"11",X"04",X"36",X"00",
		X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",
		X"44",X"01",X"FF",X"FF",X"13",X"04",X"37",X"00",X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",
		X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",X"44",X"01",X"FF",X"FF",X"15",X"04",X"38",X"00",
		X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",
		X"44",X"01",X"FF",X"FF",X"17",X"04",X"39",X"00",X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",
		X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",X"01",X"44",X"01",X"FF",X"FF",X"19",X"03",X"31",X"00",
		X"30",X"00",X"54",X"00",X"48",X"00",X"0F",X"FF",X"00",X"00",X"52",X"01",X"4F",X"01",X"55",X"01",
		X"4E",X"01",X"44",X"01",X"FF",X"FF",X"00",X"00",X"00",X"20",X"21",X"0E",X"FC",X"C3",X"04",X"C4",
		X"DE",X"F1",X"00",X"20",X"00",X"40",X"7C",X"0E",X"44",X"C4",X"4C",X"C4",X"83",X"F1",X"00",X"40",
		X"00",X"60",X"21",X"0C",X"8C",X"C4",X"94",X"C4",X"DE",X"F3",X"00",X"60",X"00",X"80",X"57",X"0C",
		X"D4",X"C4",X"DC",X"C4",X"A8",X"F3",X"00",X"C0",X"00",X"E0",X"2F",X"0B",X"1C",X"C5",X"24",X"C5",
		X"E0",X"F4",X"FF",X"FF",X"00",X"80",X"00",X"84",X"20",X"C4",X"28",X"C4",X"00",X"84",X"00",X"88",
		X"68",X"C4",X"70",X"C4",X"00",X"88",X"00",X"8C",X"B0",X"C4",X"B8",X"C4",X"00",X"8C",X"00",X"90",
		X"F8",X"C4",X"00",X"C5",X"00",X"90",X"00",X"98",X"40",X"C5",X"48",X"C5",X"FF",X"FF",X"01",X"03",
		X"50",X"01",X"55",X"01",X"53",X"01",X"48",X"01",X"00",X"00",X"42",X"01",X"55",X"01",X"54",X"01",
		X"54",X"01",X"4F",X"01",X"4E",X"01",X"00",X"00",X"46",X"01",X"4F",X"01",X"52",X"01",X"00",X"00",
		X"00",X"00",X"43",X"08",X"48",X"08",X"45",X"08",X"43",X"08",X"4B",X"08",X"FF",X"FF",X"03",X"03",
		X"52",X"03",X"4F",X"03",X"4D",X"03",X"00",X"00",X"30",X"03",X"FF",X"FF",X"03",X"0A",X"4F",X"03",
		X"4B",X"03",X"FF",X"FF",X"03",X"0A",X"45",X"02",X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",
		X"FF",X"FF",X"03",X"11",X"52",X"03",X"41",X"03",X"4D",X"03",X"00",X"00",X"30",X"03",X"FF",X"FF",
		X"03",X"18",X"4F",X"03",X"4B",X"03",X"FF",X"FF",X"03",X"18",X"45",X"02",X"52",X"02",X"52",X"02",
		X"4F",X"02",X"52",X"02",X"FF",X"FF",X"04",X"03",X"52",X"03",X"4F",X"03",X"4D",X"03",X"00",X"00",
		X"31",X"03",X"FF",X"FF",X"04",X"0A",X"4F",X"03",X"4B",X"03",X"FF",X"FF",X"04",X"0A",X"45",X"02",
		X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",X"FF",X"FF",X"04",X"11",X"52",X"03",X"41",X"03",
		X"4D",X"03",X"00",X"00",X"31",X"03",X"FF",X"FF",X"04",X"18",X"4F",X"03",X"4B",X"03",X"FF",X"FF",
		X"04",X"18",X"45",X"02",X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",X"FF",X"FF",X"05",X"03",
		X"52",X"03",X"4F",X"03",X"4D",X"03",X"00",X"00",X"32",X"03",X"FF",X"FF",X"05",X"0A",X"4F",X"03",
		X"4B",X"03",X"FF",X"FF",X"05",X"0A",X"45",X"02",X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",
		X"FF",X"FF",X"05",X"11",X"52",X"03",X"41",X"03",X"4D",X"03",X"00",X"00",X"32",X"03",X"FF",X"FF",
		X"05",X"18",X"4F",X"03",X"4B",X"03",X"FF",X"FF",X"05",X"18",X"45",X"02",X"52",X"02",X"52",X"02",
		X"4F",X"02",X"52",X"02",X"FF",X"FF",X"06",X"03",X"52",X"03",X"4F",X"03",X"4D",X"03",X"00",X"00",
		X"33",X"03",X"FF",X"FF",X"06",X"0A",X"4F",X"03",X"4B",X"03",X"FF",X"FF",X"06",X"0A",X"45",X"02",
		X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",X"FF",X"FF",X"06",X"11",X"52",X"03",X"41",X"03",
		X"4D",X"03",X"00",X"00",X"33",X"03",X"FF",X"FF",X"06",X"18",X"4F",X"03",X"4B",X"03",X"FF",X"FF",
		X"06",X"18",X"45",X"02",X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",X"FF",X"FF",X"07",X"03",
		X"52",X"03",X"4F",X"03",X"4D",X"03",X"00",X"00",X"34",X"03",X"FF",X"FF",X"07",X"0A",X"4F",X"03",
		X"4B",X"03",X"FF",X"FF",X"07",X"0A",X"45",X"02",X"52",X"02",X"52",X"02",X"4F",X"02",X"52",X"02",
		X"FF",X"FF",X"07",X"11",X"52",X"03",X"41",X"03",X"4D",X"03",X"00",X"00",X"34",X"03",X"FF",X"FF",
		X"07",X"18",X"4F",X"03",X"4B",X"03",X"FF",X"FF",X"07",X"18",X"45",X"02",X"52",X"02",X"52",X"02",
		X"4F",X"02",X"52",X"02",X"FF",X"FF",X"08",X"03",X"43",X"01",X"4F",X"01",X"4C",X"01",X"4F",X"01",
		X"52",X"01",X"28",X"01",X"52",X"01",X"47",X"01",X"42",X"01",X"57",X"01",X"29",X"01",X"FF",X"FF",
		X"16",X"03",X"31",X"03",X"50",X"03",X"FF",X"FF",X"18",X"03",X"32",X"03",X"50",X"03",X"FF",X"FF",
		X"1A",X"03",X"43",X"03",X"4F",X"03",X"49",X"03",X"4E",X"03",X"FF",X"FF",X"1C",X"03",X"44",X"03",
		X"49",X"03",X"50",X"03",X"00",X"00",X"53",X"03",X"57",X"03",X"28",X"03",X"31",X"03",X"29",X"03",
		X"FF",X"FF",X"1E",X"03",X"44",X"03",X"49",X"03",X"50",X"03",X"00",X"00",X"53",X"03",X"57",X"03",
		X"28",X"03",X"32",X"03",X"29",X"03",X"FF",X"FF",X"BE",X"C3",X"EE",X"C3",X"36",X"C4",X"7E",X"C4",
		X"C6",X"C4",X"0E",X"C5",X"12",X"C4",X"5A",X"C4",X"A2",X"C4",X"EA",X"C4",X"32",X"C5",X"56",X"C5",
		X"80",X"C5",X"70",X"C5",X"78",X"C5",X"8C",X"C5",X"A2",X"C5",X"E4",X"C5",X"F8",X"C5",X"0C",X"C6",
		X"20",X"C6",X"34",X"C6",X"16",X"0E",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",
		X"30",X"02",X"30",X"02",X"30",X"02",X"FF",X"FF",X"18",X"0E",X"30",X"05",X"30",X"05",X"30",X"05",
		X"30",X"05",X"30",X"05",X"30",X"02",X"30",X"02",X"30",X"02",X"FF",X"FF",X"1A",X"0E",X"30",X"05",
		X"30",X"05",X"30",X"05",X"30",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"FF",X"FF",
		X"1C",X"0E",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",
		X"30",X"05",X"FF",X"FF",X"1E",X"0E",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",X"30",X"05",
		X"30",X"05",X"30",X"05",X"30",X"05",X"FF",X"FF",X"01",X"13",X"43",X"08",X"48",X"08",X"41",X"08",
		X"4E",X"08",X"47",X"08",X"45",X"08",X"00",X"00",X"44",X"08",X"49",X"08",X"53",X"08",X"50",X"08",
		X"FF",X"FF",X"00",X"00",X"0F",X"00",X"0D",X"00",X"0B",X"00",X"09",X"00",X"07",X"00",X"05",X"00",
		X"03",X"00",X"00",X"00",X"F0",X"00",X"D0",X"00",X"B0",X"00",X"90",X"00",X"70",X"00",X"50",X"00",
		X"30",X"00",X"00",X"00",X"00",X"0F",X"00",X"0D",X"00",X"0B",X"00",X"09",X"00",X"07",X"00",X"05",
		X"00",X"03",X"00",X"00",X"FF",X"0F",X"DD",X"0D",X"BB",X"0B",X"99",X"09",X"77",X"07",X"55",X"05",
		X"33",X"03",X"B2",X"C6",X"DE",X"C6",X"0A",X"C7",X"36",X"C7",X"62",X"C7",X"8E",X"C7",X"BA",X"C7",
		X"E6",X"C7",X"0A",X"03",X"03",X"FF",X"05",X"0C",X"00",X"00",X"03",X"FF",X"06",X"0C",X"00",X"00",
		X"03",X"FF",X"07",X"0C",X"00",X"00",X"03",X"FF",X"08",X"0C",X"00",X"00",X"03",X"FF",X"09",X"0C",
		X"00",X"00",X"03",X"FF",X"0A",X"0C",X"00",X"00",X"03",X"FF",X"0B",X"0C",X"FF",X"FF",X"0B",X"03",
		X"03",X"FF",X"05",X"0C",X"00",X"00",X"03",X"FF",X"06",X"0C",X"00",X"00",X"03",X"FF",X"07",X"0C",
		X"00",X"00",X"03",X"FF",X"08",X"0C",X"00",X"00",X"03",X"FF",X"09",X"0C",X"00",X"00",X"03",X"FF",
		X"0A",X"0C",X"00",X"00",X"03",X"FF",X"0B",X"0C",X"FF",X"FF",X"0D",X"03",X"03",X"FF",X"05",X"0D",
		X"00",X"00",X"03",X"FF",X"06",X"0D",X"00",X"00",X"03",X"FF",X"07",X"0D",X"00",X"00",X"03",X"FF",
		X"08",X"0D",X"00",X"00",X"03",X"FF",X"09",X"0D",X"00",X"00",X"03",X"FF",X"0A",X"0D",X"00",X"00",
		X"03",X"FF",X"0B",X"0D",X"FF",X"FF",X"0E",X"03",X"03",X"FF",X"05",X"0D",X"00",X"00",X"03",X"FF",
		X"06",X"0D",X"00",X"00",X"03",X"FF",X"07",X"0D",X"00",X"00",X"03",X"FF",X"08",X"0D",X"00",X"00",
		X"03",X"FF",X"09",X"0D",X"00",X"00",X"03",X"FF",X"0A",X"0D",X"00",X"00",X"03",X"FF",X"0B",X"0D",
		X"FF",X"FF",X"10",X"03",X"03",X"FF",X"05",X"0E",X"00",X"00",X"03",X"FF",X"06",X"0E",X"00",X"00",
		X"03",X"FF",X"07",X"0E",X"00",X"00",X"03",X"FF",X"08",X"0E",X"00",X"00",X"03",X"FF",X"09",X"0E",
		X"00",X"00",X"03",X"FF",X"0A",X"0E",X"00",X"00",X"03",X"FF",X"0B",X"0E",X"FF",X"FF",X"11",X"03",
		X"03",X"FF",X"05",X"0E",X"00",X"00",X"03",X"FF",X"06",X"0E",X"00",X"00",X"03",X"FF",X"07",X"0E",
		X"00",X"00",X"03",X"FF",X"08",X"0E",X"00",X"00",X"03",X"FF",X"09",X"0E",X"00",X"00",X"03",X"FF",
		X"0A",X"0E",X"00",X"00",X"03",X"FF",X"0B",X"0E",X"FF",X"FF",X"13",X"03",X"03",X"FF",X"05",X"0F",
		X"00",X"00",X"03",X"FF",X"06",X"0F",X"00",X"00",X"03",X"FF",X"07",X"0F",X"00",X"00",X"03",X"FF",
		X"08",X"0F",X"00",X"00",X"03",X"FF",X"09",X"0F",X"00",X"00",X"03",X"FF",X"0A",X"0F",X"00",X"00",
		X"03",X"FF",X"0B",X"0F",X"FF",X"FF",X"14",X"03",X"03",X"FF",X"05",X"0F",X"00",X"00",X"03",X"FF",
		X"06",X"0F",X"00",X"00",X"03",X"FF",X"07",X"0F",X"00",X"00",X"03",X"FF",X"08",X"0F",X"00",X"00",
		X"03",X"FF",X"09",X"0F",X"00",X"00",X"03",X"FF",X"0A",X"0F",X"00",X"00",X"03",X"FF",X"0B",X"0F",
		X"FF",X"FF",X"1C",X"0C",X"43",X"06",X"52",X"06",X"45",X"06",X"44",X"06",X"49",X"06",X"54",X"06",
		X"FF",X"FF",X"1C",X"12",X"17",X"80",X"05",X"02",X"48",X"C8",X"60",X"C8",X"78",X"C8",X"90",X"C8",
		X"A8",X"C8",X"C0",X"C8",X"D8",X"C8",X"F0",X"C8",X"08",X"C9",X"20",X"C9",X"38",X"C9",X"50",X"C9",
		X"68",X"C9",X"80",X"C9",X"98",X"C9",X"B0",X"C9",X"42",X"52",X"62",X"72",X"83",X"84",X"85",X"86",
		X"03",X"04",X"05",X"06",X"10",X"20",X"30",X"77",X"67",X"57",X"38",X"28",X"18",X"80",X"70",X"60",
		X"32",X"42",X"52",X"73",X"74",X"75",X"76",X"77",X"25",X"24",X"23",X"13",X"14",X"15",X"16",X"17",
		X"63",X"64",X"65",X"71",X"51",X"41",X"31",X"11",X"23",X"13",X"03",X"04",X"05",X"06",X"07",X"87",
		X"86",X"85",X"84",X"83",X"73",X"63",X"66",X"56",X"36",X"26",X"51",X"41",X"10",X"00",X"70",X"80",
		X"51",X"52",X"53",X"68",X"67",X"66",X"85",X"75",X"65",X"25",X"15",X"05",X"28",X"27",X"26",X"31",
		X"32",X"33",X"10",X"11",X"12",X"70",X"71",X"72",X"71",X"72",X"73",X"75",X"76",X"77",X"51",X"52",
		X"53",X"35",X"36",X"37",X"11",X"12",X"13",X"15",X"16",X"17",X"55",X"56",X"57",X"31",X"32",X"33",
		X"81",X"71",X"61",X"21",X"11",X"01",X"23",X"33",X"53",X"63",X"85",X"75",X"65",X"25",X"15",X"05",
		X"27",X"37",X"57",X"67",X"78",X"88",X"18",X"08",X"56",X"57",X"58",X"54",X"64",X"74",X"36",X"37",
		X"38",X"34",X"24",X"14",X"11",X"21",X"31",X"51",X"61",X"71",X"06",X"07",X"08",X"86",X"87",X"88",
		X"56",X"66",X"76",X"36",X"26",X"16",X"64",X"74",X"84",X"24",X"14",X"04",X"61",X"71",X"81",X"21",
		X"11",X"01",X"08",X"18",X"28",X"68",X"78",X"88",X"06",X"16",X"26",X"35",X"34",X"33",X"53",X"54",
		X"55",X"66",X"76",X"86",X"51",X"61",X"70",X"80",X"31",X"21",X"10",X"00",X"28",X"38",X"58",X"68",
		X"51",X"61",X"71",X"02",X"03",X"04",X"15",X"16",X"17",X"31",X"21",X"11",X"82",X"83",X"84",X"75",
		X"76",X"77",X"55",X"54",X"53",X"33",X"34",X"35",X"23",X"22",X"21",X"11",X"12",X"13",X"16",X"26",
		X"36",X"54",X"64",X"74",X"66",X"67",X"68",X"82",X"72",X"62",X"86",X"87",X"88",X"70",X"60",X"50",
		X"01",X"11",X"21",X"14",X"24",X"34",X"16",X"26",X"36",X"56",X"66",X"76",X"54",X"64",X"74",X"61",
		X"71",X"81",X"52",X"42",X"32",X"50",X"40",X"30",X"51",X"52",X"53",X"64",X"65",X"66",X"22",X"23",
		X"24",X"35",X"36",X"37",X"70",X"71",X"72",X"86",X"87",X"88",X"10",X"11",X"12",X"06",X"07",X"08",
		X"72",X"73",X"74",X"14",X"15",X"16",X"26",X"27",X"28",X"43",X"42",X"41",X"22",X"12",X"02",X"57",
		X"67",X"77",X"84",X"83",X"82",X"60",X"61",X"62",X"00",X"01",X"02",X"13",X"14",X"15",X"74",X"75",
		X"76",X"86",X"87",X"88",X"28",X"18",X"08",X"60",X"70",X"80",X"73",X"83",X"82",X"52",X"42",X"32",
		X"55",X"56",X"57",X"24",X"23",X"22",X"85",X"84",X"83",X"70",X"60",X"50",X"30",X"20",X"10",X"03",
		X"04",X"05",X"62",X"63",X"64",X"37",X"36",X"35",X"18",X"30",X"48",X"60",X"78",X"90",X"A8",X"C0",
		X"D8",X"00",X"03",X"53",X"00",X"49",X"00",X"44",X"00",X"45",X"00",X"2D",X"00",X"4F",X"00",X"4E",
		X"00",X"45",X"00",X"FF",X"FF",X"1E",X"16",X"48",X"00",X"49",X"00",X"2D",X"00",X"53",X"00",X"43",
		X"00",X"4F",X"00",X"52",X"00",X"45",X"00",X"FF",X"FF",X"00",X"15",X"53",X"00",X"49",X"00",X"44",
		X"00",X"45",X"00",X"2D",X"00",X"54",X"00",X"57",X"00",X"4F",X"00",X"FF",X"FF",X"00",X"03",X"53",
		X"0F",X"49",X"0F",X"44",X"0F",X"45",X"0F",X"2D",X"0F",X"4F",X"0F",X"4E",X"0F",X"45",X"0F",X"FF",
		X"FF",X"1E",X"16",X"48",X"0F",X"49",X"0F",X"2D",X"0F",X"53",X"0F",X"43",X"0F",X"4F",X"0F",X"52",
		X"0F",X"45",X"0F",X"FF",X"FF",X"00",X"15",X"53",X"0F",X"49",X"0F",X"44",X"0F",X"45",X"0F",X"2D",
		X"0F",X"54",X"0F",X"57",X"0F",X"30",X"0F",X"FF",X"FF",X"01",X"03",X"B5",X"81",X"05",X"08",X"01",
		X"03",X"9C",X"81",X"05",X"08",X"1F",X"16",X"E2",X"80",X"05",X"08",X"01",X"15",X"CE",X"81",X"05",
		X"08",X"01",X"15",X"9C",X"81",X"05",X"08",X"D1",X"C9",X"E5",X"C9",X"F9",X"C9",X"D1",X"C9",X"E5",
		X"C9",X"97",X"CA",X"9F",X"CA",X"49",X"CA",X"55",X"CA",X"5B",X"CA",X"49",X"CA",X"55",X"CA",X"97",
		X"CA",X"9F",X"CA",X"0D",X"CA",X"E5",X"C9",X"F9",X"C9",X"0D",X"CA",X"E5",X"C9",X"97",X"CA",X"9F",
		X"CA",X"D1",X"C9",X"E5",X"C9",X"35",X"CA",X"00",X"15",X"08",X"FF",X"24",X"00",X"FF",X"FF",X"01",
		X"15",X"08",X"FF",X"24",X"00",X"FF",X"FF",X"1E",X"10",X"52",X"01",X"4F",X"01",X"55",X"01",X"4E",
		X"01",X"44",X"01",X"FF",X"FF",X"1F",X"11",X"B9",X"81",X"03",X"02",X"1F",X"11",X"D2",X"81",X"03",
		X"02",X"1F",X"11",X"AF",X"81",X"03",X"02",X"1F",X"10",X"00",X"00",X"2D",X"03",X"FF",X"FF",X"1F",
		X"10",X"2D",X"03",X"FF",X"FF",X"1F",X"13",X"2D",X"03",X"FF",X"FF",X"FB",X"CA",X"03",X"CB",X"0B",
		X"CB",X"17",X"CB",X"23",X"CB",X"33",X"CB",X"43",X"CB",X"57",X"CB",X"6B",X"CB",X"83",X"CB",X"9B",
		X"CB",X"B7",X"CB",X"D3",X"CB",X"F3",X"CB",X"13",X"CC",X"33",X"CC",X"1E",X"02",X"0E",X"FF",X"24",
		X"00",X"FF",X"FF",X"1F",X"02",X"0E",X"FF",X"24",X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",
		X"00",X"0C",X"FF",X"24",X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0C",X"FF",X"24",
		X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0A",X"FF",X"24",
		X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0A",X"FF",X"24",
		X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",
		X"00",X"08",X"FF",X"24",X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",
		X"00",X"0F",X"00",X"0D",X"00",X"08",X"FF",X"24",X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",
		X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"06",X"FF",X"24",
		X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",
		X"00",X"0F",X"00",X"0D",X"00",X"06",X"FF",X"24",X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",
		X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",
		X"00",X"04",X"FF",X"24",X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",
		X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"04",X"FF",X"24",
		X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",
		X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"02",X"FF",X"24",
		X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",
		X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"02",X"FF",X"24",
		X"00",X"FF",X"FF",X"1E",X"02",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",
		X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0C",
		X"00",X"FF",X"FF",X"1F",X"02",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",
		X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"00",X"6D",X"00",X"6E",X"00",X"6F",
		X"18",X"08",X"06",X"10",X"1E",X"00",X"02",X"05",X"05",X"15",X"02",X"11",X"03",X"01",X"04",X"11",
		X"05",X"01",X"05",X"11",X"04",X"05",X"03",X"15",X"0A",X"05",X"04",X"15",X"04",X"05",X"05",X"15",
		X"06",X"05",X"03",X"01",X"42",X"09",X"01",X"08",X"01",X"00",X"06",X"10",X"03",X"00",X"0C",X"04",
		X"0C",X"06",X"0C",X"02",X"06",X"12",X"05",X"02",X"04",X"12",X"04",X"02",X"07",X"12",X"03",X"02",
		X"0C",X"12",X"05",X"02",X"0B",X"0A",X"0C",X"00",X"08",X"10",X"04",X"04",X"04",X"00",X"01",X"08",
		X"0F",X"09",X"03",X"01",X"11",X"00",X"03",X"10",X"01",X"12",X"02",X"16",X"37",X"06",X"06",X"16",
		X"06",X"06",X"05",X"16",X"02",X"02",X"33",X"00",X"03",X"10",X"05",X"11",X"01",X"01",X"08",X"11",
		X"04",X"01",X"09",X"11",X"01",X"19",X"21",X"09",X"0C",X"00",X"04",X"10",X"02",X"12",X"17",X"06",
		X"02",X"04",X"05",X"05",X"01",X"01",X"05",X"09",X"14",X"19",X"02",X"09",X"03",X"08",X"02",X"0A",
		X"01",X"02",X"07",X"00",X"04",X"10",X"08",X"00",X"06",X"10",X"04",X"18",X"0B",X"08",X"03",X"00",
		X"05",X"10",X"08",X"00",X"01",X"10",X"0B",X"18",X"0A",X"08",X"05",X"00",X"05",X"10",X"07",X"00",
		X"0A",X"18",X"08",X"08",X"07",X"00",X"04",X"10",X"06",X"00",X"03",X"08",X"0B",X"18",X"09",X"08",
		X"0C",X"00",X"20",X"00",X"0C",X"0A",X"0A",X"09",X"6B",X"00",X"12",X"02",X"05",X"12",X"0A",X"06",
		X"03",X"04",X"03",X"05",X"04",X"04",X"0C",X"06",X"04",X"16",X"09",X"12",X"04",X"10",X"1D",X"01",
		X"01",X"00",X"01",X"08",X"11",X"0A",X"01",X"08",X"21",X"00",X"02",X"01",X"03",X"11",X"01",X"10",
		X"02",X"12",X"06",X"02",X"06",X"12",X"0E",X"02",X"06",X"12",X"04",X"02",X"05",X"12",X"01",X"1A",
		X"0C",X"0A",X"57",X"00",X"05",X"10",X"03",X"00",X"38",X"04",X"15",X"05",X"1E",X"01",X"1B",X"09",
		X"05",X"08",X"0D",X"00",X"0C",X"01",X"08",X"11",X"05",X"01",X"06",X"11",X"04",X"01",X"07",X"11",
		X"04",X"01",X"07",X"11",X"06",X"01",X"03",X"09",X"05",X"00",X"05",X"02",X"0A",X"00",X"33",X"02",
		X"57",X"0A",X"05",X"02",X"02",X"12",X"05",X"16",X"3F",X"06",X"04",X"04",X"07",X"05",X"1A",X"01",
		X"A0",X"00",X"12",X"01",X"15",X"00",X"15",X"06",X"10",X"00",X"05",X"05",X"03",X"15",X"03",X"05",
		X"05",X"15",X"03",X"05",X"03",X"15",X"A0",X"05",X"03",X"10",X"5A",X"05",X"03",X"16",X"03",X"06",
		X"03",X"16",X"03",X"06",X"03",X"16",X"03",X"06",X"03",X"16",X"03",X"16",X"03",X"06",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"D0",X"6E",X"D0",X"84",X"D0",X"8C",X"D0",X"0F",X"0E",X"50",X"0F",X"55",X"0F",X"53",X"0F",
		X"48",X"0F",X"FF",X"FF",X"11",X"06",X"31",X"05",X"00",X"00",X"50",X"05",X"4C",X"05",X"41",X"05",
		X"59",X"05",X"45",X"05",X"52",X"05",X"00",X"00",X"42",X"05",X"55",X"05",X"54",X"05",X"54",X"05",
		X"4F",X"05",X"4E",X"05",X"00",X"00",X"4F",X"05",X"4E",X"05",X"4C",X"05",X"59",X"05",X"FF",X"FF",
		X"11",X"06",X"31",X"05",X"00",X"00",X"4F",X"05",X"52",X"05",X"00",X"00",X"32",X"05",X"00",X"00",
		X"50",X"05",X"4C",X"05",X"41",X"05",X"59",X"05",X"45",X"05",X"52",X"05",X"53",X"05",X"00",X"00",
		X"42",X"05",X"55",X"05",X"54",X"05",X"54",X"05",X"4F",X"05",X"4E",X"05",X"FF",X"FF",X"14",X"0B",
		X"50",X"05",X"52",X"05",X"45",X"05",X"53",X"05",X"45",X"05",X"4E",X"05",X"54",X"05",X"45",X"05",
		X"44",X"05",X"FF",X"FF",X"16",X"0F",X"42",X"05",X"59",X"05",X"FF",X"FF",X"18",X"0B",X"54",X"01",
		X"45",X"01",X"48",X"01",X"4B",X"01",X"41",X"01",X"4E",X"01",X"00",X"00",X"4C",X"05",X"54",X"05",
		X"44",X"05",X"2E",X"05",X"FF",X"FF",X"D6",X"D0",X"F0",X"D0",X"D6",X"D0",X"00",X"D1",X"D6",X"D0",
		X"10",X"D1",X"20",X"D1",X"2E",X"D1",X"20",X"D1",X"3E",X"D1",X"4E",X"D1",X"6A",X"D1",X"86",X"D1",
		X"A6",X"D1",X"4E",X"D1",X"6A",X"D1",X"96",X"D1",X"B6",X"D1",X"C6",X"D1",X"E2",X"D1",X"FE",X"D1",
		X"1A",X"D2",X"2A",X"D2",X"3A",X"D2",X"18",X"05",X"45",X"00",X"56",X"00",X"45",X"00",X"52",X"00",
		X"59",X"00",X"00",X"00",X"42",X"00",X"4F",X"00",X"4E",X"00",X"55",X"00",X"53",X"00",X"FF",X"FF",
		X"18",X"12",X"35",X"05",X"04",X"FF",X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",
		X"18",X"11",X"31",X"05",X"05",X"FF",X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",
		X"18",X"12",X"33",X"05",X"04",X"FF",X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",
		X"18",X"08",X"42",X"00",X"4F",X"00",X"4E",X"00",X"55",X"00",X"53",X"00",X"FF",X"FF",X"18",X"0F",
		X"35",X"05",X"04",X"FF",X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"18",X"0E",
		X"31",X"05",X"05",X"FF",X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"17",X"05",
		X"46",X"00",X"49",X"00",X"52",X"00",X"53",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"42",X"00",
		X"4F",X"00",X"4E",X"00",X"55",X"00",X"53",X"00",X"FF",X"FF",X"19",X"05",X"53",X"00",X"45",X"00",
		X"43",X"00",X"4F",X"00",X"4E",X"00",X"44",X"00",X"00",X"00",X"42",X"00",X"4F",X"00",X"4E",X"00",
		X"55",X"00",X"53",X"00",X"FF",X"FF",X"17",X"13",X"35",X"05",X"04",X"FF",X"30",X"05",X"00",X"00",
		X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"17",X"12",X"31",X"05",X"05",X"FF",X"30",X"05",X"00",X"00",
		X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"19",X"12",X"31",X"05",X"05",X"FF",X"30",X"05",X"00",X"00",
		X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"19",X"12",X"33",X"05",X"05",X"FF",X"30",X"05",X"00",X"00",
		X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"16",X"05",X"46",X"00",X"49",X"00",X"52",X"00",X"53",X"00",
		X"54",X"00",X"00",X"00",X"00",X"00",X"42",X"00",X"4F",X"00",X"4E",X"00",X"55",X"00",X"53",X"00",
		X"FF",X"FF",X"18",X"05",X"53",X"00",X"45",X"00",X"43",X"00",X"4F",X"00",X"4E",X"00",X"44",X"00",
		X"00",X"00",X"42",X"00",X"4F",X"00",X"4E",X"00",X"55",X"00",X"53",X"00",X"FF",X"FF",X"1A",X"05",
		X"54",X"00",X"48",X"00",X"49",X"00",X"52",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"42",X"00",
		X"4F",X"00",X"4E",X"00",X"55",X"00",X"53",X"00",X"FF",X"FF",X"16",X"13",X"35",X"05",X"04",X"FF",
		X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"18",X"12",X"31",X"05",X"05",X"FF",
		X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"1A",X"12",X"33",X"05",X"05",X"FF",
		X"30",X"05",X"00",X"00",X"3E",X"05",X"3C",X"05",X"FF",X"FF",X"0A",X"09",X"59",X"0F",X"4F",X"0F",
		X"55",X"0F",X"00",X"00",X"41",X"0F",X"52",X"0F",X"45",X"0F",X"00",X"00",X"4C",X"0F",X"55",X"0F",
		X"43",X"0F",X"4B",X"0F",X"59",X"0F",X"FF",X"FF",X"59",X"05",X"4F",X"05",X"55",X"05",X"00",X"0A",
		X"43",X"05",X"41",X"05",X"4E",X"05",X"00",X"0A",X"45",X"05",X"4E",X"05",X"4A",X"05",X"4F",X"05",
		X"59",X"05",X"FF",X"59",X"05",X"41",X"05",X"4C",X"05",X"50",X"05",X"00",X"0A",X"45",X"05",X"52",
		X"05",X"4F",X"05",X"4D",X"05",X"00",X"0A",X"45",X"05",X"4E",X"05",X"4F",X"05",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0F",X"CE",X"08",X"FF",X"0F",X"0F",X"00",X"A0",X"0F",X"FF",X"00",
		X"00",X"00",X"2A",X"00",X"50",X"00",X"A0",X"00",X"88",X"08",X"66",X"06",X"44",X"04",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"44",X"04",X"88",X"08",X"CC",X"0C",X"FF",X"0F",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"44",X"04",X"88",X"08",X"CC",X"0C",X"FF",X"0F",X"F0",X"0F",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"55",X"05",X"88",X"08",X"BB",X"0B",X"DD",X"0D",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"DD",X"00",X"AA",X"0A",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"44",X"04",X"88",X"08",X"CC",X"0C",X"FF",X"0F",X"8F",X"00",
		X"00",X"00",X"88",X"00",X"FF",X"0F",X"FF",X"0F",X"F6",X"06",X"FF",X"0F",X"FF",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"0F",X"6F",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"0F",X"FF",X"0F",X"AF",X"0C",
		X"00",X"00",X"88",X"08",X"AA",X"08",X"CC",X"0C",X"80",X"00",X"A0",X"00",X"C0",X"00",X"0A",X"0F",
		X"00",X"00",X"88",X"08",X"88",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"DD",X"00",X"AA",X"0A",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"44",X"04",X"66",X"06",X"88",X"08",X"AA",X"0A",X"FF",X"0F",X"CC",X"0C",X"47",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"07",X"00",X"17",X"00",X"27",X"00",X"37",X"00",X"47",X"00",X"57",X"00",X"67",X"00",
		X"00",X"00",X"77",X"00",X"77",X"01",X"77",X"02",X"77",X"03",X"77",X"04",X"77",X"05",X"77",X"06",
		X"00",X"00",X"3F",X"00",X"5F",X"00",X"7F",X"00",X"9F",X"00",X"BF",X"00",X"DF",X"00",X"FF",X"00",
		X"00",X"00",X"40",X"00",X"60",X"00",X"80",X"00",X"A0",X"00",X"C0",X"00",X"E0",X"00",X"F0",X"00",
		X"00",X"00",X"3F",X"00",X"5F",X"00",X"7F",X"00",X"9F",X"00",X"BF",X"00",X"DF",X"00",X"FF",X"00",
		X"00",X"00",X"55",X"00",X"77",X"00",X"99",X"00",X"BB",X"00",X"DD",X"00",X"FF",X"00",X"FF",X"04",
		X"00",X"00",X"00",X"08",X"00",X"0C",X"00",X"0F",X"80",X"0F",X"A0",X"0F",X"C0",X"0F",X"F0",X"0F",
		X"00",X"00",X"00",X"0F",X"C0",X"00",X"F0",X"00",X"F8",X"00",X"F0",X"00",X"FF",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"0F",X"5C",X"00",X"8F",X"00",X"FF",X"00",X"8F",X"00",X"FF",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"0F",X"0F",X"00",X"4F",X"04",X"8F",X"08",X"4F",X"04",X"CF",X"0C",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"0C",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"0C",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"0C",X"FF",X"0F",
		X"00",X"00",X"58",X"0B",X"45",X"00",X"67",X"02",X"89",X"04",X"AB",X"06",X"CD",X"08",X"EF",X"0A",
		X"00",X"00",X"00",X"0C",X"00",X"0B",X"00",X"0A",X"00",X"09",X"00",X"08",X"00",X"07",X"00",X"06",
		X"00",X"00",X"00",X"0C",X"45",X"00",X"67",X"02",X"89",X"04",X"AB",X"06",X"CD",X"08",X"EF",X"0A",
		X"00",X"00",X"88",X"0C",X"50",X"00",X"A0",X"00",X"88",X"08",X"66",X"06",X"44",X"04",X"22",X"02",
		X"00",X"00",X"00",X"0C",X"00",X"0B",X"00",X"0A",X"00",X"09",X"00",X"08",X"88",X"08",X"AA",X"0A",
		X"00",X"00",X"44",X"04",X"44",X"04",X"00",X"00",X"30",X"03",X"50",X"05",X"70",X"07",X"05",X"07",
		X"00",X"00",X"44",X"04",X"44",X"04",X"00",X"00",X"33",X"00",X"55",X"00",X"77",X"00",X"05",X"07",
		X"00",X"00",X"44",X"04",X"44",X"04",X"00",X"00",X"33",X"03",X"55",X"05",X"77",X"07",X"05",X"07",
		X"00",X"00",X"05",X"00",X"50",X"00",X"80",X"00",X"28",X"00",X"4A",X"00",X"06",X"00",X"45",X"00",
		X"00",X"00",X"27",X"00",X"08",X"0C",X"40",X"00",X"CC",X"0C",X"0D",X"00",X"80",X"00",X"CC",X"00",
		X"00",X"00",X"0F",X"00",X"55",X"05",X"77",X"07",X"99",X"09",X"BB",X"0B",X"DD",X"0D",X"00",X"0F",
		X"00",X"00",X"88",X"0C",X"2A",X"00",X"AA",X"0A",X"88",X"08",X"66",X"06",X"44",X"04",X"22",X"02",
		X"00",X"00",X"60",X"0C",X"55",X"05",X"77",X"07",X"99",X"09",X"BB",X"0B",X"DD",X"0D",X"A0",X"00",
		X"00",X"00",X"00",X"07",X"37",X"00",X"77",X"00",X"10",X"01",X"30",X"03",X"50",X"05",X"57",X"06",
		X"00",X"00",X"00",X"07",X"37",X"00",X"77",X"00",X"11",X"00",X"33",X"00",X"55",X"00",X"57",X"06",
		X"00",X"00",X"00",X"07",X"37",X"00",X"77",X"00",X"11",X"01",X"33",X"03",X"55",X"05",X"57",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"77",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"04",X"66",X"06",X"88",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"66",X"00",X"77",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",
		X"00",X"00",X"44",X"04",X"55",X"05",X"66",X"06",X"77",X"07",X"77",X"07",X"77",X"07",X"77",X"07",
		X"CC",X"CD",X"CE",X"CF",X"15",X"94",X"95",X"96",X"97",X"0D",X"CC",X"CD",X"CE",X"CF",X"15",X"94",
		X"95",X"96",X"97",X"0D",X"CC",X"CD",X"CE",X"CF",X"15",X"94",X"95",X"96",X"97",X"0D",X"CC",X"CD",
		X"CE",X"CF",X"15",X"94",X"95",X"96",X"97",X"0D",X"CC",X"CD",X"CE",X"CF",X"15",X"94",X"95",X"96",
		X"97",X"0D",X"CC",X"CD",X"CE",X"CF",X"15",X"94",X"95",X"96",X"97",X"0D",X"D8",X"D9",X"DA",X"DB",
		X"15",X"90",X"91",X"92",X"93",X"0D",X"DC",X"DD",X"DE",X"DF",X"15",X"90",X"91",X"92",X"93",X"0D",
		X"04",X"00",X"00",X"01",X"C0",X"00",X"00",X"02",X"05",X"00",X"00",X"01",X"C0",X"00",X"00",X"02",
		X"06",X"00",X"C0",X"00",X"80",X"00",X"00",X"02",X"07",X"00",X"C0",X"00",X"80",X"00",X"00",X"01",
		X"07",X"00",X"80",X"00",X"60",X"00",X"00",X"02",X"04",X"00",X"80",X"00",X"40",X"00",X"00",X"01",
		X"05",X"00",X"60",X"00",X"60",X"00",X"00",X"01",X"06",X"00",X"60",X"00",X"40",X"00",X"00",X"01",
		X"07",X"00",X"60",X"00",X"40",X"00",X"00",X"01",X"07",X"00",X"20",X"00",X"40",X"00",X"00",X"01",
		X"04",X"00",X"80",X"00",X"30",X"00",X"00",X"01",X"05",X"00",X"80",X"00",X"30",X"00",X"00",X"01",
		X"06",X"00",X"60",X"00",X"30",X"00",X"00",X"01",X"07",X"00",X"60",X"00",X"30",X"00",X"00",X"01",
		X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",X"04",X"00",X"60",X"00",X"20",X"00",X"00",X"01",
		X"05",X"00",X"60",X"00",X"20",X"00",X"00",X"01",X"06",X"00",X"40",X"00",X"20",X"00",X"00",X"01",
		X"07",X"00",X"40",X"00",X"20",X"00",X"00",X"01",X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",
		X"04",X"00",X"40",X"00",X"20",X"00",X"00",X"01",X"05",X"00",X"40",X"00",X"20",X"00",X"00",X"01",
		X"06",X"00",X"40",X"00",X"20",X"00",X"00",X"01",X"07",X"00",X"40",X"00",X"20",X"00",X"00",X"01",
		X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",X"04",X"00",X"20",X"00",X"20",X"00",X"00",X"01",
		X"05",X"00",X"20",X"00",X"20",X"00",X"00",X"01",X"06",X"00",X"20",X"00",X"20",X"00",X"00",X"01",
		X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",
		X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",
		X"07",X"00",X"20",X"00",X"20",X"00",X"00",X"01",X"01",X"00",X"20",X"00",X"44",X"00",X"80",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"30",X"00",X"55",X"00",X"80",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"38",X"00",X"66",X"00",X"80",X"00",X"03",X"00",X"00",X"00",X"01",X"00",X"40",X"00",
		X"55",X"00",X"70",X"00",X"03",X"00",X"00",X"00",X"01",X"00",X"40",X"00",X"66",X"00",X"70",X"00",
		X"04",X"00",X"00",X"00",X"01",X"00",X"40",X"00",X"77",X"00",X"70",X"00",X"04",X"00",X"00",X"00",
		X"01",X"00",X"48",X"00",X"66",X"00",X"60",X"00",X"05",X"00",X"00",X"00",X"01",X"00",X"48",X"00",
		X"77",X"00",X"60",X"00",X"05",X"00",X"00",X"00",X"01",X"00",X"48",X"00",X"88",X"00",X"60",X"00",
		X"06",X"00",X"00",X"00",X"02",X"00",X"40",X"00",X"55",X"00",X"80",X"00",X"06",X"00",X"00",X"00",
		X"02",X"00",X"40",X"00",X"66",X"00",X"80",X"00",X"07",X"00",X"00",X"00",X"02",X"00",X"40",X"00",
		X"77",X"00",X"80",X"00",X"07",X"00",X"00",X"00",X"02",X"00",X"48",X"00",X"66",X"00",X"70",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"48",X"00",X"77",X"00",X"70",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"48",X"00",X"88",X"00",X"70",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"50",X"00",
		X"77",X"00",X"60",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"50",X"00",X"88",X"00",X"60",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"50",X"00",X"99",X"00",X"60",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"58",X"00",X"88",X"00",X"60",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"50",X"00",
		X"77",X"00",X"80",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"50",X"00",X"88",X"00",X"80",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"58",X"00",X"77",X"00",X"80",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"58",X"00",X"88",X"00",X"70",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"58",X"00",
		X"99",X"00",X"70",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"60",X"00",X"88",X"00",X"70",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"60",X"00",X"99",X"00",X"60",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"60",X"00",X"A2",X"00",X"60",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"68",X"00",
		X"99",X"00",X"60",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"68",X"00",X"A2",X"00",X"50",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"68",X"00",X"AA",X"00",X"50",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"70",X"00",X"A2",X"00",X"50",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"70",X"00",
		X"AA",X"00",X"48",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"70",X"00",X"B3",X"00",X"48",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"78",X"00",X"AA",X"00",X"48",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"78",X"00",X"B3",X"00",X"40",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"78",X"00",
		X"BB",X"00",X"40",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"80",X"00",X"B3",X"00",X"40",X"00",
		X"08",X"00",X"00",X"00",X"02",X"00",X"80",X"00",X"BB",X"00",X"38",X"00",X"08",X"00",X"00",X"00",
		X"02",X"00",X"80",X"00",X"C4",X"00",X"38",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"80",X"00",
		X"BB",X"00",X"38",X"00",X"08",X"00",X"00",X"00",X"80",X"00",X"00",X"01",X"01",X"00",X"00",X"02",
		X"01",X"00",X"00",X"04",X"B3",X"B3",X"B3",X"B4",X"B3",X"B3",X"B3",X"B4",X"91",X"00",X"C0",X"00",
		X"02",X"00",X"80",X"01",X"01",X"00",X"00",X"03",X"B1",X"B1",X"B1",X"B4",X"B1",X"B1",X"B1",X"B4",
		X"A2",X"00",X"C0",X"00",X"03",X"00",X"00",X"01",X"01",X"00",X"00",X"02",X"B2",X"B2",X"B2",X"B4",
		X"B2",X"B2",X"B2",X"B4",X"AE",X"00",X"80",X"00",X"04",X"00",X"C0",X"00",X"01",X"00",X"80",X"01",
		X"B0",X"B0",X"B0",X"B4",X"B0",X"B0",X"B0",X"B4",X"C0",X"00",X"80",X"00",X"05",X"00",X"C0",X"00",
		X"04",X"00",X"00",X"03",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"D1",X"00",X"80",X"00",
		X"06",X"00",X"C0",X"00",X"03",X"00",X"80",X"01",X"B2",X"B2",X"B1",X"B1",X"B2",X"B2",X"B3",X"B3",
		X"80",X"01",X"80",X"00",X"07",X"00",X"C0",X"00",X"03",X"00",X"80",X"01",X"B0",X"B1",X"B2",X"B3",
		X"B4",X"B3",X"B2",X"B1",X"EE",X"00",X"80",X"00",X"08",X"00",X"C0",X"00",X"03",X"00",X"80",X"01",
		X"B0",X"B0",X"B1",X"B1",X"B0",X"B0",X"B1",X"B1",X"00",X"01",X"80",X"00",X"09",X"00",X"C0",X"00",
		X"03",X"00",X"80",X"01",X"B3",X"B3",X"B4",X"B4",X"B3",X"B3",X"B4",X"B4",X"00",X"01",X"80",X"00",
		X"0A",X"00",X"C0",X"00",X"03",X"00",X"80",X"01",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",
		X"00",X"01",X"80",X"00",X"0B",X"00",X"C0",X"00",X"04",X"00",X"80",X"01",X"B4",X"B3",X"B4",X"B3",
		X"B0",X"B1",X"B0",X"B1",X"00",X"01",X"80",X"00",X"0C",X"00",X"C0",X"00",X"04",X"00",X"80",X"01",
		X"B1",X"B2",X"B1",X"B2",X"B1",X"B2",X"B1",X"B2",X"00",X"01",X"80",X"00",X"0D",X"00",X"C0",X"00",
		X"04",X"00",X"80",X"01",X"B3",X"B0",X"B3",X"B0",X"B3",X"B0",X"B3",X"B0",X"00",X"01",X"80",X"00",
		X"0E",X"00",X"C0",X"00",X"05",X"00",X"80",X"01",X"B4",X"B4",X"B4",X"B1",X"B4",X"B4",X"B4",X"B1",
		X"00",X"02",X"80",X"00",X"0F",X"00",X"C0",X"00",X"05",X"00",X"80",X"01",X"B0",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"B0",X"B0",X"00",X"01",X"80",X"00",X"10",X"00",X"C0",X"00",X"05",X"00",X"80",X"01",
		X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"80",X"01",X"80",X"00",X"11",X"00",X"C0",X"00",
		X"05",X"00",X"80",X"01",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"80",X"01",X"80",X"00",
		X"12",X"00",X"C0",X"00",X"05",X"00",X"80",X"01",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",
		X"80",X"01",X"80",X"00",X"13",X"00",X"C0",X"00",X"06",X"00",X"80",X"01",X"B4",X"B4",X"B4",X"B4",
		X"B4",X"B4",X"B4",X"B4",X"80",X"01",X"80",X"00",X"14",X"00",X"C0",X"00",X"06",X"00",X"80",X"01",
		X"B0",X"B0",X"B4",X"B4",X"B2",X"B2",X"B4",X"B4",X"80",X"01",X"80",X"00",X"15",X"00",X"C0",X"00",
		X"06",X"00",X"80",X"01",X"B0",X"B0",X"B0",X"B0",X"B1",X"B1",X"B1",X"B1",X"80",X"01",X"80",X"00",
		X"16",X"00",X"C0",X"00",X"06",X"00",X"80",X"01",X"B1",X"B1",X"B1",X"B1",X"B2",X"B2",X"B2",X"B2",
		X"80",X"01",X"80",X"00",X"17",X"00",X"C0",X"00",X"06",X"00",X"80",X"01",X"B2",X"B2",X"B2",X"B2",
		X"B3",X"B3",X"B3",X"B3",X"80",X"01",X"80",X"00",X"18",X"00",X"C0",X"00",X"07",X"00",X"80",X"01",
		X"B3",X"B3",X"B3",X"B3",X"B4",X"B4",X"B4",X"B4",X"00",X"02",X"80",X"00",X"19",X"00",X"C0",X"00",
		X"07",X"00",X"80",X"01",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"00",X"02",X"80",X"00",
		X"1A",X"00",X"C0",X"00",X"07",X"00",X"80",X"01",X"B4",X"B4",X"B4",X"B4",X"B0",X"B0",X"B0",X"B0",
		X"00",X"02",X"80",X"00",X"1B",X"00",X"C0",X"00",X"07",X"00",X"80",X"01",X"B3",X"B3",X"B3",X"B3",
		X"B1",X"B1",X"B1",X"B1",X"00",X"02",X"80",X"00",X"1C",X"00",X"C0",X"00",X"08",X"00",X"80",X"01",
		X"B2",X"B2",X"B2",X"B2",X"B4",X"B4",X"B4",X"B4",X"00",X"02",X"80",X"00",X"1D",X"00",X"C0",X"00",
		X"08",X"00",X"80",X"01",X"B0",X"B0",X"B0",X"B0",X"B3",X"B3",X"B3",X"B3",X"00",X"02",X"80",X"00",
		X"1E",X"00",X"C0",X"00",X"09",X"00",X"80",X"01",X"B4",X"B3",X"B4",X"B2",X"B4",X"B1",X"B4",X"B0",
		X"00",X"02",X"80",X"00",X"1F",X"00",X"C0",X"00",X"09",X"00",X"80",X"01",X"B0",X"B1",X"B2",X"B3",
		X"B4",X"B0",X"B1",X"B2",X"00",X"02",X"80",X"00",X"20",X"00",X"C0",X"00",X"09",X"00",X"80",X"01",
		X"B3",X"B4",X"B0",X"B1",X"B2",X"B3",X"B4",X"B0",X"00",X"00",X"02",X"00",X"00",X"00",X"0B",X"01",
		X"00",X"0B",X"01",X"01",X"08",X"02",X"03",X"08",X"02",X"02",X"07",X"03",X"04",X"07",X"03",X"00",
		X"04",X"04",X"01",X"04",X"04",X"01",X"02",X"00",X"02",X"02",X"00",X"02",X"06",X"01",X"00",X"06",
		X"01",X"00",X"03",X"02",X"03",X"03",X"02",X"01",X"0A",X"03",X"04",X"0A",X"03",X"02",X"04",X"04",
		X"01",X"00",X"04",X"00",X"0C",X"00",X"02",X"0C",X"00",X"01",X"0E",X"01",X"00",X"0E",X"01",X"02",
		X"09",X"02",X"03",X"09",X"02",X"00",X"0F",X"03",X"04",X"0F",X"03",X"01",X"04",X"04",X"01",X"04",
		X"04",X"02",X"0D",X"00",X"02",X"0D",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"01",X"05",X"02",
		X"03",X"05",X"02",X"02",X"0B",X"03",X"04",X"0B",X"03",X"00",X"04",X"04",X"01",X"0D",X"04",X"01",
		X"0E",X"00",X"02",X"0E",X"00",X"02",X"06",X"01",X"00",X"06",X"01",X"00",X"07",X"02",X"03",X"07",
		X"02",X"01",X"09",X"03",X"04",X"09",X"03",X"02",X"04",X"04",X"01",X"0F",X"04",X"00",X"05",X"00",
		X"02",X"05",X"00",X"01",X"03",X"01",X"00",X"03",X"01",X"02",X"01",X"02",X"03",X"01",X"02",X"00",
		X"0C",X"03",X"04",X"0C",X"03",X"01",X"04",X"04",X"01",X"00",X"04",X"02",X"02",X"00",X"02",X"02",
		X"00",X"00",X"08",X"01",X"00",X"08",X"01",X"01",X"0F",X"02",X"03",X"0F",X"02",X"02",X"0D",X"03",
		X"04",X"0D",X"03",X"00",X"04",X"04",X"01",X"06",X"04",X"01",X"0A",X"00",X"02",X"0A",X"00",X"02",
		X"09",X"01",X"00",X"09",X"01",X"00",X"01",X"02",X"03",X"01",X"02",X"01",X"02",X"03",X"04",X"02",
		X"03",X"02",X"04",X"04",X"01",X"02",X"04",X"00",X"03",X"00",X"02",X"03",X"00",X"01",X"05",X"01",
		X"00",X"05",X"01",X"02",X"06",X"02",X"03",X"06",X"02",X"00",X"07",X"00",X"04",X"07",X"03",X"01",
		X"04",X"01",X"01",X"0E",X"04",X"02",X"08",X"02",X"02",X"08",X"00",X"00",X"09",X"03",X"00",X"09",
		X"01",X"01",X"0A",X"04",X"03",X"0A",X"02",X"02",X"0B",X"00",X"04",X"0B",X"03",X"00",X"04",X"01",
		X"01",X"0A",X"04",X"01",X"0C",X"02",X"02",X"0C",X"00",X"02",X"0D",X"03",X"00",X"0D",X"01",X"00",
		X"0E",X"04",X"03",X"0E",X"02",X"01",X"0F",X"00",X"04",X"0F",X"03",X"02",X"04",X"01",X"01",X"06",
		X"04",X"00",X"00",X"02",X"02",X"00",X"00",X"01",X"01",X"03",X"00",X"01",X"01",X"02",X"02",X"04",
		X"03",X"02",X"02",X"00",X"03",X"00",X"04",X"03",X"03",X"01",X"04",X"01",X"01",X"08",X"04",X"02",
		X"05",X"02",X"02",X"05",X"00",X"00",X"06",X"03",X"00",X"06",X"01",X"01",X"07",X"04",X"03",X"07",
		X"02",X"02",X"08",X"00",X"04",X"08",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CB",X"01",X"E1",X"E1",X"E1",X"E1",X"08",X"80",X"02",X"E0",X"02",X"08",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
