library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"34",X"00",X"86",X"15",X"E5",X"14",X"51",X"34",X"46",X"B9",X"08",X"BA",X"04",X"BB",X"00",X"23",
		X"AA",X"AF",X"AE",X"B8",X"40",X"B0",X"02",X"94",X"10",X"94",X"10",X"FA",X"97",X"A7",X"F7",X"AA",
		X"94",X"10",X"94",X"10",X"FA",X"97",X"F7",X"AA",X"E9",X"17",X"86",X"2A",X"B9",X"0E",X"BA",X"30",
		X"B8",X"22",X"27",X"A0",X"18",X"A0",X"B8",X"40",X"A0",X"F4",X"00",X"F4",X"00",X"F4",X"69",X"F4",
		X"0D",X"F4",X"0D",X"F4",X"69",X"F4",X"1A",X"F4",X"1A",X"F4",X"69",X"E9",X"39",X"05",X"34",X"13",
		X"24",X"93",X"BA",X"30",X"B8",X"22",X"B0",X"00",X"18",X"B0",X"00",X"BB",X"00",X"B8",X"40",X"B0",
		X"01",X"34",X"55",X"14",X"6F",X"80",X"92",X"63",X"14",X"6F",X"80",X"92",X"52",X"04",X"68",X"34",
		X"55",X"B8",X"23",X"F0",X"03",X"1C",X"A0",X"F6",X"A5",X"83",X"B9",X"0C",X"BA",X"10",X"27",X"B8",
		X"22",X"A0",X"18",X"A0",X"AB",X"85",X"95",X"A5",X"F4",X"00",X"14",X"A8",X"E9",X"88",X"F4",X"00",
		X"14",X"A8",X"80",X"B2",X"8E",X"1A",X"F4",X"00",X"14",X"A8",X"80",X"B2",X"7A",X"B8",X"23",X"F0",
		X"03",X"08",X"A0",X"E6",X"95",X"34",X"13",X"B3",X"80",X"F2",X"A5",X"D2",X"A5",X"09",X"53",X"0F",
		X"96",X"A5",X"36",X"A5",X"56",X"A5",X"83",X"BA",X"0A",X"B8",X"22",X"B0",X"01",X"18",X"B0",X"00",
		X"85",X"95",X"A5",X"F4",X"64",X"F6",X"A5",X"B8",X"23",X"F0",X"03",X"14",X"F6",X"A5",X"F4",X"00",
		X"80",X"F2",X"A5",X"F4",X"00",X"80",X"F2",X"A5",X"F4",X"00",X"80",X"F2",X"A5",X"14",X"C3",X"F6",
		X"A5",X"C6",X"B9",X"60",X"BA",X"FF",X"BB",X"00",X"27",X"AE",X"AF",X"B8",X"40",X"B0",X"02",X"85",
		X"94",X"10",X"C9",X"F9",X"C6",X"A5",X"53",X"0F",X"96",X"F0",X"FA",X"97",X"67",X"AA",X"04",X"F0",
		X"F6",X"55",X"27",X"B8",X"20",X"A0",X"B8",X"21",X"A0",X"B8",X"24",X"A0",X"D5",X"AE",X"AF",X"C5",
		X"34",X"13",X"E9",X"34",X"45",X"36",X"6B",X"56",X"C5",X"09",X"12",X"37",X"32",X"F2",X"52",X"39",
		X"72",X"3B",X"80",X"F2",X"43",X"D2",X"41",X"B2",X"3F",X"92",X"3D",X"53",X"0F",X"03",X"F9",X"C6",
		X"35",X"94",X"10",X"24",X"13",X"44",X"3D",X"44",X"2A",X"44",X"00",X"24",X"8D",X"04",X"52",X"04",
		X"7A",X"04",X"B7",X"04",X"E2",X"05",X"C5",X"27",X"AE",X"AF",X"85",X"A5",X"B8",X"40",X"A0",X"B8",
		X"22",X"A0",X"18",X"A0",X"83",X"85",X"95",X"A5",X"B5",X"F4",X"0D",X"F4",X"0D",X"83",X"85",X"95",
		X"A5",X"B5",X"F4",X"0D",X"36",X"6B",X"F4",X"0D",X"36",X"6B",X"83",X"B9",X"02",X"BA",X"60",X"B8",
		X"22",X"B0",X"00",X"18",X"B0",X"00",X"B8",X"40",X"B0",X"01",X"34",X"55",X"E9",X"7A",X"BA",X"80",
		X"34",X"5E",X"B8",X"23",X"F0",X"03",X"0D",X"A0",X"E6",X"80",X"34",X"13",X"E9",X"B9",X"04",X"BA",
		X"40",X"B8",X"22",X"B0",X"00",X"18",X"B0",X"00",X"B8",X"40",X"B0",X"01",X"34",X"B6",X"B9",X"04",
		X"B8",X"23",X"B0",X"00",X"BB",X"00",X"F4",X"58",X"34",X"B6",X"B9",X"40",X"B8",X"23",X"B0",X"00",
		X"BB",X"00",X"F4",X"58",X"34",X"B6",X"F4",X"64",X"34",X"5E",X"B8",X"23",X"F0",X"03",X"10",X"A0",
		X"F6",X"13",X"E9",X"B6",X"83",X"B9",X"06",X"BA",X"20",X"B8",X"22",X"B0",X"00",X"18",X"B0",X"00",
		X"85",X"95",X"A5",X"F4",X"00",X"E9",X"D3",X"F4",X"69",X"B8",X"23",X"F0",X"03",X"08",X"A0",X"F6",
		X"13",X"F4",X"00",X"F4",X"00",X"E6",X"D7",X"C6",X"D7",X"17",X"C6",X"D7",X"F9",X"E3",X"96",X"D7",
		X"24",X"D5",X"B9",X"10",X"BA",X"40",X"BB",X"00",X"F4",X"69",X"F4",X"00",X"E9",X"F8",X"24",X"13",
		X"B9",X"30",X"BA",X"20",X"BB",X"40",X"B8",X"38",X"B0",X"04",X"F4",X"58",X"F4",X"1A",X"B8",X"38",
		X"F0",X"07",X"A0",X"C6",X"19",X"E9",X"0A",X"24",X"13",X"B0",X"04",X"F4",X"5D",X"F4",X"1A",X"B8",
		X"38",X"F0",X"07",X"A0",X"C6",X"06",X"E9",X"1B",X"24",X"13",X"B9",X"10",X"BA",X"30",X"B8",X"22",
		X"B0",X"E8",X"18",X"B0",X"E0",X"F4",X"58",X"F4",X"0D",X"E9",X"35",X"24",X"13",X"B8",X"30",X"B0",
		X"45",X"18",X"B0",X"0C",X"B8",X"40",X"B0",X"04",X"A5",X"27",X"62",X"44",X"68",X"80",X"F2",X"54",
		X"53",X"0F",X"96",X"56",X"24",X"13",X"94",X"10",X"E5",X"B8",X"23",X"F0",X"03",X"08",X"E6",X"65",
		X"27",X"AE",X"AF",X"44",X"66",X"A0",X"E9",X"4D",X"D4",X"9F",X"F8",X"C6",X"3D",X"44",X"4D",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"04",X"08",X"0C",X"10",X"14",X"18",X"1C",X"20",X"24",X"28",X"2C",X"30",X"34",X"38",X"3C",
		X"40",X"44",X"48",X"4C",X"50",X"54",X"58",X"5C",X"60",X"64",X"68",X"6C",X"70",X"74",X"78",X"7C",
		X"60",X"03",X"06",X"09",X"0C",X"0F",X"12",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",
		X"30",X"33",X"36",X"39",X"3C",X"3F",X"42",X"45",X"48",X"4B",X"4E",X"51",X"54",X"57",X"5A",X"5D",
		X"40",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0E",X"10",X"12",X"14",X"16",X"18",X"1A",X"1C",X"1E",
		X"20",X"22",X"24",X"26",X"28",X"2A",X"2C",X"2E",X"30",X"32",X"34",X"36",X"38",X"3A",X"3C",X"3E",
		X"30",X"01",X"03",X"04",X"06",X"07",X"09",X"0A",X"0C",X"0D",X"0F",X"10",X"12",X"13",X"15",X"16",
		X"18",X"19",X"1B",X"1C",X"1E",X"1F",X"21",X"22",X"24",X"25",X"27",X"28",X"2A",X"2B",X"2D",X"2E",
		X"20",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",
		X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"18",X"00",X"01",X"02",X"03",X"03",X"04",X"05",X"06",X"06",X"07",X"08",X"09",X"09",X"0A",X"0B",
		X"0C",X"0C",X"0D",X"0E",X"0F",X"0F",X"10",X"11",X"12",X"12",X"13",X"14",X"15",X"15",X"16",X"17",
		X"10",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"06",X"07",X"07",
		X"08",X"08",X"09",X"09",X"0A",X"0A",X"0B",X"0B",X"0C",X"0C",X"0D",X"0D",X"0E",X"0E",X"0F",X"0F",
		X"0C",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"03",X"04",X"04",X"04",X"05",X"05",
		X"06",X"06",X"06",X"07",X"07",X"07",X"08",X"08",X"09",X"09",X"09",X"0A",X"0A",X"0A",X"0B",X"0B",
		X"00",X"E0",X"01",X"80",X"20",X"40",X"C0",X"00",X"04",X"10",X"09",X"12",X"13",X"60",X"05",X"A0",
		X"D5",X"B8",X"20",X"80",X"53",X"0F",X"20",X"37",X"17",X"60",X"96",X"55",X"B8",X"21",X"F0",X"C6",
		X"3C",X"F2",X"E2",X"D2",X"E4",X"B2",X"E6",X"52",X"D2",X"E9",X"3C",X"FF",X"96",X"31",X"FE",X"C6",
		X"91",X"FA",X"03",X"F8",X"A9",X"F6",X"39",X"B9",X"01",X"27",X"AE",X"AF",X"B8",X"40",X"F0",X"12",
		X"48",X"32",X"4B",X"52",X"4E",X"F5",X"24",X"6F",X"F5",X"44",X"00",X"F5",X"44",X"7E",X"F5",X"24",
		X"00",X"B8",X"21",X"B0",X"00",X"B8",X"21",X"F0",X"03",X"FC",X"C6",X"D2",X"B8",X"20",X"F0",X"A3",
		X"92",X"E8",X"72",X"EA",X"F2",X"DC",X"D2",X"DE",X"B2",X"E0",X"52",X"AA",X"B8",X"21",X"F0",X"F2",
		X"E2",X"D2",X"E4",X"B2",X"E6",X"52",X"D2",X"12",X"29",X"B0",X"00",X"B8",X"20",X"F0",X"A3",X"52",
		X"AC",X"C6",X"EC",X"B8",X"21",X"A0",X"E7",X"43",X"F0",X"A8",X"B9",X"30",X"B1",X"03",X"19",X"B1",
		X"0B",X"B8",X"30",X"D4",X"36",X"B8",X"20",X"F9",X"C6",X"51",X"B9",X"08",X"B8",X"24",X"B0",X"00",
		X"FA",X"03",X"F8",X"F6",X"3C",X"FA",X"07",X"A9",X"84",X"3C",X"12",X"6C",X"B8",X"21",X"A0",X"12",
		X"BA",X"B9",X"32",X"B1",X"14",X"19",X"B1",X"0B",X"84",X"C1",X"B9",X"32",X"B1",X"27",X"19",X"B1",
		X"0B",X"B8",X"32",X"D4",X"36",X"B8",X"20",X"F9",X"C6",X"51",X"B8",X"24",X"B0",X"00",X"FA",X"A9",
		X"84",X"3C",X"B8",X"24",X"F0",X"03",X"10",X"A0",X"E9",X"3C",X"84",X"C1",X"A4",X"00",X"A4",X"2B",
		X"A4",X"4B",X"A4",X"0F",X"A4",X"38",X"A4",X"56",X"C4",X"5F",X"C4",X"B7",X"27",X"AE",X"AF",X"84",
		X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D2",X"6D",X"B8",X"21",X"A0",X"B2",X"9D",X"B9",X"18",X"BA",X"20",X"B8",X"24",X"B0",X"20",X"D2",
		X"80",X"B2",X"A5",X"F4",X"3F",X"6A",X"AA",X"F6",X"F2",X"F9",X"12",X"E5",X"FA",X"03",X"80",X"E6",
		X"E5",X"B8",X"24",X"F0",X"03",X"20",X"A0",X"A4",X"E5",X"84",X"3C",X"B8",X"21",X"A0",X"B2",X"B9",
		X"B9",X"18",X"BA",X"40",X"B8",X"24",X"B0",X"00",X"B2",X"C1",X"F4",X"58",X"F6",X"F2",X"F9",X"03",
		X"F2",X"F6",X"58",X"B8",X"24",X"F0",X"03",X"10",X"A0",X"A4",X"58",X"B8",X"21",X"A0",X"B9",X"28",
		X"BA",X"60",X"B8",X"24",X"B0",X"00",X"F4",X"69",X"F9",X"53",X"03",X"C6",X"69",X"12",X"64",X"F4",
		X"31",X"6A",X"A4",X"E6",X"F4",X"37",X"6A",X"A4",X"E6",X"F4",X"69",X"A4",X"E5",X"37",X"B2",X"74",
		X"C5",X"F5",X"04",X"05",X"B8",X"21",X"B0",X"C0",X"B9",X"28",X"BA",X"30",X"B8",X"24",X"B0",X"00",
		X"F9",X"03",X"E0",X"96",X"89",X"BA",X"48",X"A4",X"96",X"F6",X"E5",X"F9",X"53",X"03",X"96",X"96",
		X"B8",X"24",X"F0",X"03",X"20",X"A0",X"F9",X"12",X"E5",X"F4",X"69",X"A4",X"E5",X"B9",X"80",X"BA",
		X"E0",X"B8",X"24",X"B0",X"00",X"F9",X"12",X"AC",X"F4",X"69",X"E6",X"F2",X"F9",X"03",X"F0",X"F6",
		X"E5",X"B8",X"24",X"F0",X"03",X"10",X"A0",X"A4",X"E5",X"B9",X"B0",X"BA",X"80",X"B8",X"24",X"B0",
		X"00",X"F9",X"47",X"53",X"0F",X"03",X"FA",X"E6",X"D0",X"C6",X"E1",X"A8",X"E8",X"E1",X"A4",X"D0",
		X"F4",X"64",X"F6",X"F2",X"F9",X"03",X"F0",X"F6",X"58",X"B8",X"24",X"F0",X"03",X"10",X"A0",X"A4",
		X"58",X"F4",X"69",X"A4",X"58",X"FA",X"47",X"E7",X"AE",X"53",X"1F",X"AF",X"FE",X"53",X"E0",X"AE",
		X"E9",X"29",X"B8",X"21",X"B0",X"00",X"84",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2D",X"24",X"2F",X"D3",X"32",X"AB",X"35",X"AF",X"38",X"E0",X"00",X"00",X"3C",X"42",X"3F",X"D7",
		X"43",X"A3",X"47",X"A9",X"4B",X"EB",X"50",X"6F",X"55",X"38",X"F0",X"96",X"20",X"18",X"10",X"C8",
		X"18",X"F0",X"37",X"17",X"03",X"0B",X"C6",X"2A",X"C4",X"30",X"C8",X"F0",X"10",X"F5",X"64",X"00",
		X"C8",X"F0",X"10",X"F5",X"84",X"5A",X"D4",X"1A",X"A9",X"F2",X"41",X"C6",X"5E",X"AA",X"D4",X"1A",
		X"A9",X"F9",X"53",X"0F",X"E7",X"A8",X"A3",X"AF",X"F8",X"17",X"A3",X"AE",X"F9",X"53",X"30",X"47",
		X"A8",X"FF",X"97",X"67",X"AF",X"FE",X"67",X"AE",X"18",X"F8",X"03",X"FB",X"96",X"51",X"83",X"F4",
		X"70",X"D4",X"9F",X"D4",X"AA",X"27",X"62",X"F5",X"34",X"00",X"E5",X"80",X"53",X"0F",X"03",X"F6",
		X"96",X"74",X"84",X"10",X"B8",X"23",X"F0",X"03",X"08",X"E6",X"80",X"27",X"AE",X"AF",X"C4",X"81",
		X"A0",X"E9",X"88",X"D4",X"9F",X"F8",X"C6",X"DC",X"D5",X"B8",X"24",X"F0",X"03",X"08",X"E6",X"95",
		X"27",X"AE",X"AF",X"C4",X"96",X"A0",X"E9",X"67",X"D4",X"AA",X"F8",X"C6",X"DC",X"C4",X"67",X"B8",
		X"23",X"B0",X"00",X"C5",X"B8",X"30",X"D4",X"36",X"C4",X"B3",X"B8",X"24",X"B0",X"00",X"D5",X"B8",
		X"32",X"D4",X"36",X"FA",X"29",X"A8",X"83",X"F4",X"70",X"85",X"A5",X"D4",X"A3",X"B8",X"23",X"B0",
		X"20",X"D4",X"AE",X"B8",X"24",X"B0",X"20",X"27",X"62",X"F5",X"34",X"00",X"E5",X"E9",X"D4",X"D4",
		X"9F",X"F8",X"C6",X"DC",X"D5",X"E9",X"C9",X"D4",X"AA",X"F8",X"96",X"C9",X"27",X"D5",X"AE",X"AF",
		X"C5",X"AE",X"AF",X"24",X"13",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"47",X"E7",X"AE",X"53",X"1F",X"AF",X"FE",X"53",X"E0",X"AE",X"84",X"10",X"FA",X"77",X"77",
		X"AE",X"53",X"3F",X"AF",X"FE",X"53",X"C0",X"AE",X"84",X"10",X"FA",X"77",X"AE",X"53",X"7F",X"AF",
		X"FE",X"53",X"80",X"AE",X"84",X"10",X"FE",X"6F",X"E6",X"2B",X"1F",X"6F",X"E6",X"2F",X"1F",X"AE",
		X"83",X"FA",X"97",X"67",X"C6",X"56",X"83",X"FA",X"77",X"77",X"53",X"3F",X"C6",X"56",X"83",X"FA",
		X"47",X"E7",X"53",X"1F",X"C6",X"56",X"83",X"FA",X"47",X"53",X"0F",X"C6",X"56",X"83",X"FA",X"47",
		X"77",X"53",X"07",X"C6",X"56",X"83",X"17",X"83",X"F4",X"47",X"6A",X"AA",X"83",X"F4",X"47",X"37",
		X"17",X"6A",X"AA",X"83",X"F4",X"4E",X"6A",X"AA",X"83",X"F4",X"4E",X"37",X"17",X"6A",X"AA",X"83",
		X"53",X"07",X"E7",X"E7",X"43",X"F0",X"A8",X"B9",X"30",X"A3",X"A1",X"18",X"19",X"F8",X"A3",X"A1",
		X"18",X"19",X"F8",X"A3",X"A1",X"18",X"19",X"F8",X"A3",X"A1",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2A",X"0B",X"35",X"0B",X"43",X"0B",X"60",X"0B",X"78",X"0B",X"9E",X"0B",X"EB",X"0B",X"F7",X"0B",
		X"9A",X"DF",X"E5",X"34",X"01",X"15",X"B9",X"08",X"BA",X"18",X"B8",X"23",X"B0",X"00",X"18",X"B0",
		X"00",X"14",X"2A",X"B9",X"80",X"BA",X"18",X"B8",X"23",X"B0",X"00",X"18",X"B0",X"00",X"14",X"2A",
		X"D5",X"BE",X"00",X"BF",X"00",X"C5",X"05",X"E5",X"34",X"13",X"FA",X"47",X"E7",X"AE",X"53",X"1F",
		X"AF",X"FE",X"53",X"E0",X"AE",X"D5",X"AE",X"C5",X"FF",X"D5",X"AF",X"E5",X"F4",X"26",X"F4",X"26",
		X"F5",X"C5",X"14",X"5E",X"E5",X"F4",X"4E",X"F5",X"37",X"17",X"6A",X"AA",X"E6",X"20",X"B8",X"23",
		X"F0",X"03",X"10",X"A0",X"18",X"F0",X"03",X"10",X"A0",X"F6",X"20",X"E9",X"2A",X"83",X"C5",X"16",
		X"61",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"E6",X"70",X"B8",X"23",X"F0",X"53",X"E0",X"AB",X"FD",
		X"77",X"77",X"53",X"3F",X"B2",X"79",X"27",X"04",X"7B",X"FB",X"E3",X"A8",X"D5",X"FC",X"6E",X"AC",
		X"FD",X"7F",X"AD",X"E6",X"8C",X"B8",X"24",X"F0",X"53",X"E0",X"AB",X"FD",X"77",X"77",X"53",X"3F",
		X"B2",X"95",X"27",X"04",X"97",X"FB",X"E3",X"C5",X"68",X"90",X"16",X"9E",X"04",X"61",X"83",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"15",X"C5",X"16",X"04",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"F6",X"13",X"8A",X"20",X"00",X"9A",
		X"DF",X"24",X"1A",X"B8",X"23",X"F0",X"53",X"E0",X"AB",X"FD",X"77",X"77",X"53",X"3F",X"96",X"28",
		X"8A",X"20",X"A3",X"9A",X"DF",X"27",X"24",X"34",X"B2",X"2E",X"00",X"00",X"24",X"32",X"37",X"17",
		X"53",X"1F",X"6B",X"E3",X"A8",X"D5",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"F6",X"45",X"8A",X"20",
		X"00",X"9A",X"DF",X"24",X"4C",X"B8",X"24",X"F0",X"53",X"E0",X"AB",X"FD",X"77",X"77",X"53",X"3F",
		X"96",X"5A",X"8A",X"20",X"A3",X"9A",X"DF",X"27",X"24",X"66",X"B2",X"60",X"00",X"00",X"24",X"64",
		X"37",X"17",X"53",X"1F",X"6B",X"E3",X"C5",X"68",X"90",X"16",X"6D",X"24",X"04",X"05",X"83",X"15",
		X"C5",X"16",X"73",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"E6",X"D8",X"B6",X"DA",X"B8",X"22",X"F0",
		X"18",X"60",X"A0",X"53",X"E0",X"AB",X"FD",X"77",X"77",X"53",X"3F",X"96",X"95",X"8A",X"20",X"A3",
		X"9A",X"DF",X"27",X"24",X"A1",X"B2",X"9B",X"00",X"00",X"24",X"9F",X"37",X"17",X"53",X"1F",X"6B",
		X"E3",X"A8",X"D5",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"F6",X"AD",X"24",X"B4",X"B8",X"24",X"F0",
		X"53",X"E0",X"AB",X"FD",X"77",X"77",X"53",X"3F",X"96",X"C2",X"8A",X"20",X"A3",X"9A",X"DF",X"27",
		X"24",X"CE",X"B2",X"C8",X"00",X"00",X"24",X"CC",X"37",X"17",X"53",X"1F",X"6B",X"E3",X"C5",X"68",
		X"90",X"16",X"D5",X"24",X"73",X"05",X"E5",X"83",X"24",X"87",X"B5",X"76",X"E6",X"FE",X"97",X"F7",
		X"AE",X"FF",X"F7",X"AF",X"24",X"7D",X"FF",X"97",X"67",X"AF",X"FE",X"67",X"AE",X"24",X"7D",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"15",X"C5",X"16",X"04",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"E6",X"66",X"B6",X"68",X"B8",X"23",
		X"F0",X"53",X"E0",X"AB",X"FD",X"77",X"77",X"53",X"3F",X"96",X"23",X"8A",X"20",X"A3",X"9A",X"DF",
		X"27",X"44",X"2F",X"B2",X"29",X"00",X"00",X"44",X"2D",X"37",X"17",X"53",X"1F",X"6B",X"E3",X"A8",
		X"D5",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"F6",X"3B",X"44",X"42",X"B8",X"24",X"F0",X"53",X"E0",
		X"AB",X"FD",X"77",X"77",X"53",X"3F",X"96",X"50",X"8A",X"20",X"A3",X"9A",X"DF",X"27",X"44",X"5C",
		X"B2",X"56",X"00",X"00",X"44",X"5A",X"37",X"17",X"53",X"1F",X"6B",X"E3",X"C5",X"68",X"90",X"16",
		X"63",X"44",X"04",X"05",X"E5",X"83",X"44",X"15",X"76",X"74",X"FE",X"97",X"F7",X"AE",X"FF",X"F7",
		X"AF",X"85",X"44",X"0E",X"FF",X"97",X"67",X"AF",X"FE",X"67",X"AE",X"A5",X"44",X"0E",X"C5",X"16",
		X"81",X"FF",X"96",X"85",X"1F",X"FE",X"6C",X"AC",X"FF",X"5A",X"7D",X"AD",X"B6",X"90",X"E6",X"A7",
		X"FF",X"77",X"AF",X"FE",X"67",X"AE",X"FF",X"F6",X"A1",X"12",X"A3",X"53",X"7F",X"AF",X"FD",X"44",
		X"A7",X"12",X"9B",X"43",X"80",X"AF",X"FD",X"77",X"77",X"53",X"3F",X"96",X"B3",X"A3",X"A3",X"A3",
		X"27",X"44",X"BF",X"B2",X"B9",X"00",X"00",X"44",X"BD",X"37",X"17",X"53",X"1F",X"6B",X"E3",X"A8",
		X"D5",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"F6",X"CB",X"44",X"D2",X"B8",X"24",X"F0",X"53",X"E0",
		X"AB",X"FD",X"77",X"77",X"53",X"3F",X"96",X"DE",X"A3",X"A3",X"A3",X"27",X"44",X"EA",X"B2",X"E4",
		X"00",X"00",X"44",X"E8",X"37",X"17",X"53",X"1F",X"6B",X"E3",X"C5",X"68",X"90",X"16",X"F1",X"44",
		X"85",X"E5",X"83",X"44",X"A7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A3",X"E5",X"83",X"0C",X"A0",X"A0",X"A4",X"18",X"A8",X"0C",X"A4",X"06",X"A8",X"A9",X"AA",X"AB",
		X"AC",X"0C",X"B0",X"00",X"08",X"BC",X"B7",X"BC",X"B7",X"BC",X"B7",X"BC",X"B7",X"BC",X"B7",X"BC",
		X"B7",X"BC",X"B7",X"BC",X"10",X"B7",X"00",X"08",X"BA",X"00",X"0A",X"AC",X"AA",X"14",X"A8",X"A8",
		X"A8",X"AC",X"50",X"B0",X"00",X"14",X"86",X"98",X"92",X"8C",X"88",X"0A",X"80",X"82",X"84",X"88",
		X"28",X"90",X"00",X"2A",X"B0",X"0E",X"A8",X"2A",X"B0",X"0E",X"A8",X"B0",X"A8",X"B0",X"B4",X"38",
		X"B8",X"2A",X"B6",X"0E",X"B2",X"2A",X"B6",X"0E",X"B2",X"B6",X"B2",X"AC",X"B2",X"38",X"A8",X"00",
		X"2A",X"90",X"0E",X"88",X"2A",X"90",X"0E",X"88",X"70",X"90",X"2A",X"92",X"0E",X"8C",X"2A",X"92",
		X"0E",X"8C",X"1C",X"92",X"8C",X"38",X"88",X"00",X"03",X"AC",X"15",X"B0",X"18",X"AC",X"0C",X"AA",
		X"24",X"A8",X"03",X"A9",X"15",X"AA",X"18",X"A8",X"0C",X"A6",X"24",X"A4",X"18",X"A2",X"A6",X"0C",
		X"AA",X"24",X"B0",X"03",X"B1",X"2D",X"B2",X"03",X"B3",X"2D",X"B4",X"60",X"B0",X"00",X"18",X"A0",
		X"98",X"94",X"90",X"98",X"90",X"8A",X"86",X"92",X"8A",X"86",X"82",X"06",X"98",X"96",X"98",X"96",
		X"18",X"98",X"06",X"94",X"92",X"94",X"92",X"18",X"94",X"06",X"90",X"8C",X"90",X"8C",X"90",X"8C",
		X"90",X"8C",X"30",X"90",X"00",X"0E",X"AA",X"A8",X"AA",X"AC",X"B0",X"B2",X"B4",X"B2",X"B0",X"AC",
		X"AA",X"A8",X"1C",X"AA",X"0E",X"B6",X"B4",X"AC",X"B2",X"54",X"B0",X"00",X"1C",X"96",X"90",X"8A",
		X"90",X"88",X"84",X"96",X"90",X"88",X"1C",X"90",X"38",X"90",X"00",X"0A",X"A8",X"AC",X"B2",X"B6",
		X"B8",X"B6",X"B2",X"AC",X"28",X"A8",X"00",X"28",X"98",X"92",X"88",X"00",X"10",X"90",X"20",X"90",
		X"10",X"88",X"90",X"80",X"80",X"80",X"10",X"90",X"20",X"90",X"10",X"90",X"08",X"98",X"10",X"96",
		X"18",X"94",X"10",X"92",X"10",X"90",X"20",X"90",X"10",X"88",X"90",X"80",X"80",X"80",X"10",X"90",
		X"20",X"90",X"10",X"90",X"08",X"98",X"10",X"96",X"18",X"94",X"10",X"92",X"10",X"94",X"20",X"94",
		X"10",X"8C",X"94",X"84",X"84",X"84",X"10",X"94",X"20",X"94",X"10",X"94",X"08",X"9A",X"10",X"98",
		X"18",X"96",X"10",X"94",X"00",X"1C",X"A0",X"0E",X"A4",X"1C",X"9B",X"0E",X"A2",X"1C",X"A0",X"0E",
		X"A0",X"A4",X"A2",X"1C",X"99",X"0E",X"A4",X"1C",X"A2",X"00",X"A3",X"E5",X"83",X"A3",X"E5",X"83",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
