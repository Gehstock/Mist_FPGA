library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity loc_prg_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of loc_prg_rom is
	type rom is array(0 to  20479) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"00",X"32",X"81",X"A1",X"C3",X"A5",X"02",X"E1",X"87",X"E7",X"5E",X"23",X"56",X"EB",X"E9",
		X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",X"35",X"34",X"C8",X"35",X"C9",X"FF",X"FF",X"FF",
		X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",X"19",X"7C",X"E6",X"03",X"F6",X"80",X"67",X"C9",
		X"EB",X"4E",X"23",X"46",X"EB",X"09",X"C9",X"FF",X"3A",X"C0",X"98",X"26",X"98",X"6F",X"7E",X"B7",
		X"C0",X"72",X"2C",X"73",X"2C",X"7D",X"20",X"02",X"3E",X"C2",X"32",X"C0",X"98",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",X"E1",X"D1",X"C1",X"3E",
		X"01",X"32",X"81",X"A1",X"F1",X"C9",X"F5",X"AF",X"32",X"81",X"A1",X"C5",X"D5",X"E5",X"08",X"D9",
		X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"58",X"01",X"CD",X"2E",X"01",X"21",X"1E",
		X"98",X"11",X"1F",X"98",X"ED",X"A8",X"3A",X"00",X"A1",X"2F",X"12",X"1D",X"2D",X"ED",X"A8",X"3A",
		X"80",X"A0",X"2F",X"12",X"1D",X"2D",X"ED",X"A8",X"ED",X"A8",X"ED",X"A8",X"3A",X"00",X"A0",X"2F",
		X"12",X"32",X"80",X"A0",X"21",X"07",X"98",X"35",X"CD",X"C0",X"1F",X"CD",X"BE",X"00",X"21",X"52",
		X"00",X"E5",X"3A",X"00",X"98",X"CF",X"18",X"02",X"4F",X"09",X"04",X"21",X"92",X"15",X"21",X"10",
		X"98",X"7E",X"B7",X"28",X"05",X"35",X"07",X"32",X"84",X"A1",X"2E",X"14",X"7E",X"B7",X"28",X"05",
		X"35",X"07",X"32",X"86",X"A1",X"21",X"18",X"98",X"7E",X"2C",X"B6",X"2C",X"2F",X"A6",X"E6",X"C4",
		X"C8",X"47",X"E6",X"84",X"28",X"30",X"B8",X"28",X"04",X"01",X"16",X"01",X"C5",X"07",X"30",X"08",
		X"3E",X"82",X"32",X"10",X"98",X"CD",X"8C",X"20",X"3A",X"15",X"98",X"47",X"21",X"11",X"98",X"7E",
		X"C6",X"10",X"B8",X"77",X"D8",X"36",X"00",X"78",X"E6",X"0F",X"21",X"12",X"98",X"86",X"FE",X"63",
		X"38",X"02",X"3E",X"63",X"77",X"C9",X"CD",X"8C",X"20",X"3E",X"86",X"32",X"14",X"98",X"3A",X"16",
		X"98",X"47",X"21",X"13",X"98",X"7E",X"C6",X"10",X"B8",X"77",X"D8",X"C3",X"05",X"01",X"21",X"40",
		X"98",X"11",X"14",X"80",X"AF",X"CD",X"3E",X"01",X"21",X"42",X"98",X"11",X"14",X"88",X"01",X"0C",
		X"00",X"ED",X"A0",X"ED",X"A0",X"2C",X"2C",X"B9",X"38",X"F7",X"0E",X"04",X"1E",X"00",X"ED",X"A0",
		X"ED",X"A0",X"2C",X"2C",X"B9",X"38",X"F7",X"C9",X"AF",X"21",X"20",X"88",X"01",X"01",X"04",X"D7",
		X"21",X"60",X"98",X"11",X"34",X"80",X"CD",X"72",X"01",X"11",X"04",X"A0",X"CD",X"72",X"01",X"11",
		X"34",X"88",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",
		X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"11",X"04",X"00",X"19",X"C9",X"21",
		X"0E",X"99",X"34",X"5E",X"16",X"4E",X"1A",X"2C",X"86",X"77",X"C9",X"26",X"98",X"3A",X"C1",X"98",
		X"6F",X"7E",X"87",X"20",X"0F",X"26",X"9C",X"3A",X"21",X"9C",X"6F",X"7E",X"87",X"20",X"22",X"CD",
		X"C0",X"03",X"18",X"E7",X"4F",X"06",X"00",X"70",X"23",X"5E",X"2C",X"7D",X"20",X"02",X"3E",X"C2",
		X"32",X"C1",X"98",X"7B",X"21",X"EF",X"01",X"09",X"5E",X"23",X"56",X"21",X"9B",X"01",X"E5",X"EB",
		X"E9",X"4F",X"06",X"00",X"70",X"23",X"5E",X"2C",X"7D",X"FE",X"20",X"38",X"01",X"AF",X"32",X"21",
		X"9C",X"7B",X"21",X"EF",X"01",X"09",X"5E",X"23",X"56",X"21",X"9B",X"01",X"E5",X"EB",X"E9",X"FF",
		X"03",X"2C",X"03",X"84",X"04",X"DB",X"04",X"A6",X"08",X"E9",X"08",X"03",X"09",X"1E",X"09",X"00",
		X"04",X"3A",X"20",X"9C",X"6F",X"26",X"9C",X"7E",X"B7",X"C0",X"72",X"2C",X"73",X"2C",X"7D",X"FE",
		X"20",X"38",X"01",X"AF",X"32",X"20",X"9C",X"C9",X"3A",X"80",X"A1",X"47",X"E6",X"0F",X"20",X"01",
		X"47",X"4F",X"A8",X"0F",X"0F",X"0F",X"0F",X"21",X"21",X"09",X"E7",X"46",X"79",X"21",X"21",X"09",
		X"E7",X"4E",X"ED",X"43",X"15",X"98",X"3A",X"00",X"A1",X"EE",X"33",X"47",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"03",X"C6",X"03",X"FE",X"06",X"20",X"02",X"3E",X"FF",X"32",X"0C",X"98",X"78",X"21",X"00",
		X"00",X"54",X"5C",X"44",X"4C",X"0F",X"CB",X"14",X"0F",X"CB",X"11",X"0F",X"CB",X"12",X"0F",X"CB",
		X"10",X"3A",X"80",X"A1",X"E6",X"0F",X"20",X"01",X"2C",X"ED",X"53",X"BC",X"98",X"22",X"BE",X"98",
		X"21",X"0B",X"98",X"70",X"2E",X"0F",X"71",X"3E",X"0A",X"06",X"00",X"21",X"31",X"09",X"11",X"00",
		X"9F",X"0E",X"03",X"ED",X"B0",X"EB",X"01",X"3E",X"09",X"71",X"2C",X"10",X"FC",X"EB",X"3D",X"20",
		X"F0",X"21",X"31",X"09",X"11",X"C6",X"99",X"0E",X"03",X"ED",X"B0",X"3E",X"01",X"32",X"0D",X"98",
		X"21",X"00",X"98",X"34",X"C9",X"3A",X"00",X"50",X"FE",X"55",X"CA",X"01",X"50",X"21",X"00",X"98",
		X"11",X"01",X"98",X"01",X"FF",X"07",X"36",X"00",X"ED",X"B0",X"32",X"80",X"A0",X"31",X"00",X"A0",
		X"21",X"C2",X"C2",X"22",X"C0",X"98",X"21",X"D0",X"99",X"01",X"01",X"30",X"3E",X"FF",X"D7",X"21",
		X"D0",X"D0",X"22",X"CD",X"99",X"32",X"80",X"A0",X"AF",X"32",X"84",X"A1",X"32",X"86",X"A1",X"32",
		X"87",X"A1",X"3C",X"32",X"83",X"A1",X"CD",X"E5",X"1F",X"3E",X"0B",X"21",X"00",X"80",X"01",X"04",
		X"00",X"D7",X"32",X"80",X"A0",X"01",X"04",X"00",X"D7",X"3E",X"80",X"32",X"80",X"A0",X"01",X"04",
		X"00",X"D7",X"3E",X"80",X"32",X"80",X"A0",X"01",X"04",X"00",X"D7",X"CD",X"D1",X"1C",X"32",X"80",
		X"A0",X"CD",X"22",X"03",X"CD",X"EB",X"1F",X"CD",X"22",X"03",X"3E",X"01",X"32",X"81",X"A1",X"C3",
		X"9B",X"01",X"0B",X"32",X"80",X"A0",X"78",X"B1",X"20",X"F8",X"37",X"C9",X"47",X"3A",X"08",X"98",
		X"B7",X"C8",X"3A",X"09",X"98",X"B7",X"20",X"63",X"11",X"00",X"02",X"CD",X"01",X"02",X"11",X"C0",
		X"99",X"78",X"87",X"20",X"06",X"21",X"C9",X"99",X"C3",X"50",X"03",X"80",X"21",X"48",X"04",X"E7",
		X"B7",X"06",X"03",X"1A",X"8E",X"27",X"12",X"1C",X"23",X"10",X"F8",X"47",X"30",X"04",X"AF",X"32",
		X"3F",X"99",X"3A",X"01",X"99",X"B8",X"DC",X"A7",X"03",X"3A",X"3F",X"99",X"B7",X"20",X"1A",X"06",
		X"03",X"21",X"C8",X"99",X"1D",X"1A",X"BE",X"D8",X"20",X"04",X"2D",X"10",X"F7",X"C9",X"3E",X"01",
		X"32",X"3F",X"99",X"3E",X"04",X"90",X"EB",X"E7",X"EB",X"EB",X"2D",X"11",X"C8",X"99",X"ED",X"A8",
		X"ED",X"A8",X"ED",X"A8",X"11",X"02",X"02",X"CD",X"01",X"02",X"C9",X"11",X"01",X"02",X"CD",X"01",
		X"02",X"11",X"C3",X"99",X"C3",X"41",X"03",X"D5",X"C6",X"07",X"27",X"30",X"02",X"3E",X"99",X"21",
		X"01",X"99",X"77",X"2D",X"34",X"11",X"00",X"05",X"CD",X"01",X"02",X"CD",X"73",X"20",X"D1",X"C9",
		X"CD",X"59",X"2A",X"CD",X"87",X"2C",X"CD",X"2F",X"2E",X"CD",X"33",X"2B",X"21",X"19",X"98",X"CB",
		X"46",X"C8",X"C9",X"0E",X"30",X"1A",X"91",X"77",X"13",X"3E",X"20",X"E7",X"10",X"F7",X"C9",X"81",
		X"8C",X"9A",X"81",X"8C",X"8E",X"8E",X"8E",X"8E",X"90",X"90",X"90",X"90",X"90",X"90",X"91",X"91",
		X"91",X"91",X"91",X"91",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"93",X"93",X"93",X"C9",
		X"3C",X"28",X"06",X"21",X"DF",X"03",X"CD",X"C4",X"11",X"01",X"10",X"0B",X"79",X"C5",X"CD",X"DB",
		X"04",X"C1",X"0C",X"10",X"F7",X"21",X"98",X"85",X"DD",X"21",X"02",X"9F",X"06",X"0A",X"C5",X"11",
		X"20",X"00",X"CD",X"A2",X"04",X"11",X"60",X"00",X"19",X"DD",X"E5",X"D1",X"13",X"13",X"13",X"13",
		X"06",X"03",X"CD",X"D3",X"03",X"11",X"0F",X"00",X"DD",X"19",X"11",X"7E",X"FE",X"19",X"C1",X"10",
		X"DD",X"11",X"0F",X"03",X"CD",X"01",X"02",X"C9",X"00",X"00",X"00",X"10",X"00",X"00",X"20",X"00",
		X"00",X"30",X"00",X"00",X"40",X"00",X"00",X"50",X"00",X"00",X"60",X"00",X"00",X"70",X"00",X"00",
		X"80",X"00",X"00",X"90",X"00",X"00",X"00",X"01",X"00",X"10",X"01",X"00",X"20",X"01",X"00",X"30",
		X"01",X"00",X"40",X"01",X"00",X"50",X"01",X"00",X"00",X"02",X"00",X"00",X"04",X"00",X"00",X"10",
		X"00",X"00",X"50",X"00",X"DD",X"21",X"C2",X"99",X"21",X"85",X"80",X"A7",X"28",X"11",X"DD",X"21",
		X"C5",X"99",X"21",X"C5",X"82",X"3D",X"28",X"07",X"DD",X"21",X"C8",X"99",X"21",X"A5",X"81",X"11",
		X"20",X"00",X"06",X"03",X"DD",X"7E",X"00",X"4F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"20",X"1F",
		X"36",X"10",X"19",X"79",X"E6",X"0F",X"20",X"1C",X"36",X"10",X"19",X"DD",X"2B",X"10",X"E5",X"AF",
		X"ED",X"52",X"77",X"19",X"C9",X"DD",X"7E",X"00",X"4F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"77",
		X"19",X"79",X"E6",X"0F",X"77",X"19",X"DD",X"2B",X"10",X"EB",X"C9",X"47",X"E6",X"3F",X"FE",X"03",
		X"20",X"0A",X"78",X"E6",X"C0",X"F6",X"31",X"C5",X"CD",X"ED",X"04",X"C1",X"78",X"87",X"F5",X"21",
		X"2B",X"05",X"E6",X"7F",X"85",X"6F",X"30",X"01",X"24",X"F1",X"5E",X"23",X"56",X"EB",X"5E",X"23",
		X"56",X"23",X"EB",X"01",X"20",X"00",X"38",X"15",X"1A",X"FE",X"2E",X"28",X"0B",X"FE",X"2F",X"C8",
		X"D6",X"30",X"77",X"13",X"09",X"18",X"F1",X"37",X"EB",X"23",X"C3",X"FE",X"04",X"1A",X"FE",X"2E",
		X"28",X"F5",X"FE",X"2F",X"C8",X"36",X"10",X"13",X"09",X"18",X"F2",X"9B",X"05",X"A2",X"05",X"A9",
		X"05",X"B0",X"05",X"DC",X"05",X"F3",X"05",X"09",X"06",X"12",X"06",X"2A",X"06",X"3C",X"06",X"51",
		X"06",X"5B",X"06",X"68",X"06",X"75",X"06",X"81",X"06",X"92",X"06",X"A3",X"06",X"B9",X"06",X"BF",
		X"06",X"C5",X"06",X"CB",X"06",X"D1",X"06",X"D7",X"06",X"DD",X"06",X"E3",X"06",X"E9",X"06",X"EF",
		X"06",X"F6",X"06",X"00",X"07",X"07",X"07",X"07",X"07",X"37",X"07",X"37",X"07",X"66",X"07",X"73",
		X"07",X"81",X"07",X"90",X"07",X"98",X"07",X"A8",X"07",X"B4",X"07",X"CC",X"07",X"E6",X"07",X"F7",
		X"07",X"FD",X"07",X"0F",X"08",X"19",X"08",X"26",X"08",X"33",X"08",X"43",X"08",X"51",X"08",X"66",
		X"08",X"A3",X"08",X"A3",X"08",X"A3",X"08",X"A3",X"08",X"A3",X"08",X"C6",X"81",X"48",X"49",X"47",
		X"48",X"2F",X"A6",X"80",X"31",X"5B",X"55",X"50",X"2F",X"E6",X"82",X"32",X"5B",X"55",X"50",X"2F",
		X"D9",X"84",X"3F",X"3F",X"40",X"40",X"4C",X"4F",X"43",X"4F",X"5B",X"4D",X"4F",X"54",X"49",X"4F",
		X"4E",X"40",X"40",X"3F",X"3F",X"2F",X"D9",X"84",X"5B",X"40",X"47",X"55",X"54",X"54",X"41",X"4E",
		X"47",X"40",X"47",X"4F",X"54",X"54",X"4F",X"4E",X"47",X"40",X"5B",X"2F",X"B2",X"84",X"50",X"4C",
		X"45",X"41",X"53",X"45",X"40",X"44",X"45",X"50",X"4F",X"53",X"49",X"54",X"40",X"43",X"4F",X"49",
		X"4E",X"53",X"2F",X"CC",X"84",X"48",X"41",X"56",X"45",X"40",X"41",X"40",X"4E",X"49",X"43",X"45",
		X"40",X"54",X"52",X"49",X"50",X"40",X"3C",X"3C",X"2F",X"95",X"85",X"50",X"4C",X"45",X"41",X"53",
		X"45",X"2F",X"A4",X"84",X"50",X"55",X"53",X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"40",X"46",X"4F",X"52",X"2F",X"02",X"85",X"4F",X"4E",X"45",X"40",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"4C",X"59",X"2F",X"C2",X"84",X"4F",X"4E",
		X"45",X"40",X"4F",X"52",X"40",X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",
		X"2F",X"84",X"82",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"2F",X"75",X"85",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"2F",X"75",X"85",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"40",X"54",X"57",X"4F",X"2F",X"71",X"85",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",
		X"2F",X"22",X"85",X"3A",X"40",X"43",X"45",X"4E",X"54",X"55",X"52",X"49",X"40",X"31",X"39",X"38",
		X"32",X"2F",X"20",X"85",X"3A",X"40",X"43",X"45",X"4E",X"54",X"55",X"52",X"49",X"40",X"31",X"39",
		X"38",X"32",X"2F",X"DA",X"84",X"5B",X"40",X"40",X"53",X"43",X"4F",X"52",X"45",X"40",X"52",X"41",
		X"4E",X"4B",X"49",X"4E",X"47",X"40",X"40",X"5B",X"2F",X"B8",X"84",X"31",X"53",X"54",X"2F",X"B6",
		X"84",X"32",X"4E",X"44",X"2F",X"B4",X"84",X"33",X"52",X"44",X"2F",X"B2",X"84",X"34",X"54",X"48",
		X"2F",X"B0",X"84",X"35",X"54",X"48",X"2F",X"AE",X"84",X"36",X"54",X"48",X"2F",X"AC",X"84",X"37",
		X"54",X"48",X"2F",X"AA",X"84",X"38",X"54",X"48",X"2F",X"A8",X"84",X"39",X"54",X"48",X"2F",X"86",
		X"84",X"31",X"30",X"54",X"48",X"2F",X"A7",X"85",X"53",X"54",X"41",X"54",X"49",X"4F",X"4E",X"2F",
		X"A8",X"84",X"31",X"35",X"30",X"30",X"2F",X"D7",X"84",X"3F",X"3F",X"40",X"40",X"4C",X"4F",X"43",
		X"4F",X"5B",X"4D",X"4F",X"54",X"49",X"4F",X"4E",X"40",X"40",X"3F",X"3F",X"2F",X"78",X"85",X"12",
		X"10",X"16",X"14",X"1A",X"18",X"1E",X"1C",X"22",X"20",X"2F",X"77",X"85",X"13",X"11",X"17",X"15",
		X"1B",X"19",X"1F",X"1D",X"23",X"21",X"2F",X"00",X"85",X"4C",X"49",X"43",X"45",X"4E",X"53",X"45",
		X"44",X"40",X"42",X"59",X"40",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"2F",X"B6",X"85",X"12",X"10",
		X"26",X"24",X"1A",X"2A",X"28",X"1C",X"22",X"20",X"2F",X"B5",X"85",X"13",X"11",X"27",X"25",X"1B",
		X"2B",X"29",X"1D",X"23",X"21",X"2F",X"67",X"85",X"42",X"4F",X"4E",X"55",X"53",X"40",X"4C",X"49",
		X"4E",X"45",X"2F",X"67",X"85",X"43",X"52",X"41",X"5A",X"59",X"40",X"54",X"52",X"41",X"49",X"4E",
		X"2F",X"47",X"85",X"4C",X"4F",X"4F",X"50",X"40",X"53",X"57",X"45",X"45",X"50",X"45",X"52",X"2F",
		X"74",X"85",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"47",X"85",X"42",X"4F",X"4E",X"55",X"53",X"40",
		X"53",X"54",X"41",X"54",X"49",X"4F",X"4E",X"2F",X"84",X"82",X"46",X"52",X"45",X"45",X"40",X"50",
		X"4C",X"41",X"59",X"2F",X"D9",X"84",X"41",X"44",X"4A",X"55",X"53",X"54",X"40",X"52",X"41",X"49",
		X"4C",X"40",X"57",X"41",X"59",X"40",X"4C",X"49",X"4E",X"45",X"53",X"2F",X"B7",X"84",X"53",X"4F",
		X"40",X"41",X"53",X"40",X"54",X"4F",X"40",X"4C",X"45",X"54",X"40",X"59",X"4F",X"55",X"52",X"40",
		X"54",X"52",X"41",X"49",X"4E",X"2F",X"B5",X"84",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"40",
		X"53",X"41",X"46",X"45",X"4C",X"59",X"2F",X"CF",X"85",X"41",X"4E",X"44",X"2F",X"11",X"85",X"40",
		X"50",X"45",X"52",X"46",X"45",X"43",X"54",X"40",X"43",X"4C",X"45",X"41",X"52",X"40",X"2F",X"91",
		X"85",X"40",X"43",X"4C",X"45",X"41",X"52",X"40",X"2F",X"6E",X"85",X"40",X"35",X"30",X"30",X"30",
		X"40",X"50",X"54",X"53",X"40",X"2F",X"6E",X"85",X"40",X"31",X"30",X"30",X"30",X"40",X"50",X"54",
		X"53",X"40",X"2F",X"31",X"8D",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"C3",X"C3",X"2F",X"8E",X"8D",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"2F",X"00",X"84",
		X"2F",X"00",X"85",X"4C",X"49",X"43",X"45",X"4E",X"53",X"45",X"44",X"40",X"42",X"59",X"40",X"4B",
		X"4F",X"4E",X"41",X"4D",X"49",X"2F",X"44",X"84",X"4D",X"4F",X"56",X"45",X"40",X"54",X"48",X"45",
		X"40",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"40",X"54",X"4F",X"40",X"53",X"45",X"4C",
		X"45",X"43",X"54",X"2E",X"42",X"84",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"40",X"41",X"4E",
		X"44",X"40",X"50",X"52",X"45",X"53",X"53",X"40",X"46",X"49",X"52",X"45",X"42",X"55",X"54",X"54",
		X"4F",X"4E",X"2F",X"00",X"80",X"2F",X"3A",X"BE",X"98",X"B7",X"28",X"05",X"3E",X"26",X"C3",X"DB",
		X"04",X"3E",X"0A",X"CD",X"DB",X"04",X"3A",X"12",X"98",X"FE",X"63",X"38",X"02",X"3E",X"63",X"CD",
		X"CD",X"08",X"21",X"64",X"83",X"11",X"20",X"00",X"06",X"01",X"C3",X"A7",X"04",X"4F",X"0F",X"0F",
		X"0F",X"0F",X"E6",X"0F",X"47",X"04",X"AF",X"81",X"27",X"0E",X"00",X"C6",X"06",X"27",X"30",X"01",
		X"0C",X"10",X"F8",X"D6",X"06",X"27",X"D0",X"0D",X"C9",X"3A",X"00",X"99",X"01",X"C4",X"06",X"11",
		X"E0",X"FF",X"21",X"04",X"81",X"B8",X"38",X"05",X"71",X"19",X"10",X"F9",X"C9",X"36",X"10",X"19",
		X"10",X"F3",X"C9",X"3A",X"02",X"99",X"3C",X"01",X"C5",X"10",X"11",X"20",X"00",X"21",X"A4",X"81",
		X"B8",X"38",X"05",X"71",X"19",X"10",X"F9",X"C9",X"36",X"10",X"19",X"10",X"F3",X"C9",X"C3",X"CD",
		X"30",X"00",X"11",X"22",X"04",X"31",X"06",X"15",X"02",X"33",X"07",X"21",X"03",X"24",X"05",X"13",
		X"01",X"00",X"00",X"01",X"30",X"85",X"00",X"90",X"76",X"00",X"30",X"70",X"00",X"80",X"62",X"00",
		X"00",X"54",X"00",X"90",X"39",X"00",X"00",X"36",X"00",X"50",X"28",X"00",X"10",X"24",X"00",X"3A",
		X"BE",X"98",X"B7",X"28",X"08",X"21",X"C0",X"21",X"E5",X"11",X"26",X"03",X"FF",X"21",X"7B",X"09",
		X"E5",X"3A",X"01",X"98",X"CF",X"AF",X"15",X"8A",X"09",X"FB",X"09",X"29",X"0C",X"38",X"0D",X"43",
		X"0E",X"41",X"10",X"75",X"22",X"49",X"10",X"72",X"10",X"A6",X"10",X"3A",X"12",X"98",X"B7",X"C8",
		X"AF",X"21",X"00",X"98",X"34",X"2C",X"77",X"2C",X"77",X"C9",X"3A",X"03",X"98",X"CF",X"94",X"09",
		X"34",X"0B",X"9D",X"10",X"3A",X"07",X"98",X"0F",X"D8",X"CD",X"91",X"11",X"3A",X"2C",X"98",X"FE",
		X"20",X"D8",X"AF",X"32",X"2C",X"98",X"21",X"DB",X"09",X"CD",X"C4",X"11",X"21",X"40",X"98",X"01",
		X"01",X"50",X"D7",X"3C",X"CD",X"61",X"11",X"1E",X"2A",X"FF",X"1E",X"04",X"FF",X"1C",X"FF",X"1E",
		X"1D",X"FF",X"1C",X"FF",X"1C",X"FF",X"1C",X"FF",X"1E",X"4E",X"FF",X"3E",X"04",X"32",X"3E",X"98",
		X"CD",X"6F",X"11",X"21",X"02",X"98",X"36",X"00",X"2C",X"34",X"C9",X"81",X"8C",X"9A",X"81",X"8C",
		X"8C",X"8C",X"8C",X"95",X"95",X"95",X"95",X"90",X"90",X"91",X"91",X"91",X"91",X"91",X"91",X"91",
		X"8E",X"8E",X"8E",X"8E",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"3A",X"03",X"98",X"CF",X"15",
		X"0A",X"A7",X"0A",X"D3",X"0A",X"11",X"0B",X"47",X"0B",X"50",X"0B",X"79",X"0B",X"A1",X"0B",X"0F",
		X"0C",X"18",X"0C",X"9D",X"10",X"3A",X"07",X"98",X"0F",X"D8",X"CD",X"91",X"11",X"3A",X"2C",X"98",
		X"FE",X"20",X"D8",X"AF",X"32",X"2C",X"98",X"CD",X"61",X"11",X"CD",X"6F",X"11",X"21",X"83",X"0A",
		X"CD",X"C4",X"11",X"11",X"03",X"03",X"FF",X"1E",X"0E",X"FF",X"21",X"A3",X"0A",X"11",X"40",X"98",
		X"01",X"04",X"00",X"ED",X"B0",X"CD",X"7D",X"11",X"11",X"6E",X"85",X"21",X"1B",X"42",X"CD",X"31",
		X"11",X"21",X"BB",X"44",X"CD",X"31",X"11",X"21",X"BB",X"43",X"3E",X"02",X"CD",X"1F",X"11",X"11",
		X"6A",X"85",X"21",X"BB",X"44",X"CD",X"31",X"11",X"21",X"BB",X"44",X"CD",X"31",X"11",X"21",X"DB",
		X"43",X"3E",X"02",X"CD",X"1F",X"11",X"3E",X"80",X"32",X"21",X"98",X"21",X"02",X"98",X"36",X"02",
		X"2C",X"34",X"C9",X"81",X"8C",X"9A",X"81",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"9A",X"8C",
		X"9A",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"9A",X"9A",X"9A",X"9A",X"93",
		X"93",X"93",X"93",X"C1",X"98",X"58",X"01",X"3A",X"07",X"98",X"0F",X"D0",X"21",X"42",X"98",X"34",
		X"7E",X"FE",X"70",X"21",X"00",X"FF",X"28",X"06",X"FE",X"90",X"C0",X"21",X"80",X"FF",X"11",X"6A",
		X"86",X"19",X"EB",X"21",X"DB",X"3C",X"CD",X"31",X"11",X"21",X"02",X"98",X"35",X"C0",X"36",X"40",
		X"2C",X"34",X"C9",X"3A",X"07",X"98",X"0F",X"D0",X"3A",X"02",X"98",X"DD",X"21",X"40",X"98",X"01",
		X"90",X"88",X"FD",X"21",X"02",X"98",X"21",X"FD",X"10",X"22",X"1B",X"99",X"CD",X"AB",X"10",X"FD",
		X"35",X"00",X"C0",X"FD",X"34",X"01",X"11",X"6E",X"86",X"21",X"BB",X"42",X"3E",X"02",X"CD",X"1F",
		X"11",X"11",X"6A",X"86",X"21",X"DB",X"42",X"3E",X"02",X"CD",X"1F",X"11",X"11",X"1B",X"03",X"FF",
		X"C9",X"3A",X"02",X"98",X"C6",X"1F",X"E6",X"20",X"20",X"14",X"3E",X"20",X"21",X"48",X"04",X"E7",
		X"E5",X"DD",X"E1",X"21",X"F4",X"85",X"CD",X"9F",X"04",X"CD",X"01",X"0C",X"18",X"06",X"21",X"F4",
		X"85",X"CD",X"3C",X"0B",X"21",X"02",X"98",X"35",X"C0",X"2C",X"34",X"C9",X"11",X"20",X"00",X"01",
		X"10",X"0A",X"71",X"19",X"10",X"FC",X"C9",X"11",X"9B",X"03",X"FF",X"21",X"03",X"98",X"34",X"C9",
		X"3A",X"07",X"98",X"0F",X"D0",X"3A",X"02",X"98",X"DD",X"21",X"40",X"98",X"01",X"90",X"88",X"FD",
		X"21",X"02",X"98",X"21",X"FD",X"10",X"22",X"1B",X"99",X"CD",X"AB",X"10",X"FD",X"35",X"00",X"FD",
		X"7E",X"00",X"E6",X"3F",X"C0",X"FD",X"34",X"01",X"C9",X"3A",X"07",X"98",X"0F",X"D0",X"21",X"42",
		X"98",X"35",X"7E",X"FE",X"70",X"28",X"11",X"FE",X"6C",X"C0",X"3E",X"03",X"32",X"17",X"98",X"11",
		X"21",X"03",X"FF",X"21",X"03",X"98",X"34",X"C9",X"11",X"EE",X"85",X"21",X"DB",X"3C",X"C3",X"31",
		X"11",X"3A",X"02",X"98",X"C6",X"1F",X"E6",X"20",X"20",X"43",X"3E",X"2F",X"21",X"48",X"04",X"E7",
		X"E5",X"DD",X"E1",X"21",X"14",X"85",X"CD",X"9F",X"04",X"CD",X"01",X"0C",X"CD",X"34",X"0B",X"3A",
		X"07",X"98",X"E6",X"0F",X"C0",X"21",X"17",X"98",X"35",X"7E",X"20",X"02",X"36",X"03",X"87",X"F5",
		X"21",X"F5",X"0B",X"E7",X"5E",X"23",X"56",X"EB",X"11",X"6E",X"85",X"CD",X"43",X"11",X"F1",X"21",
		X"FB",X"0B",X"E7",X"5E",X"23",X"56",X"EB",X"11",X"6A",X"85",X"C3",X"43",X"11",X"21",X"14",X"85",
		X"CD",X"3C",X"0B",X"18",X"C7",X"FB",X"41",X"3B",X"42",X"5B",X"42",X"DB",X"3C",X"DB",X"40",X"DB",
		X"3C",X"01",X"20",X"00",X"11",X"0B",X"0C",X"09",X"C3",X"08",X"05",X"50",X"54",X"53",X"2F",X"11",
		X"A1",X"03",X"FF",X"21",X"03",X"98",X"34",X"C9",X"21",X"40",X"98",X"01",X"01",X"40",X"AF",X"D7",
		X"21",X"03",X"98",X"34",X"AF",X"32",X"17",X"98",X"C9",X"3A",X"03",X"98",X"CF",X"9A",X"0C",X"D2",
		X"0C",X"08",X"0D",X"3F",X"0C",X"45",X"0C",X"8B",X"0C",X"34",X"0B",X"18",X"0C",X"9D",X"10",X"CD",
		X"4B",X"0C",X"C3",X"A7",X"0A",X"CD",X"4B",X"0C",X"C3",X"D3",X"0A",X"3A",X"07",X"98",X"E6",X"1F",
		X"C0",X"DD",X"21",X"1F",X"99",X"DD",X"7E",X"FE",X"D6",X"10",X"27",X"DD",X"77",X"FE",X"DD",X"7E",
		X"FF",X"DE",X"00",X"27",X"DD",X"77",X"FF",X"21",X"F4",X"85",X"CD",X"9F",X"04",X"CD",X"01",X"0C",
		X"21",X"1E",X"99",X"11",X"6F",X"86",X"7E",X"CD",X"7C",X"0C",X"2D",X"7E",X"0F",X"0F",X"0F",X"0F",
		X"CD",X"84",X"0C",X"7E",X"E6",X"0F",X"C6",X"2C",X"12",X"1D",X"C9",X"CD",X"7D",X"11",X"11",X"25",
		X"03",X"FF",X"1E",X"24",X"FF",X"21",X"03",X"98",X"34",X"C9",X"3A",X"07",X"98",X"0F",X"D8",X"CD",
		X"91",X"11",X"3A",X"2C",X"98",X"FE",X"20",X"D8",X"AF",X"32",X"2C",X"98",X"CD",X"61",X"11",X"CD",
		X"6F",X"11",X"21",X"83",X"0A",X"CD",X"C4",X"11",X"11",X"03",X"03",X"FF",X"1E",X"0E",X"FF",X"21",
		X"A3",X"0A",X"11",X"40",X"98",X"01",X"04",X"00",X"ED",X"B0",X"CD",X"7D",X"11",X"21",X"03",X"98",
		X"34",X"C9",X"11",X"6E",X"85",X"21",X"BB",X"3C",X"CD",X"31",X"11",X"21",X"FB",X"40",X"CD",X"31",
		X"11",X"21",X"BB",X"43",X"3E",X"02",X"CD",X"1F",X"11",X"11",X"6A",X"85",X"21",X"BB",X"44",X"CD",
		X"31",X"11",X"21",X"7B",X"41",X"CD",X"31",X"11",X"21",X"DB",X"43",X"3E",X"02",X"CD",X"1F",X"11",
		X"21",X"02",X"98",X"36",X"02",X"2C",X"34",X"C9",X"11",X"30",X"0D",X"21",X"00",X"15",X"22",X"1D",
		X"99",X"21",X"9A",X"9A",X"22",X"6C",X"8E",X"22",X"6E",X"8E",X"EB",X"11",X"6C",X"86",X"01",X"04",
		X"00",X"ED",X"B0",X"21",X"03",X"98",X"34",X"C9",X"11",X"34",X"0D",X"21",X"40",X"00",X"18",X"DE",
		X"2C",X"2C",X"31",X"2D",X"2C",X"30",X"2C",X"2C",X"3A",X"03",X"98",X"CF",X"9A",X"0C",X"4E",X"0D",
		X"28",X"0D",X"94",X"0D",X"A6",X"0D",X"BD",X"0D",X"E1",X"0F",X"18",X"0C",X"9D",X"10",X"FD",X"21",
		X"00",X"9D",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"1F",X"01",X"11",X"6E",
		X"85",X"21",X"9B",X"44",X"CD",X"31",X"11",X"21",X"FB",X"44",X"CD",X"31",X"11",X"21",X"BB",X"43",
		X"3E",X"02",X"CD",X"1F",X"11",X"11",X"6A",X"85",X"21",X"9B",X"40",X"CD",X"31",X"11",X"21",X"1B",
		X"45",X"CD",X"31",X"11",X"21",X"DB",X"43",X"3E",X"02",X"CD",X"1F",X"11",X"21",X"02",X"98",X"36",
		X"02",X"2C",X"34",X"C9",X"CD",X"4B",X"0C",X"CD",X"C6",X"0D",X"21",X"1D",X"99",X"7E",X"2C",X"B6",
		X"C0",X"21",X"03",X"98",X"34",X"C9",X"21",X"18",X"02",X"22",X"20",X"9D",X"7C",X"32",X"47",X"98",
		X"0F",X"32",X"3F",X"9D",X"11",X"22",X"03",X"FF",X"21",X"03",X"98",X"34",X"C9",X"CD",X"09",X"0F",
		X"CD",X"C6",X"0D",X"C3",X"7A",X"0F",X"21",X"ED",X"0D",X"E5",X"DD",X"21",X"40",X"98",X"FD",X"21",
		X"00",X"9D",X"21",X"FD",X"10",X"22",X"1B",X"99",X"FD",X"7E",X"01",X"FD",X"77",X"1E",X"CF",X"B9",
		X"0F",X"C3",X"0F",X"C3",X"0F",X"A0",X"0F",X"C3",X"0F",X"C3",X"0F",X"C3",X"0F",X"FD",X"7E",X"1E",
		X"FD",X"BE",X"01",X"C8",X"FE",X"05",X"C8",X"B7",X"20",X"08",X"FD",X"36",X"1F",X"FF",X"FD",X"36",
		X"00",X"C0",X"FE",X"04",X"20",X"07",X"CD",X"0D",X"0E",X"FD",X"7E",X"1E",X"3C",X"87",X"87",X"21",
		X"27",X"0E",X"E7",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"FD",X"7E",X"1E",X"FE",X"04",
		X"C2",X"31",X"11",X"0F",X"C3",X"1F",X"11",X"EE",X"85",X"9B",X"44",X"6E",X"85",X"BB",X"3C",X"6A",
		X"85",X"9B",X"3C",X"EA",X"85",X"DB",X"40",X"6A",X"86",X"DB",X"42",X"6E",X"86",X"BB",X"42",X"EE",
		X"85",X"BB",X"3C",X"3A",X"03",X"98",X"CF",X"51",X"0E",X"CD",X"0E",X"E1",X"0F",X"18",X"0C",X"9D",
		X"10",X"3A",X"07",X"98",X"0F",X"D8",X"CD",X"91",X"11",X"3A",X"2C",X"98",X"FE",X"20",X"D8",X"AF",
		X"32",X"2C",X"98",X"CD",X"61",X"11",X"CD",X"6F",X"11",X"21",X"83",X"0A",X"CD",X"C4",X"11",X"11",
		X"03",X"03",X"FF",X"1E",X"0E",X"FF",X"21",X"C5",X"0E",X"11",X"40",X"98",X"01",X"08",X"00",X"ED",
		X"B0",X"3E",X"FF",X"32",X"1F",X"9D",X"32",X"3F",X"9D",X"ED",X"43",X"20",X"9D",X"21",X"C0",X"04",
		X"22",X"00",X"9D",X"11",X"6E",X"85",X"21",X"9B",X"44",X"CD",X"31",X"11",X"21",X"BB",X"44",X"CD",
		X"31",X"11",X"21",X"7B",X"44",X"CD",X"31",X"11",X"11",X"6A",X"85",X"21",X"FB",X"40",X"CD",X"31",
		X"11",X"21",X"BB",X"44",X"CD",X"31",X"11",X"21",X"BB",X"40",X"CD",X"31",X"11",X"21",X"02",X"98",
		X"36",X"40",X"2C",X"34",X"C9",X"E1",X"78",X"78",X"01",X"D4",X"98",X"8C",X"07",X"CD",X"1E",X"0F",
		X"3A",X"1F",X"99",X"B7",X"28",X"06",X"CD",X"43",X"0F",X"C3",X"7A",X"0F",X"3A",X"07",X"98",X"E6",
		X"04",X"21",X"00",X"00",X"28",X"03",X"2A",X"CA",X"0E",X"22",X"45",X"98",X"3A",X"42",X"98",X"FE",
		X"7C",X"D8",X"3E",X"03",X"32",X"22",X"9D",X"32",X"1F",X"99",X"3C",X"32",X"47",X"98",X"2A",X"CA",
		X"0E",X"22",X"45",X"98",X"11",X"23",X"03",X"FF",X"C9",X"3A",X"07",X"98",X"0F",X"D8",X"DD",X"21",
		X"44",X"98",X"FD",X"21",X"20",X"9D",X"21",X"ED",X"10",X"22",X"1B",X"99",X"18",X"13",X"3A",X"07",
		X"98",X"0F",X"D0",X"21",X"FD",X"10",X"22",X"1B",X"99",X"DD",X"21",X"40",X"98",X"FD",X"21",X"00",
		X"9D",X"FD",X"7E",X"01",X"CF",X"A0",X"0F",X"BE",X"0F",X"BE",X"0F",X"A9",X"0F",X"C3",X"0F",X"C3",
		X"0F",X"DC",X"0F",X"DD",X"21",X"44",X"98",X"FD",X"21",X"20",X"9D",X"3A",X"07",X"98",X"0F",X"30",
		X"14",X"FD",X"35",X"02",X"FD",X"7E",X"02",X"20",X"04",X"FD",X"36",X"02",X"03",X"21",X"74",X"0F",
		X"E7",X"7E",X"DD",X"77",X"00",X"FD",X"7E",X"01",X"B7",X"28",X"C6",X"FE",X"03",X"28",X"C2",X"FD",
		X"35",X"00",X"18",X"BD",X"CC",X"D0",X"D4",X"05",X"06",X"07",X"DD",X"21",X"40",X"98",X"DD",X"7E",
		X"01",X"DD",X"96",X"05",X"30",X"02",X"ED",X"44",X"FE",X"0C",X"D0",X"DD",X"7E",X"02",X"DD",X"96",
		X"06",X"30",X"02",X"ED",X"44",X"FE",X"0C",X"D0",X"21",X"02",X"98",X"36",X"80",X"2C",X"34",X"C9",
		X"11",X"01",X"90",X"FD",X"36",X"00",X"40",X"18",X"03",X"11",X"FF",X"70",X"DD",X"7E",X"02",X"83",
		X"DD",X"77",X"02",X"BA",X"C0",X"FD",X"34",X"01",X"C9",X"01",X"70",X"68",X"18",X"08",X"01",X"90",
		X"88",X"18",X"03",X"01",X"70",X"88",X"FD",X"7E",X"00",X"CD",X"AB",X"10",X"FD",X"7E",X"1F",X"FD",
		X"86",X"00",X"FD",X"77",X"00",X"E6",X"3F",X"C0",X"FD",X"34",X"01",X"C9",X"FD",X"36",X"01",X"00",
		X"C9",X"DD",X"21",X"40",X"98",X"CD",X"EF",X"0F",X"DD",X"21",X"44",X"98",X"C3",X"12",X"10",X"11",
		X"31",X"10",X"21",X"02",X"98",X"35",X"7E",X"20",X"02",X"2C",X"34",X"0F",X"0F",X"E6",X"03",X"EB",
		X"E7",X"7E",X"DD",X"77",X"00",X"3E",X"04",X"E7",X"7E",X"DD",X"77",X"03",X"C9",X"11",X"39",X"10",
		X"18",X"E0",X"3A",X"3F",X"9D",X"07",X"30",X"F5",X"21",X"22",X"9D",X"35",X"7E",X"20",X"02",X"36",
		X"03",X"21",X"74",X"0F",X"E7",X"7E",X"DD",X"77",X"00",X"3E",X"03",X"E7",X"7E",X"DD",X"77",X"03",
		X"C9",X"F1",X"E1",X"D1",X"C1",X"10",X"0C",X"04",X"08",X"83",X"81",X"93",X"91",X"1A",X"09",X"08",
		X"07",X"CD",X"6D",X"22",X"21",X"01",X"98",X"34",X"C9",X"CD",X"55",X"11",X"CD",X"92",X"15",X"CD",
		X"55",X"11",X"FE",X"03",X"20",X"17",X"11",X"0E",X"03",X"FF",X"1E",X"03",X"FF",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"05",X"C0",
		X"34",X"C9",X"3A",X"03",X"98",X"CF",X"7C",X"10",X"34",X"0B",X"9D",X"10",X"3A",X"07",X"98",X"0F",
		X"D8",X"CD",X"91",X"11",X"3A",X"2C",X"98",X"FE",X"20",X"D8",X"AF",X"32",X"2C",X"98",X"CD",X"61",
		X"11",X"CD",X"6F",X"11",X"11",X"01",X"08",X"FF",X"21",X"03",X"98",X"34",X"C9",X"21",X"03",X"98",
		X"36",X"00",X"2D",X"2D",X"34",X"C9",X"AF",X"32",X"01",X"98",X"C9",X"6F",X"CB",X"3F",X"AD",X"ED",
		X"47",X"11",X"7A",X"4D",X"26",X"00",X"29",X"19",X"CD",X"0D",X"11",X"80",X"DD",X"77",X"01",X"EB",
		X"23",X"CD",X"0D",X"11",X"81",X"DD",X"77",X"02",X"FD",X"7E",X"00",X"E6",X"0F",X"FE",X"08",X"C0",
		X"FD",X"AE",X"00",X"0F",X"0F",X"0F",X"0F",X"FD",X"CB",X"1F",X"7E",X"20",X"04",X"C6",X"09",X"E6",
		X"0F",X"4F",X"06",X"00",X"2A",X"1B",X"99",X"09",X"7E",X"DD",X"77",X"00",X"C9",X"91",X"8D",X"89",
		X"85",X"81",X"9D",X"99",X"95",X"91",X"8D",X"89",X"85",X"81",X"9D",X"99",X"95",X"D1",X"CD",X"C9",
		X"C5",X"C1",X"FD",X"F9",X"F5",X"F1",X"ED",X"E9",X"E5",X"E1",X"DD",X"D9",X"D5",X"5E",X"16",X"00",
		X"EB",X"29",X"29",X"29",X"29",X"ED",X"57",X"07",X"ED",X"47",X"7C",X"D0",X"ED",X"44",X"C9",X"ED",
		X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"01",X"1C",X"00",X"EB",X"09",X"EB",X"3D",X"20",X"EF",
		X"C9",X"D5",X"3E",X"04",X"CD",X"1F",X"11",X"EB",X"E3",X"EB",X"CB",X"DA",X"3E",X"04",X"CD",X"1F",
		X"11",X"D1",X"C9",X"D5",X"3E",X"04",X"CD",X"1F",X"11",X"EB",X"E3",X"EB",X"CB",X"DA",X"3E",X"04",
		X"CD",X"1F",X"11",X"D1",X"C9",X"11",X"01",X"98",X"21",X"17",X"98",X"4E",X"1A",X"EB",X"71",X"12",
		X"C9",X"11",X"00",X"03",X"FF",X"1C",X"FF",X"1C",X"3A",X"0A",X"98",X"B7",X"20",X"FF",X"C9",X"11",
		X"00",X"02",X"FF",X"1C",X"3A",X"0A",X"98",X"B7",X"20",X"FF",X"1C",X"FF",X"C9",X"21",X"6A",X"8E",
		X"11",X"18",X"00",X"0E",X"02",X"06",X"08",X"36",X"C0",X"23",X"10",X"FB",X"0D",X"19",X"20",X"F5",
		X"C9",X"21",X"B7",X"11",X"E5",X"3A",X"2C",X"98",X"3C",X"32",X"2C",X"98",X"6F",X"26",X"00",X"E6",
		X"1E",X"BD",X"20",X"03",X"25",X"ED",X"44",X"6F",X"29",X"29",X"29",X"29",X"11",X"00",X"86",X"19",
		X"3E",X"10",X"01",X"01",X"1C",X"D7",X"C9",X"7D",X"E6",X"E0",X"6F",X"CB",X"94",X"01",X"01",X"08",
		X"3E",X"10",X"D7",X"C9",X"22",X"30",X"98",X"11",X"04",X"88",X"01",X"04",X"00",X"CD",X"DC",X"11",
		X"2A",X"30",X"98",X"3E",X"04",X"E7",X"11",X"00",X"8C",X"01",X"1C",X"00",X"D9",X"06",X"20",X"D9",
		X"C5",X"ED",X"B0",X"C1",X"B7",X"ED",X"42",X"EB",X"ED",X"42",X"3E",X"20",X"E7",X"EB",X"D9",X"10",
		X"EE",X"C9",X"21",X"10",X"39",X"10",X"1C",X"01",X"0A",X"01",X"2B",X"01",X"09",X"20",X"0C",X"20",
		X"40",X"02",X"30",X"20",X"36",X"01",X"25",X"10",X"08",X"10",X"50",X"02",X"20",X"20",X"20",X"02",
		X"50",X"10",X"40",X"02",X"40",X"20",X"40",X"20",X"40",X"20",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"01",X"40",X"20",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"02",X"40",X"20",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"01",X"40",X"01",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"10",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"10",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"20",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"3A",X"09",X"99",X"B7",X"C8",X"FD",
		X"E5",X"E1",X"4F",X"06",X"03",X"2C",X"AF",X"86",X"86",X"2C",X"10",X"FB",X"06",X"06",X"86",X"2C",
		X"10",X"FC",X"FE",X"1E",X"D8",X"41",X"3E",X"F0",X"A5",X"6F",X"D9",X"CD",X"8F",X"01",X"E6",X"1E",
		X"21",X"FE",X"12",X"E7",X"7E",X"B7",X"28",X"F3",X"23",X"08",X"7E",X"D9",X"B5",X"6F",X"7E",X"B7",
		X"28",X"E4",X"35",X"3E",X"F0",X"A5",X"6F",X"08",X"B5",X"6F",X"34",X"10",X"D9",X"C9",X"00",X"00",
		X"04",X"01",X"06",X"02",X"08",X"03",X"0B",X"04",X"0B",X"05",X"0B",X"06",X"0B",X"07",X"0B",X"08",
		X"0B",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"07",X"02",X"09",X"03",X"06",X"40",
		X"1A",X"E6",X"3F",X"FE",X"10",X"30",X"06",X"B5",X"6F",X"34",X"E6",X"F0",X"6F",X"13",X"10",X"F0",
		X"3E",X"0F",X"B5",X"6F",X"06",X"03",X"7E",X"36",X"00",X"2D",X"86",X"36",X"00",X"10",X"FA",X"77",
		X"C9",X"21",X"02",X"99",X"3E",X"03",X"BE",X"38",X"01",X"7E",X"87",X"87",X"87",X"ED",X"44",X"C6",
		X"80",X"2C",X"77",X"2E",X"07",X"36",X"04",X"3A",X"02",X"99",X"FE",X"08",X"38",X"02",X"3E",X"07",
		X"87",X"21",X"9F",X"13",X"E7",X"4E",X"23",X"46",X"ED",X"43",X"0C",X"99",X"3A",X"02",X"99",X"47",
		X"E6",X"0F",X"4F",X"A8",X"0F",X"47",X"0F",X"0F",X"80",X"81",X"E6",X"07",X"21",X"96",X"13",X"E7",
		X"7E",X"32",X"06",X"99",X"47",X"E6",X"0E",X"4F",X"A8",X"0F",X"0F",X"0F",X"0F",X"E6",X"0E",X"81",
		X"6F",X"67",X"22",X"09",X"99",X"C9",X"44",X"54",X"64",X"45",X"56",X"55",X"65",X"66",X"46",X"18",
		X"00",X"10",X"01",X"0C",X"02",X"0A",X"03",X"08",X"04",X"06",X"05",X"05",X"06",X"04",X"07",X"11",
		X"A0",X"99",X"21",X"C2",X"13",X"01",X"10",X"00",X"ED",X"B0",X"21",X"C2",X"13",X"0E",X"10",X"ED",
		X"B0",X"C9",X"01",X"08",X"08",X"08",X"01",X"02",X"02",X"01",X"02",X"02",X"00",X"00",X"01",X"00",
		X"00",X"00",X"3A",X"02",X"99",X"87",X"87",X"87",X"6F",X"67",X"22",X"0E",X"99",X"01",X"01",X"40",
		X"3E",X"FF",X"DD",X"E5",X"E1",X"D7",X"CD",X"C4",X"14",X"CD",X"65",X"14",X"CD",X"53",X"15",X"CD",
		X"3C",X"14",X"C9",X"3A",X"08",X"99",X"D6",X"04",X"2E",X"00",X"67",X"22",X"06",X"9D",X"E6",X"F0",
		X"6F",X"AC",X"87",X"87",X"87",X"87",X"67",X"11",X"10",X"10",X"19",X"22",X"04",X"9D",X"3A",X"07",
		X"9D",X"6F",X"26",X"9A",X"6E",X"26",X"00",X"29",X"29",X"29",X"3E",X"04",X"E7",X"11",X"3B",X"45",
		X"19",X"5E",X"23",X"56",X"ED",X"53",X"08",X"9D",X"11",X"82",X"99",X"3A",X"09",X"98",X"B7",X"28",
		X"02",X"1E",X"92",X"01",X"08",X"00",X"21",X"02",X"9D",X"ED",X"B0",X"C9",X"DD",X"E5",X"E1",X"FD",
		X"E5",X"D1",X"01",X"00",X"10",X"1A",X"B7",X"28",X"17",X"7D",X"E6",X"C0",X"6F",X"D9",X"CD",X"8F",
		X"01",X"D9",X"E6",X"3F",X"B5",X"6F",X"7E",X"3C",X"20",X"EF",X"71",X"EB",X"35",X"EB",X"20",X"E9",
		X"0C",X"13",X"10",X"E1",X"C9",X"3A",X"06",X"99",X"4F",X"E6",X"0F",X"47",X"A9",X"0F",X"0F",X"0F",
		X"0F",X"4F",X"ED",X"43",X"24",X"98",X"0E",X"24",X"11",X"18",X"19",X"DD",X"E5",X"E1",X"CD",X"B1",
		X"14",X"ED",X"4B",X"24",X"98",X"58",X"41",X"16",X"00",X"4A",X"1C",X"CB",X"38",X"30",X"01",X"0C",
		X"36",X"1E",X"19",X"36",X"1C",X"2C",X"36",X"1F",X"19",X"36",X"1D",X"2C",X"10",X"F2",X"CB",X"41",
		X"28",X"06",X"36",X"23",X"19",X"36",X"22",X"2C",X"3A",X"25",X"98",X"47",X"0E",X"21",X"11",X"1A",
		X"1B",X"36",X"20",X"2C",X"CB",X"38",X"30",X"02",X"71",X"2C",X"72",X"2C",X"73",X"2C",X"10",X"FA",
		X"36",X"20",X"2C",X"C9",X"3A",X"06",X"99",X"47",X"E6",X"03",X"4F",X"A8",X"0F",X"0F",X"E6",X"0C",
		X"B1",X"87",X"21",X"3D",X"15",X"E7",X"7E",X"32",X"08",X"99",X"23",X"7E",X"5F",X"AF",X"57",X"DD",
		X"E5",X"E1",X"19",X"77",X"FD",X"35",X"00",X"CD",X"13",X"15",X"23",X"D9",X"FD",X"E5",X"C1",X"CD",
		X"8F",X"01",X"E6",X"07",X"28",X"F9",X"21",X"0B",X"15",X"E7",X"7E",X"57",X"60",X"69",X"E7",X"35",
		X"F2",X"07",X"15",X"34",X"C3",X"EF",X"14",X"7A",X"D9",X"77",X"C9",X"00",X"01",X"02",X"03",X"05",
		X"07",X"09",X"0C",X"2B",X"2B",X"FD",X"7E",X"03",X"B7",X"28",X"06",X"36",X"03",X"FD",X"35",X"03",
		X"C9",X"FD",X"7E",X"09",X"B7",X"28",X"06",X"36",X"09",X"FD",X"35",X"09",X"C9",X"36",X"09",X"AF",
		X"06",X"0F",X"FD",X"E5",X"D1",X"EB",X"23",X"B6",X"28",X"FC",X"35",X"EB",X"C9",X"8A",X"16",X"89",
		X"19",X"8A",X"1D",X"00",X"00",X"7A",X"16",X"79",X"19",X"7A",X"1D",X"00",X"00",X"8A",X"1C",X"89",
		X"20",X"8A",X"25",X"3A",X"06",X"99",X"C6",X"11",X"47",X"E6",X"0F",X"4F",X"A8",X"0F",X"0F",X"0F",
		X"0F",X"81",X"87",X"ED",X"44",X"C6",X"1C",X"C8",X"47",X"36",X"20",X"2C",X"10",X"FB",X"7D",X"E6",
		X"3F",X"2F",X"C6",X"40",X"47",X"04",X"FD",X"E5",X"D1",X"EB",X"7D",X"6F",X"D9",X"CD",X"8F",X"01",
		X"D9",X"E6",X"0F",X"12",X"B5",X"6F",X"E6",X"F0",X"35",X"34",X"28",X"EF",X"35",X"6F",X"13",X"10",
		X"EA",X"C9",X"CD",X"01",X"17",X"3A",X"01",X"98",X"CF",X"AF",X"15",X"E3",X"15",X"BE",X"16",X"7D",
		X"17",X"6C",X"18",X"DC",X"18",X"30",X"19",X"A8",X"19",X"F1",X"19",X"D9",X"1A",X"54",X"1D",X"AF",
		X"21",X"40",X"98",X"01",X"01",X"50",X"D7",X"21",X"00",X"9D",X"01",X"02",X"00",X"D7",X"21",X"00",
		X"9A",X"01",X"02",X"00",X"D7",X"21",X"00",X"99",X"01",X"01",X"80",X"D7",X"21",X"01",X"98",X"34",
		X"AF",X"32",X"2C",X"98",X"32",X"03",X"98",X"3A",X"08",X"98",X"47",X"3A",X"BE",X"98",X"A0",X"32",
		X"20",X"98",X"C9",X"CD",X"1E",X"16",X"3A",X"0A",X"98",X"B7",X"C4",X"4E",X"16",X"3A",X"08",X"98",
		X"B7",X"28",X"1A",X"11",X"0B",X"03",X"ED",X"53",X"24",X"98",X"21",X"01",X"98",X"34",X"2C",X"36",
		X"00",X"3A",X"08",X"98",X"B7",X"C4",X"91",X"20",X"AF",X"32",X"2C",X"98",X"C9",X"21",X"01",X"98",
		X"34",X"2C",X"36",X"01",X"AF",X"32",X"2C",X"98",X"3E",X"25",X"32",X"20",X"99",X"C9",X"11",X"80",
		X"99",X"21",X"6D",X"17",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"0C",X"98",X"32",X"00",X"99",X"CD",
		X"AF",X"13",X"CD",X"41",X"13",X"DD",X"21",X"00",X"9B",X"FD",X"21",X"A0",X"99",X"CD",X"D2",X"13",
		X"DD",X"21",X"00",X"99",X"21",X"00",X"9B",X"CD",X"0D",X"1C",X"CD",X"F3",X"13",X"C9",X"21",X"00",
		X"99",X"11",X"60",X"99",X"01",X"20",X"00",X"ED",X"B0",X"21",X"80",X"99",X"11",X"90",X"99",X"0E",
		X"10",X"ED",X"B0",X"11",X"40",X"9B",X"21",X"00",X"9B",X"0E",X"40",X"ED",X"B0",X"C9",X"81",X"8C",
		X"9A",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"3A",X"08",
		X"98",X"B7",X"28",X"0B",X"ED",X"5B",X"24",X"98",X"FF",X"3A",X"0A",X"98",X"B7",X"28",X"08",X"11",
		X"01",X"02",X"FF",X"11",X"02",X"03",X"FF",X"11",X"00",X"02",X"FF",X"1E",X"02",X"FF",X"11",X"01",
		X"03",X"FF",X"1D",X"FF",X"21",X"2C",X"98",X"34",X"21",X"6E",X"16",X"C3",X"C4",X"11",X"3A",X"2C",
		X"98",X"FE",X"21",X"30",X"16",X"3A",X"07",X"98",X"0F",X"D8",X"3E",X"10",X"CD",X"91",X"11",X"3A",
		X"2C",X"98",X"FE",X"20",X"D8",X"11",X"0E",X"03",X"FF",X"18",X"B3",X"21",X"02",X"98",X"35",X"28",
		X"11",X"3E",X"07",X"A6",X"C0",X"3E",X"18",X"A6",X"ED",X"5B",X"24",X"98",X"20",X"02",X"CB",X"FB",
		X"FF",X"C9",X"36",X"40",X"2D",X"34",X"11",X"CB",X"03",X"FF",X"1E",X"8E",X"FF",X"CD",X"20",X"17",
		X"C9",X"3A",X"08",X"98",X"0F",X"D0",X"3A",X"07",X"98",X"47",X"E6",X"07",X"C0",X"11",X"01",X"03",
		X"3A",X"09",X"98",X"0F",X"30",X"01",X"1C",X"3E",X"18",X"A0",X"20",X"02",X"CB",X"FB",X"FF",X"C9",
		X"3A",X"06",X"99",X"ED",X"44",X"C6",X"66",X"32",X"38",X"98",X"C9",X"3A",X"06",X"99",X"47",X"3A",
		X"38",X"98",X"ED",X"44",X"C6",X"66",X"B8",X"3A",X"38",X"98",X"CD",X"CD",X"30",X"3A",X"38",X"98",
		X"CD",X"47",X"17",X"32",X"38",X"98",X"C9",X"4F",X"E6",X"F0",X"47",X"A9",X"4F",X"3A",X"06",X"99",
		X"C6",X"88",X"5F",X"E6",X"F0",X"57",X"AB",X"5F",X"B9",X"20",X"0A",X"78",X"BA",X"30",X"0B",X"7B",
		X"2F",X"C6",X"2F",X"80",X"C9",X"3E",X"02",X"80",X"81",X"C9",X"3E",X"FF",X"C9",X"01",X"00",X"90",
		X"50",X"A0",X"30",X"F0",X"84",X"00",X"02",X"00",X"00",X"D1",X"01",X"01",X"C1",X"3A",X"38",X"98",
		X"3C",X"28",X"3A",X"CD",X"2B",X"17",X"3A",X"38",X"98",X"3C",X"C0",X"11",X"00",X"9D",X"21",X"80",
		X"99",X"01",X"10",X"00",X"3A",X"09",X"98",X"B7",X"28",X"02",X"2E",X"90",X"ED",X"B0",X"21",X"00",
		X"99",X"35",X"CD",X"15",X"18",X"CD",X"EF",X"24",X"CD",X"E9",X"17",X"11",X"00",X"06",X"FF",X"11",
		X"00",X"05",X"FF",X"3A",X"0C",X"99",X"32",X"9B",X"9C",X"C3",X"D1",X"1C",X"C9",X"21",X"02",X"98",
		X"35",X"C0",X"3A",X"0A",X"99",X"B7",X"28",X"16",X"21",X"01",X"98",X"34",X"2C",X"2C",X"36",X"00",
		X"3E",X"10",X"32",X"98",X"9C",X"CD",X"82",X"20",X"CD",X"7B",X"2E",X"C3",X"13",X"20",X"21",X"08",
		X"C0",X"22",X"01",X"98",X"AF",X"32",X"2C",X"98",X"C9",X"3A",X"08",X"9D",X"21",X"F5",X"17",X"E7",
		X"7E",X"32",X"0C",X"9D",X"C9",X"D1",X"F1",X"C1",X"E1",X"F1",X"C1",X"F1",X"E1",X"C1",X"D1",X"D1",
		X"E1",X"F1",X"C1",X"D1",X"E1",X"F1",X"F1",X"C1",X"C1",X"F1",X"F1",X"E1",X"E1",X"C1",X"C1",X"D1",
		X"D1",X"D1",X"D1",X"E1",X"E1",X"11",X"30",X"9D",X"21",X"2C",X"18",X"3E",X"04",X"01",X"10",X"00",
		X"EB",X"09",X"EB",X"ED",X"B0",X"3D",X"20",X"F5",X"CD",X"58",X"24",X"C9",X"00",X"00",X"10",X"70",
		X"A0",X"30",X"F0",X"06",X"00",X"02",X"00",X"00",X"81",X"03",X"01",X"81",X"00",X"00",X"10",X"B0",
		X"A0",X"30",X"F0",X"0A",X"00",X"02",X"00",X"00",X"81",X"02",X"01",X"81",X"00",X"00",X"F0",X"30",
		X"A0",X"30",X"F0",X"E2",X"00",X"02",X"00",X"00",X"81",X"02",X"01",X"81",X"00",X"00",X"F0",X"70",
		X"A0",X"30",X"F0",X"E6",X"00",X"02",X"00",X"00",X"81",X"02",X"01",X"81",X"CD",X"AE",X"33",X"CD",
		X"C1",X"3B",X"CD",X"D1",X"1C",X"CD",X"CE",X"26",X"CD",X"7E",X"2A",X"3A",X"07",X"98",X"E6",X"0F",
		X"CC",X"22",X"20",X"3A",X"00",X"9D",X"B7",X"C0",X"CD",X"EF",X"1F",X"DD",X"21",X"00",X"9D",X"DD",
		X"36",X"06",X"F0",X"CD",X"3F",X"35",X"CD",X"B3",X"32",X"CD",X"98",X"35",X"3E",X"01",X"32",X"0D",
		X"9D",X"11",X"80",X"99",X"21",X"00",X"9D",X"36",X"01",X"01",X"10",X"00",X"3A",X"09",X"98",X"B7",
		X"28",X"02",X"1E",X"90",X"ED",X"B0",X"AF",X"32",X"2C",X"98",X"21",X"40",X"98",X"01",X"01",X"50",
		X"D7",X"21",X"A0",X"99",X"01",X"01",X"12",X"D7",X"21",X"98",X"9C",X"01",X"01",X"68",X"D7",X"21",
		X"80",X"9B",X"01",X"01",X"08",X"D7",X"21",X"01",X"98",X"36",X"05",X"C9",X"CD",X"95",X"11",X"3A",
		X"2C",X"98",X"FE",X"20",X"D8",X"21",X"6E",X"16",X"CD",X"C4",X"11",X"AF",X"21",X"20",X"99",X"01",
		X"01",X"20",X"D7",X"21",X"00",X"9D",X"01",X"02",X"00",X"D7",X"3E",X"08",X"32",X"89",X"9B",X"3A",
		X"00",X"99",X"B7",X"20",X"0A",X"3E",X"0A",X"32",X"01",X"98",X"AF",X"32",X"03",X"98",X"C9",X"CD",
		X"20",X"17",X"CD",X"FF",X"1B",X"28",X"06",X"3E",X"06",X"32",X"01",X"98",X"C9",X"21",X"03",X"40",
		X"22",X"01",X"98",X"11",X"00",X"9B",X"CD",X"44",X"1C",X"21",X"00",X"9B",X"CD",X"0D",X"1C",X"C9",
		X"3A",X"09",X"98",X"EE",X"01",X"32",X"09",X"98",X"20",X"47",X"21",X"00",X"99",X"11",X"60",X"99",
		X"01",X"20",X"00",X"ED",X"B0",X"11",X"40",X"9B",X"CD",X"44",X"1C",X"21",X"40",X"99",X"11",X"00",
		X"99",X"01",X"20",X"00",X"ED",X"B0",X"21",X"00",X"9B",X"CD",X"0D",X"1C",X"11",X"0B",X"03",X"ED",
		X"53",X"24",X"98",X"11",X"01",X"03",X"FF",X"1C",X"FF",X"21",X"0B",X"98",X"3A",X"09",X"98",X"A6",
		X"32",X"0E",X"98",X"EE",X"01",X"32",X"83",X"A1",X"21",X"01",X"98",X"36",X"02",X"2C",X"36",X"80",
		X"C9",X"21",X"00",X"99",X"11",X"40",X"99",X"01",X"20",X"00",X"ED",X"B0",X"11",X"00",X"9B",X"CD",
		X"44",X"1C",X"21",X"60",X"99",X"11",X"00",X"99",X"01",X"20",X"00",X"ED",X"B0",X"21",X"40",X"9B",
		X"CD",X"0D",X"1C",X"11",X"0C",X"03",X"18",X"B7",X"3A",X"06",X"99",X"47",X"E6",X"0F",X"4F",X"A8",
		X"47",X"87",X"81",X"ED",X"44",X"16",X"FF",X"87",X"5F",X"38",X"01",X"15",X"21",X"0E",X"86",X"19",
		X"79",X"87",X"87",X"4F",X"2F",X"C6",X"21",X"5F",X"16",X"00",X"78",X"0F",X"0F",X"D9",X"47",X"3E",
		X"10",X"D9",X"41",X"77",X"2C",X"10",X"FC",X"19",X"D9",X"10",X"F6",X"C9",X"3A",X"09",X"99",X"B7",
		X"11",X"13",X"01",X"28",X"01",X"1D",X"FF",X"3A",X"09",X"99",X"B7",X"CA",X"CD",X"20",X"C3",X"AA",
		X"20",X"3A",X"00",X"9D",X"0F",X"D2",X"88",X"18",X"3A",X"07",X"98",X"0F",X"D8",X"AF",X"21",X"44",
		X"98",X"01",X"01",X"60",X"D7",X"3A",X"02",X"98",X"FE",X"BF",X"CC",X"A8",X"19",X"3A",X"02",X"98",
		X"FE",X"B0",X"CC",X"DC",X"19",X"3A",X"02",X"98",X"47",X"E6",X"07",X"20",X"17",X"11",X"2B",X"03",
		X"3A",X"09",X"99",X"B7",X"28",X"01",X"1C",X"3E",X"18",X"A0",X"20",X"02",X"CB",X"FB",X"FF",X"1E",
		X"2F",X"FF",X"1C",X"FF",X"3A",X"09",X"99",X"B7",X"11",X"2D",X"03",X"28",X"01",X"1C",X"FF",X"21",
		X"02",X"98",X"35",X"C0",X"34",X"11",X"AD",X"03",X"FF",X"AF",X"21",X"40",X"98",X"01",X"01",X"60",
		X"D7",X"3E",X"10",X"CD",X"95",X"11",X"3A",X"2C",X"98",X"FE",X"20",X"D8",X"21",X"6E",X"16",X"CD",
		X"C4",X"11",X"CD",X"B3",X"32",X"11",X"00",X"9B",X"3A",X"09",X"98",X"0F",X"30",X"02",X"1E",X"40",
		X"CD",X"44",X"1C",X"3A",X"09",X"98",X"0F",X"38",X"57",X"11",X"00",X"9B",X"21",X"A0",X"99",X"D5",
		X"DD",X"E1",X"E5",X"FD",X"E1",X"CD",X"1E",X"13",X"CD",X"BA",X"12",X"21",X"02",X"99",X"34",X"CD",
		X"41",X"13",X"CD",X"D2",X"13",X"DD",X"E5",X"E1",X"CD",X"0D",X"1C",X"CD",X"F3",X"13",X"CD",X"20",
		X"17",X"AF",X"21",X"20",X"99",X"01",X"01",X"20",X"D7",X"21",X"80",X"9B",X"01",X"01",X"10",X"D7",
		X"21",X"98",X"9C",X"01",X"01",X"70",X"D7",X"21",X"20",X"9D",X"06",X"0B",X"11",X"20",X"00",X"77",
		X"19",X"10",X"FC",X"21",X"00",X"99",X"34",X"21",X"01",X"98",X"34",X"AF",X"32",X"03",X"98",X"C9",
		X"11",X"40",X"9B",X"21",X"A0",X"99",X"C3",X"7F",X"1A",X"3A",X"00",X"A1",X"CB",X"4F",X"28",X"15",
		X"3A",X"02",X"99",X"C6",X"02",X"E6",X"03",X"20",X"0C",X"3A",X"03",X"98",X"CF",X"FC",X"1A",X"1D",
		X"1B",X"4A",X"1B",X"69",X"1B",X"21",X"03",X"40",X"22",X"01",X"98",X"C9",X"21",X"03",X"98",X"34",
		X"11",X"13",X"00",X"21",X"4F",X"84",X"3E",X"64",X"CD",X"10",X"1B",X"3E",X"C0",X"21",X"4F",X"8C",
		X"0E",X"1C",X"06",X"0D",X"77",X"2C",X"10",X"FC",X"19",X"0D",X"20",X"F6",X"C9",X"21",X"40",X"02",
		X"22",X"02",X"98",X"AF",X"21",X"30",X"98",X"06",X"04",X"77",X"2C",X"10",X"FC",X"11",X"67",X"85",
		X"21",X"43",X"47",X"CD",X"39",X"1B",X"11",X"67",X"8D",X"3E",X"0A",X"01",X"0D",X"00",X"ED",X"B0",
		X"EB",X"01",X"13",X"00",X"09",X"EB",X"3D",X"20",X"F2",X"C9",X"21",X"02",X"98",X"2C",X"34",X"21",
		X"30",X"98",X"34",X"7E",X"EB",X"FE",X"06",X"30",X"9C",X"87",X"21",X"F5",X"1B",X"E7",X"4E",X"23",
		X"46",X"ED",X"43",X"32",X"98",X"1C",X"AF",X"12",X"C9",X"3A",X"07",X"98",X"0F",X"D8",X"21",X"31",
		X"98",X"7E",X"34",X"FE",X"15",X"38",X"06",X"3E",X"02",X"32",X"03",X"98",X"C9",X"11",X"20",X"00",
		X"47",X"04",X"21",X"47",X"84",X"E7",X"3A",X"30",X"98",X"FE",X"05",X"28",X"47",X"3E",X"07",X"B8",
		X"DC",X"DD",X"1B",X"E5",X"21",X"F0",X"1B",X"3A",X"30",X"98",X"E7",X"46",X"E1",X"7D",X"E6",X"1F",
		X"21",X"60",X"85",X"B5",X"6F",X"3A",X"31",X"98",X"90",X"38",X"23",X"FE",X"0D",X"D0",X"D9",X"2A",
		X"32",X"98",X"23",X"22",X"32",X"98",X"2B",X"11",X"0D",X"00",X"CD",X"C3",X"1B",X"D9",X"01",X"C0",
		X"06",X"09",X"D9",X"06",X"0A",X"7E",X"19",X"D9",X"77",X"19",X"D9",X"10",X"F8",X"C9",X"06",X"0A",
		X"3E",X"10",X"18",X"04",X"3E",X"10",X"06",X"1C",X"77",X"19",X"10",X"FC",X"C9",X"3E",X"71",X"CD",
		X"D6",X"1B",X"01",X"80",X"04",X"09",X"3E",X"C0",X"C3",X"D6",X"1B",X"08",X"07",X"05",X"01",X"00",
		X"00",X"01",X"03",X"07",X"08",X"43",X"47",X"47",X"48",X"4B",X"49",X"4F",X"4A",X"53",X"4B",X"21",
		X"40",X"99",X"3A",X"09",X"98",X"B7",X"20",X"02",X"2E",X"60",X"7E",X"B7",X"C9",X"3A",X"06",X"99",
		X"C6",X"22",X"47",X"4F",X"E6",X"0F",X"5F",X"A8",X"0F",X"0F",X"0F",X"0F",X"57",X"3E",X"88",X"91",
		X"ED",X"53",X"2C",X"98",X"32",X"2E",X"98",X"16",X"9A",X"5F",X"D9",X"3A",X"2D",X"98",X"47",X"D9",
		X"3A",X"2C",X"98",X"01",X"10",X"00",X"ED",X"A0",X"1C",X"3D",X"20",X"FA",X"EB",X"09",X"09",X"EB",
		X"D9",X"10",X"EC",X"C9",X"3A",X"06",X"99",X"C6",X"22",X"47",X"4F",X"E6",X"0F",X"6F",X"A8",X"0F",
		X"0F",X"0F",X"0F",X"67",X"3E",X"88",X"91",X"22",X"2C",X"98",X"32",X"2E",X"98",X"26",X"9A",X"6F",
		X"D9",X"3A",X"2D",X"98",X"47",X"D9",X"3A",X"2C",X"98",X"01",X"10",X"00",X"08",X"7E",X"E6",X"3F",
		X"12",X"23",X"13",X"08",X"0D",X"2C",X"3D",X"20",X"F3",X"09",X"09",X"D9",X"10",X"E7",X"21",X"00",
		X"9A",X"AF",X"01",X"01",X"00",X"D7",X"C9",X"21",X"60",X"98",X"3A",X"00",X"9E",X"B7",X"28",X"38",
		X"EB",X"3A",X"0E",X"98",X"0F",X"30",X"1B",X"01",X"06",X"00",X"21",X"14",X"9E",X"ED",X"B0",X"CD",
		X"BE",X"1C",X"21",X"0E",X"9E",X"11",X"80",X"98",X"06",X"06",X"7E",X"2F",X"12",X"23",X"13",X"10",
		X"F9",X"C9",X"21",X"14",X"9E",X"CD",X"A8",X"1C",X"CD",X"BE",X"1C",X"21",X"0E",X"9E",X"0E",X"0A",
		X"EB",X"09",X"EB",X"0E",X"06",X"ED",X"B0",X"C9",X"21",X"80",X"98",X"01",X"01",X"10",X"AF",X"D7",
		X"C9",X"CD",X"87",X"1C",X"06",X"08",X"11",X"20",X"00",X"21",X"40",X"98",X"DD",X"21",X"00",X"9D",
		X"3A",X"0E",X"98",X"0F",X"38",X"35",X"0E",X"07",X"DD",X"7E",X"00",X"B7",X"28",X"22",X"DD",X"7E",
		X"0C",X"77",X"2C",X"2C",X"DD",X"7E",X"02",X"D6",X"08",X"77",X"2D",X"DD",X"7E",X"03",X"C6",X"27",
		X"2F",X"C6",X"20",X"77",X"DD",X"7E",X"0D",X"2C",X"2C",X"77",X"2C",X"DD",X"19",X"10",X"D9",X"C9",
		X"2C",X"77",X"2C",X"77",X"2C",X"2C",X"DD",X"19",X"10",X"CE",X"C9",X"DD",X"7E",X"00",X"B7",X"28",
		X"28",X"0E",X"00",X"DD",X"7E",X"0C",X"EE",X"02",X"77",X"2C",X"DD",X"7E",X"03",X"D6",X"08",X"30",
		X"02",X"0E",X"80",X"77",X"2C",X"DD",X"7E",X"02",X"ED",X"44",X"D6",X"07",X"77",X"2C",X"DD",X"7E",
		X"0D",X"B1",X"77",X"2C",X"DD",X"19",X"10",X"D3",X"C9",X"2C",X"77",X"2C",X"77",X"2C",X"2C",X"DD",
		X"19",X"10",X"C8",X"C9",X"CD",X"FF",X"1B",X"20",X"04",X"21",X"C0",X"21",X"E5",X"3A",X"03",X"98",
		X"CF",X"69",X"1D",X"7F",X"1D",X"95",X"1D",X"D2",X"1D",X"11",X"0D",X"03",X"FF",X"3A",X"09",X"98",
		X"B7",X"1E",X"0B",X"28",X"01",X"1C",X"FF",X"21",X"03",X"98",X"34",X"2D",X"36",X"60",X"C9",X"21",
		X"02",X"98",X"35",X"C0",X"2C",X"34",X"CD",X"22",X"1E",X"11",X"8C",X"03",X"FF",X"1C",X"FF",X"16",
		X"08",X"FF",X"C3",X"F0",X"20",X"3A",X"28",X"98",X"B7",X"C4",X"8F",X"1E",X"21",X"02",X"98",X"35",
		X"C0",X"11",X"A0",X"03",X"FF",X"21",X"29",X"98",X"36",X"0A",X"2D",X"7E",X"B7",X"20",X"01",X"34",
		X"3A",X"28",X"98",X"B7",X"C4",X"38",X"1F",X"21",X"28",X"98",X"7E",X"B7",X"36",X"00",X"28",X"02",
		X"3E",X"80",X"3C",X"21",X"03",X"98",X"34",X"2D",X"77",X"11",X"FF",X"08",X"FF",X"AF",X"32",X"2C",
		X"98",X"C9",X"21",X"02",X"98",X"35",X"C0",X"34",X"3E",X"10",X"CD",X"95",X"11",X"3A",X"2C",X"98",
		X"FE",X"20",X"D8",X"CD",X"FF",X"1B",X"28",X"1B",X"21",X"05",X"80",X"01",X"20",X"1A",X"11",X"06",
		X"00",X"3E",X"10",X"2C",X"77",X"10",X"FC",X"19",X"06",X"1A",X"0D",X"20",X"F6",X"3E",X"06",X"32",
		X"01",X"98",X"C9",X"21",X"17",X"1E",X"11",X"00",X"98",X"01",X"0A",X"00",X"ED",X"B0",X"AF",X"32",
		X"0E",X"98",X"3C",X"32",X"83",X"A1",X"C9",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AF",X"32",X"28",X"98",X"DD",X"21",X"C0",X"99",X"3A",X"09",X"98",X"B7",X"28",X"04",
		X"DD",X"21",X"C3",X"99",X"06",X"0A",X"21",X"02",X"9F",X"11",X"0E",X"00",X"7E",X"DD",X"BE",X"02",
		X"20",X"11",X"2B",X"7E",X"DD",X"BE",X"01",X"20",X"0B",X"2B",X"7E",X"DD",X"BE",X"00",X"20",X"05",
		X"C3",X"57",X"1E",X"2B",X"2B",X"38",X"04",X"19",X"10",X"E2",X"C9",X"E5",X"21",X"28",X"98",X"70",
		X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"05",X"28",X"11",X"21",X"6B",X"9F",X"11",
		X"77",X"9F",X"78",X"87",X"87",X"4F",X"87",X"81",X"4F",X"06",X"00",X"ED",X"B8",X"DD",X"E5",X"E1",
		X"D1",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"EB",X"01",X"01",X"09",X"3E",X"40",X"D7",X"C9",X"21",
		X"02",X"98",X"34",X"EB",X"21",X"04",X"99",X"DF",X"20",X"04",X"36",X"08",X"EB",X"35",X"3A",X"02",
		X"98",X"47",X"E6",X"03",X"20",X"0A",X"11",X"32",X"03",X"CB",X"50",X"28",X"02",X"CB",X"FB",X"FF",
		X"21",X"2B",X"98",X"DF",X"CD",X"0D",X"3B",X"B7",X"C4",X"D8",X"1E",X"C3",X"38",X"1F",X"21",X"2A",
		X"98",X"34",X"28",X"06",X"2D",X"34",X"3E",X"04",X"BE",X"C0",X"21",X"29",X"98",X"36",X"10",X"21",
		X"02",X"98",X"36",X"01",X"E1",X"C3",X"38",X"1F",X"21",X"2B",X"98",X"DF",X"C0",X"36",X"10",X"2D",
		X"47",X"E6",X"33",X"28",X"D9",X"E6",X"30",X"28",X"19",X"34",X"28",X"DE",X"2D",X"CB",X"68",X"3E",
		X"01",X"28",X"02",X"ED",X"44",X"86",X"FE",X"FF",X"20",X"02",X"3E",X"03",X"FE",X"04",X"28",X"CA",
		X"77",X"2C",X"78",X"E6",X"03",X"C8",X"4F",X"2D",X"7E",X"FE",X"03",X"D0",X"2D",X"46",X"21",X"7B",
		X"9F",X"11",X"F4",X"FF",X"19",X"10",X"FD",X"E7",X"CB",X"49",X"28",X"0E",X"34",X"3E",X"5B",X"BE",
		X"D0",X"36",X"3B",X"21",X"2A",X"98",X"34",X"28",X"A1",X"C9",X"35",X"7E",X"FE",X"3B",X"D0",X"36",
		X"5B",X"21",X"2A",X"98",X"34",X"28",X"93",X"C9",X"CD",X"8D",X"1F",X"DD",X"21",X"7B",X"9F",X"21",
		X"A4",X"86",X"11",X"02",X"00",X"01",X"F4",X"FF",X"3A",X"28",X"98",X"DD",X"09",X"19",X"3D",X"20",
		X"FA",X"DD",X"E5",X"D1",X"06",X"03",X"CD",X"D3",X"03",X"2B",X"3A",X"29",X"98",X"D6",X"03",X"5F",
		X"3E",X"8E",X"16",X"2B",X"01",X"10",X"04",X"20",X"0B",X"36",X"37",X"CD",X"B5",X"1F",X"16",X"36",
		X"05",X"CD",X"83",X"1F",X"1D",X"71",X"1C",X"20",X"01",X"72",X"CD",X"B5",X"1F",X"CD",X"83",X"1F",
		X"10",X"F3",X"C9",X"08",X"7D",X"D6",X"20",X"6F",X"30",X"01",X"25",X"08",X"C9",X"3A",X"07",X"98",
		X"47",X"E6",X"07",X"C0",X"3E",X"18",X"A0",X"28",X"22",X"FE",X"08",X"C0",X"21",X"84",X"84",X"3A",
		X"28",X"98",X"87",X"85",X"6F",X"3E",X"8E",X"01",X"10",X"18",X"11",X"20",X"00",X"71",X"CD",X"B5",
		X"1F",X"19",X"10",X"F9",X"C9",X"CB",X"DC",X"77",X"CB",X"9C",X"C9",X"11",X"FF",X"08",X"FF",X"C9",
		X"21",X"CE",X"99",X"5E",X"16",X"99",X"1A",X"3C",X"C8",X"3D",X"47",X"3E",X"FF",X"12",X"1C",X"20",
		X"02",X"1E",X"D0",X"73",X"3E",X"10",X"B8",X"28",X"17",X"3A",X"BF",X"98",X"21",X"08",X"98",X"B6",
		X"C8",X"78",X"C3",X"F0",X"1F",X"3E",X"01",X"32",X"82",X"A1",X"C9",X"AF",X"32",X"82",X"A1",X"AF",
		X"32",X"00",X"A1",X"3E",X"00",X"32",X"80",X"A1",X"00",X"00",X"00",X"00",X"3E",X"01",X"32",X"80",
		X"A1",X"C9",X"47",X"11",X"CD",X"99",X"1A",X"6F",X"26",X"99",X"70",X"2C",X"20",X"02",X"2E",X"D0",
		X"EB",X"73",X"C9",X"3E",X"1E",X"CD",X"02",X"20",X"3E",X"04",X"C3",X"02",X"20",X"3E",X"84",X"C3",
		X"02",X"20",X"2A",X"30",X"99",X"29",X"29",X"7C",X"E6",X"0F",X"C8",X"C6",X"1D",X"C3",X"02",X"20",
		X"3E",X"01",X"CD",X"02",X"20",X"3E",X"02",X"CD",X"02",X"20",X"3E",X"03",X"C3",X"02",X"20",X"3E",
		X"05",X"C3",X"02",X"20",X"3E",X"85",X"C3",X"02",X"20",X"3E",X"85",X"CD",X"02",X"20",X"3E",X"06",
		X"C3",X"02",X"20",X"3E",X"85",X"3E",X"86",X"C3",X"02",X"20",X"3E",X"07",X"C3",X"02",X"20",X"3E",
		X"08",X"C3",X"02",X"20",X"3E",X"87",X"C3",X"02",X"20",X"3E",X"09",X"CD",X"02",X"20",X"3E",X"0A",
		X"C3",X"02",X"20",X"3E",X"0B",X"C3",X"02",X"20",X"3E",X"0C",X"C3",X"02",X"20",X"3E",X"0D",X"C3",
		X"02",X"20",X"3E",X"0E",X"C3",X"02",X"20",X"3E",X"0F",X"C3",X"02",X"20",X"3E",X"10",X"C3",X"02",
		X"20",X"3E",X"00",X"CD",X"02",X"20",X"3E",X"11",X"CD",X"02",X"20",X"3E",X"12",X"CD",X"02",X"20",
		X"3E",X"13",X"CD",X"02",X"20",X"3E",X"14",X"C3",X"02",X"20",X"3E",X"84",X"CD",X"02",X"20",X"3E",
		X"85",X"CD",X"02",X"20",X"3E",X"86",X"CD",X"02",X"20",X"3E",X"87",X"CD",X"02",X"20",X"3E",X"15",
		X"CD",X"02",X"20",X"3E",X"16",X"CD",X"02",X"20",X"3E",X"17",X"C3",X"02",X"20",X"3E",X"84",X"CD",
		X"02",X"20",X"3E",X"85",X"CD",X"02",X"20",X"3E",X"86",X"CD",X"02",X"20",X"3E",X"87",X"CD",X"02",
		X"20",X"3E",X"18",X"CD",X"02",X"20",X"3E",X"19",X"CD",X"02",X"20",X"3E",X"1A",X"C3",X"02",X"20",
		X"3E",X"00",X"CD",X"02",X"20",X"3E",X"1B",X"CD",X"02",X"20",X"3E",X"1C",X"CD",X"02",X"20",X"3E",
		X"1D",X"C3",X"02",X"20",X"3A",X"BE",X"98",X"B7",X"28",X"0B",X"AF",X"32",X"12",X"98",X"21",X"00",
		X"00",X"22",X"00",X"98",X"C9",X"21",X"C0",X"21",X"E5",X"3A",X"01",X"98",X"CF",X"25",X"21",X"38",
		X"21",X"8E",X"21",X"BB",X"21",X"21",X"40",X"98",X"01",X"01",X"50",X"AF",X"D7",X"32",X"2C",X"98",
		X"21",X"02",X"98",X"36",X"10",X"2D",X"34",X"C9",X"3A",X"07",X"98",X"0F",X"D8",X"3E",X"10",X"CD",
		X"91",X"11",X"3A",X"2C",X"98",X"FE",X"20",X"D8",X"11",X"01",X"02",X"FF",X"11",X"02",X"03",X"FF",
		X"11",X"00",X"02",X"FF",X"1E",X"02",X"FF",X"11",X"01",X"03",X"FF",X"1D",X"FF",X"CD",X"EF",X"1F",
		X"21",X"01",X"98",X"34",X"2C",X"36",X"FF",X"2C",X"AF",X"77",X"32",X"09",X"98",X"32",X"2C",X"98",
		X"3C",X"32",X"83",X"A1",X"11",X"00",X"04",X"FF",X"11",X"07",X"03",X"FF",X"16",X"08",X"FF",X"3A",
		X"0D",X"98",X"47",X"E6",X"0F",X"78",X"E6",X"F0",X"C8",X"0F",X"0F",X"0F",X"0F",X"C9",X"21",X"02",
		X"98",X"DF",X"CC",X"75",X"22",X"3A",X"12",X"98",X"A7",X"C8",X"3D",X"11",X"08",X"03",X"28",X"01",
		X"1C",X"0E",X"07",X"3A",X"07",X"98",X"47",X"E6",X"0F",X"C0",X"78",X"E6",X"30",X"20",X"04",X"CB",
		X"FB",X"CB",X"F9",X"FF",X"59",X"FF",X"11",X"00",X"04",X"FF",X"C9",X"AF",X"32",X"01",X"98",X"C9",
		X"3A",X"1C",X"98",X"E6",X"C0",X"C8",X"07",X"38",X"3B",X"3A",X"BE",X"98",X"B7",X"20",X"0B",X"3A",
		X"12",X"98",X"FE",X"02",X"D8",X"D6",X"02",X"32",X"12",X"98",X"AF",X"21",X"C3",X"99",X"01",X"01",
		X"03",X"D7",X"21",X"00",X"01",X"22",X"09",X"98",X"AF",X"21",X"C0",X"99",X"01",X"01",X"03",X"D7",
		X"AF",X"32",X"01",X"98",X"32",X"0E",X"98",X"3C",X"32",X"83",X"A1",X"32",X"08",X"98",X"21",X"00",
		X"98",X"36",X"03",X"C9",X"3A",X"BE",X"98",X"B7",X"20",X"09",X"3A",X"12",X"98",X"A7",X"C8",X"3D",
		X"32",X"12",X"98",X"21",X"00",X"00",X"C3",X"E5",X"21",X"81",X"8C",X"9A",X"81",X"8C",X"8C",X"8E",
		X"8E",X"8E",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"92",X"92",X"92",X"92",X"92",X"93",X"93",X"93",X"24",X"01",X"30",X"10",X"3C",X"02",X"30",
		X"20",X"24",X"01",X"60",X"02",X"48",X"10",X"24",X"01",X"3C",X"20",X"24",X"02",X"30",X"20",X"21",
		X"01",X"2A",X"01",X"21",X"10",X"1E",X"02",X"1E",X"02",X"3C",X"20",X"24",X"01",X"24",X"01",X"2A",
		X"10",X"24",X"10",X"24",X"02",X"30",X"20",X"24",X"20",X"54",X"01",X"A8",X"FF",X"AF",X"32",X"2C",
		X"98",X"32",X"03",X"98",X"C9",X"3A",X"03",X"98",X"CF",X"81",X"22",X"97",X"22",X"E7",X"22",X"5A",
		X"23",X"3E",X"10",X"CD",X"95",X"11",X"3A",X"2C",X"98",X"FE",X"20",X"D8",X"21",X"19",X"22",X"CD",
		X"C4",X"11",X"21",X"03",X"98",X"34",X"C9",X"21",X"03",X"98",X"34",X"11",X"27",X"03",X"FF",X"1C",
		X"FF",X"1C",X"FF",X"1E",X"0F",X"FF",X"AF",X"21",X"00",X"9D",X"01",X"01",X"20",X"D7",X"21",X"00",
		X"99",X"01",X"01",X"40",X"D7",X"21",X"90",X"9C",X"01",X"01",X"70",X"D7",X"21",X"2E",X"23",X"11",
		X"00",X"9D",X"01",X"10",X"00",X"ED",X"B0",X"11",X"00",X"99",X"0E",X"10",X"ED",X"B0",X"11",X"54",
		X"9A",X"CD",X"D7",X"22",X"CD",X"D7",X"22",X"3E",X"04",X"01",X"20",X"00",X"ED",X"A0",X"1C",X"0D",
		X"3D",X"20",X"F9",X"EB",X"09",X"EB",X"C9",X"3E",X"C0",X"21",X"52",X"8D",X"11",X"20",X"00",X"06",
		X"0C",X"77",X"19",X"10",X"FC",X"21",X"53",X"8D",X"06",X"0C",X"77",X"19",X"10",X"FC",X"01",X"03",
		X"04",X"21",X"54",X"9A",X"E5",X"C5",X"7D",X"CD",X"CD",X"30",X"C1",X"E1",X"23",X"23",X"10",X"F4",
		X"06",X"04",X"11",X"18",X"00",X"19",X"0D",X"20",X"EB",X"AF",X"32",X"08",X"98",X"21",X"01",X"00",
		X"22",X"28",X"98",X"21",X"39",X"22",X"22",X"2A",X"98",X"21",X"03",X"98",X"34",X"C9",X"01",X"00",
		X"80",X"38",X"80",X"30",X"18",X"74",X"00",X"02",X"00",X"00",X"D1",X"01",X"01",X"C1",X"00",X"00",
		X"00",X"90",X"00",X"00",X"34",X"04",X"78",X"00",X"02",X"00",X"08",X"FF",X"00",X"00",X"02",X"03",
		X"01",X"1C",X"03",X"0B",X"00",X"1D",X"01",X"02",X"08",X"22",X"CD",X"71",X"23",X"3A",X"07",X"98",
		X"0F",X"DC",X"6E",X"32",X"CD",X"A7",X"34",X"CD",X"63",X"2E",X"CD",X"D1",X"1C",X"CD",X"7E",X"2A",
		X"C9",X"21",X"28",X"98",X"35",X"28",X"57",X"7E",X"FE",X"12",X"C0",X"2C",X"7E",X"3D",X"F8",X"3A",
		X"08",X"99",X"CD",X"27",X"24",X"3A",X"29",X"98",X"FE",X"10",X"38",X"1F",X"21",X"4E",X"24",X"CB",
		X"67",X"28",X"03",X"21",X"53",X"24",X"46",X"23",X"4E",X"23",X"EB",X"09",X"EB",X"ED",X"A0",X"ED",
		X"A0",X"CB",X"DA",X"3E",X"80",X"AE",X"1D",X"12",X"1D",X"12",X"C9",X"21",X"44",X"24",X"0F",X"38",
		X"03",X"21",X"49",X"24",X"46",X"23",X"4E",X"23",X"EB",X"09",X"01",X"20",X"00",X"1A",X"77",X"09",
		X"13",X"1A",X"77",X"13",X"CB",X"DC",X"1A",X"EE",X"80",X"77",X"ED",X"42",X"77",X"C9",X"3A",X"29",
		X"98",X"FE",X"FF",X"28",X"40",X"EB",X"2A",X"2A",X"98",X"ED",X"A0",X"ED",X"A0",X"22",X"2A",X"98",
		X"B7",X"C8",X"47",X"3A",X"2A",X"99",X"F6",X"28",X"6F",X"26",X"99",X"70",X"3E",X"01",X"AD",X"32",
		X"2A",X"99",X"3A",X"08",X"99",X"CD",X"27",X"24",X"21",X"21",X"00",X"19",X"01",X"1F",X"00",X"3E",
		X"FF",X"77",X"2C",X"77",X"09",X"77",X"2C",X"77",X"CB",X"DC",X"3E",X"80",X"77",X"2D",X"77",X"ED",
		X"42",X"77",X"2D",X"77",X"C9",X"CD",X"F2",X"23",X"AF",X"32",X"00",X"9D",X"32",X"03",X"98",X"32",
		X"2C",X"98",X"21",X"01",X"98",X"34",X"C9",X"3D",X"4F",X"E6",X"0F",X"47",X"A9",X"16",X"00",X"87",
		X"CB",X"12",X"87",X"CB",X"12",X"80",X"80",X"5F",X"47",X"FE",X"0F",X"20",X"02",X"CB",X"EB",X"3E",
		X"84",X"B2",X"57",X"C9",X"00",X"21",X"86",X"84",X"00",X"00",X"22",X"84",X"86",X"80",X"00",X"41",
		X"87",X"85",X"80",X"00",X"21",X"85",X"87",X"00",X"3A",X"02",X"99",X"FE",X"0E",X"38",X"02",X"3E",
		X"0A",X"C6",X"02",X"0F",X"0F",X"E6",X"03",X"C8",X"4F",X"06",X"0C",X"11",X"20",X"00",X"21",X"A2",
		X"24",X"DD",X"21",X"40",X"9D",X"7E",X"32",X"80",X"9B",X"D9",X"CD",X"72",X"29",X"3A",X"80",X"9B",
		X"B7",X"28",X"13",X"DD",X"E5",X"E1",X"CD",X"2A",X"28",X"CD",X"31",X"2C",X"38",X"08",X"D9",X"AF",
		X"0D",X"28",X"0B",X"DD",X"19",X"D9",X"D9",X"23",X"10",X"DB",X"AF",X"DD",X"77",X"00",X"32",X"80",
		X"9B",X"C9",X"01",X"0A",X"1B",X"11",X"03",X"19",X"09",X"13",X"02",X"0B",X"1A",X"12",X"3A",X"07",
		X"9D",X"5F",X"16",X"9A",X"1A",X"E6",X"3F",X"C6",X"F0",X"FE",X"FC",X"D8",X"21",X"38",X"99",X"7E",
		X"BB",X"28",X"07",X"73",X"2C",X"36",X"00",X"C3",X"44",X"20",X"2C",X"34",X"7E",X"FE",X"03",X"CA",
		X"3F",X"20",X"FE",X"04",X"D8",X"36",X"00",X"C3",X"B6",X"2D",X"3A",X"08",X"9D",X"21",X"E3",X"24",
		X"E7",X"6E",X"C9",X"03",X"03",X"03",X"03",X"02",X"02",X"01",X"01",X"01",X"01",X"02",X"02",X"AF",
		X"32",X"01",X"9D",X"3A",X"07",X"9D",X"6F",X"26",X"9A",X"7E",X"EB",X"E6",X"3F",X"6F",X"C6",X"F0",
		X"FE",X"FC",X"D4",X"DA",X"24",X"26",X"00",X"29",X"29",X"29",X"01",X"3C",X"45",X"09",X"3A",X"09",
		X"9D",X"FE",X"04",X"20",X"07",X"3A",X"08",X"9D",X"E6",X"03",X"EE",X"02",X"47",X"EE",X"02",X"87",
		X"E7",X"7E",X"FE",X"04",X"20",X"01",X"78",X"EE",X"02",X"87",X"21",X"E0",X"25",X"E7",X"4E",X"23",
		X"46",X"7B",X"E6",X"F0",X"6F",X"AB",X"87",X"87",X"87",X"87",X"67",X"09",X"22",X"02",X"9D",X"22",
		X"04",X"9D",X"3A",X"07",X"9D",X"2A",X"08",X"9D",X"22",X"28",X"98",X"32",X"2A",X"98",X"7D",X"C6",
		X"F0",X"FE",X"FC",X"30",X"04",X"CD",X"24",X"26",X"D8",X"AF",X"32",X"2C",X"98",X"3A",X"07",X"9D",
		X"6F",X"26",X"9A",X"7E",X"B7",X"28",X"5F",X"FE",X"0B",X"28",X"5B",X"CB",X"6F",X"20",X"57",X"C6",
		X"F0",X"FE",X"FC",X"30",X"51",X"7D",X"32",X"07",X"9D",X"7E",X"E6",X"3F",X"EB",X"6F",X"26",X"00",
		X"29",X"29",X"29",X"01",X"3B",X"45",X"09",X"06",X"00",X"7E",X"C6",X"F0",X"FE",X"FC",X"38",X"06",
		X"04",X"23",X"23",X"C3",X"89",X"25",X"78",X"FE",X"04",X"30",X"25",X"4E",X"23",X"46",X"ED",X"43",
		X"08",X"9D",X"87",X"21",X"E0",X"25",X"E7",X"4E",X"23",X"46",X"7B",X"E6",X"F0",X"6F",X"AB",X"87",
		X"87",X"87",X"87",X"67",X"09",X"22",X"02",X"9D",X"22",X"04",X"9D",X"AF",X"32",X"06",X"9D",X"C9",
		X"3A",X"07",X"9D",X"6F",X"26",X"9A",X"D9",X"21",X"2C",X"98",X"7E",X"34",X"E6",X"07",X"21",X"D8",
		X"25",X"E7",X"7E",X"D9",X"85",X"C3",X"60",X"25",X"02",X"DE",X"1E",X"22",X"C2",X"FC",X"40",X"24",
		X"10",X"10",X"20",X"00",X"10",X"F0",X"00",X"00",X"3A",X"07",X"9D",X"2A",X"08",X"9D",X"22",X"28",
		X"98",X"32",X"2A",X"98",X"7D",X"FE",X"0C",X"30",X"09",X"CD",X"24",X"26",X"30",X"04",X"CD",X"24",
		X"26",X"D8",X"3A",X"07",X"9D",X"6F",X"26",X"9A",X"4E",X"EB",X"21",X"00",X"9A",X"3E",X"03",X"06",
		X"00",X"BE",X"28",X"07",X"2C",X"10",X"FA",X"3D",X"20",X"F5",X"C9",X"71",X"12",X"CD",X"0E",X"14",
		X"C9",X"C3",X"E8",X"25",X"ED",X"4B",X"29",X"98",X"79",X"21",X"83",X"35",X"E7",X"7E",X"80",X"32",
		X"2A",X"98",X"6F",X"26",X"9A",X"7E",X"E6",X"3F",X"6F",X"C6",X"F0",X"FE",X"FC",X"30",X"25",X"26",
		X"00",X"29",X"29",X"29",X"11",X"3B",X"45",X"19",X"79",X"FE",X"04",X"20",X"07",X"3A",X"28",X"98",
		X"E6",X"03",X"EE",X"02",X"57",X"87",X"E7",X"4E",X"23",X"46",X"ED",X"43",X"28",X"98",X"3E",X"F0",
		X"81",X"FE",X"FC",X"C9",X"37",X"C9",X"21",X"00",X"00",X"54",X"06",X"08",X"0F",X"30",X"01",X"19",
		X"CB",X"23",X"CB",X"12",X"10",X"F6",X"C9",X"87",X"5F",X"16",X"00",X"30",X"01",X"14",X"21",X"7A",
		X"4D",X"19",X"7E",X"C9",X"87",X"3C",X"5F",X"16",X"00",X"30",X"01",X"14",X"21",X"7A",X"4D",X"19",
		X"7E",X"C9",X"DD",X"66",X"06",X"3A",X"03",X"99",X"57",X"AF",X"06",X"80",X"5F",X"6F",X"ED",X"52",
		X"D0",X"19",X"CB",X"3A",X"CB",X"1B",X"ED",X"52",X"30",X"02",X"B0",X"19",X"CB",X"38",X"30",X"F2",
		X"2F",X"37",X"C9",X"87",X"5F",X"16",X"00",X"30",X"01",X"14",X"21",X"7A",X"4D",X"19",X"5E",X"23",
		X"56",X"63",X"7C",X"AA",X"E6",X"01",X"4F",X"CD",X"99",X"26",X"E6",X"FE",X"B1",X"C9",X"21",X"80",
		X"9B",X"7E",X"B7",X"28",X"09",X"2C",X"7E",X"CF",X"4A",X"29",X"1F",X"27",X"6A",X"27",X"3A",X"07",
		X"98",X"E6",X"0F",X"C0",X"21",X"89",X"9B",X"DF",X"C0",X"CD",X"8F",X"01",X"E6",X"1B",X"6F",X"26",
		X"00",X"22",X"80",X"9B",X"C9",X"1E",X"F3",X"3A",X"02",X"99",X"FE",X"08",X"38",X"04",X"87",X"2F",
		X"83",X"5F",X"3A",X"82",X"9B",X"B7",X"C8",X"CD",X"66",X"26",X"7C",X"32",X"82",X"9B",X"B7",X"CA",
		X"99",X"27",X"FE",X"0A",X"CA",X"5F",X"20",X"C6",X"D8",X"FE",X"FC",X"D8",X"C3",X"5A",X"20",X"CD",
		X"9A",X"28",X"3A",X"07",X"98",X"E6",X"1F",X"CC",X"F5",X"26",X"ED",X"4B",X"85",X"9B",X"ED",X"5B",
		X"02",X"9D",X"78",X"92",X"C6",X"05",X"FE",X"0B",X"D0",X"79",X"93",X"C6",X"05",X"FE",X"0B",X"D0",
		X"3A",X"82",X"9B",X"CD",X"31",X"29",X"78",X"87",X"87",X"87",X"87",X"81",X"47",X"7A",X"87",X"87",
		X"87",X"87",X"4F",X"ED",X"43",X"C9",X"99",X"AF",X"32",X"CB",X"99",X"11",X"00",X"01",X"FF",X"21",
		X"81",X"9B",X"34",X"2D",X"36",X"40",X"CD",X"64",X"20",X"C9",X"21",X"80",X"9B",X"35",X"C2",X"9A",
		X"28",X"21",X"0D",X"99",X"7E",X"34",X"FE",X"07",X"38",X"02",X"3E",X"07",X"21",X"91",X"27",X"E7",
		X"7E",X"32",X"89",X"9B",X"CD",X"64",X"28",X"21",X"00",X"00",X"22",X"80",X"9B",X"CD",X"64",X"20",
		X"C9",X"30",X"20",X"18",X"14",X"10",X"0C",X"0A",X"08",X"E1",X"21",X"71",X"27",X"E5",X"CD",X"8F",
		X"01",X"E6",X"03",X"28",X"0F",X"06",X"04",X"11",X"20",X"00",X"21",X"40",X"9D",X"7E",X"B7",X"28",
		X"79",X"19",X"10",X"F9",X"CD",X"69",X"20",X"3A",X"88",X"9B",X"6F",X"26",X"9A",X"3E",X"01",X"32",
		X"94",X"9C",X"7E",X"08",X"7E",X"0F",X"E6",X"03",X"20",X"02",X"3E",X"04",X"C6",X"20",X"77",X"08",
		X"EB",X"21",X"09",X"99",X"34",X"E6",X"1F",X"FE",X"18",X"38",X"13",X"2C",X"35",X"20",X"0F",X"F5",
		X"D9",X"AF",X"32",X"2C",X"98",X"01",X"08",X"C0",X"ED",X"43",X"01",X"98",X"D9",X"F1",X"E6",X"07",
		X"87",X"21",X"D3",X"36",X"E7",X"7E",X"83",X"4F",X"42",X"08",X"02",X"16",X"07",X"FF",X"43",X"59",
		X"FF",X"60",X"69",X"DD",X"21",X"00",X"9D",X"06",X"06",X"11",X"20",X"00",X"DD",X"7E",X"00",X"0F",
		X"30",X"0B",X"DD",X"7E",X"07",X"BC",X"CC",X"22",X"28",X"BD",X"CC",X"22",X"28",X"DD",X"19",X"10",
		X"EB",X"C9",X"DD",X"34",X"00",X"DD",X"36",X"01",X"04",X"C9",X"3E",X"01",X"77",X"2C",X"77",X"2C",
		X"ED",X"4B",X"85",X"9B",X"71",X"2C",X"70",X"2C",X"71",X"2C",X"70",X"2C",X"36",X"F0",X"2C",X"3A",
		X"87",X"9B",X"57",X"78",X"0F",X"0F",X"0F",X"0F",X"B1",X"CB",X"4A",X"20",X"02",X"D6",X"11",X"77",
		X"2C",X"36",X"00",X"2C",X"7A",X"FE",X"02",X"3E",X"01",X"30",X"01",X"3C",X"77",X"CB",X"D5",X"36",
		X"02",X"C3",X"7D",X"20",X"3A",X"87",X"9B",X"CF",X"70",X"28",X"70",X"28",X"87",X"28",X"87",X"28",
		X"2A",X"85",X"9B",X"11",X"F0",X"EF",X"19",X"7C",X"0F",X"0F",X"0F",X"0F",X"85",X"F5",X"C6",X"02",
		X"CD",X"CD",X"30",X"F1",X"C3",X"CD",X"30",X"2A",X"85",X"9B",X"7C",X"0F",X"0F",X"0F",X"0F",X"85",
		X"F5",X"D6",X"20",X"CD",X"CD",X"30",X"F1",X"C3",X"CD",X"30",X"3A",X"81",X"9B",X"B7",X"C8",X"01",
		X"18",X"00",X"FE",X"02",X"28",X"18",X"3A",X"82",X"9B",X"FE",X"28",X"30",X"02",X"0E",X"0C",X"FE",
		X"0A",X"30",X"02",X"0E",X"04",X"3A",X"07",X"98",X"2F",X"A1",X"20",X"02",X"06",X"04",X"3A",X"87",
		X"9B",X"80",X"CF",X"F7",X"28",X"F7",X"28",X"15",X"29",X"15",X"29",X"D3",X"28",X"D3",X"28",X"D9",
		X"28",X"D9",X"28",X"11",X"FF",X"FF",X"C3",X"DC",X"28",X"11",X"20",X"00",X"2A",X"83",X"9B",X"3E",
		X"10",X"CD",X"F0",X"28",X"7A",X"2F",X"57",X"7B",X"2F",X"5F",X"13",X"19",X"3E",X"88",X"CB",X"DC",
		X"06",X"04",X"77",X"19",X"10",X"FC",X"C9",X"3A",X"82",X"9B",X"CD",X"31",X"29",X"2A",X"83",X"9B",
		X"1E",X"2C",X"78",X"83",X"77",X"2D",X"79",X"83",X"77",X"2D",X"7A",X"83",X"77",X"2D",X"73",X"11",
		X"01",X"00",X"C3",X"EC",X"28",X"3A",X"82",X"9B",X"CD",X"31",X"29",X"2A",X"83",X"9B",X"1E",X"20",
		X"7B",X"70",X"E7",X"71",X"7B",X"E7",X"72",X"7B",X"E7",X"36",X"00",X"11",X"E0",X"FF",X"C3",X"EC",
		X"28",X"01",X"00",X"00",X"D6",X"64",X"38",X"04",X"04",X"C3",X"34",X"29",X"C6",X"64",X"D6",X"0A",
		X"38",X"04",X"0C",X"C3",X"3E",X"29",X"C6",X"0A",X"57",X"C9",X"CD",X"72",X"29",X"11",X"FF",X"80",
		X"E6",X"08",X"20",X"0C",X"D9",X"CD",X"8F",X"01",X"D9",X"E6",X"07",X"20",X"4B",X"11",X"3F",X"30",
		X"D9",X"CD",X"8F",X"01",X"D9",X"A3",X"B2",X"32",X"82",X"9B",X"21",X"81",X"9B",X"34",X"CD",X"7D",
		X"20",X"C9",X"CD",X"DA",X"29",X"38",X"31",X"22",X"83",X"9B",X"3A",X"80",X"9B",X"E6",X"18",X"0F",
		X"0F",X"0F",X"32",X"87",X"9B",X"CD",X"AD",X"29",X"3A",X"87",X"9B",X"ED",X"4B",X"85",X"9B",X"57",
		X"78",X"0F",X"0F",X"0F",X"0F",X"B1",X"CB",X"4A",X"20",X"02",X"D6",X"11",X"6F",X"26",X"9A",X"32",
		X"88",X"9B",X"7E",X"E6",X"18",X"28",X"01",X"C9",X"AF",X"32",X"80",X"9B",X"C9",X"3A",X"87",X"9B",
		X"87",X"21",X"D2",X"29",X"E7",X"5E",X"23",X"56",X"2A",X"83",X"9B",X"19",X"7D",X"87",X"87",X"87",
		X"E6",X"F8",X"57",X"7D",X"CB",X"1C",X"1F",X"CB",X"1C",X"1F",X"E6",X"F8",X"5F",X"ED",X"53",X"85",
		X"9B",X"C9",X"DF",X"FF",X"3F",X"00",X"3F",X"00",X"42",X"00",X"3A",X"80",X"9B",X"CB",X"67",X"20",
		X"38",X"0E",X"00",X"61",X"CB",X"5F",X"20",X"01",X"0C",X"E6",X"07",X"28",X"2A",X"87",X"47",X"3A",
		X"06",X"99",X"57",X"E6",X"F0",X"6F",X"AA",X"B8",X"D8",X"87",X"C6",X"13",X"CB",X"20",X"CB",X"20",
		X"90",X"47",X"29",X"29",X"CB",X"E5",X"EB",X"21",X"F0",X"85",X"CB",X"41",X"28",X"05",X"ED",X"52",
		X"78",X"E7",X"C9",X"19",X"78",X"E7",X"C9",X"37",X"C9",X"0E",X"00",X"61",X"CB",X"5F",X"20",X"01",
		X"0C",X"E6",X"07",X"28",X"F2",X"47",X"3A",X"06",X"99",X"57",X"E6",X"F0",X"6F",X"AA",X"87",X"CB",
		X"41",X"28",X"01",X"2F",X"C6",X"0E",X"4F",X"29",X"29",X"54",X"5D",X"29",X"7C",X"B8",X"D8",X"21",
		X"40",X"85",X"ED",X"52",X"78",X"84",X"67",X"06",X"00",X"09",X"C9",X"3E",X"C0",X"06",X"04",X"11",
		X"20",X"00",X"CB",X"DC",X"77",X"19",X"10",X"FC",X"C9",X"21",X"94",X"9C",X"7E",X"B7",X"C8",X"34",
		X"3D",X"CA",X"4D",X"2E",X"3D",X"28",X"0A",X"D6",X"04",X"C0",X"77",X"3E",X"10",X"32",X"98",X"9C",
		X"C9",X"AF",X"32",X"98",X"9C",X"32",X"93",X"9C",X"3E",X"10",X"32",X"9C",X"9C",X"C9",X"3A",X"07",
		X"98",X"E6",X"03",X"C0",X"3A",X"9D",X"9C",X"B7",X"C0",X"21",X"98",X"9C",X"7E",X"B7",X"C0",X"21",
		X"93",X"9C",X"7E",X"B7",X"FA",X"D5",X"2A",X"C8",X"3A",X"34",X"99",X"B7",X"C0",X"36",X"A1",X"CD",
		X"4D",X"2E",X"3A",X"90",X"9C",X"47",X"3A",X"07",X"9D",X"B8",X"20",X"6F",X"3A",X"92",X"9C",X"32",
		X"99",X"9C",X"3A",X"A0",X"9C",X"6F",X"26",X"9A",X"3A",X"91",X"9C",X"47",X"AE",X"E6",X"3F",X"28",
		X"0F",X"78",X"E6",X"3F",X"C6",X"F0",X"FE",X"FC",X"38",X"50",X"78",X"AE",X"E6",X"3C",X"20",X"4A",
		X"70",X"7D",X"C3",X"CD",X"30",X"34",X"6F",X"7E",X"B7",X"28",X"3A",X"5F",X"16",X"9A",X"1A",X"E6",
		X"3F",X"6F",X"C6",X"F0",X"FE",X"FC",X"30",X"23",X"26",X"00",X"29",X"29",X"E5",X"29",X"01",X"3C",
		X"45",X"09",X"3A",X"99",X"9C",X"4F",X"87",X"E7",X"7E",X"32",X"99",X"9C",X"E1",X"06",X"00",X"09",
		X"01",X"63",X"46",X"09",X"1A",X"B6",X"12",X"7B",X"C3",X"CD",X"30",X"3A",X"99",X"9C",X"C6",X"4C",
		X"12",X"7B",X"CD",X"CD",X"30",X"AF",X"32",X"93",X"9C",X"C9",X"00",X"AF",X"32",X"93",X"9C",X"3E",
		X"10",X"32",X"98",X"9C",X"C9",X"3A",X"09",X"9D",X"EE",X"02",X"C6",X"4C",X"77",X"32",X"91",X"9C",
		X"C3",X"78",X"20",X"21",X"98",X"9C",X"7E",X"B7",X"C8",X"FA",X"9B",X"2B",X"3A",X"00",X"9D",X"0F",
		X"D0",X"3A",X"34",X"99",X"B7",X"C0",X"3E",X"10",X"32",X"93",X"9C",X"36",X"A0",X"2C",X"3A",X"09",
		X"9D",X"77",X"32",X"92",X"9C",X"2C",X"36",X"00",X"EE",X"02",X"47",X"3A",X"07",X"9D",X"32",X"A0",
		X"9C",X"32",X"90",X"9C",X"6F",X"26",X"9A",X"7E",X"E6",X"3F",X"C6",X"F0",X"FE",X"FC",X"30",X"B5",
		X"7E",X"EB",X"87",X"87",X"21",X"63",X"46",X"80",X"E7",X"7E",X"EB",X"B6",X"77",X"32",X"91",X"9C",
		X"7D",X"C9",X"6F",X"26",X"9A",X"7E",X"22",X"96",X"9C",X"32",X"95",X"9C",X"7D",X"CD",X"CD",X"30",
		X"2A",X"96",X"9C",X"3A",X"95",X"9C",X"BE",X"C8",X"C3",X"85",X"2B",X"5E",X"34",X"3A",X"99",X"9C",
		X"21",X"83",X"35",X"E7",X"16",X"9C",X"1A",X"86",X"13",X"12",X"5F",X"16",X"9A",X"1A",X"E6",X"3F",
		X"6F",X"C6",X"F0",X"FE",X"FC",X"30",X"4C",X"26",X"00",X"29",X"29",X"E5",X"29",X"01",X"3B",X"45",
		X"09",X"3A",X"99",X"9C",X"4F",X"87",X"E7",X"7E",X"C6",X"F0",X"FE",X"FC",X"30",X"2A",X"23",X"7E",
		X"32",X"99",X"9C",X"E1",X"06",X"00",X"09",X"01",X"63",X"46",X"09",X"1A",X"B6",X"EB",X"BE",X"20",
		X"14",X"3A",X"A0",X"9C",X"BD",X"20",X"0F",X"21",X"98",X"9C",X"5E",X"16",X"9C",X"AF",X"12",X"77",
		X"2C",X"2C",X"36",X"01",X"C9",X"77",X"7D",X"C9",X"E1",X"21",X"98",X"9C",X"5E",X"16",X"9C",X"AF",
		X"12",X"77",X"C9",X"1A",X"FE",X"40",X"38",X"1E",X"21",X"38",X"99",X"7B",X"BE",X"20",X"13",X"2C",
		X"34",X"7E",X"D6",X"03",X"38",X"10",X"01",X"3F",X"20",X"28",X"03",X"01",X"B6",X"2D",X"C5",X"28",
		X"05",X"2D",X"73",X"2C",X"36",X"00",X"3A",X"99",X"9C",X"C6",X"4C",X"12",X"AF",X"32",X"98",X"9C",
		X"C9",X"3A",X"07",X"9D",X"47",X"DD",X"7E",X"07",X"B8",X"28",X"4A",X"DD",X"66",X"09",X"32",X"30",
		X"98",X"22",X"31",X"98",X"CD",X"56",X"2C",X"D8",X"C6",X"F0",X"FE",X"FC",X"D0",X"CD",X"56",X"2C",
		X"D8",X"C6",X"F0",X"FE",X"FC",X"D0",X"3A",X"32",X"98",X"21",X"83",X"35",X"E7",X"3A",X"30",X"98",
		X"86",X"32",X"30",X"98",X"B8",X"28",X"1E",X"6F",X"26",X"9A",X"7E",X"E6",X"3F",X"6F",X"26",X"00",
		X"29",X"29",X"29",X"11",X"3B",X"45",X"19",X"3A",X"32",X"98",X"87",X"E7",X"7E",X"23",X"4E",X"ED",
		X"43",X"32",X"98",X"B7",X"C9",X"37",X"C9",X"21",X"9D",X"9C",X"7E",X"B7",X"C8",X"3A",X"9A",X"9C",
		X"B7",X"20",X"51",X"21",X"A0",X"9C",X"7E",X"B7",X"28",X"45",X"5F",X"16",X"9A",X"1A",X"87",X"87",
		X"47",X"3A",X"9E",X"9C",X"EE",X"02",X"80",X"21",X"63",X"46",X"E7",X"7E",X"2F",X"EB",X"A6",X"77",
		X"7D",X"CD",X"82",X"2B",X"21",X"98",X"9C",X"DF",X"2E",X"9C",X"DF",X"2E",X"93",X"DF",X"21",X"A0",
		X"9C",X"11",X"9F",X"9C",X"01",X"60",X"00",X"ED",X"B0",X"EB",X"70",X"3A",X"9B",X"9C",X"FE",X"04",
		X"30",X"02",X"3E",X"04",X"32",X"9B",X"9C",X"3A",X"39",X"99",X"FE",X"03",X"C4",X"44",X"20",X"21",
		X"9D",X"9C",X"35",X"C9",X"21",X"98",X"9C",X"DF",X"2E",X"9C",X"DF",X"2E",X"93",X"DF",X"21",X"A0",
		X"9C",X"11",X"9F",X"9C",X"ED",X"A0",X"1A",X"08",X"ED",X"A0",X"7E",X"B7",X"20",X"FA",X"08",X"12",
		X"21",X"9D",X"9C",X"35",X"21",X"9B",X"9C",X"DF",X"CA",X"98",X"2D",X"7E",X"FE",X"03",X"C0",X"CD",
		X"3F",X"20",X"3A",X"20",X"9D",X"B7",X"C0",X"ED",X"4B",X"A3",X"9C",X"78",X"B7",X"20",X"04",X"3A",
		X"A0",X"9C",X"47",X"91",X"38",X"17",X"D6",X"02",X"20",X"08",X"0E",X"02",X"11",X"10",X"F0",X"C3",
		X"51",X"2D",X"D6",X"1E",X"C0",X"0E",X"03",X"11",X"00",X"00",X"C3",X"51",X"2D",X"C6",X"02",X"20",
		X"08",X"0E",X"00",X"11",X"10",X"10",X"C3",X"51",X"2D",X"C6",X"1E",X"C0",X"0E",X"01",X"11",X"20",
		X"00",X"78",X"E6",X"F0",X"6F",X"A8",X"87",X"87",X"87",X"87",X"67",X"19",X"22",X"22",X"9D",X"22",
		X"24",X"9D",X"ED",X"43",X"26",X"9D",X"68",X"26",X"9A",X"7E",X"E6",X"3F",X"6F",X"26",X"00",X"29",
		X"29",X"29",X"11",X"3B",X"45",X"19",X"79",X"87",X"E7",X"5E",X"23",X"56",X"ED",X"53",X"28",X"9D",
		X"21",X"8F",X"34",X"22",X"2A",X"9D",X"21",X"02",X"01",X"22",X"20",X"9D",X"21",X"D4",X"07",X"22",
		X"2C",X"9D",X"3E",X"01",X"32",X"2E",X"9D",X"C9",X"3A",X"20",X"9D",X"0F",X"30",X"12",X"21",X"A0",
		X"9C",X"06",X"60",X"3A",X"27",X"9D",X"4F",X"7E",X"B7",X"28",X"05",X"B9",X"C8",X"2C",X"10",X"F7",
		X"3A",X"0C",X"99",X"32",X"9B",X"9C",X"ED",X"4B",X"A0",X"9C",X"78",X"91",X"38",X"17",X"D6",X"02",
		X"20",X"08",X"0E",X"02",X"11",X"10",X"F0",X"C3",X"E9",X"2D",X"D6",X"1E",X"C0",X"0E",X"03",X"11",
		X"00",X"00",X"C3",X"E9",X"2D",X"C6",X"02",X"20",X"08",X"0E",X"00",X"11",X"10",X"10",X"C3",X"E9",
		X"2D",X"C6",X"1E",X"C0",X"0E",X"01",X"11",X"20",X"00",X"78",X"E6",X"F0",X"6F",X"A8",X"87",X"87",
		X"87",X"87",X"67",X"19",X"22",X"22",X"9D",X"22",X"24",X"9D",X"ED",X"43",X"26",X"9D",X"68",X"26",
		X"9A",X"7E",X"E6",X"3F",X"6F",X"26",X"00",X"29",X"29",X"29",X"11",X"3B",X"45",X"19",X"79",X"87",
		X"E7",X"5E",X"23",X"56",X"ED",X"53",X"28",X"9D",X"21",X"8F",X"34",X"22",X"2A",X"9D",X"21",X"01",
		X"03",X"22",X"20",X"9D",X"3E",X"01",X"32",X"2E",X"9D",X"CD",X"44",X"20",X"C3",X"49",X"20",X"21",
		X"9C",X"9C",X"7E",X"B7",X"C8",X"FA",X"3A",X"2E",X"36",X"9F",X"34",X"6E",X"7E",X"B7",X"C8",X"36",
		X"00",X"5F",X"16",X"9A",X"1A",X"B7",X"C8",X"7B",X"C3",X"82",X"2B",X"77",X"C9",X"AF",X"32",X"98",
		X"9C",X"06",X"3F",X"26",X"9A",X"11",X"A0",X"9C",X"1A",X"B7",X"C8",X"6F",X"7E",X"A0",X"77",X"1C",
		X"20",X"F6",X"C9",X"DD",X"21",X"00",X"9E",X"3A",X"00",X"9E",X"B7",X"28",X"08",X"3A",X"01",X"9E",
		X"CF",X"75",X"2E",X"C2",X"2E",X"21",X"1F",X"9E",X"DF",X"C0",X"C9",X"DD",X"21",X"00",X"9E",X"DD",
		X"36",X"00",X"01",X"DD",X"36",X"01",X"01",X"3A",X"0C",X"9D",X"D6",X"C0",X"0F",X"0F",X"E6",X"0F",
		X"21",X"B4",X"30",X"E7",X"11",X"74",X"30",X"3A",X"0E",X"98",X"B7",X"28",X"03",X"11",X"94",X"30",
		X"7E",X"DD",X"77",X"04",X"EB",X"E7",X"11",X"1A",X"9E",X"01",X"06",X"00",X"ED",X"B0",X"56",X"23",
		X"5E",X"2A",X"02",X"9D",X"19",X"22",X"02",X"9E",X"AF",X"DD",X"77",X"05",X"3C",X"DD",X"77",X"06",
		X"C9",X"C9",X"DD",X"35",X"06",X"C0",X"06",X"06",X"DD",X"70",X"06",X"D9",X"DD",X"34",X"05",X"DD",
		X"7E",X"05",X"21",X"11",X"2F",X"E7",X"7E",X"B7",X"FA",X"0D",X"2F",X"87",X"87",X"4F",X"87",X"81",
		X"4F",X"06",X"00",X"DD",X"7E",X"04",X"0F",X"0F",X"21",X"1C",X"2F",X"E7",X"5E",X"23",X"56",X"EB",
		X"09",X"ED",X"4B",X"02",X"9E",X"11",X"0E",X"9E",X"CD",X"FF",X"2E",X"3A",X"03",X"9E",X"4F",X"06",
		X"06",X"7E",X"FE",X"FF",X"28",X"01",X"81",X"12",X"23",X"1C",X"10",X"F5",X"C9",X"DD",X"36",X"00",
		X"00",X"C9",X"00",X"01",X"02",X"03",X"02",X"03",X"04",X"05",X"06",X"FF",X"24",X"2F",X"78",X"2F",
		X"CC",X"2F",X"20",X"30",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"02",X"FF",X"FF",X"00",X"02",X"00",X"00",X"FF",X"FF",X"FD",X"FD",X"00",X"03",X"00",X"03",
		X"00",X"03",X"00",X"00",X"FD",X"FD",X"FA",X"FA",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"00",
		X"FC",X"FC",X"F8",X"F8",X"01",X"04",X"01",X"04",X"01",X"04",X"FE",X"FE",X"FB",X"FB",X"F8",X"F8",
		X"02",X"04",X"FF",X"FF",X"02",X"04",X"FC",X"FC",X"FF",X"FF",X"F9",X"F9",X"03",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"FF",X"FF",X"00",X"02",X"00",X"00",X"FF",X"FF",X"03",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"03",X"03",X"06",X"06",X"00",X"04",X"00",X"04",
		X"00",X"04",X"00",X"00",X"04",X"04",X"08",X"08",X"01",X"04",X"01",X"04",X"01",X"04",X"02",X"02",
		X"05",X"05",X"08",X"08",X"02",X"04",X"FF",X"FF",X"02",X"04",X"04",X"04",X"FF",X"FF",X"07",X"07",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FD",X"FD",X"00",X"02",
		X"FF",X"FF",X"00",X"02",X"00",X"00",X"FD",X"FD",X"FA",X"FA",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"FC",X"FC",X"F8",X"F8",X"00",X"04",X"00",X"04",X"00",X"04",X"FE",X"FE",X"FB",X"FB",
		X"F8",X"F8",X"01",X"04",X"01",X"04",X"01",X"04",X"FC",X"FC",X"FF",X"FF",X"F9",X"F9",X"02",X"04",
		X"02",X"04",X"02",X"04",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"03",X"03",X"00",X"02",X"FF",X"FF",X"00",X"02",X"00",X"00",X"03",X"03",X"06",X"06",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"00",X"04",X"04",X"08",X"08",X"00",X"04",X"00",X"04",X"00",X"04",
		X"02",X"02",X"05",X"05",X"08",X"08",X"01",X"04",X"01",X"04",X"01",X"04",X"04",X"04",X"FF",X"FF",
		X"07",X"07",X"02",X"04",X"02",X"04",X"02",X"04",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0B",X"0E",X"0C",X"0D",X"0C",X"0A",X"07",X"06",X"09",X"0A",X"0C",X"0D",
		X"0C",X"0E",X"FE",X"08",X"0F",X"0E",X"0F",X"0D",X"0C",X"0B",X"0B",X"03",X"0A",X"09",X"0F",X"0D",
		X"0A",X"0E",X"0B",X"FA",X"0E",X"0C",X"0A",X"0D",X"0E",X"09",X"06",X"08",X"0A",X"09",X"0E",X"0F",
		X"0A",X"0C",X"FC",X"07",X"0E",X"08",X"0F",X"0A",X"0E",X"0A",X"07",X"05",X"09",X"0A",X"0E",X"0A",
		X"09",X"0B",X"08",X"FA",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",
		X"08",X"08",X"08",X"08",X"11",X"FE",X"83",X"3A",X"00",X"9A",X"C3",X"F0",X"30",X"B7",X"28",X"F4",
		X"6F",X"26",X"9A",X"3D",X"4F",X"E6",X"0F",X"47",X"A9",X"16",X"00",X"87",X"CB",X"12",X"87",X"CB",
		X"12",X"80",X"80",X"5F",X"78",X"FE",X"0F",X"20",X"02",X"CB",X"EB",X"3E",X"84",X"B2",X"57",X"7E",
		X"6F",X"26",X"00",X"29",X"29",X"7C",X"E5",X"87",X"21",X"73",X"3C",X"E7",X"4E",X"23",X"46",X"E1",
		X"29",X"29",X"3E",X"03",X"A4",X"20",X"21",X"29",X"09",X"3E",X"04",X"CD",X"16",X"31",X"EB",X"01",
		X"80",X"07",X"09",X"EB",X"3E",X"04",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"EB",X"01",
		X"1C",X"00",X"09",X"EB",X"3D",X"20",X"EF",X"C9",X"3D",X"28",X"3A",X"7D",X"B7",X"28",X"06",X"2E",
		X"00",X"87",X"C3",X"66",X"31",X"29",X"09",X"13",X"13",X"23",X"23",X"CB",X"63",X"28",X"04",X"1B",
		X"1B",X"2B",X"2B",X"CB",X"4A",X"20",X"0A",X"01",X"08",X"00",X"09",X"EB",X"01",X"40",X"00",X"09",
		X"EB",X"3E",X"02",X"CD",X"A8",X"31",X"01",X"08",X"00",X"09",X"EB",X"01",X"C0",X"07",X"09",X"EB",
		X"3E",X"02",X"C3",X"A8",X"31",X"7D",X"29",X"09",X"D9",X"07",X"07",X"07",X"E6",X"03",X"CF",X"77",
		X"31",X"96",X"31",X"9A",X"31",X"B8",X"31",X"D9",X"01",X"08",X"00",X"09",X"01",X"40",X"00",X"EB",
		X"09",X"EB",X"3E",X"02",X"CD",X"16",X"31",X"01",X"08",X"00",X"09",X"EB",X"01",X"C0",X"07",X"09",
		X"EB",X"3E",X"02",X"C3",X"16",X"31",X"D9",X"C3",X"82",X"31",X"D9",X"3E",X"04",X"CD",X"A8",X"31",
		X"EB",X"01",X"80",X"07",X"09",X"EB",X"3E",X"04",X"ED",X"A0",X"ED",X"A0",X"23",X"23",X"EB",X"01",
		X"1E",X"00",X"09",X"EB",X"3D",X"20",X"F1",X"C9",X"D9",X"23",X"23",X"13",X"13",X"C3",X"9B",X"31",
		X"3A",X"35",X"99",X"CB",X"4F",X"0E",X"05",X"20",X"01",X"0D",X"21",X"2C",X"99",X"06",X"04",X"D9",
		X"21",X"07",X"9D",X"11",X"20",X"00",X"06",X"06",X"3A",X"36",X"99",X"4F",X"3A",X"08",X"99",X"BE",
		X"20",X"0B",X"08",X"71",X"7D",X"D9",X"91",X"77",X"2C",X"05",X"C8",X"D9",X"08",X"19",X"10",X"EF",
		X"D9",X"36",X"00",X"C9",X"3A",X"08",X"99",X"5F",X"D6",X"02",X"0E",X"01",X"C3",X"41",X"32",X"3A",
		X"08",X"99",X"5F",X"D6",X"20",X"0E",X"02",X"C3",X"41",X"32",X"3A",X"08",X"99",X"5F",X"C6",X"20",
		X"0E",X"03",X"C3",X"41",X"32",X"3A",X"2B",X"99",X"F6",X"28",X"6F",X"26",X"99",X"7E",X"B7",X"C8",
		X"36",X"00",X"08",X"7D",X"EE",X"01",X"32",X"2B",X"99",X"08",X"0F",X"38",X"C7",X"0F",X"38",X"09",
		X"0F",X"0F",X"0F",X"38",X"CA",X"0F",X"38",X"D2",X"C9",X"3A",X"08",X"99",X"5F",X"C6",X"02",X"0E",
		X"00",X"6F",X"26",X"9A",X"54",X"7E",X"E6",X"3F",X"FE",X"10",X"D0",X"32",X"37",X"99",X"3E",X"01",
		X"32",X"94",X"9C",X"D9",X"CD",X"4D",X"2E",X"D9",X"36",X"00",X"43",X"ED",X"43",X"35",X"99",X"7D",
		X"32",X"08",X"99",X"CD",X"87",X"20",X"CD",X"C0",X"31",X"3E",X"04",X"C3",X"74",X"32",X"3A",X"34",
		X"99",X"B7",X"28",X"A1",X"3D",X"32",X"34",X"99",X"47",X"D9",X"CC",X"B3",X"32",X"CD",X"90",X"32",
		X"D9",X"CD",X"32",X"33",X"3A",X"35",X"99",X"CF",X"CF",X"32",X"EF",X"32",X"FB",X"32",X"1F",X"33",
		X"21",X"AF",X"32",X"3A",X"35",X"99",X"E7",X"4E",X"11",X"2C",X"99",X"06",X"04",X"26",X"9D",X"1A",
		X"B7",X"C8",X"6F",X"7E",X"81",X"77",X"2C",X"2C",X"7E",X"81",X"77",X"1C",X"10",X"F1",X"C9",X"F8",
		X"08",X"08",X"F8",X"2A",X"36",X"99",X"7C",X"B7",X"C8",X"26",X"9A",X"77",X"ED",X"4B",X"38",X"99",
		X"78",X"BD",X"C0",X"79",X"FE",X"03",X"C0",X"3D",X"32",X"39",X"99",X"C3",X"44",X"20",X"C9",X"D9",
		X"68",X"26",X"00",X"19",X"E5",X"11",X"04",X"00",X"19",X"3E",X"FF",X"06",X"04",X"11",X"20",X"00",
		X"CB",X"DC",X"36",X"80",X"CB",X"9C",X"77",X"19",X"10",X"F6",X"D1",X"79",X"C3",X"F0",X"30",X"D9",
		X"78",X"ED",X"44",X"83",X"6F",X"62",X"E5",X"2B",X"C3",X"D9",X"32",X"D9",X"EB",X"11",X"E0",X"FF",
		X"AF",X"B0",X"28",X"03",X"19",X"10",X"FD",X"E5",X"19",X"3E",X"FF",X"06",X"04",X"11",X"01",X"00",
		X"CB",X"DC",X"36",X"80",X"CB",X"9C",X"77",X"19",X"10",X"F6",X"D1",X"79",X"C3",X"F0",X"30",X"D9",
		X"EB",X"11",X"20",X"00",X"AF",X"B0",X"28",X"03",X"19",X"10",X"FD",X"E5",X"1E",X"80",X"19",X"C3",
		X"09",X"33",X"2A",X"36",X"99",X"4C",X"7D",X"3D",X"57",X"E6",X"0F",X"67",X"AA",X"16",X"00",X"87",
		X"CB",X"12",X"87",X"CB",X"12",X"84",X"84",X"5F",X"7C",X"FE",X"0F",X"20",X"02",X"CB",X"EB",X"3E",
		X"84",X"B2",X"57",X"D9",X"C9",X"26",X"00",X"11",X"96",X"33",X"3A",X"0D",X"9D",X"DD",X"BE",X"0D",
		X"28",X"03",X"11",X"7E",X"33",X"DD",X"7E",X"1F",X"C6",X"08",X"0F",X"0F",X"0F",X"0F",X"84",X"E6",
		X"0F",X"DD",X"AE",X"11",X"EB",X"E7",X"7E",X"DD",X"86",X"0F",X"DD",X"77",X"0C",X"C9",X"00",X"1E",
		X"1A",X"16",X"12",X"0E",X"0A",X"06",X"02",X"1C",X"18",X"14",X"10",X"0C",X"08",X"04",X"00",X"1E",
		X"1A",X"16",X"12",X"0E",X"0A",X"06",X"00",X"3C",X"38",X"34",X"30",X"2C",X"28",X"24",X"20",X"1C",
		X"18",X"14",X"10",X"0C",X"08",X"04",X"00",X"3C",X"38",X"34",X"30",X"2C",X"28",X"24",X"3A",X"00",
		X"9D",X"0F",X"30",X"06",X"CD",X"A5",X"3A",X"CD",X"6E",X"32",X"CD",X"A7",X"34",X"CD",X"63",X"2E",
		X"C9",X"DD",X"7E",X"06",X"C6",X"04",X"DD",X"77",X"06",X"C9",X"3A",X"0D",X"9D",X"DD",X"BE",X"0D",
		X"20",X"EF",X"3A",X"06",X"9D",X"32",X"33",X"99",X"3A",X"3B",X"99",X"CB",X"5F",X"28",X"24",X"ED",
		X"4B",X"30",X"99",X"3E",X"04",X"81",X"4F",X"30",X"09",X"04",X"3E",X"03",X"B8",X"30",X"03",X"01",
		X"FF",X"03",X"ED",X"43",X"30",X"99",X"2A",X"32",X"99",X"04",X"09",X"22",X"32",X"99",X"7C",X"32",
		X"06",X"9D",X"C9",X"ED",X"4B",X"30",X"99",X"3E",X"F8",X"81",X"4F",X"38",X"E5",X"05",X"78",X"3C",
		X"20",X"E0",X"01",X"00",X"00",X"C3",X"F2",X"33",X"3A",X"20",X"9D",X"B7",X"C8",X"3A",X"21",X"9D",
		X"CF",X"2D",X"34",X"2D",X"34",X"52",X"34",X"52",X"34",X"6D",X"34",X"81",X"34",X"3A",X"9B",X"9C",
		X"FE",X"04",X"38",X"07",X"21",X"00",X"00",X"22",X"20",X"9D",X"C9",X"06",X"0C",X"3D",X"20",X"02",
		X"06",X"04",X"2A",X"24",X"9D",X"3A",X"07",X"98",X"A0",X"28",X"03",X"21",X"00",X"00",X"22",X"22",
		X"9D",X"C9",X"3A",X"26",X"9D",X"C6",X"09",X"32",X"26",X"9D",X"3A",X"2C",X"9D",X"32",X"3D",X"9D",
		X"CD",X"36",X"35",X"3A",X"3D",X"9D",X"32",X"2C",X"9D",X"CD",X"C4",X"3A",X"C9",X"CD",X"53",X"20",
		X"21",X"9B",X"34",X"22",X"2A",X"9D",X"DD",X"36",X"0E",X"01",X"DD",X"36",X"10",X"40",X"DD",X"34",
		X"01",X"CD",X"C4",X"3A",X"DD",X"35",X"10",X"C0",X"21",X"00",X"00",X"22",X"20",X"9D",X"C9",X"D4",
		X"04",X"02",X"D0",X"04",X"02",X"CC",X"04",X"02",X"FF",X"8F",X"34",X"D4",X"05",X"01",X"D0",X"06",
		X"01",X"CC",X"07",X"01",X"FF",X"9B",X"34",X"DD",X"21",X"00",X"9D",X"CD",X"D6",X"34",X"DD",X"21",
		X"20",X"9D",X"CD",X"18",X"34",X"11",X"20",X"00",X"DD",X"19",X"3A",X"07",X"98",X"0F",X"30",X"02",
		X"DD",X"19",X"06",X"02",X"1E",X"40",X"DD",X"7E",X"00",X"B7",X"28",X"05",X"D9",X"CD",X"D6",X"34",
		X"D9",X"DD",X"19",X"10",X"F1",X"C9",X"DD",X"7E",X"01",X"CF",X"33",X"35",X"33",X"35",X"33",X"35",
		X"33",X"35",X"E6",X"34",X"06",X"35",X"3A",X"0D",X"9D",X"DD",X"BE",X"0D",X"21",X"15",X"35",X"28",
		X"03",X"21",X"24",X"35",X"11",X"40",X"01",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"72",X"0E",
		X"DD",X"73",X"10",X"DD",X"34",X"01",X"CD",X"C4",X"3A",X"DD",X"35",X"10",X"C0",X"AF",X"DD",X"77",
		X"00",X"DD",X"77",X"01",X"C9",X"C1",X"08",X"04",X"D1",X"04",X"04",X"E1",X"0C",X"04",X"F1",X"10",
		X"04",X"FF",X"15",X"35",X"91",X"07",X"03",X"81",X"08",X"03",X"93",X"09",X"03",X"83",X"1A",X"03",
		X"FF",X"24",X"35",X"CD",X"CA",X"33",X"3A",X"03",X"99",X"3D",X"DD",X"BE",X"06",X"38",X"59",X"DD",
		X"7E",X"08",X"CF",X"E2",X"36",X"EC",X"36",X"F8",X"36",X"02",X"37",X"0E",X"37",X"2A",X"37",X"48",
		X"37",X"66",X"37",X"82",X"37",X"9E",X"37",X"BC",X"37",X"D8",X"37",X"F6",X"37",X"F6",X"37",X"F6",
		X"37",X"F6",X"37",X"0E",X"38",X"2D",X"38",X"4C",X"38",X"6D",X"38",X"8E",X"38",X"AF",X"38",X"D0",
		X"38",X"EF",X"38",X"0E",X"39",X"2D",X"39",X"4C",X"39",X"6D",X"39",X"8E",X"39",X"AD",X"39",X"CC",
		X"39",X"ED",X"39",X"FE",X"E0",X"02",X"20",X"00",X"3A",X"34",X"99",X"B7",X"C8",X"3A",X"36",X"99",
		X"95",X"3E",X"00",X"C0",X"3A",X"37",X"99",X"C9",X"3A",X"34",X"99",X"B7",X"28",X"14",X"3A",X"36",
		X"99",X"DD",X"BE",X"07",X"20",X"0C",X"DD",X"7E",X"02",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"C3",
		X"C3",X"35",X"DD",X"7E",X"02",X"C6",X"06",X"E6",X"F0",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"C6",
		X"06",X"E6",X"F0",X"DD",X"77",X"05",X"DD",X"7E",X"09",X"21",X"83",X"35",X"E7",X"7E",X"DD",X"4E",
		X"07",X"81",X"DD",X"77",X"07",X"6F",X"26",X"9A",X"7E",X"E6",X"3F",X"CC",X"88",X"35",X"6F",X"C6",
		X"F0",X"FE",X"FC",X"D4",X"B5",X"36",X"26",X"00",X"29",X"29",X"29",X"11",X"3B",X"45",X"19",X"DD",
		X"7E",X"09",X"FE",X"04",X"20",X"05",X"DD",X"7E",X"08",X"E6",X"03",X"57",X"87",X"E7",X"46",X"23",
		X"DD",X"7E",X"08",X"C6",X"F0",X"38",X"11",X"A0",X"C6",X"F0",X"FE",X"FC",X"38",X"0A",X"DD",X"34",
		X"00",X"DD",X"36",X"01",X"04",X"C3",X"69",X"20",X"DD",X"70",X"08",X"7E",X"DD",X"77",X"09",X"DD",
		X"36",X"06",X"00",X"FE",X"04",X"20",X"03",X"DD",X"71",X"07",X"3A",X"2D",X"9D",X"DD",X"BE",X"0D",
		X"C8",X"3A",X"0D",X"9D",X"DD",X"BE",X"0D",X"20",X"75",X"D9",X"11",X"01",X"01",X"FF",X"D9",X"21",
		X"9D",X"9C",X"34",X"7A",X"2C",X"77",X"DD",X"7E",X"08",X"C6",X"F0",X"30",X"55",X"DD",X"6E",X"07",
		X"26",X"9A",X"7E",X"E6",X"3F",X"FE",X"18",X"D8",X"E6",X"07",X"87",X"EB",X"21",X"D2",X"36",X"E7",
		X"3A",X"08",X"9D",X"BE",X"C0",X"1A",X"D6",X"08",X"12",X"23",X"6E",X"26",X"00",X"CB",X"7D",X"28",
		X"01",X"25",X"19",X"7E",X"D6",X"08",X"77",X"16",X"07",X"45",X"FF",X"58",X"FF",X"CD",X"82",X"20",
		X"CD",X"7B",X"2E",X"11",X"0A",X"01",X"FF",X"21",X"09",X"99",X"35",X"2C",X"35",X"C0",X"AF",X"32",
		X"2C",X"98",X"01",X"08",X"C0",X"ED",X"43",X"01",X"98",X"21",X"80",X"9B",X"7E",X"B7",X"C8",X"36",
		X"01",X"C9",X"FE",X"FC",X"D8",X"21",X"02",X"04",X"22",X"00",X"9D",X"C3",X"30",X"20",X"CD",X"31",
		X"2C",X"D0",X"C3",X"7D",X"20",X"3A",X"0D",X"9D",X"DD",X"BE",X"0D",X"20",X"0C",X"11",X"0F",X"01",
		X"FF",X"CD",X"78",X"20",X"3E",X"01",X"32",X"94",X"9C",X"CD",X"8F",X"01",X"E6",X"03",X"28",X"F9",
		X"6F",X"C9",X"1D",X"FE",X"15",X"02",X"1B",X"FE",X"11",X"02",X"1E",X"20",X"18",X"E0",X"16",X"20",
		X"12",X"E0",X"CD",X"20",X"3A",X"DD",X"86",X"05",X"DD",X"77",X"03",X"C9",X"CD",X"20",X"3A",X"ED",
		X"44",X"DD",X"86",X"05",X"DD",X"77",X"03",X"C9",X"CD",X"20",X"3A",X"DD",X"86",X"04",X"DD",X"77",
		X"02",X"C9",X"CD",X"20",X"3A",X"ED",X"44",X"DD",X"86",X"04",X"DD",X"77",X"02",X"C9",X"CD",X"92",
		X"26",X"01",X"00",X"40",X"CD",X"37",X"3A",X"CD",X"6D",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"02",
		X"CD",X"96",X"3A",X"DD",X"74",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",X"01",X"01",X"40",
		X"CD",X"37",X"3A",X"CD",X"6D",X"3A",X"DD",X"74",X"02",X"CD",X"96",X"3A",X"7C",X"C6",X"10",X"DD",
		X"77",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",X"26",X"01",X"01",X"80",X"CD",X"37",
		X"3A",X"CD",X"7A",X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"02",X"CD",X"96",X"3A",X"DD",X"74",X"03",
		X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",X"26",X"01",X"00",X"80",X"CD",X"37",X"3A",X"CD",
		X"7A",X"3A",X"DD",X"74",X"02",X"CD",X"96",X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"03",X"CD",X"55",
		X"33",X"C9",X"CD",X"92",X"26",X"01",X"00",X"00",X"CD",X"37",X"3A",X"CD",X"6D",X"3A",X"DD",X"74",
		X"02",X"CD",X"89",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",
		X"26",X"01",X"01",X"00",X"CD",X"37",X"3A",X"CD",X"6D",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"02",
		X"CD",X"89",X"3A",X"DD",X"74",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",X"26",X"01",
		X"00",X"C0",X"CD",X"37",X"3A",X"CD",X"7A",X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"02",X"CD",X"89",
		X"3A",X"DD",X"74",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",X"01",X"01",X"C0",X"CD",X"37",
		X"3A",X"CD",X"7A",X"3A",X"DD",X"74",X"02",X"CD",X"89",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"03",
		X"26",X"08",X"CD",X"57",X"33",X"C9",X"DD",X"34",X"06",X"DD",X"34",X"06",X"3A",X"03",X"99",X"D6",
		X"02",X"DD",X"BE",X"06",X"D0",X"3E",X"08",X"DD",X"AE",X"11",X"DD",X"77",X"11",X"C9",X"CD",X"92",
		X"26",X"01",X"00",X"40",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"6D",X"3A",X"7C",X"D6",X"10",
		X"DD",X"77",X"02",X"CD",X"96",X"3A",X"DD",X"74",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",
		X"01",X"00",X"40",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"6D",X"3A",X"7C",X"D6",X"10",X"DD",
		X"77",X"02",X"CD",X"96",X"3A",X"DD",X"74",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",X"01",
		X"01",X"40",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"6D",X"3A",X"DD",X"74",X"02",X"CD",X"96",
		X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",X"26",
		X"01",X"01",X"40",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"6D",X"3A",X"DD",X"74",X"02",X"CD",
		X"96",X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",
		X"26",X"01",X"01",X"80",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"7A",X"3A",X"7C",X"C6",X"10",
		X"DD",X"77",X"02",X"CD",X"96",X"3A",X"DD",X"74",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",
		X"92",X"26",X"01",X"01",X"80",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"7A",X"3A",X"7C",X"C6",
		X"10",X"DD",X"77",X"02",X"CD",X"96",X"3A",X"DD",X"74",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",
		X"CD",X"92",X"26",X"01",X"00",X"80",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"7A",X"3A",X"DD",
		X"74",X"02",X"CD",X"96",X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"03",X"CD",X"55",X"33",X"C9",X"CD",
		X"92",X"26",X"01",X"00",X"80",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"7A",X"3A",X"DD",X"74",
		X"02",X"CD",X"96",X"3A",X"7C",X"C6",X"10",X"DD",X"77",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",
		X"26",X"01",X"00",X"00",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"6D",X"3A",X"DD",X"74",X"02",
		X"CD",X"89",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",
		X"01",X"00",X"00",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"6D",X"3A",X"DD",X"74",X"02",X"CD",
		X"89",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",X"01",
		X"01",X"00",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"6D",X"3A",X"7C",X"D6",X"10",X"DD",X"77",
		X"02",X"CD",X"89",X"3A",X"DD",X"74",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",X"26",
		X"01",X"01",X"00",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"6D",X"3A",X"7C",X"D6",X"10",X"DD",
		X"77",X"02",X"CD",X"89",X"3A",X"DD",X"74",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",
		X"26",X"01",X"00",X"C0",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"7A",X"3A",X"7C",X"C6",X"10",
		X"DD",X"77",X"02",X"CD",X"89",X"3A",X"DD",X"74",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",
		X"01",X"00",X"C0",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"7A",X"3A",X"7C",X"C6",X"10",X"DD",
		X"77",X"02",X"CD",X"89",X"3A",X"DD",X"74",X"03",X"CD",X"55",X"33",X"C9",X"CD",X"92",X"26",X"01",
		X"01",X"C0",X"CD",X"37",X"3A",X"CD",X"0E",X"3A",X"CD",X"7A",X"3A",X"DD",X"74",X"02",X"CD",X"89",
		X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"CD",X"92",X"26",
		X"01",X"01",X"C0",X"CD",X"37",X"3A",X"CD",X"17",X"3A",X"CD",X"7A",X"3A",X"DD",X"74",X"02",X"CD",
		X"89",X"3A",X"7C",X"D6",X"10",X"DD",X"77",X"03",X"26",X"08",X"CD",X"57",X"33",X"C9",X"21",X"00",
		X"FD",X"19",X"D0",X"11",X"00",X"03",X"C9",X"21",X"00",X"FD",X"09",X"D0",X"01",X"00",X"03",X"C9",
		X"CD",X"92",X"26",X"DD",X"77",X"1F",X"5F",X"3A",X"07",X"99",X"87",X"87",X"87",X"CD",X"66",X"26",
		X"7C",X"CB",X"15",X"30",X"01",X"3C",X"C9",X"C6",X"02",X"30",X"02",X"3E",X"FF",X"CB",X"41",X"28",
		X"02",X"ED",X"44",X"E6",X"FC",X"0F",X"0F",X"80",X"DD",X"77",X"1F",X"87",X"21",X"7A",X"4D",X"5F",
		X"16",X"00",X"30",X"01",X"14",X"19",X"4E",X"23",X"5E",X"16",X"00",X"42",X"CB",X"21",X"CB",X"10",
		X"CB",X"21",X"CB",X"10",X"CB",X"23",X"CB",X"12",X"CB",X"23",X"CB",X"12",X"C9",X"3A",X"07",X"99",
		X"DD",X"66",X"04",X"2E",X"80",X"09",X"3D",X"20",X"FC",X"C9",X"3A",X"07",X"99",X"DD",X"66",X"04",
		X"2E",X"80",X"B7",X"ED",X"42",X"3D",X"20",X"FB",X"C9",X"3A",X"07",X"99",X"47",X"DD",X"66",X"05",
		X"2E",X"80",X"19",X"10",X"FD",X"C9",X"3A",X"07",X"99",X"47",X"DD",X"66",X"05",X"2E",X"80",X"B7",
		X"ED",X"52",X"10",X"FC",X"C9",X"CD",X"0D",X"3B",X"3A",X"3B",X"99",X"E6",X"33",X"C8",X"47",X"21",
		X"3A",X"99",X"AE",X"A0",X"C8",X"47",X"11",X"2A",X"99",X"1A",X"F6",X"28",X"6F",X"26",X"99",X"70",
		X"EE",X"01",X"12",X"C9",X"DD",X"35",X"0E",X"C0",X"DD",X"E5",X"E1",X"11",X"0A",X"00",X"19",X"5E",
		X"2C",X"56",X"2C",X"EB",X"7E",X"3C",X"28",X"0D",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"DD",X"75",
		X"0A",X"DD",X"74",X"0B",X"C9",X"23",X"4E",X"23",X"46",X"60",X"69",X"C3",X"D8",X"3A",X"21",X"20",
		X"99",X"35",X"20",X"0F",X"23",X"7E",X"34",X"2B",X"EB",X"21",X"F2",X"11",X"87",X"E7",X"ED",X"A0",
		X"7E",X"18",X"4F",X"3A",X"A8",X"9C",X"B7",X"28",X"49",X"3E",X"08",X"18",X"45",X"3A",X"3B",X"99",
		X"32",X"3A",X"99",X"3A",X"08",X"98",X"0F",X"30",X"D5",X"3A",X"0E",X"98",X"B7",X"28",X"10",X"3A",
		X"18",X"98",X"E6",X"01",X"47",X"3A",X"1C",X"98",X"E6",X"3E",X"B0",X"32",X"3B",X"99",X"C9",X"3A",
		X"1C",X"98",X"E6",X"01",X"4F",X"3A",X"18",X"98",X"87",X"E6",X"74",X"47",X"0F",X"E6",X"08",X"ED",
		X"44",X"80",X"CB",X"77",X"28",X"02",X"D6",X"30",X"B1",X"47",X"3A",X"1E",X"98",X"07",X"07",X"E6",
		X"02",X"B0",X"32",X"3B",X"99",X"C9",X"DD",X"6E",X"07",X"26",X"9A",X"7E",X"E6",X"3F",X"BE",X"28",
		X"05",X"3E",X"01",X"32",X"94",X"9C",X"7E",X"E6",X"3F",X"FE",X"04",X"30",X"15",X"EB",X"47",X"87",
		X"87",X"4F",X"DD",X"7E",X"09",X"EE",X"02",X"81",X"21",X"B1",X"3B",X"E7",X"7E",X"12",X"16",X"07",
		X"FF",X"C9",X"FE",X"0C",X"30",X"07",X"36",X"0B",X"EB",X"16",X"07",X"FF",X"C9",X"CB",X"67",X"C8",
		X"3A",X"80",X"9B",X"B7",X"CA",X"BD",X"27",X"EB",X"1A",X"E6",X"07",X"87",X"21",X"D3",X"36",X"E7",
		X"7E",X"83",X"4F",X"EB",X"3A",X"88",X"9B",X"B9",X"28",X"04",X"BD",X"C2",X"BD",X"27",X"11",X"71",
		X"27",X"D5",X"C3",X"BD",X"27",X"05",X"05",X"04",X"04",X"07",X"06",X"06",X"07",X"08",X"09",X"08",
		X"09",X"CD",X"C8",X"3B",X"CD",X"F4",X"3B",X"C9",X"3A",X"00",X"9D",X"0F",X"D0",X"ED",X"5B",X"02",
		X"9D",X"2A",X"07",X"9D",X"D9",X"06",X"05",X"11",X"20",X"00",X"DD",X"21",X"20",X"9D",X"D9",X"CD",
		X"3E",X"3C",X"38",X"06",X"D9",X"DD",X"19",X"10",X"F5",X"C9",X"CD",X"33",X"3C",X"21",X"02",X"04",
		X"22",X"00",X"9D",X"C9",X"0E",X"04",X"11",X"20",X"00",X"FD",X"21",X"20",X"9D",X"FD",X"7E",X"00",
		X"0F",X"30",X"20",X"FD",X"E5",X"DD",X"E1",X"DD",X"19",X"41",X"D9",X"FD",X"56",X"03",X"FD",X"5E",
		X"02",X"FD",X"66",X"08",X"FD",X"6E",X"07",X"D9",X"D9",X"CD",X"3E",X"3C",X"38",X"0B",X"D9",X"DD",
		X"19",X"10",X"F5",X"FD",X"19",X"0D",X"20",X"D5",X"C9",X"CD",X"56",X"3B",X"FD",X"34",X"00",X"FD",
		X"36",X"01",X"04",X"CD",X"69",X"20",X"DD",X"34",X"00",X"DD",X"36",X"01",X"04",X"C9",X"DD",X"7E",
		X"00",X"0F",X"D0",X"DD",X"7E",X"02",X"93",X"C6",X"08",X"FE",X"11",X"D0",X"DD",X"7E",X"03",X"92",
		X"C6",X"08",X"FE",X"11",X"D0",X"DD",X"7E",X"07",X"BD",X"20",X"14",X"7C",X"D6",X"08",X"FE",X"08",
		X"30",X"0D",X"C6",X"08",X"E6",X"FE",X"67",X"DD",X"7E",X"08",X"E6",X"FE",X"BC",X"20",X"02",X"37",
		X"C9",X"B7",X"C9",X"7B",X"3C",X"7B",X"38",X"5B",X"34",X"BB",X"2C",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"5B",X"5A",X"82",X"63",
		X"53",X"52",X"62",X"61",X"51",X"50",X"60",X"81",X"59",X"58",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"43",X"42",X"82",X"4B",
		X"3B",X"3A",X"4A",X"49",X"39",X"38",X"48",X"81",X"41",X"40",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"AD",X"AF",X"82",X"AE",
		X"6B",X"6A",X"7A",X"AC",X"69",X"68",X"78",X"81",X"79",X"7B",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"97",
		X"82",X"38",X"62",X"95",X"38",X"50",X"60",X"81",X"59",X"58",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"5B",X"5A",X"82",X"63",
		X"53",X"38",X"96",X"61",X"38",X"82",X"94",X"81",X"99",X"98",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"43",X"42",X"82",X"97",
		X"38",X"3A",X"4A",X"95",X"82",X"38",X"48",X"81",X"99",X"98",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"9B",X"9A",X"82",X"4B",
		X"38",X"82",X"96",X"49",X"39",X"38",X"94",X"81",X"41",X"40",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"AD",X"AF",X"82",X"97",
		X"AD",X"AF",X"96",X"95",X"AD",X"AF",X"94",X"81",X"79",X"7B",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"AE",
		X"7A",X"7A",X"7A",X"AC",X"78",X"78",X"78",X"81",X"99",X"98",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"97",
		X"8F",X"8E",X"7A",X"95",X"8D",X"8C",X"78",X"81",X"79",X"7B",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"97",
		X"82",X"82",X"96",X"95",X"82",X"82",X"94",X"81",X"99",X"98",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"BF",
		X"8B",X"8A",X"BE",X"BD",X"89",X"88",X"BC",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"BF",
		X"8B",X"8A",X"BE",X"BD",X"89",X"88",X"BC",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"BF",
		X"8B",X"8A",X"BE",X"BD",X"89",X"88",X"BC",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"BF",
		X"8B",X"8A",X"BE",X"BD",X"89",X"88",X"BC",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"65",X"63",X"53",X"5B",X"5B",X"5D",X"51",X"50",X"5D",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"65",X"5B",X"5B",X"5A",X"63",X"5D",X"59",X"58",X"5D",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"52",X"57",X"56",X"52",X"6F",
		X"55",X"54",X"54",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"52",X"5F",X"5E",X"52",X"54",
		X"54",X"5C",X"6F",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"4B",X"42",X"65",X"65",X"43",
		X"42",X"65",X"65",X"41",X"40",X"65",X"65",X"4B",X"62",X"65",X"65",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"4B",X"62",X"65",X"65",X"47",
		X"46",X"65",X"65",X"45",X"42",X"65",X"65",X"4B",X"42",X"65",X"65",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"65",X"65",X"4B",X"44",X"65",
		X"65",X"4B",X"4A",X"65",X"65",X"49",X"48",X"65",X"65",X"6E",X"44",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"65",X"65",X"6E",X"44",X"65",
		X"65",X"4F",X"4E",X"65",X"65",X"4B",X"4C",X"65",X"65",X"4B",X"44",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"64",X"64",X"64",X"64",X"64",
		X"64",X"64",X"64",X"67",X"33",X"3B",X"3B",X"6A",X"31",X"30",X"3D",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"64",X"64",X"64",X"64",X"64",
		X"64",X"64",X"64",X"3B",X"3B",X"3A",X"67",X"3D",X"39",X"38",X"6B",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"6A",X"37",X"36",X"32",X"73",
		X"35",X"34",X"34",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"32",X"3F",X"3E",X"6B",X"34",
		X"34",X"3C",X"73",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2B",X"22",X"64",X"64",X"23",
		X"22",X"64",X"64",X"21",X"20",X"64",X"64",X"76",X"66",X"64",X"64",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"74",X"66",X"64",X"64",X"27",
		X"26",X"64",X"64",X"25",X"22",X"64",X"64",X"2B",X"22",X"64",X"64",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"64",X"64",X"2B",X"24",X"64",
		X"64",X"2B",X"2A",X"64",X"64",X"29",X"28",X"64",X"64",X"72",X"76",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"64",X"64",X"72",X"74",X"64",
		X"64",X"2F",X"2E",X"64",X"64",X"2B",X"2C",X"64",X"64",X"2B",X"24",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"7B",X"7A",X"7A",X"7A",X"7B",
		X"7A",X"7A",X"7A",X"7B",X"7A",X"7A",X"7A",X"79",X"78",X"78",X"78",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"83",X"5B",X"5A",X"82",X"63",
		X"53",X"B6",X"66",X"61",X"B5",X"54",X"64",X"81",X"5D",X"5C",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"47",X"46",X"82",X"4B",
		X"BB",X"3E",X"4E",X"49",X"39",X"B8",X"4C",X"81",X"41",X"40",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"AD",X"AF",X"82",X"B2",
		X"73",X"72",X"7E",X"B0",X"71",X"70",X"7C",X"81",X"79",X"7B",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"97",
		X"82",X"38",X"66",X"95",X"38",X"54",X"64",X"81",X"5D",X"5C",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"5F",X"5E",X"82",X"67",
		X"57",X"38",X"96",X"65",X"38",X"82",X"94",X"81",X"99",X"98",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"47",X"46",X"82",X"97",
		X"38",X"3E",X"4E",X"95",X"82",X"38",X"4C",X"81",X"99",X"98",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"9B",X"9A",X"82",X"4F",
		X"38",X"82",X"96",X"4D",X"3D",X"38",X"94",X"81",X"45",X"44",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"B1",X"B3",X"82",X"97",
		X"B1",X"B3",X"96",X"95",X"B1",X"B3",X"94",X"81",X"7D",X"7F",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"B2",
		X"7E",X"7E",X"7E",X"B0",X"7C",X"7C",X"7C",X"81",X"99",X"98",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"97",
		X"8F",X"8E",X"93",X"95",X"8D",X"8C",X"91",X"81",X"7D",X"7F",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"9B",X"9A",X"82",X"97",
		X"82",X"82",X"96",X"95",X"82",X"82",X"94",X"81",X"99",X"98",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"BF",
		X"8B",X"8A",X"DA",X"BD",X"89",X"88",X"D8",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"BF",
		X"8B",X"8A",X"BE",X"BD",X"89",X"88",X"BC",X"81",X"DD",X"DC",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"C3",X"C2",X"82",X"DB",
		X"8B",X"8A",X"BE",X"D9",X"89",X"88",X"BC",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"DF",X"DE",X"82",X"BF",
		X"8B",X"8A",X"BE",X"BD",X"89",X"88",X"BC",X"81",X"C1",X"C0",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"65",X"63",X"53",X"5B",X"5B",X"54",X"51",X"50",X"54",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"65",X"5B",X"5B",X"5A",X"63",X"54",X"59",X"58",X"54",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"52",X"57",X"56",X"52",X"6F",
		X"55",X"54",X"54",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"52",X"5F",X"5E",X"52",X"54",
		X"54",X"5C",X"6F",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"4B",X"42",X"65",X"65",X"43",
		X"42",X"65",X"65",X"41",X"40",X"65",X"65",X"4B",X"62",X"65",X"65",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"4B",X"62",X"65",X"65",X"47",
		X"46",X"65",X"65",X"45",X"42",X"65",X"65",X"4B",X"42",X"65",X"65",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"65",X"65",X"4B",X"44",X"65",
		X"65",X"4B",X"4A",X"65",X"65",X"49",X"48",X"65",X"65",X"6E",X"42",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"65",X"65",X"6E",X"42",X"65",
		X"65",X"4F",X"4E",X"65",X"65",X"4B",X"4C",X"65",X"65",X"4B",X"44",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"64",X"64",X"64",X"64",X"64",
		X"64",X"64",X"64",X"61",X"13",X"1B",X"1B",X"68",X"11",X"70",X"1D",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"64",X"64",X"64",X"64",X"64",
		X"64",X"64",X"64",X"1B",X"1B",X"1A",X"61",X"1D",X"19",X"18",X"69",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"68",X"17",X"16",X"12",X"6D",
		X"15",X"14",X"14",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"12",X"1F",X"1E",X"69",X"14",
		X"14",X"1C",X"6D",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0B",X"02",X"64",X"64",X"03",
		X"02",X"64",X"64",X"01",X"00",X"64",X"64",X"77",X"60",X"64",X"64",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"75",X"60",X"64",X"64",X"07",
		X"06",X"64",X"64",X"05",X"02",X"64",X"64",X"0B",X"02",X"64",X"64",X"C0",X"C0",X"10",X"10",X"C0",
		X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"64",X"64",X"0B",X"04",X"64",
		X"64",X"0B",X"0A",X"64",X"64",X"09",X"08",X"64",X"64",X"6C",X"77",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"64",X"64",X"6C",X"75",X"64",
		X"64",X"0F",X"0E",X"64",X"64",X"0B",X"0C",X"64",X"64",X"0B",X"04",X"10",X"10",X"C0",X"C0",X"10",
		X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"10",X"10",X"C0",X"C0",X"83",X"5F",X"5E",X"82",X"67",
		X"57",X"BA",X"62",X"65",X"B9",X"50",X"60",X"81",X"59",X"58",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"43",X"42",X"82",X"4F",
		X"B7",X"3A",X"4A",X"4D",X"3D",X"B4",X"48",X"81",X"45",X"44",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"B1",X"B3",X"82",X"AE",
		X"6F",X"6E",X"7A",X"AC",X"6D",X"6C",X"78",X"81",X"7D",X"7F",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"83",X"5F",X"5E",X"82",X"67",
		X"57",X"56",X"66",X"65",X"55",X"54",X"64",X"81",X"5D",X"5C",X"80",X"9C",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"83",X"47",X"46",X"82",X"4F",
		X"3F",X"3E",X"4E",X"4D",X"3D",X"3C",X"4C",X"81",X"45",X"44",X"80",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"9D",X"83",X"B1",X"B3",X"82",X"B2",
		X"77",X"76",X"7E",X"B0",X"75",X"74",X"7C",X"81",X"7D",X"7F",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"0E",X"04",X"0F",X"04",X"0C",
		X"04",X"0D",X"04",X"06",X"03",X"07",X"02",X"09",X"01",X"08",X"00",X"04",X"01",X"0B",X"00",X"0A",
		X"03",X"05",X"02",X"01",X"00",X"03",X"01",X"00",X"02",X"02",X"03",X"06",X"03",X"07",X"02",X"0C",
		X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"09",X"01",X"08",X"00",X"04",X"01",X"0F",X"04",X"0C",
		X"04",X"05",X"02",X"0E",X"04",X"0B",X"00",X"0A",X"03",X"0D",X"04",X"0E",X"04",X"03",X"01",X"0C",
		X"04",X"02",X"03",X"01",X"00",X"0F",X"04",X"00",X"02",X"0D",X"04",X"06",X"03",X"07",X"02",X"0C",
		X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"0C",X"04",X"0D",X"04",X"06",X"03",X"07",X"02",X"09",
		X"01",X"08",X"00",X"04",X"01",X"0B",X"00",X"0A",X"03",X"05",X"02",X"01",X"00",X"03",X"01",X"00",
		X"02",X"02",X"03",X"0E",X"04",X"0F",X"04",X"0C",X"04",X"0D",X"04",X"0E",X"04",X"1F",X"00",X"1D",
		X"03",X"0D",X"04",X"15",X"03",X"17",X"02",X"0C",X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"1B",
		X"01",X"19",X"00",X"11",X"01",X"0F",X"04",X"0C",X"04",X"13",X"02",X"0E",X"04",X"1E",X"00",X"1C",
		X"03",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"1A",X"01",X"18",X"00",X"14",X"03",X"16",X"02",X"0C",
		X"04",X"0D",X"04",X"10",X"01",X"0F",X"04",X"0C",X"04",X"12",X"02",X"0E",X"04",X"1F",X"00",X"1D",
		X"03",X"0D",X"04",X"15",X"03",X"17",X"02",X"0C",X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"1B",
		X"01",X"19",X"00",X"11",X"01",X"0F",X"04",X"0C",X"04",X"13",X"02",X"0E",X"04",X"1E",X"00",X"1C",
		X"03",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"1A",X"01",X"18",X"00",X"14",X"03",X"16",X"02",X"0C",
		X"04",X"0D",X"04",X"10",X"01",X"0F",X"04",X"0C",X"04",X"12",X"02",X"0E",X"04",X"0F",X"04",X"0C",
		X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"0C",X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"0C",
		X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"0C",X"04",X"0D",X"04",X"0E",X"04",X"0F",X"04",X"0C",
		X"04",X"0D",X"04",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"80",X"40",X"80",X"80",X"40",X"40",
		X"80",X"40",X"80",X"40",X"40",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"40",X"00",
		X"40",X"40",X"00",X"00",X"40",X"00",X"40",X"40",X"00",X"40",X"00",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"00",X"40",X"40",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"40",X"40",X"40",
		X"00",X"00",X"40",X"00",X"40",X"40",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"00",X"00",X"40",
		X"00",X"00",X"40",X"00",X"40",X"40",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"40",X"40",X"40",
		X"00",X"00",X"40",X"00",X"40",X"40",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"00",X"00",X"40",
		X"00",X"00",X"40",X"C1",X"01",X"00",X"C1",X"00",X"00",X"FD",X"01",X"00",X"FD",X"00",X"00",X"F9",
		X"01",X"00",X"F9",X"00",X"00",X"F5",X"01",X"00",X"F5",X"00",X"00",X"F1",X"00",X"00",X"F1",X"01",
		X"00",X"ED",X"00",X"00",X"ED",X"00",X"00",X"E9",X"00",X"00",X"E9",X"00",X"00",X"E5",X"00",X"00",
		X"E5",X"00",X"00",X"E1",X"00",X"00",X"E1",X"00",X"00",X"DD",X"00",X"00",X"DD",X"00",X"00",X"D9",
		X"00",X"00",X"D9",X"00",X"00",X"D5",X"00",X"00",X"D5",X"00",X"00",X"D1",X"00",X"00",X"D1",X"01",
		X"00",X"CD",X"00",X"00",X"CD",X"00",X"00",X"C9",X"00",X"00",X"C9",X"00",X"00",X"C5",X"00",X"00",
		X"C5",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"64",X"64",X"64",X"64",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"64",X"64",X"64",X"64",X"A3",X"A2",X"10",
		X"10",X"10",X"10",X"10",X"10",X"93",X"92",X"64",X"64",X"64",X"FE",X"FE",X"A6",X"A3",X"A2",X"10",
		X"10",X"10",X"71",X"71",X"8F",X"64",X"64",X"CB",X"CA",X"FD",X"FC",X"A9",X"A8",X"A3",X"A2",X"71",
		X"71",X"71",X"8E",X"64",X"C9",X"C8",X"C7",X"C6",X"A5",X"A4",X"A1",X"A0",X"A5",X"71",X"71",X"8C",
		X"64",X"FE",X"FE",X"A7",X"A1",X"A0",X"A4",X"10",X"10",X"71",X"71",X"8D",X"64",X"64",X"A1",X"A0",
		X"A4",X"10",X"10",X"10",X"10",X"10",X"91",X"90",X"64",X"64",X"64",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"64",X"64",X"64",X"64",X"64",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"64",X"64",X"64",X"64",X"64",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",
		X"C0",X"80",X"80",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"C0",X"C0",X"C0",X"80",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",
		X"C0",X"80",X"C0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"80",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"71",X"71",
		X"71",X"71",X"71",X"71",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",
		X"71",X"A3",X"A2",X"10",X"10",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"FE",X"FE",
		X"A6",X"A3",X"A2",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"CB",X"CA",X"FD",X"FC",X"A9",
		X"A8",X"A3",X"AB",X"AA",X"71",X"71",X"71",X"71",X"C9",X"C8",X"C7",X"C6",X"A5",X"A4",X"A1",X"A9",
		X"A8",X"71",X"71",X"71",X"71",X"FE",X"FE",X"A7",X"A1",X"A0",X"A4",X"10",X"71",X"71",X"71",X"71",
		X"71",X"71",X"A1",X"A0",X"A4",X"10",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",
		X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"10",X"10",X"10",X"10",X"10",X"71",X"71",X"71",
		X"71",X"71",X"71",X"71",X"71",X"A3",X"A2",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",
		X"71",X"71",X"FE",X"FE",X"A6",X"A3",X"A2",X"AB",X"AB",X"AF",X"71",X"71",X"71",X"71",X"71",X"CB",
		X"CA",X"FD",X"FC",X"A9",X"10",X"10",X"10",X"AE",X"71",X"71",X"71",X"71",X"C9",X"C8",X"C7",X"C6",
		X"A5",X"10",X"10",X"10",X"AC",X"71",X"71",X"71",X"71",X"FE",X"FE",X"A7",X"A1",X"A0",X"A9",X"A9",
		X"AD",X"71",X"71",X"71",X"71",X"71",X"A1",X"A0",X"A4",X"10",X"10",X"71",X"71",X"71",X"71",X"71",
		X"71",X"71",X"71",X"10",X"10",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",
		X"10",X"10",X"10",X"10",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"80",X"80",X"80",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"10",
		X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"10",X"71",X"71",X"71",
		X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"A3",X"10",X"10",X"10",X"10",X"B7",X"B6",
		X"71",X"71",X"71",X"71",X"71",X"71",X"FE",X"10",X"10",X"10",X"10",X"10",X"B3",X"71",X"71",X"71",
		X"71",X"71",X"71",X"CB",X"10",X"10",X"10",X"10",X"10",X"B2",X"71",X"71",X"71",X"71",X"71",X"71",
		X"C9",X"10",X"10",X"10",X"10",X"10",X"B0",X"71",X"71",X"71",X"71",X"71",X"71",X"FE",X"10",X"10",
		X"10",X"10",X"10",X"B1",X"71",X"71",X"71",X"71",X"71",X"71",X"A1",X"10",X"10",X"10",X"10",X"B5",
		X"B4",X"71",X"71",X"71",X"71",X"71",X"71",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",
		X"71",X"71",X"71",X"71",X"10",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",
		X"71",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"B7",X"B6",X"71",X"71",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"BF",X"71",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"BE",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"BB",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"BA",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"B8",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"B9",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"BC",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"BD",X"71",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"B5",X"B4",X"71",X"71",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"06",X"FF",X"0D",X"FF",
		X"13",X"FF",X"19",X"FF",X"1F",X"FE",X"26",X"FD",X"2C",X"FC",X"32",X"FB",X"38",X"FA",X"3E",X"F8",
		X"44",X"F7",X"4A",X"F5",X"50",X"F3",X"56",X"F1",X"5C",X"EF",X"62",X"ED",X"68",X"EA",X"6D",X"E7",
		X"73",X"E5",X"79",X"E2",X"7E",X"DF",X"84",X"DC",X"89",X"D8",X"8E",X"D5",X"93",X"D1",X"99",X"CE",
		X"9E",X"CA",X"A2",X"C6",X"A7",X"C2",X"AC",X"BE",X"B1",X"B9",X"B5",X"B5",X"B9",X"B1",X"BE",X"AC",
		X"C2",X"A7",X"C6",X"A2",X"CA",X"9E",X"CE",X"99",X"D1",X"93",X"D5",X"8E",X"D8",X"89",X"DC",X"84",
		X"DF",X"7E",X"E2",X"79",X"E5",X"73",X"E7",X"6D",X"EA",X"68",X"ED",X"62",X"EF",X"5C",X"F1",X"56",
		X"F3",X"50",X"F5",X"4A",X"F7",X"44",X"F8",X"3E",X"FA",X"38",X"FB",X"32",X"FC",X"2C",X"FD",X"26",
		X"FE",X"1F",X"FF",X"19",X"FF",X"13",X"FF",X"0D",X"FF",X"06",X"FF",X"00",X"FF",X"06",X"FF",X"0D",
		X"FF",X"13",X"FF",X"19",X"FE",X"1F",X"FD",X"26",X"FC",X"2C",X"FB",X"32",X"FA",X"38",X"F8",X"3E",
		X"F7",X"44",X"F5",X"4A",X"F3",X"50",X"F1",X"56",X"EF",X"5C",X"ED",X"62",X"EA",X"68",X"E7",X"6D",
		X"E5",X"73",X"E2",X"79",X"DF",X"7E",X"DC",X"84",X"D8",X"89",X"D5",X"8E",X"D1",X"93",X"CE",X"99",
		X"CA",X"9E",X"C6",X"A2",X"C2",X"A7",X"BE",X"AC",X"B9",X"B1",X"B5",X"B5",X"B1",X"B9",X"AC",X"BE",
		X"A7",X"C2",X"A2",X"C6",X"9E",X"CA",X"99",X"CE",X"93",X"D1",X"8E",X"D5",X"89",X"D8",X"84",X"DC",
		X"7E",X"DF",X"79",X"E2",X"73",X"E5",X"6D",X"E7",X"68",X"EA",X"62",X"ED",X"5C",X"EF",X"56",X"F1",
		X"50",X"F3",X"4A",X"F5",X"44",X"F7",X"3E",X"F8",X"38",X"FA",X"32",X"FB",X"2C",X"FC",X"26",X"FD",
		X"1F",X"FE",X"19",X"FF",X"13",X"FF",X"0D",X"FF",X"06",X"FF",X"00",X"FF",X"06",X"FF",X"0D",X"FF",
		X"13",X"FF",X"19",X"FF",X"1F",X"FE",X"26",X"FD",X"2C",X"FC",X"32",X"FB",X"38",X"FA",X"3E",X"F8",
		X"44",X"F7",X"4A",X"F5",X"50",X"F3",X"56",X"F1",X"5C",X"EF",X"62",X"ED",X"68",X"EA",X"6D",X"E7",
		X"73",X"E5",X"79",X"E2",X"7E",X"DF",X"84",X"DC",X"89",X"D8",X"8E",X"D5",X"93",X"D1",X"99",X"CE",
		X"9E",X"CA",X"A2",X"C6",X"A7",X"C2",X"AC",X"BE",X"B1",X"B9",X"B5",X"B5",X"B9",X"B1",X"BE",X"AC",
		X"C2",X"A7",X"C6",X"A2",X"CA",X"9E",X"CE",X"99",X"D1",X"93",X"D5",X"8E",X"D8",X"89",X"DC",X"84",
		X"DF",X"7E",X"E2",X"79",X"E5",X"73",X"E7",X"6D",X"EA",X"68",X"ED",X"62",X"EF",X"5C",X"F1",X"56",
		X"F3",X"50",X"F5",X"4A",X"F7",X"44",X"F8",X"3E",X"FA",X"38",X"FB",X"32",X"FC",X"2C",X"FD",X"26",
		X"FE",X"1F",X"FF",X"19",X"FF",X"13",X"FF",X"0D",X"FF",X"06",X"FF",X"00",X"FF",X"06",X"FF",X"0D",
		X"FF",X"13",X"FF",X"19",X"FE",X"1F",X"FD",X"26",X"FC",X"2C",X"FB",X"32",X"FA",X"38",X"F8",X"3E",
		X"F7",X"44",X"F5",X"4A",X"F3",X"50",X"F1",X"56",X"EF",X"5C",X"ED",X"62",X"EA",X"68",X"E7",X"6D",
		X"E5",X"73",X"E2",X"79",X"DF",X"7E",X"DC",X"84",X"D8",X"89",X"D5",X"8E",X"D1",X"93",X"CE",X"99",
		X"CA",X"9E",X"C6",X"A2",X"C2",X"A7",X"BE",X"AC",X"B9",X"B1",X"B5",X"B5",X"B1",X"B9",X"AC",X"BE",
		X"A7",X"C2",X"A2",X"C6",X"9E",X"CA",X"99",X"CE",X"93",X"D1",X"8E",X"D5",X"89",X"D8",X"84",X"DC",
		X"7E",X"DF",X"79",X"E2",X"73",X"E5",X"6D",X"E7",X"68",X"EA",X"62",X"ED",X"5C",X"EF",X"56",X"F1",
		X"50",X"F3",X"4A",X"F5",X"44",X"F7",X"3E",X"F8",X"38",X"FA",X"32",X"FB",X"2C",X"FC",X"26",X"FD",
		X"1F",X"FE",X"19",X"FF",X"13",X"FF",X"0D",X"FF",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
