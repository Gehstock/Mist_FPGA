library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity wacko_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of wacko_sp_bits is
	type rom is array(0 to 32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"99",X"99",X"00",X"90",X"A9",X"93",X"00",X"99",X"9F",X"93",X"00",X"33",X"9F",X"9B",
		X"00",X"93",X"FF",X"9B",X"00",X"93",X"F9",X"93",X"00",X"B9",X"99",X"9B",X"00",X"B9",X"33",X"9B",
		X"00",X"39",X"39",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"93",X"33",X"00",X"09",X"99",X"33",
		X"00",X"00",X"99",X"33",X"00",X"90",X"33",X"39",X"00",X"99",X"99",X"99",X"00",X"39",X"B9",X"90",
		X"00",X"33",X"99",X"99",X"00",X"93",X"9B",X"39",X"90",X"99",X"93",X"33",X"09",X"00",X"33",X"33",
		X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"99",X"00",X"99",X"93",X"33",X"09",X"33",X"93",X"33",
		X"00",X"33",X"33",X"33",X"00",X"99",X"33",X"33",X"00",X"99",X"39",X"33",X"09",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"99",X"99",X"9D",
		X"99",X"99",X"99",X"DD",X"9D",X"22",X"99",X"DD",X"99",X"DD",X"99",X"DD",X"49",X"9D",X"22",X"DD",
		X"9D",X"9D",X"22",X"9D",X"92",X"D2",X"99",X"9D",X"99",X"22",X"99",X"99",X"00",X"99",X"95",X"22",
		X"00",X"59",X"95",X"29",X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"92",X"00",X"99",X"59",X"22",
		X"00",X"99",X"99",X"22",X"00",X"99",X"29",X"29",X"00",X"D2",X"22",X"99",X"00",X"22",X"99",X"22",
		X"00",X"22",X"99",X"22",X"00",X"29",X"99",X"22",X"00",X"99",X"9A",X"22",X"00",X"29",X"99",X"29",
		X"00",X"22",X"99",X"2A",X"00",X"99",X"22",X"29",X"00",X"9A",X"22",X"29",X"00",X"99",X"22",X"22",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"99",X"99",X"9D",X"99",X"99",X"99",X"DD",
		X"9D",X"22",X"99",X"DD",X"99",X"DD",X"99",X"DD",X"99",X"9D",X"22",X"DD",X"9D",X"9D",X"22",X"9D",
		X"92",X"D2",X"99",X"9D",X"99",X"22",X"99",X"99",X"00",X"99",X"95",X"22",X"09",X"59",X"95",X"29",
		X"09",X"99",X"99",X"22",X"09",X"22",X"22",X"92",X"00",X"29",X"22",X"22",X"00",X"22",X"92",X"22",
		X"00",X"99",X"22",X"29",X"00",X"D9",X"22",X"99",X"00",X"D9",X"99",X"22",X"00",X"29",X"DD",X"22",
		X"00",X"29",X"99",X"22",X"00",X"29",X"9A",X"22",X"00",X"29",X"99",X"29",X"00",X"22",X"99",X"2A",
		X"00",X"99",X"22",X"29",X"00",X"9A",X"22",X"29",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"22",
		X"00",X"99",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"99",X"22",X"00",X"22",X"9A",X"22",X"00",X"22",X"99",X"22",
		X"00",X"22",X"99",X"99",X"99",X"92",X"22",X"A9",X"92",X"99",X"22",X"99",X"92",X"22",X"22",X"99",
		X"92",X"99",X"99",X"22",X"92",X"00",X"91",X"29",X"92",X"00",X"92",X"29",X"99",X"99",X"99",X"29",
		X"09",X"29",X"09",X"29",X"00",X"29",X"09",X"29",X"00",X"99",X"09",X"19",X"00",X"90",X"09",X"99",
		X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"99",X"00",X"00",X"90",X"92",X"00",X"00",X"90",
		X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"99",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"99",
		X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"A9",X"00",X"22",X"22",X"99",X"00",X"22",X"29",X"92",
		X"00",X"22",X"99",X"29",X"00",X"22",X"92",X"29",X"00",X"22",X"22",X"99",X"00",X"22",X"99",X"99",
		X"00",X"92",X"9A",X"22",X"00",X"99",X"99",X"22",X"00",X"2D",X"29",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"29",X"00",X"22",X"99",X"99",X"00",X"22",X"90",X"99",X"00",X"29",X"00",X"92",
		X"00",X"99",X"00",X"22",X"00",X"90",X"00",X"22",X"00",X"90",X"00",X"22",X"00",X"90",X"00",X"22",
		X"00",X"99",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"D2",X"00",X"22",
		X"00",X"DD",X"00",X"22",X"00",X"2D",X"00",X"22",X"99",X"22",X"00",X"22",X"92",X"2D",X"00",X"99",
		X"92",X"2D",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"09",X"09",X"09",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"44",X"9B",X"99",X"09",X"99",X"BB",X"9B",X"9B",X"BB",X"BB",X"9B",X"B9",X"BB",X"BB",
		X"99",X"B9",X"BB",X"BB",X"99",X"B9",X"99",X"BB",X"09",X"BB",X"99",X"BB",X"09",X"99",X"99",X"BB",
		X"00",X"95",X"99",X"BB",X"00",X"95",X"99",X"BB",X"00",X"4F",X"99",X"BB",X"00",X"99",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"B9",X"44",X"BB",X"99",X"90",X"04",X"99",X"BB",X"90",
		X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"99",X"00",X"09",X"99",X"BB",
		X"00",X"99",X"77",X"BB",X"00",X"9B",X"77",X"BB",X"00",X"BB",X"77",X"BB",X"00",X"B9",X"99",X"BB",
		X"00",X"99",X"11",X"BB",X"00",X"99",X"77",X"BB",X"00",X"19",X"97",X"BB",X"00",X"71",X"11",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"43",X"9B",X"99",X"09",X"99",X"BB",X"9B",X"9B",X"BB",X"BB",
		X"9B",X"B9",X"BB",X"BB",X"94",X"B9",X"BB",X"BB",X"99",X"B9",X"BB",X"BB",X"09",X"BB",X"99",X"BB",
		X"09",X"BB",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",X"95",X"99",X"BB",X"00",X"4F",X"99",X"BB",
		X"00",X"49",X"99",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"B9",X"00",X"BB",X"99",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"99",
		X"00",X"09",X"99",X"B9",X"00",X"99",X"77",X"B9",X"00",X"9B",X"77",X"BB",X"00",X"BB",X"77",X"BB",
		X"00",X"B9",X"99",X"BB",X"00",X"99",X"11",X"BB",X"00",X"99",X"77",X"BB",X"00",X"19",X"97",X"BB",
		X"00",X"77",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",X"11",X"17",X"BB",X"00",X"77",X"77",X"BB",
		X"00",X"77",X"79",X"BB",X"00",X"99",X"79",X"BB",X"00",X"11",X"99",X"B9",X"00",X"77",X"9B",X"B9",
		X"00",X"77",X"BB",X"B9",X"00",X"99",X"B9",X"B9",X"00",X"11",X"99",X"B9",X"00",X"77",X"1B",X"BB",
		X"00",X"77",X"99",X"BB",X"00",X"77",X"BB",X"9B",X"00",X"99",X"BB",X"9B",X"00",X"11",X"BB",X"99",
		X"00",X"77",X"BB",X"19",X"09",X"77",X"BB",X"99",X"09",X"99",X"9B",X"BB",X"09",X"B9",X"99",X"BB",
		X"09",X"99",X"9B",X"99",X"09",X"90",X"9B",X"99",X"00",X"B9",X"9B",X"90",X"00",X"BB",X"9B",X"99",
		X"00",X"BB",X"99",X"9B",X"00",X"BB",X"09",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",
		X"09",X"99",X"00",X"99",X"99",X"90",X"00",X"09",X"9B",X"90",X"00",X"9B",X"99",X"00",X"00",X"99",
		X"00",X"71",X"11",X"BB",X"00",X"79",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",X"BB",X"99",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"99",X"BB",X"B9",X"00",X"99",X"BB",X"99",X"00",X"19",X"BB",X"00",
		X"00",X"79",X"99",X"00",X"00",X"77",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"11",X"BB",X"00",
		X"00",X"77",X"BB",X"00",X"00",X"77",X"BB",X"09",X"00",X"77",X"BB",X"99",X"00",X"99",X"BB",X"9B",
		X"00",X"11",X"BB",X"BB",X"00",X"77",X"BB",X"BB",X"00",X"77",X"BB",X"BB",X"00",X"99",X"9B",X"BB",
		X"00",X"09",X"99",X"BB",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"99",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"9B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"90",
		X"99",X"99",X"66",X"99",X"9E",X"9E",X"66",X"69",X"9E",X"E9",X"66",X"66",X"9E",X"E9",X"99",X"99",
		X"99",X"E9",X"9C",X"66",X"09",X"EE",X"CC",X"66",X"09",X"EE",X"CC",X"66",X"99",X"EE",X"CC",X"66",
		X"99",X"E9",X"99",X"66",X"99",X"99",X"99",X"66",X"99",X"99",X"CC",X"66",X"99",X"99",X"9C",X"66",
		X"99",X"49",X"9C",X"66",X"99",X"99",X"9C",X"66",X"9C",X"CC",X"CC",X"66",X"9C",X"C9",X"CC",X"66",
		X"9C",X"99",X"CC",X"66",X"99",X"99",X"CC",X"66",X"09",X"99",X"C9",X"66",X"09",X"99",X"99",X"66",
		X"09",X"F9",X"9D",X"66",X"00",X"99",X"DD",X"66",X"00",X"CC",X"D6",X"66",X"00",X"99",X"66",X"66",
		X"00",X"99",X"99",X"00",X"00",X"96",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"90",X"00",X"99",X"66",X"99",X"09",X"9E",X"66",X"69",
		X"09",X"E9",X"66",X"66",X"09",X"E9",X"99",X"99",X"09",X"E9",X"9C",X"66",X"00",X"EE",X"CC",X"66",
		X"09",X"EE",X"CC",X"66",X"99",X"EE",X"CC",X"66",X"9C",X"E9",X"99",X"66",X"99",X"99",X"99",X"66",
		X"99",X"99",X"CC",X"66",X"99",X"99",X"9C",X"66",X"99",X"49",X"9C",X"66",X"99",X"99",X"9C",X"66",
		X"9C",X"CC",X"CC",X"66",X"9C",X"C9",X"CC",X"66",X"9C",X"99",X"CC",X"66",X"99",X"99",X"CC",X"66",
		X"09",X"99",X"C9",X"66",X"09",X"99",X"99",X"66",X"09",X"99",X"9D",X"66",X"00",X"CC",X"DD",X"66",
		X"00",X"99",X"D6",X"66",X"00",X"DD",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"99",X"66",X"66",X"00",X"55",X"99",X"66",
		X"00",X"99",X"9D",X"66",X"00",X"99",X"DD",X"66",X"00",X"99",X"DD",X"66",X"00",X"55",X"D9",X"66",
		X"00",X"99",X"99",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"D6",X"66",X"66",X"00",X"DD",X"99",X"66",X"99",X"66",X"99",X"66",X"99",X"66",X"9D",X"66",
		X"99",X"66",X"DD",X"66",X"97",X"66",X"D6",X"99",X"97",X"66",X"D6",X"CC",X"97",X"66",X"96",X"CC",
		X"97",X"69",X"96",X"C9",X"97",X"99",X"99",X"CC",X"97",X"00",X"97",X"CC",X"99",X"00",X"97",X"9C",
		X"99",X"00",X"99",X"9C",X"09",X"00",X"79",X"99",X"09",X"00",X"77",X"9C",X"09",X"00",X"99",X"99",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"99",X"66",X"66",X"00",X"55",X"99",X"66",X"00",X"99",X"9D",X"66",X"00",X"99",X"DD",X"66",
		X"00",X"99",X"DD",X"66",X"00",X"55",X"D9",X"66",X"00",X"99",X"99",X"66",X"00",X"66",X"66",X"66",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"69",X"66",
		X"00",X"99",X"69",X"66",X"00",X"DD",X"69",X"66",X"00",X"6D",X"69",X"66",X"09",X"66",X"69",X"99",
		X"09",X"66",X"69",X"CC",X"09",X"66",X"69",X"CC",X"09",X"99",X"69",X"CC",X"00",X"77",X"69",X"CC",
		X"00",X"99",X"99",X"CC",X"00",X"99",X"79",X"CC",X"00",X"97",X"99",X"CC",X"00",X"77",X"99",X"9C",
		X"00",X"77",X"99",X"9C",X"00",X"77",X"00",X"9C",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"90",X"00",X"09",X"9E",X"99",X"00",X"09",X"99",X"E9",
		X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"99",X"E9",
		X"00",X"EE",X"9E",X"99",X"00",X"99",X"99",X"B9",X"00",X"EE",X"97",X"B9",X"00",X"9E",X"99",X"99",
		X"00",X"99",X"99",X"B9",X"00",X"E9",X"99",X"99",X"00",X"9B",X"E9",X"EE",X"00",X"9B",X"99",X"E9",
		X"00",X"9E",X"9E",X"E9",X"00",X"9E",X"9E",X"E9",X"00",X"9E",X"9E",X"99",X"00",X"9B",X"99",X"B9",
		X"00",X"9B",X"99",X"E9",X"09",X"99",X"E9",X"EB",X"09",X"E9",X"E9",X"EB",X"09",X"49",X"E9",X"B9",
		X"00",X"00",X"B9",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"90",
		X"00",X"09",X"9E",X"99",X"00",X"09",X"99",X"E9",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"9E",X"99",X"E9",X"00",X"9E",X"99",X"E9",X"00",X"E9",X"9E",X"99",X"00",X"99",X"99",X"B9",
		X"00",X"E9",X"97",X"B9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"B9",X"00",X"E9",X"99",X"99",
		X"00",X"9B",X"99",X"EE",X"00",X"9B",X"99",X"E9",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"9E",X"E9",
		X"00",X"9E",X"9E",X"99",X"00",X"9B",X"99",X"B9",X"00",X"9B",X"9E",X"E9",X"09",X"99",X"EE",X"EB",
		X"09",X"E9",X"EE",X"EB",X"09",X"49",X"9E",X"B9",X"00",X"9E",X"99",X"EE",X"00",X"9E",X"E9",X"EE",
		X"09",X"99",X"99",X"EE",X"09",X"9E",X"9E",X"EE",X"00",X"9E",X"9E",X"9E",X"09",X"9E",X"99",X"99",
		X"09",X"99",X"E9",X"99",X"09",X"EB",X"E9",X"9E",X"09",X"BE",X"99",X"99",X"09",X"B9",X"9E",X"EE",
		X"00",X"99",X"9E",X"99",X"00",X"E9",X"E9",X"99",X"00",X"E9",X"49",X"99",X"00",X"E9",X"E9",X"E9",
		X"00",X"E9",X"9E",X"9E",X"00",X"9E",X"9E",X"99",X"00",X"E9",X"9E",X"EE",X"00",X"E9",X"9E",X"99",
		X"00",X"99",X"9E",X"99",X"00",X"B9",X"99",X"00",X"00",X"B9",X"EE",X"00",X"00",X"E9",X"9E",X"00",
		X"00",X"EE",X"9E",X"90",X"00",X"EE",X"9E",X"90",X"00",X"9E",X"99",X"90",X"00",X"99",X"9E",X"99",
		X"00",X"E9",X"9E",X"B9",X"00",X"E9",X"9E",X"99",X"00",X"E9",X"99",X"EE",X"09",X"99",X"E9",X"9E",
		X"09",X"EE",X"EE",X"99",X"09",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9E",X"E9",X"99",X"09",X"9E",X"E9",X"EE",X"09",X"99",X"99",X"EE",X"09",X"9E",X"99",X"E9",
		X"00",X"9E",X"99",X"99",X"00",X"9E",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"EB",X"E9",X"99",
		X"00",X"B9",X"99",X"99",X"00",X"B9",X"9E",X"E9",X"00",X"99",X"9E",X"99",X"00",X"E9",X"EE",X"99",
		X"00",X"E9",X"4E",X"90",X"00",X"E9",X"99",X"90",X"00",X"EB",X"E9",X"99",X"09",X"BB",X"E9",X"E9",
		X"09",X"B9",X"99",X"EE",X"99",X"99",X"EE",X"99",X"9E",X"99",X"EE",X"E9",X"99",X"90",X"99",X"E9",
		X"99",X"00",X"00",X"9B",X"9E",X"00",X"00",X"9E",X"99",X"99",X"00",X"99",X"09",X"E9",X"00",X"E9",
		X"00",X"EE",X"00",X"E9",X"09",X"9E",X"00",X"E9",X"09",X"9E",X"00",X"E9",X"99",X"9E",X"00",X"99",
		X"9E",X"99",X"00",X"E9",X"99",X"B9",X"00",X"99",X"9E",X"B9",X"00",X"9B",X"99",X"99",X"00",X"99",
		X"99",X"00",X"09",X"00",X"9A",X"00",X"99",X"00",X"99",X"00",X"79",X"99",X"09",X"00",X"79",X"77",
		X"09",X"99",X"77",X"77",X"00",X"97",X"79",X"77",X"00",X"97",X"79",X"97",X"00",X"97",X"97",X"99",
		X"00",X"97",X"97",X"44",X"00",X"77",X"99",X"99",X"00",X"79",X"49",X"77",X"00",X"99",X"04",X"77",
		X"09",X"F9",X"00",X"97",X"09",X"99",X"00",X"99",X"09",X"99",X"00",X"E9",X"09",X"99",X"40",X"E9",
		X"09",X"97",X"90",X"79",X"00",X"97",X"94",X"79",X"00",X"97",X"99",X"79",X"00",X"79",X"79",X"79",
		X"00",X"99",X"77",X"79",X"00",X"90",X"77",X"79",X"00",X"09",X"77",X"79",X"00",X"99",X"77",X"79",
		X"00",X"97",X"77",X"79",X"00",X"77",X"77",X"79",X"00",X"77",X"77",X"79",X"00",X"77",X"77",X"99",
		X"00",X"99",X"97",X"77",X"00",X"91",X"99",X"77",X"00",X"91",X"99",X"77",X"00",X"99",X"11",X"77",
		X"00",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"9A",X"00",X"77",X"99",X"9A",X"00",X"79",X"99",
		X"9A",X"00",X"79",X"77",X"9A",X"90",X"77",X"97",X"99",X"99",X"77",X"99",X"09",X"79",X"99",X"99",
		X"09",X"77",X"97",X"99",X"09",X"77",X"99",X"99",X"09",X"77",X"00",X"77",X"09",X"99",X"00",X"79",
		X"09",X"99",X"00",X"79",X"99",X"99",X"00",X"79",X"97",X"97",X"00",X"79",X"97",X"77",X"00",X"79",
		X"97",X"77",X"00",X"79",X"97",X"79",X"00",X"79",X"97",X"99",X"00",X"79",X"99",X"99",X"90",X"79",
		X"00",X"09",X"90",X"79",X"00",X"09",X"90",X"79",X"00",X"99",X"99",X"79",X"00",X"97",X"79",X"79",
		X"00",X"97",X"79",X"79",X"00",X"97",X"77",X"79",X"00",X"97",X"77",X"79",X"00",X"77",X"77",X"99",
		X"00",X"99",X"97",X"77",X"00",X"91",X"99",X"77",X"00",X"91",X"99",X"77",X"00",X"99",X"11",X"77",
		X"00",X"49",X"99",X"77",X"00",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"77",
		X"00",X"94",X"49",X"77",X"00",X"94",X"49",X"77",X"00",X"19",X"44",X"77",X"00",X"19",X"99",X"77",
		X"00",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"77",
		X"00",X"49",X"49",X"77",X"00",X"99",X"49",X"77",X"00",X"99",X"49",X"77",X"00",X"99",X"99",X"77",
		X"00",X"94",X"97",X"77",X"00",X"94",X"97",X"99",X"00",X"94",X"97",X"00",X"00",X"99",X"77",X"00",
		X"00",X"91",X"77",X"00",X"00",X"91",X"77",X"00",X"00",X"99",X"77",X"00",X"00",X"11",X"77",X"00",
		X"00",X"99",X"77",X"00",X"00",X"11",X"77",X"90",X"00",X"11",X"77",X"99",X"00",X"99",X"77",X"77",
		X"00",X"94",X"99",X"77",X"00",X"79",X"19",X"77",X"00",X"79",X"91",X"77",X"00",X"99",X"99",X"99",
		X"00",X"49",X"99",X"77",X"00",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"77",
		X"00",X"94",X"49",X"77",X"09",X"94",X"49",X"77",X"09",X"19",X"44",X"77",X"09",X"19",X"99",X"77",
		X"09",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"97",
		X"00",X"49",X"49",X"97",X"00",X"99",X"49",X"99",X"00",X"99",X"49",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"97",X"00",X"00",X"94",X"97",X"00",X"00",X"94",X"97",X"00",X"00",X"99",X"77",X"00",
		X"00",X"91",X"77",X"00",X"00",X"91",X"77",X"99",X"00",X"99",X"77",X"97",X"00",X"11",X"77",X"77",
		X"00",X"99",X"77",X"77",X"00",X"11",X"77",X"77",X"00",X"11",X"77",X"77",X"00",X"99",X"77",X"79",
		X"00",X"94",X"99",X"99",X"00",X"79",X"19",X"90",X"00",X"99",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"92",X"99",X"09",X"00",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"92",X"22",X"99",
		X"99",X"92",X"29",X"99",X"99",X"92",X"99",X"99",X"09",X"92",X"94",X"99",X"09",X"99",X"94",X"99",
		X"00",X"99",X"44",X"99",X"90",X"99",X"49",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"99",
		X"99",X"99",X"92",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"29",X"99",X"09",X"99",X"22",X"99",
		X"09",X"99",X"29",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"92",X"99",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",X"92",X"22",X"99",
		X"99",X"99",X"29",X"99",X"99",X"99",X"99",X"99",X"09",X"99",X"94",X"99",X"09",X"99",X"94",X"99",
		X"00",X"99",X"44",X"99",X"90",X"99",X"49",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"99",
		X"99",X"99",X"92",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"59",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"29",X"99",X"09",X"99",X"22",X"99",
		X"09",X"99",X"29",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"D9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"09",X"99",X"22",X"99",X"09",X"99",X"22",X"99",X"09",X"99",X"22",X"99",
		X"09",X"99",X"22",X"9D",X"09",X"99",X"29",X"D9",X"09",X"99",X"99",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"E9",X"99",X"00",X"09",X"EE",X"93",X"00",X"99",X"3E",X"39",X"00",X"39",X"99",X"39",
		X"00",X"99",X"FF",X"99",X"00",X"99",X"99",X"90",X"00",X"9F",X"99",X"90",X"00",X"9F",X"99",X"90",
		X"00",X"99",X"AA",X"99",X"00",X"39",X"F9",X"39",X"00",X"33",X"99",X"39",X"00",X"33",X"33",X"99",
		X"00",X"33",X"99",X"90",X"00",X"33",X"39",X"00",X"00",X"93",X"39",X"00",X"99",X"93",X"94",X"00",
		X"93",X"99",X"99",X"99",X"93",X"09",X"99",X"39",X"93",X"09",X"B3",X"39",X"99",X"99",X"33",X"39",
		X"00",X"33",X"33",X"39",X"00",X"99",X"39",X"99",X"00",X"00",X"39",X"90",X"00",X"00",X"39",X"00",
		X"00",X"00",X"39",X"00",X"00",X"90",X"33",X"00",X"00",X"99",X"93",X"00",X"00",X"39",X"93",X"00",
		X"00",X"39",X"93",X"00",X"00",X"33",X"93",X"00",X"00",X"33",X"93",X"00",X"00",X"99",X"99",X"00",
		X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"9D",
		X"09",X"99",X"00",X"D9",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",X"99",
		X"99",X"D9",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"D9",X"94",X"99",X"99",X"9D",X"44",X"99",
		X"99",X"99",X"44",X"99",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"F9",X"99",
		X"99",X"99",X"D9",X"99",X"90",X"99",X"D9",X"09",X"90",X"99",X"D9",X"09",X"90",X"90",X"99",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"9D",X"00",X"90",X"99",X"D9",X"00",X"99",X"99",X"99",X"09",X"99",X"94",X"99",
		X"99",X"D9",X"49",X"99",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"FD",X"99",X"99",X"99",X"3D",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"D9",X"99",
		X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"9D",X"90",X"99",X"99",X"99",X"00",X"99",X"90",X"90",X"00",
		X"99",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"90",X"99",X"90",X"00",X"99",X"95",X"99",X"00",X"99",X"95",X"99",
		X"00",X"99",X"59",X"99",X"00",X"99",X"99",X"99",X"00",X"D9",X"99",X"99",X"00",X"D9",X"FD",X"99",
		X"00",X"DD",X"3D",X"99",X"00",X"9D",X"DD",X"99",X"00",X"9D",X"D9",X"99",X"00",X"9D",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"D9",X"90",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"A0",X"00",X"00",X"FF",X"FA",X"00",X"00",X"AF",X"FA",X"00",X"00",X"AA",X"FF",
		X"00",X"0A",X"FF",X"FF",X"00",X"0A",X"FA",X"FF",X"00",X"AA",X"FF",X"FF",X"00",X"FA",X"AA",X"FF",
		X"00",X"AA",X"FA",X"AF",X"00",X"AF",X"FF",X"AF",X"00",X"AF",X"FF",X"FF",X"00",X"AA",X"FF",X"FF",
		X"00",X"FA",X"AF",X"FF",X"00",X"FA",X"AA",X"FF",X"00",X"FA",X"FF",X"FF",X"00",X"FA",X"FF",X"FA",
		X"00",X"FA",X"AF",X"FF",X"00",X"AF",X"AF",X"FF",X"00",X"AF",X"AA",X"AF",X"00",X"AF",X"FA",X"AA",
		X"00",X"AF",X"AA",X"FA",X"00",X"AF",X"FF",X"FA",X"00",X"FF",X"FF",X"AA",X"00",X"FF",X"FF",X"FF",
		X"00",X"AA",X"FF",X"FF",X"00",X"FF",X"FF",X"AA",X"00",X"AF",X"FF",X"00",X"00",X"0A",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"AA",X"0A",X"00",X"00",X"FF",X"0A",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"A0",X"AF",X"00",X"00",X"AA",X"AF",
		X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"FF",X"00",X"0A",
		X"AA",X"FF",X"00",X"AA",X"AF",X"FF",X"00",X"AF",X"AF",X"FF",X"00",X"AF",X"AA",X"FF",X"00",X"FF",
		X"00",X"AF",X"00",X"AA",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"0A",X"A0",X"A0",X"00",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"0A",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"F0",X"00",X"3F",X"F3",X"30",
		X"00",X"0F",X"F0",X"00",X"AA",X"F3",X"F0",X"00",X"00",X"30",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"3F",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"F9",X"90",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"9F",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"50",
		X"00",X"99",X"0E",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"0A",X"99",X"00",X"00",X"0A",X"99",X"0A",X"00",X"0A",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"0A",X"99",X"00",X"00",X"05",X"99",X"00",X"00",X"0A",X"99",X"83",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"77",X"00",X"00",X"90",X"E9",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"77",X"00",X"00",X"00",X"E7",X"10",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"99",X"00",X"59",X"00",X"95",X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",
		X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"09",X"99",X"99",X"99",
		X"09",X"A9",X"44",X"9A",X"99",X"AA",X"99",X"AA",X"9A",X"3A",X"99",X"33",X"9A",X"33",X"99",X"5A",
		X"9A",X"33",X"99",X"35",X"9A",X"5A",X"44",X"33",X"9A",X"3A",X"44",X"AA",X"9A",X"99",X"44",X"AA",
		X"9A",X"90",X"99",X"9A",X"9A",X"90",X"99",X"99",X"93",X"90",X"99",X"09",X"93",X"90",X"99",X"09",
		X"9A",X"00",X"99",X"09",X"9A",X"00",X"99",X"09",X"9A",X"00",X"99",X"09",X"93",X"00",X"44",X"00",
		X"9A",X"00",X"99",X"00",X"9A",X"09",X"00",X"90",X"9A",X"99",X"00",X"99",X"9A",X"95",X"00",X"59",
		X"9A",X"59",X"00",X"95",X"9A",X"99",X"00",X"99",X"9A",X"99",X"00",X"99",X"99",X"00",X"00",X"00",
		X"00",X"99",X"00",X"99",X"00",X"59",X"00",X"95",X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",
		X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"99",X"99",X"99",
		X"00",X"99",X"44",X"99",X"00",X"9A",X"99",X"A9",X"00",X"9A",X"99",X"39",X"00",X"93",X"99",X"39",
		X"00",X"93",X"99",X"A9",X"00",X"9A",X"44",X"A9",X"00",X"93",X"44",X"39",X"00",X"93",X"44",X"A9",
		X"00",X"9A",X"99",X"A9",X"00",X"9A",X"99",X"39",X"00",X"9A",X"99",X"A9",X"00",X"9A",X"99",X"A9",
		X"00",X"9A",X"99",X"39",X"00",X"93",X"99",X"39",X"00",X"93",X"99",X"A9",X"00",X"93",X"44",X"99",
		X"00",X"9A",X"99",X"90",X"00",X"99",X"00",X"90",X"00",X"09",X"00",X"99",X"00",X"95",X"00",X"59",
		X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",X"00",X"A9",X"00",X"99",X"00",X"9A",X"00",X"90",
		X"00",X"99",X"00",X"99",X"00",X"59",X"00",X"95",X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",
		X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"99",X"99",X"99",
		X"00",X"99",X"44",X"90",X"00",X"9A",X"99",X"99",X"00",X"9A",X"99",X"A9",X"00",X"93",X"99",X"3A",
		X"00",X"93",X"99",X"AA",X"00",X"A3",X"44",X"A3",X"00",X"A3",X"44",X"A3",X"00",X"AA",X"44",X"A3",
		X"00",X"3A",X"99",X"AA",X"00",X"3A",X"99",X"3A",X"00",X"3A",X"99",X"3A",X"00",X"AA",X"99",X"A3",
		X"00",X"3A",X"99",X"A3",X"00",X"3A",X"99",X"A3",X"00",X"3A",X"99",X"3A",X"00",X"3A",X"44",X"3A",
		X"00",X"AA",X"99",X"AA",X"00",X"A9",X"00",X"9A",X"00",X"99",X"00",X"99",X"00",X"95",X"00",X"59",
		X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"44",X"00",
		X"00",X"94",X"99",X"99",X"00",X"44",X"22",X"49",X"00",X"49",X"99",X"44",X"00",X"99",X"AA",X"44",
		X"99",X"99",X"9A",X"11",X"91",X"59",X"99",X"51",X"9E",X"11",X"99",X"55",X"99",X"11",X"11",X"55",
		X"09",X"11",X"71",X"55",X"00",X"E9",X"79",X"EE",X"00",X"EE",X"77",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"44",X"00",
		X"00",X"94",X"99",X"99",X"00",X"44",X"22",X"49",X"00",X"49",X"99",X"44",X"00",X"92",X"AA",X"44",
		X"99",X"99",X"9A",X"11",X"91",X"79",X"99",X"71",X"9E",X"11",X"99",X"77",X"99",X"11",X"11",X"77",
		X"09",X"11",X"51",X"77",X"00",X"E9",X"59",X"EE",X"00",X"EE",X"55",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"9E",X"09",X"00",X"00",X"F9",X"09",
		X"00",X"00",X"FF",X"99",X"00",X"90",X"FF",X"93",X"00",X"99",X"F4",X"93",X"00",X"33",X"FF",X"9B",
		X"00",X"93",X"FF",X"9B",X"00",X"93",X"FF",X"93",X"00",X"B9",X"4F",X"9B",X"00",X"B9",X"99",X"9B",
		X"00",X"39",X"39",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"93",X"33",X"00",X"09",X"99",X"33",
		X"00",X"00",X"99",X"33",X"00",X"A0",X"33",X"39",X"04",X"AA",X"99",X"99",X"04",X"05",X"B9",X"90",
		X"00",X"95",X"99",X"00",X"00",X"94",X"93",X"91",X"00",X"49",X"93",X"91",X"40",X"79",X"43",X"15",
		X"00",X"99",X"44",X"11",X"00",X"5A",X"34",X"59",X"00",X"11",X"94",X"11",X"70",X"A5",X"A1",X"55",
		X"00",X"15",X"11",X"91",X"00",X"50",X"A1",X"00",X"04",X"00",X"11",X"00",X"47",X"07",X"10",X"07",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"99",X"99",X"00",X"90",X"A9",X"93",X"00",X"99",X"FF",X"93",X"00",X"33",X"FF",X"9B",
		X"00",X"93",X"9F",X"9B",X"00",X"93",X"9F",X"93",X"00",X"B9",X"F9",X"9B",X"00",X"B9",X"99",X"9B",
		X"00",X"39",X"33",X"39",X"00",X"93",X"39",X"39",X"00",X"99",X"33",X"33",X"00",X"09",X"99",X"33",
		X"00",X"00",X"B9",X"33",X"00",X"00",X"33",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"90",
		X"00",X"09",X"33",X"00",X"00",X"99",X"39",X"00",X"00",X"93",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"39",X"39",X"00",X"00",X"39",X"33",X"90",X"00",X"39",X"33",X"99",X"00",X"99",X"33",X"39",
		X"00",X"00",X"33",X"99",X"00",X"00",X"93",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"9B",X"94",X"90",
		X"09",X"99",X"99",X"99",X"09",X"E9",X"99",X"B9",X"99",X"EE",X"B9",X"BB",X"91",X"9E",X"BB",X"9B",
		X"91",X"99",X"99",X"9B",X"91",X"11",X"59",X"BB",X"91",X"EE",X"59",X"99",X"91",X"EE",X"99",X"95",
		X"91",X"EE",X"99",X"99",X"91",X"E1",X"99",X"B9",X"91",X"11",X"99",X"99",X"91",X"19",X"BB",X"9B",
		X"91",X"99",X"9B",X"B9",X"91",X"9B",X"99",X"00",X"91",X"9B",X"B7",X"00",X"91",X"BB",X"BB",X"00",
		X"91",X"B9",X"BB",X"00",X"91",X"99",X"BB",X"00",X"91",X"90",X"19",X"00",X"91",X"90",X"99",X"90",
		X"91",X"00",X"B9",X"99",X"91",X"00",X"B9",X"B9",X"91",X"00",X"B9",X"BB",X"91",X"00",X"B9",X"BB",
		X"99",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"9B",X"00",X"00",X"B9",X"9B",X"00",X"00",X"99",X"99",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"9B",X"93",X"90",
		X"00",X"99",X"99",X"99",X"00",X"19",X"99",X"B9",X"00",X"E9",X"B9",X"BB",X"00",X"E1",X"BB",X"9B",
		X"00",X"EE",X"99",X"9B",X"00",X"1E",X"59",X"BB",X"00",X"11",X"59",X"99",X"00",X"11",X"99",X"95",
		X"00",X"11",X"99",X"99",X"00",X"11",X"BB",X"B9",X"00",X"99",X"BB",X"99",X"00",X"BB",X"99",X"BB",
		X"00",X"9B",X"B7",X"B9",X"00",X"99",X"B7",X"99",X"00",X"91",X"B7",X"00",X"00",X"91",X"BB",X"00",
		X"00",X"91",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"B9",X"99",X"00",X"00",X"B9",X"B9",X"00",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"BB",
		X"00",X"00",X"B9",X"9B",X"00",X"00",X"B9",X"9B",X"00",X"00",X"B9",X"99",X"00",X"00",X"99",X"09",
		X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"99",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"EE",X"66",X"00",X"00",X"EE",X"6D",X"00",
		X"00",X"99",X"6D",X"90",X"00",X"94",X"99",X"90",X"00",X"44",X"C9",X"90",X"00",X"99",X"C9",X"90",
		X"00",X"CC",X"99",X"90",X"00",X"CC",X"9D",X"90",X"00",X"C9",X"9D",X"90",X"00",X"99",X"DD",X"90",
		X"00",X"99",X"99",X"90",X"00",X"95",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"CC",X"99",X"90",
		X"00",X"CC",X"96",X"90",X"00",X"99",X"96",X"90",X"00",X"66",X"66",X"90",X"00",X"69",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"90",X"96",X"00",X"00",X"90",X"99",X"00",X"00",X"09",X"C9",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"77",X"00",X"00",X"09",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"EE",X"66",X"90",X"00",X"EE",X"66",X"90",X"00",X"99",X"6D",X"90",
		X"00",X"94",X"99",X"90",X"00",X"94",X"C9",X"90",X"00",X"99",X"C9",X"90",X"00",X"CC",X"99",X"90",
		X"00",X"CC",X"9D",X"90",X"00",X"C9",X"9D",X"99",X"00",X"99",X"DD",X"69",X"00",X"99",X"DD",X"69",
		X"00",X"95",X"DD",X"69",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"CC",X"99",X"99",
		X"00",X"99",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"99",X"69",X"69",X"00",X"96",X"99",X"99",
		X"00",X"96",X"90",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"9C",X"99",X"00",X"99",X"99",X"66",
		X"00",X"77",X"00",X"66",X"00",X"77",X"00",X"99",X"00",X"99",X"00",X"97",X"00",X"00",X"00",X"99",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"9A",X"00",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"9E",X"00",X"E9",X"99",X"EE",X"00",X"E9",X"9E",X"9E",X"00",X"99",X"E9",X"99",
		X"99",X"9E",X"99",X"9B",X"9E",X"9E",X"99",X"9B",X"9E",X"EE",X"99",X"BB",X"99",X"EE",X"99",X"99",
		X"91",X"9E",X"99",X"9E",X"91",X"9E",X"EE",X"9E",X"99",X"99",X"99",X"9E",X"00",X"9E",X"E9",X"99",
		X"00",X"EE",X"E9",X"90",X"00",X"99",X"9E",X"00",X"00",X"19",X"9B",X"00",X"00",X"E1",X"9B",X"00",
		X"00",X"E9",X"9B",X"00",X"00",X"99",X"99",X"90",X"00",X"B9",X"EE",X"99",X"00",X"BE",X"EE",X"9E",
		X"09",X"99",X"99",X"EE",X"09",X"09",X"09",X"EE",X"09",X"09",X"09",X"99",X"09",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"9A",X"00",X"00",X"99",X"9A",X"00",
		X"00",X"91",X"99",X"00",X"00",X"E9",X"99",X"90",X"00",X"E9",X"9E",X"99",X"00",X"B9",X"E9",X"EE",
		X"09",X"9B",X"99",X"99",X"09",X"99",X"99",X"19",X"99",X"E9",X"99",X"99",X"9E",X"E9",X"99",X"E9",
		X"9E",X"99",X"99",X"EE",X"9E",X"9E",X"99",X"EE",X"99",X"99",X"99",X"99",X"9E",X"9E",X"E9",X"9B",
		X"9E",X"9E",X"E9",X"9B",X"99",X"99",X"9E",X"99",X"00",X"B9",X"9B",X"09",X"00",X"EE",X"9B",X"00",
		X"00",X"99",X"9B",X"90",X"09",X"9E",X"09",X"99",X"09",X"EE",X"00",X"E9",X"99",X"99",X"09",X"99",
		X"9E",X"E9",X"09",X"E9",X"9E",X"E9",X"09",X"E9",X"99",X"E9",X"00",X"EE",X"00",X"99",X"00",X"99",
		X"09",X"99",X"00",X"99",X"99",X"77",X"00",X"79",X"93",X"77",X"09",X"79",X"99",X"77",X"09",X"77",
		X"97",X"77",X"09",X"97",X"97",X"77",X"09",X"99",X"97",X"99",X"09",X"99",X"97",X"99",X"99",X"99",
		X"97",X"90",X"77",X"79",X"97",X"99",X"77",X"99",X"99",X"77",X"77",X"99",X"00",X"77",X"77",X"77",
		X"00",X"77",X"77",X"77",X"09",X"77",X"77",X"77",X"99",X"77",X"99",X"97",X"97",X"94",X"49",X"97",
		X"97",X"94",X"49",X"97",X"97",X"99",X"44",X"49",X"97",X"94",X"99",X"49",X"97",X"99",X"11",X"A9",
		X"97",X"09",X"11",X"99",X"94",X"00",X"11",X"79",X"94",X"00",X"99",X"77",X"0A",X"00",X"19",X"77",
		X"09",X"00",X"19",X"97",X"09",X"00",X"99",X"97",X"00",X"00",X"99",X"97",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",
		X"09",X"99",X"00",X"99",X"99",X"77",X"00",X"99",X"99",X"77",X"09",X"99",X"93",X"77",X"09",X"79",
		X"93",X"77",X"09",X"97",X"99",X"77",X"09",X"99",X"97",X"79",X"09",X"99",X"97",X"79",X"99",X"99",
		X"97",X"79",X"77",X"99",X"97",X"90",X"77",X"77",X"99",X"99",X"77",X"99",X"00",X"77",X"77",X"90",
		X"00",X"77",X"77",X"99",X"00",X"77",X"77",X"77",X"00",X"97",X"99",X"77",X"00",X"97",X"49",X"77",
		X"00",X"97",X"49",X"77",X"00",X"99",X"44",X"77",X"00",X"97",X"99",X"77",X"00",X"99",X"11",X"77",
		X"00",X"49",X"11",X"79",X"00",X"44",X"11",X"47",X"00",X"74",X"99",X"49",X"00",X"79",X"19",X"79",
		X"00",X"77",X"19",X"79",X"00",X"79",X"00",X"A9",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"92",X"09",X"99",X"00",X"92",X"99",X"99",
		X"00",X"92",X"22",X"99",X"00",X"22",X"29",X"90",X"00",X"29",X"99",X"90",X"00",X"29",X"99",X"99",
		X"00",X"92",X"94",X"99",X"00",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"95",X"90",X"09",X"99",X"99",X"90",X"09",X"99",X"95",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"D9",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"22",X"99",X"00",X"92",X"22",X"99",X"00",X"92",X"29",X"99",X"00",X"92",X"99",X"99",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"09",X"00",X"99",X"59",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"59",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"93",X"00",
		X"00",X"99",X"34",X"00",X"00",X"92",X"99",X"00",X"00",X"29",X"22",X"00",X"00",X"24",X"22",X"00",
		X"09",X"22",X"92",X"00",X"09",X"99",X"99",X"09",X"99",X"95",X"99",X"99",X"92",X"99",X"99",X"22",
		X"92",X"29",X"99",X"22",X"92",X"99",X"92",X"29",X"99",X"99",X"22",X"99",X"00",X"99",X"29",X"9D",
		X"00",X"92",X"99",X"2D",X"00",X"99",X"92",X"D2",X"00",X"D9",X"22",X"DD",X"00",X"2D",X"22",X"DD",
		X"00",X"DD",X"22",X"2D",X"00",X"DD",X"22",X"D9",X"00",X"DD",X"22",X"99",X"00",X"D2",X"22",X"00",
		X"00",X"DD",X"A2",X"00",X"00",X"99",X"22",X"99",X"00",X"09",X"99",X"22",X"00",X"09",X"99",X"22",
		X"00",X"99",X"99",X"92",X"00",X"92",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"99",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"94",X"00",
		X"00",X"99",X"44",X"00",X"00",X"92",X"99",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"22",X"00",
		X"00",X"22",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"95",X"00",
		X"00",X"29",X"99",X"00",X"00",X"22",X"92",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"99",X"90",
		X"00",X"9D",X"9D",X"90",X"00",X"9D",X"9D",X"90",X"00",X"92",X"9D",X"99",X"00",X"9D",X"9D",X"D9",
		X"00",X"9D",X"99",X"D9",X"00",X"9D",X"29",X"D9",X"00",X"99",X"29",X"D9",X"00",X"09",X"29",X"D9",
		X"00",X"09",X"99",X"99",X"00",X"09",X"22",X"90",X"00",X"09",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"99",X"99",X"00",X"90",X"F9",X"93",X"00",X"99",X"FF",X"93",X"00",X"33",X"A9",X"9B",
		X"00",X"93",X"99",X"9B",X"00",X"93",X"99",X"93",X"00",X"B9",X"99",X"9B",X"00",X"B9",X"33",X"9B",
		X"00",X"39",X"39",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"33",X"33",X"00",X"09",X"93",X"33",
		X"00",X"00",X"99",X"33",X"00",X"00",X"33",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"90",
		X"00",X"99",X"99",X"90",X"00",X"94",X"93",X"99",X"00",X"49",X"93",X"49",X"00",X"99",X"33",X"44",
		X"99",X"99",X"33",X"11",X"91",X"59",X"33",X"51",X"9E",X"11",X"99",X"55",X"99",X"11",X"11",X"55",
		X"09",X"11",X"71",X"55",X"00",X"E9",X"79",X"EE",X"00",X"EE",X"77",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",X"00",X"00",X"99",X"99",
		X"00",X"90",X"F9",X"93",X"00",X"99",X"99",X"93",X"00",X"33",X"99",X"9B",X"00",X"93",X"99",X"9B",
		X"00",X"93",X"F9",X"93",X"00",X"B9",X"99",X"9B",X"00",X"B9",X"33",X"9B",X"00",X"39",X"39",X"39",
		X"00",X"93",X"33",X"39",X"00",X"99",X"33",X"33",X"00",X"09",X"93",X"33",X"00",X"00",X"99",X"33",
		X"00",X"00",X"33",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"90",X"00",X"00",X"99",X"00",
		X"00",X"99",X"93",X"90",X"00",X"94",X"93",X"99",X"00",X"49",X"33",X"49",X"00",X"99",X"33",X"44",
		X"99",X"99",X"33",X"11",X"91",X"79",X"33",X"71",X"9E",X"11",X"99",X"77",X"99",X"11",X"11",X"77",
		X"09",X"11",X"51",X"77",X"00",X"E9",X"59",X"EE",X"00",X"EE",X"55",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"49",X"00",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"49",X"90",X"00",X"00",X"F9",X"90",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"49",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"04",X"00",X"00",X"F9",X"00",X"50",
		X"00",X"99",X"0E",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"0A",X"9A",X"00",X"00",X"0A",X"49",X"00",X"00",X"0A",X"44",X"0A",X"00",X"0A",X"4A",X"00",
		X"00",X"0A",X"A4",X"00",X"00",X"0A",X"A4",X"00",X"00",X"05",X"49",X"00",X"00",X"0A",X"9A",X"83",
		X"00",X"00",X"A4",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"74",X"00",X"00",X"90",X"E9",X"00",
		X"00",X"90",X"9A",X"00",X"00",X"90",X"77",X"00",X"00",X"00",X"E7",X"10",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"09",X"E9",X"99",X"00",X"0E",X"EE",X"93",X"00",X"09",X"EE",X"93",
		X"00",X"99",X"39",X"33",X"00",X"93",X"99",X"39",X"00",X"93",X"9A",X"39",X"00",X"93",X"9F",X"99",
		X"00",X"93",X"9F",X"90",X"00",X"99",X"99",X"90",X"00",X"39",X"39",X"90",X"00",X"99",X"33",X"90",
		X"00",X"93",X"93",X"00",X"00",X"93",X"33",X"90",X"00",X"9B",X"93",X"90",X"00",X"9B",X"33",X"90",
		X"00",X"99",X"93",X"90",X"00",X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"33",X"99",X"90",X"00",X"9B",X"33",X"90",X"09",X"09",X"B3",X"39",
		X"09",X"99",X"39",X"99",X"09",X"93",X"B9",X"90",X"00",X"99",X"39",X"90",X"00",X"33",X"33",X"90",
		X"90",X"33",X"33",X"90",X"00",X"99",X"33",X"90",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"9D",X"00",X"00",X"99",X"9D",X"00",X"99",X"94",X"DD",X"00",X"99",X"94",X"DD",
		X"00",X"99",X"94",X"DD",X"99",X"99",X"94",X"D9",X"D2",X"22",X"99",X"D9",X"D2",X"22",X"22",X"D9",
		X"D2",X"22",X"22",X"D9",X"22",X"22",X"99",X"99",X"99",X"99",X"99",X"92",X"95",X"95",X"99",X"22",
		X"99",X"95",X"99",X"22",X"09",X"99",X"99",X"29",X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"92",
		X"09",X"59",X"95",X"99",X"99",X"99",X"99",X"99",X"92",X"22",X"22",X"22",X"99",X"92",X"99",X"22",
		X"09",X"22",X"99",X"22",X"00",X"99",X"DD",X"22",X"09",X"99",X"22",X"22",X"99",X"92",X"22",X"92",
		X"9A",X"22",X"29",X"92",X"99",X"22",X"2D",X"92",X"09",X"22",X"2D",X"92",X"09",X"22",X"2D",X"22",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"9D",
		X"00",X"00",X"99",X"9D",X"00",X"99",X"94",X"DD",X"00",X"99",X"94",X"DD",X"00",X"99",X"94",X"DD",
		X"99",X"99",X"94",X"D9",X"D2",X"22",X"99",X"D9",X"D2",X"22",X"22",X"D9",X"D2",X"22",X"22",X"D9",
		X"22",X"22",X"99",X"99",X"99",X"99",X"99",X"92",X"95",X"95",X"99",X"22",X"99",X"95",X"99",X"22",
		X"29",X"99",X"99",X"29",X"92",X"22",X"29",X"22",X"9D",X"22",X"29",X"92",X"99",X"22",X"22",X"99",
		X"00",X"29",X"92",X"99",X"00",X"22",X"22",X"22",X"00",X"99",X"99",X"22",X"00",X"9D",X"DD",X"22",
		X"00",X"A2",X"DD",X"22",X"09",X"92",X"22",X"22",X"99",X"92",X"22",X"92",X"9A",X"22",X"29",X"92",
		X"99",X"22",X"2D",X"92",X"09",X"22",X"2D",X"92",X"09",X"22",X"2D",X"22",X"09",X"22",X"2D",X"22",
		X"09",X"22",X"2D",X"22",X"09",X"22",X"2D",X"22",X"09",X"22",X"2D",X"22",X"99",X"22",X"2D",X"22",
		X"9A",X"22",X"2D",X"22",X"99",X"99",X"2D",X"22",X"09",X"9A",X"2D",X"29",X"09",X"99",X"2D",X"29",
		X"99",X"99",X"2D",X"29",X"99",X"22",X"2D",X"29",X"22",X"99",X"29",X"29",X"22",X"29",X"99",X"29",
		X"22",X"90",X"92",X"2A",X"29",X"00",X"22",X"29",X"22",X"00",X"29",X"29",X"22",X"00",X"99",X"29",
		X"92",X"00",X"22",X"19",X"99",X"00",X"22",X"99",X"09",X"00",X"22",X"00",X"09",X"00",X"92",X"00",
		X"99",X"00",X"92",X"00",X"92",X"00",X"99",X"00",X"92",X"00",X"09",X"00",X"22",X"00",X"99",X"00",
		X"99",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"99",
		X"09",X"22",X"2D",X"22",X"09",X"22",X"29",X"22",X"99",X"22",X"99",X"29",X"9A",X"22",X"92",X"99",
		X"99",X"99",X"22",X"90",X"09",X"92",X"22",X"00",X"09",X"91",X"22",X"00",X"09",X"99",X"22",X"99",
		X"09",X"22",X"22",X"29",X"99",X"99",X"22",X"22",X"91",X"D9",X"29",X"22",X"92",X"D9",X"99",X"22",
		X"99",X"DD",X"90",X"22",X"00",X"29",X"90",X"22",X"00",X"99",X"00",X"22",X"00",X"90",X"00",X"22",
		X"09",X"00",X"00",X"22",X"09",X"00",X"09",X"22",X"99",X"00",X"99",X"22",X"92",X"00",X"92",X"22",
		X"92",X"90",X"92",X"29",X"99",X"90",X"92",X"99",X"09",X"99",X"99",X"90",X"00",X"29",X"00",X"99",
		X"00",X"29",X"00",X"29",X"00",X"D2",X"00",X"22",X"90",X"D2",X"00",X"22",X"99",X"D2",X"00",X"92",
		X"DD",X"D2",X"00",X"92",X"2D",X"29",X"00",X"99",X"22",X"99",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"09",X"00",X"49",X"49",X"99",X"00",X"49",X"49",X"BB",
		X"00",X"93",X"49",X"BB",X"90",X"99",X"99",X"BB",X"90",X"BB",X"BB",X"BB",X"99",X"99",X"BB",X"BB",
		X"BB",X"99",X"BB",X"99",X"BB",X"99",X"99",X"99",X"BB",X"BB",X"99",X"B9",X"9B",X"99",X"99",X"B9",
		X"99",X"99",X"99",X"B9",X"05",X"99",X"99",X"B9",X"09",X"44",X"99",X"B9",X"09",X"BB",X"99",X"99",
		X"09",X"BB",X"BB",X"90",X"09",X"BB",X"BB",X"00",X"44",X"99",X"BB",X"00",X"40",X"90",X"BB",X"00",
		X"40",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"90",X"00",X"99",X"9B",X"90",
		X"00",X"BB",X"99",X"99",X"00",X"B9",X"79",X"B9",X"00",X"99",X"77",X"BB",X"00",X"91",X"77",X"BB",
		X"09",X"77",X"17",X"BB",X"09",X"77",X"77",X"BB",X"09",X"99",X"77",X"BB",X"09",X"11",X"77",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"09",X"00",X"49",X"49",X"99",
		X"00",X"39",X"39",X"BB",X"00",X"94",X"49",X"9B",X"90",X"99",X"99",X"9B",X"90",X"BB",X"BB",X"BB",
		X"99",X"99",X"BB",X"BB",X"BB",X"49",X"BB",X"99",X"BB",X"99",X"BB",X"99",X"BB",X"BB",X"99",X"B9",
		X"9B",X"BB",X"99",X"B9",X"99",X"99",X"99",X"B9",X"05",X"99",X"99",X"B9",X"09",X"44",X"99",X"B9",
		X"09",X"BB",X"99",X"99",X"09",X"BB",X"99",X"90",X"09",X"BB",X"BB",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"90",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"99",X"9B",X"00",X"00",X"BB",X"99",X"90",X"00",X"B9",X"79",X"99",X"00",X"99",X"79",X"B9",
		X"00",X"91",X"79",X"B9",X"09",X"77",X"19",X"B9",X"09",X"77",X"79",X"B9",X"09",X"99",X"79",X"B9",
		X"09",X"77",X"77",X"BB",X"99",X"99",X"79",X"BB",X"9B",X"11",X"99",X"B9",X"9B",X"77",X"9B",X"B9",
		X"99",X"77",X"9B",X"99",X"99",X"99",X"B9",X"90",X"99",X"11",X"B9",X"90",X"09",X"77",X"99",X"00",
		X"09",X"77",X"9B",X"00",X"00",X"99",X"9B",X"00",X"00",X"11",X"BB",X"99",X"00",X"77",X"BB",X"91",
		X"00",X"77",X"9B",X"99",X"00",X"77",X"9B",X"B9",X"00",X"99",X"9B",X"19",X"00",X"77",X"9B",X"99",
		X"09",X"77",X"99",X"BB",X"99",X"77",X"B9",X"BB",X"BB",X"77",X"BB",X"BB",X"BB",X"99",X"99",X"99",
		X"BB",X"00",X"B9",X"90",X"9B",X"00",X"BB",X"00",X"99",X"99",X"BB",X"09",X"09",X"B9",X"BB",X"99",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"9B",X"BB",X"09",X"99",X"99",X"B9",X"99",X"90",X"09",X"99",
		X"9B",X"90",X"00",X"99",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"99",X"00",X"00",X"99",
		X"09",X"11",X"79",X"B9",X"09",X"99",X"79",X"B9",X"99",X"BB",X"79",X"B9",X"9B",X"BB",X"99",X"99",
		X"9B",X"BB",X"BB",X"90",X"99",X"99",X"BB",X"90",X"99",X"BB",X"BB",X"00",X"99",X"BB",X"B9",X"00",
		X"09",X"99",X"99",X"00",X"09",X"9B",X"BB",X"00",X"00",X"99",X"BB",X"09",X"00",X"11",X"BB",X"99",
		X"00",X"77",X"BB",X"9B",X"00",X"77",X"BB",X"9B",X"00",X"77",X"BB",X"BB",X"00",X"99",X"BB",X"BB",
		X"00",X"77",X"BB",X"BB",X"00",X"77",X"BB",X"BB",X"00",X"77",X"BB",X"BB",X"00",X"77",X"BB",X"BB",
		X"00",X"99",X"99",X"99",X"00",X"09",X"BB",X"90",X"00",X"09",X"BB",X"00",X"00",X"09",X"B9",X"00",
		X"00",X"99",X"B9",X"00",X"00",X"BB",X"B9",X"00",X"00",X"BB",X"B9",X"00",X"09",X"99",X"BB",X"00",
		X"09",X"BB",X"BB",X"00",X"09",X"BB",X"BB",X"00",X"09",X"BB",X"BB",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"96",X"99",X"00",
		X"00",X"66",X"66",X"00",X"00",X"69",X"66",X"00",X"00",X"69",X"66",X"00",X"00",X"66",X"66",X"00",
		X"90",X"96",X"66",X"00",X"99",X"96",X"66",X"90",X"99",X"96",X"66",X"90",X"E9",X"99",X"96",X"99",
		X"9E",X"E9",X"C9",X"69",X"EE",X"E9",X"C9",X"66",X"9E",X"EE",X"C9",X"66",X"99",X"99",X"99",X"66",
		X"CC",X"94",X"9E",X"66",X"9C",X"44",X"EE",X"66",X"49",X"94",X"9E",X"66",X"44",X"94",X"99",X"66",
		X"94",X"99",X"C9",X"66",X"99",X"9C",X"C9",X"66",X"99",X"99",X"99",X"66",X"99",X"99",X"99",X"66",
		X"99",X"F9",X"C9",X"66",X"C9",X"F9",X"99",X"66",X"C9",X"99",X"9D",X"66",X"C9",X"99",X"DD",X"66",
		X"99",X"99",X"6D",X"66",X"09",X"9C",X"2D",X"66",X"09",X"CC",X"6D",X"66",X"09",X"99",X"6D",X"66",
		X"00",X"99",X"90",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"69",X"00",X"00",X"69",X"69",X"00",
		X"00",X"69",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"96",X"66",X"00",X"99",X"96",X"66",X"90",
		X"E9",X"96",X"66",X"90",X"E9",X"66",X"96",X"99",X"9E",X"99",X"C9",X"69",X"9E",X"E9",X"C9",X"66",
		X"9E",X"EE",X"C9",X"66",X"9E",X"99",X"99",X"66",X"99",X"94",X"9E",X"66",X"CC",X"94",X"EE",X"66",
		X"99",X"94",X"9E",X"66",X"49",X"44",X"99",X"66",X"94",X"99",X"C9",X"66",X"99",X"9C",X"C9",X"66",
		X"99",X"99",X"99",X"66",X"99",X"99",X"99",X"66",X"99",X"F9",X"C9",X"66",X"C9",X"F9",X"99",X"66",
		X"C9",X"99",X"9D",X"66",X"CC",X"99",X"DD",X"66",X"99",X"9C",X"6D",X"66",X"09",X"CC",X"2D",X"66",
		X"09",X"99",X"6D",X"66",X"09",X"DD",X"6D",X"66",X"09",X"66",X"6D",X"66",X"09",X"66",X"6D",X"66",
		X"09",X"66",X"6D",X"66",X"09",X"66",X"6D",X"66",X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",
		X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",X"09",X"99",X"66",X"66",X"09",X"59",X"99",X"66",
		X"09",X"59",X"DD",X"66",X"09",X"59",X"DD",X"66",X"09",X"59",X"DD",X"66",X"09",X"59",X"99",X"66",
		X"09",X"99",X"66",X"66",X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",
		X"09",X"66",X"99",X"66",X"09",X"D6",X"99",X"66",X"09",X"66",X"D9",X"66",X"99",X"66",X"DD",X"66",
		X"99",X"69",X"66",X"66",X"99",X"69",X"66",X"99",X"99",X"99",X"66",X"CC",X"99",X"99",X"66",X"CC",
		X"79",X"99",X"69",X"9C",X"77",X"00",X"99",X"9C",X"77",X"00",X"77",X"9C",X"99",X"00",X"77",X"9C",
		X"77",X"00",X"77",X"9C",X"77",X"00",X"97",X"9C",X"97",X"00",X"77",X"CC",X"99",X"00",X"99",X"99",
		X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",
		X"09",X"99",X"66",X"66",X"09",X"59",X"99",X"66",X"09",X"59",X"DD",X"66",X"09",X"59",X"DD",X"66",
		X"09",X"59",X"DD",X"66",X"09",X"59",X"99",X"66",X"09",X"99",X"66",X"66",X"09",X"66",X"66",X"66",
		X"09",X"66",X"66",X"66",X"09",X"66",X"66",X"66",X"09",X"66",X"99",X"66",X"09",X"66",X"90",X"66",
		X"09",X"99",X"00",X"66",X"09",X"D9",X"00",X"66",X"99",X"D9",X"00",X"66",X"9C",X"D9",X"00",X"99",
		X"CC",X"96",X"00",X"CC",X"C9",X"96",X"00",X"CC",X"99",X"96",X"09",X"CC",X"99",X"96",X"99",X"CC",
		X"09",X"99",X"9C",X"CC",X"99",X"77",X"CC",X"CC",X"97",X"77",X"C9",X"9C",X"97",X"77",X"99",X"9C",
		X"99",X"77",X"00",X"99",X"00",X"99",X"99",X"90",X"00",X"90",X"9C",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"09",X"E9",X"00",X"00",X"09",X"EE",X"00",X"00",X"99",X"9E",X"00",X"00",X"9E",X"99",X"00",
		X"00",X"99",X"E9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"00",X"9E",X"99",X"00",X"00",X"EE",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9E",X"99",X"90",X"00",X"9E",X"99",X"90",X"00",X"9E",X"99",X"90",
		X"99",X"99",X"9E",X"00",X"9E",X"BB",X"9E",X"99",X"9E",X"9E",X"99",X"E9",X"09",X"9B",X"99",X"E4",
		X"99",X"99",X"99",X"9E",X"9E",X"9E",X"99",X"99",X"E9",X"EE",X"99",X"9E",X"9E",X"99",X"99",X"9E",
		X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"09",X"E9",X"00",X"00",X"09",X"EE",X"00",
		X"00",X"99",X"9E",X"00",X"00",X"9E",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"E9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"00",X"99",X"A9",X"00",
		X"00",X"9E",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"90",
		X"00",X"9E",X"99",X"90",X"00",X"9E",X"99",X"90",X"99",X"99",X"99",X"00",X"9E",X"BB",X"9E",X"99",
		X"9E",X"9E",X"99",X"E9",X"09",X"9B",X"9E",X"E4",X"99",X"99",X"EE",X"9E",X"9E",X"9E",X"E9",X"99",
		X"E9",X"EE",X"99",X"9E",X"9E",X"99",X"99",X"9E",X"99",X"E9",X"99",X"EE",X"09",X"E9",X"99",X"EE",
		X"E9",X"99",X"99",X"99",X"9E",X"E9",X"99",X"E9",X"9E",X"99",X"99",X"E9",X"99",X"9E",X"E9",X"99",
		X"E9",X"9E",X"99",X"E9",X"99",X"99",X"E9",X"EB",X"E9",X"9E",X"E9",X"9B",X"9E",X"9E",X"E9",X"9E",
		X"99",X"99",X"9B",X"E9",X"9E",X"E9",X"99",X"E9",X"9E",X"E9",X"99",X"E9",X"99",X"EE",X"99",X"9E",
		X"09",X"9E",X"99",X"E4",X"00",X"99",X"99",X"9E",X"00",X"EE",X"99",X"99",X"00",X"49",X"9B",X"EE",
		X"00",X"E9",X"99",X"99",X"00",X"E9",X"99",X"00",X"00",X"E9",X"9E",X"00",X"00",X"99",X"9E",X"00",
		X"00",X"9E",X"99",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"9E",X"00",X"00",X"99",X"9E",X"00",
		X"09",X"BB",X"99",X"00",X"99",X"BB",X"EE",X"90",X"9E",X"99",X"EE",X"99",X"9E",X"E9",X"99",X"E9",
		X"EE",X"99",X"EE",X"E9",X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"9E",X"99",X"EE",X"9E",X"99",X"99",X"9E",X"E9",X"99",X"99",X"99",X"9E",X"E9",X"99",X"99",
		X"9E",X"99",X"9E",X"E9",X"99",X"9E",X"9E",X"90",X"09",X"99",X"9E",X"00",X"09",X"9E",X"E9",X"00",
		X"09",X"9E",X"E9",X"00",X"09",X"E9",X"E9",X"00",X"99",X"99",X"EB",X"00",X"9E",X"E9",X"E9",X"00",
		X"9E",X"E9",X"99",X"00",X"9E",X"EE",X"99",X"00",X"9E",X"9E",X"EE",X"00",X"9E",X"9E",X"99",X"90",
		X"E9",X"99",X"9E",X"90",X"E9",X"00",X"9E",X"90",X"BB",X"00",X"9E",X"00",X"B9",X"00",X"9E",X"99",
		X"99",X"00",X"99",X"E9",X"E9",X"00",X"9B",X"9E",X"E9",X"00",X"99",X"9E",X"99",X"90",X"09",X"9E",
		X"09",X"90",X"09",X"EE",X"99",X"99",X"00",X"EE",X"E9",X"9E",X"00",X"9E",X"E9",X"9E",X"00",X"99",
		X"E9",X"9E",X"09",X"B9",X"99",X"EE",X"99",X"B9",X"EE",X"E9",X"9E",X"B9",X"99",X"99",X"99",X"99",
		X"90",X"00",X"99",X"00",X"99",X"00",X"49",X"99",X"A9",X"00",X"49",X"97",X"A9",X"00",X"99",X"99",
		X"9A",X"90",X"77",X"79",X"9A",X"94",X"99",X"77",X"99",X"99",X"99",X"77",X"09",X"79",X"99",X"99",
		X"09",X"77",X"99",X"99",X"09",X"77",X"77",X"99",X"99",X"97",X"97",X"99",X"97",X"97",X"99",X"77",
		X"97",X"99",X"49",X"77",X"79",X"99",X"49",X"99",X"79",X"99",X"09",X"00",X"77",X"97",X"09",X"00",
		X"97",X"77",X"09",X"00",X"99",X"99",X"09",X"00",X"09",X"99",X"09",X"00",X"09",X"99",X"99",X"00",
		X"09",X"09",X"79",X"00",X"09",X"99",X"79",X"00",X"00",X"97",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"79",X"77",X"90",
		X"00",X"99",X"77",X"99",X"09",X"11",X"77",X"79",X"09",X"11",X"97",X"77",X"09",X"99",X"99",X"77",
		X"00",X"00",X"00",X"99",X"90",X"00",X"90",X"39",X"90",X"00",X"99",X"39",X"90",X"00",X"97",X"99",
		X"99",X"00",X"97",X"77",X"A9",X"00",X"77",X"77",X"AA",X"90",X"79",X"77",X"A9",X"90",X"99",X"77",
		X"A9",X"94",X"77",X"79",X"99",X"99",X"97",X"79",X"99",X"79",X"99",X"99",X"33",X"79",X"09",X"94",
		X"99",X"77",X"09",X"40",X"77",X"77",X"00",X"40",X"77",X"77",X"00",X"40",X"77",X"77",X"00",X"40",
		X"79",X"97",X"00",X"40",X"79",X"97",X"00",X"00",X"99",X"97",X"00",X"00",X"90",X"77",X"00",X"00",
		X"00",X"77",X"09",X"00",X"00",X"77",X"09",X"00",X"00",X"77",X"99",X"00",X"00",X"77",X"97",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"79",X"77",X"90",
		X"00",X"99",X"77",X"99",X"09",X"11",X"77",X"79",X"09",X"11",X"97",X"77",X"09",X"99",X"99",X"77",
		X"09",X"19",X"99",X"77",X"99",X"19",X"94",X"77",X"97",X"11",X"94",X"77",X"97",X"99",X"94",X"97",
		X"97",X"49",X"19",X"97",X"9E",X"49",X"99",X"9E",X"9E",X"44",X"49",X"99",X"97",X"99",X"99",X"79",
		X"97",X"19",X"19",X"79",X"97",X"19",X"99",X"79",X"97",X"19",X"97",X"79",X"99",X"99",X"97",X"39",
		X"00",X"19",X"97",X"79",X"00",X"19",X"77",X"79",X"09",X"19",X"77",X"77",X"09",X"99",X"77",X"77",
		X"09",X"91",X"77",X"77",X"09",X"99",X"77",X"97",X"09",X"91",X"77",X"99",X"09",X"91",X"99",X"00",
		X"09",X"19",X"90",X"00",X"09",X"19",X"99",X"00",X"09",X"99",X"79",X"00",X"09",X"94",X"79",X"00",
		X"09",X"94",X"79",X"09",X"00",X"99",X"77",X"99",X"00",X"91",X"77",X"97",X"00",X"91",X"77",X"37",
		X"00",X"49",X"77",X"77",X"00",X"49",X"97",X"77",X"00",X"91",X"99",X"77",X"00",X"99",X"99",X"99",
		X"09",X"19",X"99",X"77",X"99",X"19",X"94",X"77",X"97",X"11",X"94",X"77",X"97",X"99",X"94",X"97",
		X"97",X"49",X"19",X"99",X"9E",X"49",X"99",X"E9",X"7E",X"44",X"49",X"EE",X"79",X"99",X"99",X"7E",
		X"99",X"19",X"19",X"77",X"00",X"19",X"99",X"77",X"00",X"19",X"97",X"77",X"00",X"99",X"97",X"77",
		X"00",X"19",X"97",X"77",X"00",X"19",X"77",X"99",X"09",X"19",X"77",X"00",X"09",X"99",X"77",X"00",
		X"09",X"91",X"77",X"00",X"09",X"99",X"77",X"00",X"09",X"91",X"77",X"00",X"09",X"91",X"99",X"09",
		X"09",X"19",X"90",X"99",X"09",X"19",X"99",X"97",X"09",X"99",X"79",X"77",X"09",X"94",X"77",X"77",
		X"09",X"94",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"91",X"77",X"79",X"00",X"91",X"77",X"99",
		X"00",X"49",X"77",X"00",X"00",X"49",X"97",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"49",X"99",X"99",X"49",X"49",X"99",X"99",X"49",X"49",X"99",X"99",X"44",X"49",X"99",
		X"99",X"94",X"99",X"99",X"99",X"99",X"92",X"99",X"09",X"29",X"22",X"99",X"99",X"22",X"22",X"99",
		X"99",X"92",X"22",X"99",X"99",X"92",X"22",X"99",X"99",X"92",X"22",X"99",X"9D",X"92",X"29",X"99",
		X"99",X"92",X"29",X"99",X"99",X"92",X"29",X"99",X"99",X"92",X"29",X"99",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"90",
		X"00",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"49",X"99",X"99",X"49",X"49",X"99",X"99",X"49",X"49",X"99",X"99",X"44",X"49",X"99",
		X"99",X"94",X"99",X"99",X"99",X"29",X"92",X"99",X"09",X"29",X"22",X"99",X"99",X"22",X"22",X"99",
		X"99",X"92",X"22",X"99",X"99",X"92",X"22",X"99",X"99",X"92",X"22",X"99",X"9D",X"92",X"29",X"99",
		X"99",X"92",X"29",X"99",X"99",X"92",X"29",X"99",X"99",X"92",X"29",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"92",X"09",X"99",X"99",X"22",
		X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"92",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"D9",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"99",X"99",X"99",X"22",X"99",X"22",X"90",
		X"22",X"99",X"22",X"00",X"29",X"99",X"22",X"00",X"29",X"99",X"22",X"00",X"99",X"99",X"22",X"00",
		X"09",X"99",X"92",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"90",X"09",X"99",X"99",X"90",X"09",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"95",X"95",X"00",X"00",X"95",X"55",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"59",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"EE",X"EE",X"90",X"09",X"9E",X"99",X"90",X"09",X"E3",X"E9",X"90",X"00",X"99",X"93",X"00",
		X"00",X"FF",X"99",X"00",X"00",X"A9",X"F9",X"00",X"00",X"A9",X"FF",X"00",X"00",X"F9",X"F9",X"00",
		X"00",X"FF",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"33",X"00",
		X"00",X"33",X"99",X"00",X"00",X"39",X"93",X"00",X"99",X"33",X"93",X"00",X"93",X"33",X"93",X"00",
		X"93",X"33",X"39",X"00",X"99",X"33",X"99",X"00",X"33",X"93",X"33",X"00",X"99",X"99",X"99",X"00",
		X"00",X"99",X"93",X"00",X"00",X"99",X"93",X"00",X"00",X"93",X"33",X"00",X"00",X"93",X"39",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"93",X"99",X"00",
		X"00",X"33",X"99",X"00",X"00",X"39",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"90",X"99",X"00",
		X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"90",X"99",X"00",X"00",X"99",
		X"99",X"00",X"00",X"99",X"99",X"09",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"D9",X"9D",X"99",
		X"99",X"D9",X"9D",X"99",X"99",X"D9",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"D9",X"9D",X"99",X"99",X"D9",X"9D",X"99",
		X"09",X"99",X"99",X"99",X"09",X"D9",X"9D",X"99",X"00",X"9D",X"D9",X"99",X"00",X"9D",X"D9",X"99",
		X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"90",X"09",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"09",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"D9",X"9D",X"99",X"99",X"99",X"9D",X"99",
		X"99",X"D9",X"99",X"99",X"99",X"D9",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"D9",X"99",
		X"99",X"D9",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",X"09",X"09",X"09",X"09",X"00",X"00",X"09",
		X"09",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"9D",X"90",X"99",X"99",X"9D",X"90",X"99",X"99",X"9D",X"90",
		X"99",X"99",X"99",X"90",X"99",X"D9",X"D9",X"90",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0A",X"FF",X"00",X"00",X"0A",X"FF",X"00",X"00",X"0A",X"AA",X"00",
		X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"0A",X"FA",X"00",X"00",X"AF",X"FA",X"AA",X"00",X"AF",X"FF",X"FF",
		X"00",X"FF",X"AA",X"FF",X"00",X"FA",X"AF",X"FF",X"00",X"FA",X"FF",X"FA",X"00",X"AA",X"FF",X"FA",
		X"00",X"FF",X"AA",X"FA",X"00",X"FF",X"FA",X"FF",X"00",X"FF",X"FA",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"AF",X"AA",X"00",X"FF",X"AF",X"AF",X"00",X"FF",X"AF",X"AF",
		X"00",X"AA",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FA",X"FF",X"00",X"AA",X"FF",X"FF",
		X"00",X"AF",X"FF",X"FF",X"00",X"FF",X"AF",X"FF",X"00",X"FF",X"AA",X"FF",X"00",X"AA",X"FF",X"FF",
		X"00",X"AF",X"FF",X"FF",X"00",X"FF",X"FF",X"AF",X"00",X"FF",X"FF",X"0A",X"00",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"0A",X"00",X"00",X"AF",X"0A",X"00",X"00",X"AF",
		X"AA",X"00",X"00",X"AF",X"FF",X"00",X"00",X"FF",X"AF",X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",
		X"AF",X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",X"00",X"00",X"00",X"AA",X"00",X"00",X"A0",X"AA",
		X"00",X"00",X"A0",X"A0",X"00",X"00",X"A0",X"00",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"AF",X"A0",X"00",X"AA",
		X"AF",X"A0",X"00",X"FA",X"FF",X"AA",X"00",X"FF",X"FF",X"FA",X"00",X"FF",X"AA",X"FA",X"00",X"FF",
		X"00",X"FA",X"00",X"FA",X"00",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"0A",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"F0",X"0A",X"00",X"0F",X"3F",X"00",
		X"00",X"0F",X"0F",X"00",X"AA",X"0F",X"0F",X"0A",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"03",X"F3",X"00",X"00",X"00",X"30",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"A0",X"00",X"0A",X"00",X"0A",
		X"0A",X"A0",X"00",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"09",X"9F",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",
		X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",
		X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"95",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"09",X"9F",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"9F",X"FF",X"00",X"00",X"99",X"9F",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"9F",X"F9",X"00",X"00",X"9F",X"99",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",
		X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"95",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"09",X"9F",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"9F",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"9F",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"F9",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"95",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9F",X"00",X"00",X"0E",X"9F",X"00",X"19",X"5E",X"9F",X"40",X"99",X"99",X"99",
		X"00",X"91",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"39",X"99",X"00",
		X"06",X"97",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9A",X"01",X"00",X"39",X"99",X"00",
		X"70",X"00",X"99",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"99",X"09",X"00",X"09",X"29",X"99",
		X"00",X"09",X"20",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"09",X"90",X"00",X"90",X"99",X"00",
		X"09",X"90",X"49",X"99",X"99",X"99",X"49",X"9A",X"9A",X"59",X"49",X"AA",X"9A",X"55",X"44",X"A3",
		X"A3",X"95",X"49",X"53",X"AA",X"99",X"9A",X"33",X"AA",X"AA",X"A9",X"3A",X"33",X"3A",X"AA",X"AA",
		X"AA",X"AA",X"99",X"53",X"A3",X"3A",X"99",X"33",X"33",X"A9",X"44",X"3A",X"3A",X"99",X"44",X"33",
		X"3A",X"94",X"99",X"A3",X"3A",X"94",X"F9",X"A3",X"AA",X"94",X"F9",X"A3",X"AA",X"94",X"F9",X"A3",
		X"A3",X"99",X"F9",X"AA",X"A3",X"99",X"A9",X"9A",X"A3",X"09",X"99",X"99",X"A3",X"09",X"49",X"09",
		X"AA",X"99",X"94",X"09",X"3A",X"95",X"99",X"09",X"3A",X"59",X"09",X"09",X"A9",X"99",X"99",X"09",
		X"99",X"95",X"95",X"90",X"90",X"99",X"99",X"90",X"90",X"95",X"00",X"00",X"90",X"99",X"00",X"00",
		X"00",X"99",X"00",X"90",X"00",X"9A",X"00",X"90",X"00",X"93",X"09",X"00",X"00",X"9A",X"99",X"00",
		X"00",X"9A",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"59",X"49",X"00",X"00",X"55",X"44",X"00",
		X"00",X"95",X"49",X"00",X"00",X"99",X"9A",X"00",X"00",X"AA",X"A9",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"3A",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"A9",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"94",X"99",X"00",X"00",X"94",X"F9",X"00",X"00",X"94",X"F9",X"00",X"00",X"94",X"F9",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"A9",X"49",X"00",
		X"00",X"99",X"94",X"00",X"00",X"95",X"99",X"00",X"00",X"59",X"09",X"00",X"00",X"95",X"99",X"00",
		X"00",X"95",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"59",X"49",X"00",X"00",X"55",X"44",X"00",
		X"00",X"9A",X"49",X"00",X"00",X"99",X"9A",X"00",X"00",X"A3",X"AA",X"90",X"00",X"AA",X"AA",X"90",
		X"00",X"3A",X"99",X"90",X"00",X"AA",X"99",X"99",X"00",X"A9",X"44",X"A9",X"00",X"99",X"44",X"A9",
		X"00",X"94",X"99",X"A9",X"00",X"94",X"F9",X"A9",X"00",X"94",X"F9",X"A9",X"00",X"94",X"F9",X"A9",
		X"00",X"99",X"A9",X"A9",X"00",X"99",X"99",X"A9",X"00",X"A9",X"99",X"99",X"00",X"A9",X"49",X"90",
		X"00",X"99",X"94",X"90",X"00",X"95",X"99",X"90",X"00",X"59",X"09",X"90",X"00",X"95",X"99",X"90",
		X"00",X"95",X"95",X"90",X"00",X"99",X"99",X"00",X"00",X"9A",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"94",X"44",X"00",
		X"00",X"49",X"99",X"00",X"00",X"99",X"22",X"90",X"00",X"92",X"92",X"99",X"99",X"22",X"99",X"49",
		X"91",X"99",X"A9",X"11",X"11",X"99",X"A2",X"11",X"91",X"99",X"9A",X"11",X"EE",X"11",X"11",X"59",
		X"9E",X"11",X"11",X"EE",X"99",X"11",X"11",X"E9",X"00",X"EE",X"EE",X"99",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"94",X"44",X"00",
		X"00",X"49",X"94",X"00",X"00",X"92",X"22",X"90",X"00",X"22",X"92",X"99",X"99",X"29",X"99",X"49",
		X"91",X"99",X"A9",X"11",X"11",X"99",X"A2",X"11",X"91",X"99",X"9A",X"11",X"EE",X"11",X"11",X"79",
		X"9E",X"11",X"11",X"EE",X"99",X"11",X"11",X"E9",X"00",X"EE",X"EE",X"99",X"00",X"99",X"99",X"00",
		X"00",X"00",X"E0",X"99",X"00",X"00",X"EE",X"93",X"00",X"00",X"E9",X"93",X"00",X"09",X"99",X"33",
		X"00",X"99",X"9F",X"33",X"00",X"93",X"9F",X"39",X"00",X"93",X"9F",X"39",X"00",X"93",X"9F",X"99",
		X"00",X"93",X"9F",X"90",X"00",X"99",X"9F",X"90",X"00",X"39",X"9F",X"90",X"00",X"99",X"99",X"90",
		X"77",X"93",X"93",X"00",X"00",X"93",X"33",X"90",X"00",X"9B",X"93",X"90",X"00",X"9B",X"33",X"90",
		X"00",X"99",X"93",X"90",X"00",X"09",X"99",X"90",X"00",X"A5",X"99",X"00",X"40",X"99",X"70",X"00",
		X"40",X"99",X"99",X"00",X"00",X"59",X"99",X"1A",X"00",X"99",X"B9",X"AA",X"0A",X"43",X"B4",X"90",
		X"00",X"44",X"34",X"95",X"55",X"A4",X"B5",X"11",X"04",X"99",X"95",X"90",X"00",X"1A",X"44",X"90",
		X"00",X"91",X"59",X"11",X"00",X"99",X"59",X"00",X"70",X"00",X"05",X"05",X"00",X"50",X"00",X"05",
		X"00",X"0E",X"00",X"00",X"00",X"09",X"E9",X"99",X"00",X"0E",X"EE",X"93",X"00",X"09",X"EE",X"93",
		X"00",X"99",X"39",X"33",X"00",X"93",X"99",X"39",X"00",X"93",X"9F",X"39",X"00",X"93",X"9F",X"99",
		X"00",X"93",X"9F",X"90",X"00",X"99",X"9F",X"90",X"00",X"39",X"99",X"90",X"00",X"99",X"39",X"90",
		X"00",X"93",X"33",X"00",X"00",X"93",X"93",X"90",X"00",X"9B",X"39",X"90",X"00",X"9B",X"33",X"90",
		X"00",X"99",X"93",X"90",X"00",X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"99",X"39",X"00",
		X"00",X"93",X"33",X"00",X"00",X"33",X"93",X"00",X"00",X"39",X"99",X"00",X"00",X"99",X"39",X"00",
		X"00",X"99",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"93",X"39",X"00",
		X"00",X"93",X"39",X"00",X"00",X"93",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",
		X"00",X"99",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",
		X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",
		X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"9F",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"95",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"99",X"00",
		X"99",X"BB",X"49",X"00",X"11",X"BB",X"49",X"99",X"11",X"9B",X"99",X"BB",X"1E",X"9B",X"BB",X"BB",
		X"1E",X"9B",X"9B",X"BB",X"1E",X"9B",X"99",X"BB",X"11",X"9B",X"95",X"99",X"1E",X"9B",X"95",X"99",
		X"1E",X"99",X"99",X"90",X"EE",X"E9",X"99",X"00",X"E1",X"99",X"94",X"99",X"E1",X"9B",X"99",X"BB",
		X"E1",X"BB",X"BB",X"99",X"E1",X"BB",X"99",X"09",X"E1",X"B9",X"77",X"00",X"E1",X"99",X"77",X"00",
		X"E1",X"9B",X"B7",X"00",X"E1",X"99",X"BB",X"00",X"E1",X"09",X"BB",X"00",X"11",X"09",X"BB",X"00",
		X"99",X"09",X"BB",X"09",X"90",X"00",X"BB",X"99",X"90",X"00",X"BB",X"9B",X"90",X"00",X"B9",X"BB",
		X"90",X"00",X"99",X"BB",X"00",X"00",X"90",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"00",X"91",X"90",X"99",X"00",X"91",X"99",X"99",X"00",X"9E",X"B9",X"99",X"00",
		X"9E",X"BB",X"49",X"00",X"9E",X"BB",X"49",X"99",X"91",X"9B",X"99",X"BB",X"91",X"9B",X"BB",X"BB",
		X"91",X"9B",X"9B",X"BB",X"91",X"9B",X"99",X"BB",X"91",X"9B",X"95",X"99",X"91",X"9B",X"95",X"99",
		X"91",X"99",X"99",X"90",X"91",X"19",X"BB",X"99",X"99",X"99",X"BB",X"BB",X"09",X"9B",X"99",X"BB",
		X"01",X"BB",X"77",X"99",X"09",X"9B",X"77",X"00",X"09",X"99",X"77",X"00",X"00",X"19",X"77",X"00",
		X"00",X"9B",X"B7",X"00",X"00",X"99",X"BB",X"00",X"00",X"09",X"BB",X"00",X"00",X"09",X"BB",X"00",
		X"00",X"09",X"BB",X"09",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B9",X"BB",
		X"00",X"00",X"99",X"BB",X"00",X"00",X"90",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"96",X"66",X"00",
		X"00",X"66",X"99",X"00",X"09",X"99",X"96",X"00",X"09",X"E9",X"66",X"00",X"09",X"EE",X"96",X"00",
		X"00",X"9E",X"96",X"00",X"00",X"99",X"96",X"00",X"09",X"99",X"96",X"00",X"09",X"9C",X"96",X"00",
		X"09",X"C9",X"96",X"00",X"09",X"99",X"96",X"00",X"09",X"95",X"96",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"9C",X"66",X"00",X"00",X"CC",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"00",X"99",X"66",X"00",X"09",X"96",X"69",X"00",X"09",X"99",X"69",X"00",
		X"09",X"09",X"96",X"00",X"00",X"09",X"96",X"00",X"00",X"09",X"96",X"00",X"00",X"99",X"66",X"00",
		X"00",X"77",X"99",X"00",X"00",X"77",X"77",X"00",X"00",X"99",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"69",X"00",X"00",X"96",X"66",X"00",
		X"09",X"99",X"99",X"00",X"09",X"E9",X"96",X"00",X"09",X"EE",X"66",X"00",X"00",X"99",X"96",X"00",
		X"00",X"49",X"96",X"00",X"09",X"99",X"96",X"00",X"09",X"9C",X"96",X"00",X"09",X"C9",X"96",X"00",
		X"09",X"99",X"96",X"00",X"09",X"95",X"96",X"00",X"09",X"99",X"96",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"96",X"00",X"00",X"CC",X"96",X"00",
		X"00",X"99",X"96",X"00",X"00",X"99",X"96",X"00",X"00",X"96",X"96",X"00",X"00",X"66",X"96",X"00",
		X"00",X"66",X"99",X"99",X"00",X"66",X"9C",X"99",X"00",X"66",X"CC",X"66",X"00",X"99",X"9C",X"66",
		X"00",X"77",X"99",X"66",X"00",X"77",X"00",X"99",X"00",X"99",X"00",X"77",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"E9",X"99",X"99",
		X"9E",X"E9",X"9E",X"E9",X"9E",X"E9",X"EE",X"99",X"99",X"99",X"EE",X"9E",X"09",X"9E",X"99",X"9E",
		X"99",X"9E",X"99",X"9E",X"E9",X"E9",X"79",X"9E",X"E9",X"99",X"99",X"99",X"9E",X"99",X"99",X"E9",
		X"19",X"99",X"99",X"E9",X"99",X"E9",X"E9",X"E9",X"90",X"99",X"E9",X"9E",X"00",X"E9",X"E9",X"99",
		X"00",X"E9",X"9E",X"09",X"00",X"EE",X"9E",X"00",X"00",X"99",X"9E",X"00",X"00",X"9E",X"99",X"00",
		X"00",X"9E",X"B9",X"00",X"09",X"E1",X"99",X"99",X"09",X"91",X"E9",X"9E",X"99",X"99",X"E9",X"EE",
		X"9E",X"E9",X"99",X"99",X"19",X"E9",X"EE",X"91",X"1E",X"99",X"99",X"94",X"99",X"00",X"09",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"E9",X"99",X"00",
		X"00",X"E9",X"9E",X"00",X"00",X"E9",X"EE",X"00",X"00",X"99",X"EE",X"90",X"00",X"9E",X"99",X"99",
		X"99",X"99",X"99",X"E9",X"EB",X"99",X"99",X"E9",X"9B",X"99",X"79",X"EE",X"9E",X"99",X"99",X"9E",
		X"99",X"99",X"99",X"99",X"19",X"99",X"99",X"E9",X"99",X"99",X"E9",X"99",X"E9",X"E9",X"E9",X"E9",
		X"11",X"E9",X"9E",X"EE",X"99",X"EE",X"9E",X"B9",X"00",X"99",X"9E",X"99",X"09",X"9E",X"99",X"09",
		X"09",X"9E",X"E9",X"09",X"99",X"EE",X"E9",X"00",X"E9",X"99",X"99",X"99",X"99",X"9E",X"9E",X"EE",
		X"9E",X"BE",X"E9",X"E9",X"9E",X"B9",X"99",X"99",X"99",X"E9",X"09",X"E9",X"00",X"99",X"00",X"99",
		X"99",X"99",X"99",X"99",X"39",X"79",X"97",X"39",X"99",X"77",X"97",X"99",X"97",X"77",X"77",X"99",
		X"77",X"77",X"77",X"77",X"79",X"77",X"77",X"77",X"79",X"77",X"77",X"99",X"99",X"97",X"77",X"99",
		X"99",X"97",X"77",X"90",X"90",X"99",X"77",X"90",X"90",X"97",X"77",X"99",X"09",X"97",X"77",X"77",
		X"99",X"97",X"77",X"77",X"97",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"79",X"97",X"77",X"77",X"79",X"97",X"77",X"77",X"79",X"97",X"79",X"74",X"79",X"97",X"49",
		X"94",X"97",X"99",X"49",X"9A",X"97",X"19",X"A9",X"99",X"09",X"99",X"99",X"99",X"09",X"44",X"79",
		X"90",X"00",X"99",X"79",X"00",X"00",X"11",X"79",X"00",X"00",X"99",X"79",X"00",X"00",X"00",X"79",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",
		X"99",X"99",X"99",X"99",X"39",X"79",X"97",X"39",X"39",X"77",X"97",X"39",X"97",X"77",X"77",X"99",
		X"97",X"77",X"77",X"79",X"79",X"77",X"79",X"77",X"79",X"77",X"79",X"99",X"99",X"97",X"79",X"99",
		X"99",X"97",X"77",X"90",X"90",X"99",X"77",X"90",X"90",X"97",X"77",X"90",X"00",X"97",X"77",X"00",
		X"00",X"97",X"77",X"90",X"00",X"77",X"77",X"90",X"00",X"77",X"77",X"99",X"00",X"77",X"77",X"79",
		X"00",X"79",X"97",X"79",X"00",X"79",X"97",X"77",X"00",X"79",X"97",X"77",X"00",X"79",X"97",X"77",
		X"00",X"97",X"99",X"77",X"00",X"97",X"19",X"77",X"00",X"99",X"99",X"49",X"00",X"79",X"44",X"49",
		X"00",X"79",X"99",X"79",X"00",X"99",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",
		X"99",X"90",X"00",X"00",X"99",X"99",X"09",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"29",X"90",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"49",X"00",
		X"99",X"99",X"99",X"90",X"92",X"99",X"99",X"99",X"92",X"99",X"99",X"90",X"92",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"22",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"99",X"09",X"99",X"09",X"99",X"09",X"29",X"99",X"99",X"00",X"29",X"92",X"90",
		X"00",X"29",X"29",X"90",X"00",X"29",X"99",X"90",X"00",X"99",X"94",X"00",X"00",X"99",X"94",X"00",
		X"00",X"29",X"44",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"22",X"00",X"99",X"59",X"92",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"59",X"99",
		X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"92",X"99",X"99",X"90",X"92",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"00",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"93",X"92",X"00",
		X"00",X"94",X"92",X"09",X"00",X"29",X"22",X"09",X"00",X"92",X"22",X"09",X"00",X"92",X"22",X"09",
		X"99",X"22",X"22",X"99",X"29",X"99",X"22",X"92",X"29",X"95",X"92",X"A2",X"29",X"99",X"92",X"22",
		X"22",X"99",X"92",X"29",X"2A",X"99",X"22",X"99",X"92",X"59",X"99",X"DD",X"99",X"99",X"92",X"22",
		X"9D",X"22",X"22",X"D2",X"9D",X"92",X"22",X"DD",X"9D",X"99",X"A2",X"2D",X"99",X"99",X"22",X"D2",
		X"09",X"92",X"22",X"D9",X"09",X"92",X"22",X"99",X"09",X"99",X"2A",X"00",X"00",X"D9",X"22",X"00",
		X"00",X"D9",X"22",X"00",X"00",X"99",X"92",X"90",X"00",X"22",X"22",X"90",X"00",X"29",X"22",X"90",
		X"00",X"29",X"92",X"90",X"00",X"29",X"99",X"90",X"00",X"22",X"00",X"90",X"00",X"99",X"00",X"90",
		X"00",X"9D",X"00",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"94",X"92",X"00",
		X"00",X"99",X"92",X"00",X"00",X"29",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"95",X"92",X"00",X"00",X"99",X"92",X"00",
		X"00",X"59",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"DD",X"00",
		X"00",X"9D",X"DD",X"00",X"00",X"99",X"DD",X"00",X"00",X"DD",X"D2",X"00",X"00",X"2D",X"2D",X"00",
		X"00",X"D2",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"2D",X"DD",X"00",X"00",X"D2",X"92",X"00",
		X"00",X"DD",X"9D",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"29",X"00",X"00",X"9D",X"22",X"00",
		X"00",X"99",X"22",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"09",X"E9",X"99",X"00",X"0E",X"EE",X"93",X"00",X"09",X"EE",X"93",
		X"00",X"99",X"39",X"33",X"00",X"93",X"99",X"39",X"00",X"93",X"9F",X"39",X"00",X"93",X"9F",X"99",
		X"00",X"93",X"9A",X"90",X"00",X"99",X"99",X"90",X"00",X"39",X"39",X"90",X"00",X"99",X"33",X"90",
		X"00",X"93",X"93",X"00",X"00",X"93",X"33",X"90",X"00",X"9B",X"93",X"90",X"00",X"9B",X"33",X"90",
		X"00",X"99",X"93",X"90",X"00",X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"B9",X"99",X"99",X"93",X"B9",X"49",
		X"91",X"9B",X"39",X"11",X"11",X"99",X"B9",X"11",X"91",X"99",X"99",X"11",X"EE",X"11",X"11",X"59",
		X"9E",X"11",X"11",X"EE",X"99",X"11",X"11",X"E9",X"00",X"EE",X"EE",X"99",X"00",X"99",X"99",X"00",
		X"00",X"09",X"E9",X"00",X"00",X"0E",X"EE",X"99",X"09",X"09",X"EE",X"93",X"09",X"99",X"39",X"33",
		X"09",X"93",X"99",X"39",X"00",X"93",X"9F",X"39",X"00",X"93",X"9F",X"99",X"00",X"93",X"9A",X"90",
		X"00",X"99",X"9A",X"90",X"00",X"39",X"39",X"90",X"00",X"99",X"33",X"90",X"00",X"93",X"93",X"00",
		X"00",X"93",X"33",X"90",X"00",X"93",X"93",X"90",X"00",X"9B",X"33",X"90",X"00",X"99",X"93",X"90",
		X"00",X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"33",X"00",X"00",X"99",X"B9",X"99",X"99",X"93",X"B9",X"49",
		X"91",X"9B",X"39",X"11",X"11",X"99",X"B9",X"11",X"91",X"99",X"99",X"11",X"EE",X"11",X"11",X"79",
		X"9E",X"11",X"11",X"EE",X"99",X"11",X"11",X"E9",X"00",X"EE",X"EE",X"99",X"00",X"99",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"09",X"9F",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"9F",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"44",X"00",X"00",X"99",X"49",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"F9",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"95",X"00",
		X"00",X"55",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9F",X"00",X"00",X"0E",X"9F",X"00",X"19",X"5E",X"9F",X"40",X"99",X"49",X"99",
		X"00",X"91",X"99",X"09",X"00",X"99",X"AA",X"09",X"00",X"A9",X"A9",X"09",X"00",X"3A",X"49",X"00",
		X"06",X"97",X"94",X"00",X"00",X"9A",X"9A",X"00",X"00",X"A9",X"4A",X"01",X"00",X"39",X"9A",X"00",
		X"70",X"00",X"A9",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"49",X"09",X"00",X"09",X"29",X"99",
		X"00",X"09",X"20",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"E0",X"00",X"99",X"E0",X"9E",X"90",X"93",X"EE",X"EE",X"90",X"93",X"99",X"E9",X"90",
		X"93",X"33",X"99",X"90",X"93",X"39",X"AA",X"90",X"93",X"99",X"FF",X"00",X"99",X"9A",X"99",X"00",
		X"09",X"9F",X"99",X"00",X"09",X"99",X"FF",X"00",X"00",X"39",X"99",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"39",X"93",X"00",X"00",X"39",X"33",X"00",X"09",X"B4",X"33",X"00",
		X"09",X"49",X"33",X"00",X"99",X"94",X"33",X"00",X"93",X"99",X"93",X"00",X"99",X"9B",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"39",X"99",X"00",X"00",X"39",X"39",X"00",X"99",X"33",X"33",X"00",
		X"33",X"33",X"99",X"00",X"93",X"33",X"00",X"09",X"93",X"33",X"90",X"90",X"99",X"33",X"99",X"00",
		X"93",X"33",X"33",X"90",X"93",X"33",X"39",X"09",X"99",X"93",X"99",X"00",X"99",X"99",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"90",X"00",X"99",X"39",X"90",X"00",X"49",X"39",X"99",
		X"09",X"49",X"99",X"99",X"99",X"99",X"92",X"92",X"22",X"22",X"92",X"22",X"29",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"22",X"92",X"99",X"99",X"22",X"99",X"99",X"59",X"29",
		X"95",X"99",X"59",X"29",X"99",X"99",X"59",X"29",X"00",X"99",X"59",X"99",X"09",X"95",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"22",X"99",X"90",X"29",X"29",X"22",X"99",X"22",X"22",X"DD",X"29",
		X"99",X"29",X"D2",X"29",X"99",X"99",X"29",X"2A",X"92",X"99",X"29",X"29",X"22",X"99",X"99",X"29",
		X"22",X"9A",X"99",X"29",X"29",X"99",X"92",X"99",X"29",X"99",X"92",X"90",X"29",X"22",X"92",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"90",
		X"00",X"00",X"99",X"90",X"00",X"99",X"49",X"90",X"00",X"49",X"49",X"99",X"09",X"49",X"99",X"99",
		X"99",X"99",X"92",X"92",X"22",X"22",X"92",X"22",X"29",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"99",X"22",X"92",X"99",X"99",X"22",X"99",X"99",X"59",X"29",X"95",X"99",X"59",X"29",
		X"99",X"99",X"59",X"29",X"29",X"22",X"59",X"99",X"DD",X"22",X"99",X"90",X"99",X"29",X"22",X"90",
		X"09",X"22",X"29",X"90",X"00",X"22",X"22",X"99",X"00",X"99",X"DD",X"29",X"09",X"DD",X"D2",X"29",
		X"99",X"22",X"29",X"2A",X"92",X"22",X"29",X"29",X"22",X"99",X"99",X"29",X"22",X"9A",X"99",X"29",
		X"29",X"99",X"92",X"99",X"29",X"99",X"92",X"90",X"29",X"22",X"92",X"90",X"29",X"22",X"92",X"90",
		X"29",X"22",X"92",X"90",X"29",X"99",X"92",X"99",X"29",X"9A",X"92",X"A9",X"99",X"99",X"92",X"99",
		X"92",X"99",X"92",X"90",X"92",X"22",X"92",X"90",X"92",X"22",X"92",X"90",X"92",X"22",X"92",X"00",
		X"99",X"22",X"92",X"00",X"29",X"22",X"92",X"00",X"22",X"99",X"92",X"00",X"22",X"00",X"22",X"90",
		X"29",X"00",X"22",X"90",X"99",X"00",X"99",X"90",X"29",X"00",X"99",X"00",X"22",X"00",X"29",X"00",
		X"22",X"00",X"29",X"00",X"22",X"00",X"99",X"00",X"22",X"00",X"92",X"00",X"22",X"00",X"91",X"00",
		X"22",X"00",X"99",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"29",X"00",X"22",X"00",
		X"99",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"29",X"92",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"99",
		X"29",X"99",X"92",X"99",X"29",X"9A",X"92",X"A9",X"99",X"99",X"22",X"99",X"92",X"99",X"29",X"00",
		X"92",X"99",X"2A",X"00",X"92",X"22",X"29",X"00",X"92",X"22",X"29",X"00",X"99",X"99",X"22",X"00",
		X"29",X"99",X"22",X"99",X"22",X"92",X"29",X"29",X"22",X"12",X"9A",X"22",X"29",X"92",X"99",X"22",
		X"99",X"12",X"00",X"22",X"09",X"99",X"00",X"22",X"99",X"09",X"00",X"22",X"92",X"00",X"09",X"22",
		X"92",X"00",X"99",X"29",X"22",X"00",X"92",X"29",X"22",X"00",X"22",X"99",X"22",X"00",X"22",X"90",
		X"22",X"00",X"22",X"90",X"22",X"00",X"22",X"00",X"92",X"00",X"92",X"00",X"99",X"00",X"92",X"00",
		X"09",X"90",X"99",X"99",X"00",X"90",X"00",X"29",X"00",X"90",X"00",X"22",X"99",X"90",X"00",X"22",
		X"22",X"90",X"00",X"22",X"22",X"90",X"00",X"92",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"9B",X"9B",X"00",X"90",X"9B",X"BB",X"00",X"99",X"9B",X"BB",
		X"00",X"9B",X"BB",X"B9",X"00",X"9B",X"BB",X"B9",X"00",X"BB",X"BB",X"99",X"99",X"BB",X"BB",X"90",
		X"BB",X"BB",X"BB",X"90",X"BB",X"BB",X"99",X"00",X"BB",X"B9",X"59",X"00",X"BB",X"99",X"59",X"00",
		X"99",X"99",X"59",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"99",X"00",X"99",X"BB",X"99",X"00",
		X"B4",X"BB",X"BB",X"00",X"44",X"BB",X"BB",X"00",X"49",X"99",X"BB",X"00",X"09",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"09",X"BB",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"99",X"B9",X"00",X"00",X"97",X"99",X"90",X"00",X"97",X"9B",X"90",X"99",X"99",X"9B",X"90",
		X"99",X"11",X"9B",X"90",X"9B",X"77",X"9B",X"90",X"BB",X"99",X"9B",X"90",X"B9",X"11",X"9B",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9B",X"9B",X"00",X"90",X"9B",X"BB",
		X"00",X"99",X"9B",X"BB",X"00",X"9B",X"BB",X"B9",X"00",X"9B",X"BB",X"B9",X"00",X"BB",X"BB",X"99",
		X"99",X"BB",X"BB",X"90",X"BB",X"BB",X"BB",X"90",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"99",X"00",
		X"BB",X"B9",X"59",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"99",X"00",
		X"99",X"B9",X"99",X"00",X"BB",X"BB",X"99",X"00",X"BB",X"BB",X"BB",X"00",X"09",X"99",X"BB",X"00",
		X"09",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"09",X"BB",X"00",
		X"00",X"99",X"B9",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"BB",X"00",X"00",X"97",X"BB",X"00",
		X"99",X"99",X"BB",X"00",X"99",X"11",X"BB",X"00",X"9B",X"77",X"BB",X"00",X"BB",X"99",X"BB",X"00",
		X"B9",X"77",X"9B",X"90",X"B9",X"99",X"9B",X"90",X"99",X"11",X"9B",X"90",X"97",X"77",X"99",X"00",
		X"99",X"77",X"99",X"00",X"19",X"99",X"9B",X"09",X"71",X"11",X"BB",X"09",X"77",X"77",X"BB",X"09",
		X"97",X"77",X"BB",X"09",X"99",X"79",X"BB",X"99",X"91",X"79",X"BB",X"91",X"97",X"79",X"BB",X"BB",
		X"99",X"79",X"B9",X"BB",X"09",X"79",X"B9",X"BB",X"09",X"79",X"B9",X"BB",X"99",X"77",X"B9",X"BB",
		X"9B",X"77",X"19",X"B9",X"BB",X"77",X"99",X"B9",X"BB",X"77",X"BB",X"99",X"B9",X"99",X"BB",X"90",
		X"B9",X"00",X"99",X"00",X"BB",X"00",X"BB",X"99",X"BB",X"00",X"BB",X"9B",X"9B",X"90",X"BB",X"BB",
		X"99",X"90",X"BB",X"BB",X"99",X"90",X"BB",X"9B",X"9B",X"90",X"BB",X"9B",X"BB",X"00",X"9B",X"9B",
		X"BB",X"00",X"99",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B9",X"99",X"00",X"00",X"99",
		X"B9",X"11",X"BB",X"00",X"B9",X"99",X"BB",X"00",X"B9",X"BB",X"9B",X"99",X"99",X"BB",X"9B",X"BB",
		X"97",X"BB",X"BB",X"99",X"99",X"BB",X"BB",X"99",X"19",X"BB",X"BB",X"9B",X"71",X"BB",X"99",X"9B",
		X"77",X"BB",X"BB",X"9B",X"97",X"BB",X"BB",X"9B",X"99",X"99",X"BB",X"9B",X"91",X"79",X"B9",X"BB",
		X"97",X"79",X"B9",X"BB",X"99",X"79",X"B9",X"BB",X"09",X"79",X"B9",X"BB",X"09",X"79",X"BB",X"BB",
		X"00",X"77",X"BB",X"BB",X"00",X"77",X"BB",X"B9",X"00",X"77",X"BB",X"B9",X"00",X"77",X"BB",X"99",
		X"00",X"99",X"BB",X"90",X"00",X"BB",X"99",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"90",X"00",
		X"00",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"9B",X"B9",X"90",X"00",X"9B",X"99",X"99",X"00",
		X"BB",X"BB",X"B9",X"00",X"BB",X"BB",X"B9",X"00",X"99",X"BB",X"B9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"96",X"69",X"00",X"00",X"96",X"66",X"00",X"00",X"66",X"66",X"00",X"09",X"66",X"66",X"00",
		X"99",X"66",X"66",X"00",X"99",X"99",X"66",X"00",X"E9",X"9E",X"66",X"00",X"9E",X"9E",X"66",X"00",
		X"9E",X"EE",X"66",X"90",X"9E",X"9E",X"66",X"90",X"EE",X"EE",X"66",X"90",X"9E",X"9E",X"96",X"90",
		X"9E",X"9E",X"99",X"90",X"C9",X"9C",X"E9",X"90",X"99",X"9C",X"E9",X"90",X"99",X"9C",X"99",X"90",
		X"99",X"C9",X"99",X"90",X"99",X"99",X"D9",X"90",X"CC",X"9F",X"D9",X"90",X"9C",X"99",X"D9",X"90",
		X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"69",X"9F",X"99",X"96",X"69",X"99",X"99",X"96",X"69",
		X"99",X"CC",X"96",X"69",X"CC",X"C9",X"96",X"69",X"99",X"99",X"96",X"69",X"69",X"96",X"96",X"69",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"99",X"00",
		X"09",X"66",X"69",X"00",X"09",X"66",X"66",X"00",X"09",X"66",X"66",X"00",X"09",X"99",X"66",X"00",
		X"09",X"9E",X"66",X"00",X"99",X"9E",X"66",X"00",X"99",X"9E",X"66",X"90",X"9E",X"9E",X"66",X"90",
		X"EE",X"EE",X"66",X"90",X"EE",X"9E",X"96",X"90",X"EE",X"9E",X"99",X"90",X"99",X"9C",X"E9",X"90",
		X"C9",X"9C",X"E9",X"90",X"99",X"9C",X"99",X"90",X"99",X"C9",X"99",X"90",X"99",X"99",X"D9",X"90",
		X"CC",X"9F",X"D9",X"90",X"9C",X"99",X"D9",X"90",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"69",
		X"9F",X"9C",X"96",X"69",X"99",X"CC",X"96",X"69",X"CC",X"CC",X"96",X"69",X"CC",X"99",X"96",X"69",
		X"99",X"9D",X"96",X"69",X"69",X"66",X"96",X"69",X"69",X"66",X"96",X"69",X"69",X"66",X"96",X"99",
		X"69",X"66",X"96",X"69",X"69",X"66",X"96",X"99",X"99",X"66",X"99",X"69",X"96",X"66",X"69",X"66",
		X"96",X"66",X"69",X"66",X"66",X"66",X"69",X"66",X"66",X"66",X"69",X"66",X"66",X"66",X"99",X"66",
		X"99",X"99",X"99",X"66",X"DD",X"DD",X"99",X"66",X"DD",X"DD",X"99",X"66",X"9D",X"DD",X"99",X"66",
		X"99",X"99",X"69",X"66",X"9D",X"66",X"99",X"66",X"D9",X"66",X"90",X"66",X"D9",X"66",X"90",X"66",
		X"69",X"66",X"90",X"66",X"6D",X"66",X"00",X"66",X"66",X"66",X"99",X"66",X"99",X"99",X"D9",X"66",
		X"C9",X"99",X"69",X"66",X"99",X"99",X"69",X"99",X"96",X"99",X"99",X"CC",X"66",X"90",X"97",X"C9",
		X"96",X"00",X"97",X"C9",X"96",X"00",X"77",X"C9",X"99",X"00",X"77",X"C9",X"99",X"00",X"79",X"C9",
		X"79",X"99",X"79",X"9C",X"79",X"97",X"99",X"99",X"77",X"97",X"90",X"CC",X"99",X"09",X"90",X"99",
		X"99",X"66",X"96",X"90",X"96",X"66",X"99",X"90",X"96",X"66",X"99",X"90",X"66",X"66",X"99",X"90",
		X"66",X"66",X"99",X"90",X"66",X"66",X"96",X"90",X"99",X"99",X"96",X"90",X"DD",X"DD",X"96",X"90",
		X"DD",X"DD",X"96",X"90",X"9D",X"DD",X"96",X"90",X"99",X"99",X"96",X"90",X"96",X"66",X"96",X"90",
		X"D9",X"66",X"96",X"90",X"D9",X"66",X"96",X"90",X"69",X"66",X"96",X"90",X"6D",X"66",X"96",X"90",
		X"66",X"66",X"96",X"90",X"99",X"66",X"96",X"90",X"CC",X"66",X"96",X"90",X"CC",X"66",X"99",X"90",
		X"9C",X"66",X"9C",X"90",X"9C",X"66",X"9C",X"99",X"CC",X"66",X"9C",X"C9",X"C9",X"66",X"CC",X"C9",
		X"99",X"99",X"C9",X"C9",X"97",X"77",X"99",X"C9",X"77",X"77",X"99",X"99",X"79",X"77",X"09",X"90",
		X"99",X"79",X"09",X"90",X"09",X"99",X"99",X"00",X"09",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"E9",X"9B",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9E",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"EE",X"99",X"00",
		X"9E",X"9E",X"E9",X"00",X"E9",X"9E",X"99",X"00",X"99",X"99",X"9E",X"99",X"E9",X"B9",X"9E",X"E9",
		X"E9",X"99",X"9E",X"99",X"9E",X"9E",X"EE",X"90",X"E9",X"99",X"9E",X"90",X"E9",X"E4",X"9E",X"90",
		X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"E9",X"9B",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"99",X"00",
		X"00",X"A9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9E",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"0E",X"79",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"9E",X"9E",X"99",X"00",X"E9",X"9E",X"99",X"00",
		X"99",X"99",X"9E",X"99",X"E9",X"B9",X"99",X"E9",X"E9",X"99",X"99",X"99",X"9E",X"9E",X"9E",X"90",
		X"E9",X"99",X"9E",X"90",X"E9",X"E4",X"9E",X"90",X"E9",X"EE",X"EE",X"90",X"E9",X"EE",X"EE",X"99",
		X"EE",X"E9",X"EE",X"E9",X"9E",X"99",X"99",X"E9",X"9E",X"E9",X"9E",X"99",X"9E",X"9E",X"9E",X"00",
		X"E4",X"9E",X"99",X"99",X"EE",X"9E",X"99",X"B9",X"EE",X"9E",X"99",X"99",X"99",X"99",X"99",X"90",
		X"99",X"EE",X"99",X"90",X"E9",X"B9",X"99",X"00",X"EE",X"9B",X"99",X"99",X"E9",X"99",X"99",X"E9",
		X"99",X"90",X"9E",X"E9",X"09",X"90",X"EE",X"99",X"99",X"90",X"9E",X"90",X"9E",X"90",X"9E",X"90",
		X"9E",X"90",X"99",X"90",X"99",X"00",X"E9",X"00",X"99",X"90",X"E9",X"00",X"09",X"99",X"9E",X"00",
		X"09",X"E9",X"9E",X"00",X"99",X"99",X"99",X"00",X"9E",X"90",X"9E",X"00",X"99",X"90",X"9E",X"00",
		X"9E",X"90",X"9E",X"00",X"EE",X"99",X"94",X"00",X"9E",X"9E",X"99",X"00",X"99",X"E9",X"E9",X"00",
		X"E9",X"EE",X"E9",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"EE",X"9E",X"99",X"E9",X"EE",X"9E",X"E9",X"EE",X"E9",X"EE",X"E9",X"9E",X"99",X"99",X"E9",
		X"9E",X"E9",X"9E",X"99",X"9E",X"9E",X"9E",X"00",X"E4",X"99",X"99",X"00",X"EE",X"99",X"E9",X"00",
		X"EE",X"9E",X"EE",X"00",X"99",X"99",X"EE",X"00",X"E9",X"EE",X"99",X"00",X"E9",X"99",X"99",X"00",
		X"9E",X"9B",X"99",X"00",X"9E",X"99",X"99",X"00",X"E9",X"9E",X"EE",X"00",X"E9",X"99",X"9E",X"00",
		X"E9",X"90",X"9E",X"00",X"99",X"00",X"9E",X"00",X"B9",X"00",X"99",X"00",X"99",X"00",X"9E",X"90",
		X"E9",X"00",X"9E",X"99",X"EE",X"00",X"B9",X"E9",X"99",X"00",X"B9",X"E9",X"E9",X"00",X"99",X"99",
		X"E9",X"00",X"9E",X"9E",X"E9",X"90",X"90",X"9E",X"EE",X"90",X"9E",X"9E",X"99",X"99",X"9E",X"99",
		X"EE",X"E9",X"9E",X"EE",X"9E",X"99",X"E9",X"E9",X"9E",X"BE",X"EE",X"E9",X"99",X"99",X"99",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"97",X"90",X"00",X"99",X"97",
		X"99",X"00",X"77",X"97",X"AA",X"00",X"99",X"77",X"A9",X"40",X"F9",X"77",X"99",X"90",X"99",X"99",
		X"49",X"90",X"99",X"00",X"49",X"94",X"77",X"00",X"99",X"94",X"77",X"90",X"77",X"79",X"77",X"90",
		X"77",X"79",X"77",X"90",X"79",X"77",X"77",X"90",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",
		X"79",X"97",X"77",X"00",X"99",X"97",X"77",X"00",X"79",X"E7",X"77",X"00",X"79",X"E7",X"77",X"00",
		X"77",X"E7",X"77",X"00",X"99",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"09",X"77",X"77",X"00",X"09",X"99",X"77",X"00",
		X"97",X"44",X"77",X"00",X"79",X"94",X"79",X"90",X"79",X"99",X"99",X"90",X"79",X"94",X"97",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"09",X"77",X"79",
		X"00",X"09",X"77",X"79",X"99",X"09",X"79",X"79",X"99",X"09",X"99",X"99",X"99",X"00",X"79",X"90",
		X"33",X"00",X"77",X"90",X"93",X"00",X"77",X"40",X"99",X"40",X"77",X"00",X"97",X"94",X"77",X"00",
		X"97",X"99",X"99",X"00",X"77",X"79",X"9E",X"00",X"79",X"99",X"9E",X"00",X"79",X"77",X"9E",X"00",
		X"99",X"77",X"97",X"00",X"77",X"77",X"97",X"00",X"77",X"77",X"97",X"00",X"97",X"77",X"97",X"00",
		X"00",X"77",X"97",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"09",X"99",X"77",X"00",
		X"97",X"44",X"77",X"00",X"79",X"94",X"79",X"90",X"79",X"99",X"99",X"90",X"79",X"94",X"97",X"90",
		X"79",X"44",X"97",X"90",X"79",X"99",X"97",X"90",X"E9",X"91",X"99",X"90",X"E9",X"91",X"99",X"90",
		X"99",X"11",X"99",X"90",X"97",X"99",X"99",X"90",X"97",X"91",X"99",X"90",X"97",X"91",X"99",X"90",
		X"97",X"11",X"E9",X"90",X"97",X"99",X"E9",X"00",X"97",X"11",X"E9",X"00",X"97",X"11",X"E9",X"00",
		X"97",X"11",X"7E",X"00",X"97",X"99",X"7E",X"90",X"97",X"19",X"7E",X"90",X"77",X"19",X"77",X"90",
		X"77",X"19",X"79",X"90",X"77",X"99",X"79",X"90",X"77",X"91",X"99",X"90",X"77",X"99",X"90",X"00",
		X"77",X"11",X"00",X"00",X"77",X"99",X"00",X"00",X"77",X"49",X"00",X"00",X"77",X"44",X"00",X"09",
		X"97",X"44",X"99",X"99",X"97",X"99",X"79",X"77",X"97",X"91",X"77",X"77",X"97",X"91",X"77",X"37",
		X"99",X"99",X"77",X"77",X"09",X"19",X"77",X"77",X"00",X"19",X"99",X"79",X"00",X"99",X"99",X"99",
		X"79",X"44",X"97",X"90",X"79",X"99",X"97",X"90",X"E9",X"91",X"99",X"90",X"E9",X"91",X"99",X"90",
		X"99",X"11",X"99",X"90",X"97",X"99",X"E9",X"99",X"97",X"91",X"E9",X"99",X"97",X"91",X"E9",X"E9",
		X"97",X"11",X"7E",X"E9",X"97",X"99",X"7E",X"79",X"97",X"11",X"7E",X"77",X"97",X"11",X"77",X"77",
		X"97",X"11",X"77",X"77",X"97",X"99",X"77",X"97",X"97",X"19",X"77",X"99",X"77",X"19",X"77",X"00",
		X"77",X"19",X"79",X"00",X"77",X"99",X"79",X"09",X"77",X"91",X"99",X"99",X"77",X"99",X"90",X"97",
		X"77",X"11",X"00",X"77",X"77",X"99",X"00",X"77",X"77",X"49",X"99",X"79",X"77",X"44",X"77",X"79",
		X"97",X"44",X"77",X"99",X"97",X"99",X"77",X"90",X"97",X"91",X"77",X"90",X"99",X"91",X"77",X"00",
		X"09",X"99",X"77",X"00",X"00",X"19",X"77",X"00",X"00",X"19",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"99",X"09",X"00",X"99",X"99",X"09",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"92",X"99",X"99",X"99",X"92",X"99",
		X"99",X"99",X"29",X"99",X"99",X"99",X"22",X"99",X"99",X"99",X"92",X"99",X"99",X"99",X"92",X"99",
		X"99",X"49",X"99",X"90",X"99",X"49",X"29",X"09",X"99",X"99",X"29",X"99",X"99",X"22",X"29",X"99",
		X"99",X"29",X"29",X"99",X"99",X"95",X"29",X"99",X"99",X"95",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"92",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"92",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"D9",X"99",X"99",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"09",X"00",X"09",X"99",X"09",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"99",X"92",X"99",X"99",X"99",X"92",X"99",
		X"99",X"99",X"29",X"99",X"99",X"99",X"22",X"99",X"99",X"99",X"92",X"99",X"99",X"99",X"92",X"99",
		X"99",X"49",X"99",X"90",X"99",X"49",X"29",X"00",X"99",X"99",X"29",X"99",X"99",X"22",X"29",X"99",
		X"99",X"29",X"29",X"99",X"99",X"95",X"29",X"99",X"99",X"95",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"95",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"92",X"99",X"90",X"99",X"22",X"99",X"00",
		X"99",X"92",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"9D",X"99",X"D9",X"90",X"9D",X"99",X"D9",X"90",X"9D",X"99",X"D9",X"90",X"D9",X"99",X"99",X"99",
		X"D9",X"99",X"D9",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"22",X"99",X"99",X"99",X"22",
		X"99",X"99",X"99",X"22",X"99",X"99",X"99",X"22",X"09",X"99",X"99",X"22",X"09",X"99",X"99",X"22",
		X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",
		X"9D",X"99",X"D9",X"90",X"9D",X"99",X"D9",X"90",X"9D",X"99",X"D9",X"90",X"DD",X"99",X"D9",X"99",
		X"D9",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"92",X"99",X"00",X"99",X"92",X"29",X"00",X"99",X"99",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"95",X"90",X"00",
		X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"E0",X"00",X"33",X"EE",X"00",X"00",X"93",X"EE",X"00",X"00",X"99",X"99",X"99",X"00",
		X"09",X"F9",X"39",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"93",X"00",X"09",X"99",X"93",X"00",
		X"99",X"A9",X"39",X"00",X"93",X"99",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"33",X"39",X"00",
		X"00",X"39",X"33",X"00",X"00",X"33",X"33",X"00",X"90",X"33",X"99",X"00",X"90",X"33",X"9B",X"00",
		X"99",X"33",X"93",X"00",X"39",X"33",X"B3",X"00",X"33",X"33",X"33",X"00",X"93",X"99",X"9B",X"00",
		X"99",X"93",X"99",X"00",X"09",X"33",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"99",X"00",
		X"00",X"33",X"B9",X"00",X"09",X"33",X"99",X"00",X"09",X"93",X"90",X"00",X"09",X"33",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"D9",X"00",X"09",X"00",
		X"9D",X"00",X"99",X"90",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"99",
		X"99",X"90",X"9D",X"99",X"99",X"90",X"9D",X"99",X"99",X"49",X"99",X"99",X"99",X"44",X"9D",X"99",
		X"99",X"44",X"D9",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"99",X"99",X"9F",X"99",X"99",
		X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"90",X"99",X"9D",X"99",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"9D",X"99",X"09",X"00",X"99",X"99",X"99",X"90",X"99",X"49",X"99",X"99",
		X"99",X"94",X"9D",X"99",X"99",X"99",X"D9",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"DF",X"99",X"99",X"99",X"D3",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"9D",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"90",X"99",X"99",X"90",X"90",
		X"99",X"00",X"90",X"90",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"09",X"99",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"59",X"99",X"00",X"99",X"59",X"99",X"00",
		X"99",X"95",X"99",X"00",X"99",X"99",X"9D",X"00",X"99",X"99",X"DD",X"00",X"99",X"DF",X"DD",X"00",
		X"99",X"D3",X"D9",X"00",X"99",X"DD",X"D9",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AF",X"A0",X"00",
		X"00",X"AF",X"A0",X"00",X"00",X"AF",X"A0",X"00",X"00",X"FF",X"A0",X"00",X"00",X"FF",X"A0",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",X"FF",X"A0",
		X"00",X"AA",X"AA",X"A0",X"00",X"AF",X"FA",X"A0",X"00",X"FF",X"FF",X"00",X"00",X"AF",X"FF",X"00",
		X"0A",X"AF",X"FF",X"AA",X"0A",X"FA",X"FF",X"FF",X"0A",X"AA",X"AA",X"FF",X"0A",X"AF",X"FA",X"FF",
		X"00",X"AF",X"FA",X"FA",X"00",X"AF",X"FF",X"A0",X"0A",X"FF",X"FF",X"AA",X"AF",X"FF",X"FF",X"FF",
		X"AF",X"FA",X"FA",X"FF",X"AF",X"AA",X"FA",X"FA",X"AF",X"AF",X"AA",X"AA",X"0A",X"AF",X"FF",X"A0",
		X"00",X"FF",X"FF",X"AA",X"00",X"FF",X"FF",X"FA",X"00",X"FF",X"AF",X"FA",X"0A",X"AA",X"AA",X"FA",
		X"0A",X"FA",X"FF",X"FA",X"00",X"FF",X"FF",X"FA",X"00",X"FA",X"FF",X"A0",X"00",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"AA",X"00",X"00",X"A0",X"FA",X"00",X"0A",X"AA",
		X"FF",X"00",X"0A",X"FA",X"FF",X"00",X"AA",X"FF",X"FF",X"00",X"AF",X"FF",X"FA",X"00",X"AF",X"FF",
		X"FA",X"00",X"AA",X"FF",X"AA",X"00",X"0A",X"FF",X"00",X"0A",X"00",X"FA",X"00",X"AA",X"00",X"AA",
		X"00",X"AF",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"AA",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"A0",X"FF",X"00",X"00",X"AA",X"AF",X"00",X"00",X"FA",X"0A",X"00",X"00",X"FA",
		X"0A",X"00",X"00",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"A0",
		X"A0",X"00",X"A0",X"00",X"0A",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A0",X"FF",X"0F",X"00",X"00",X"33",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"A0",X"00",X"0F",X"AA",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"FF",X"0F",X"00",X"A0",X"33",X"03",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"0A",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"00",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"55",X"00",X"00",X"9F",X"F5",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"9F",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"99",X"F5",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",
		X"00",X"59",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"90",X"99",X"00",
		X"09",X"90",X"95",X"00",X"09",X"90",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"55",X"00",X"00",X"9F",X"99",X"00",X"00",X"FF",X"9F",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"99",X"9F",X"00",X"00",X"FF",X"99",X"00",X"00",X"9F",X"F9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"F9",X"FF",X"00",X"00",X"FF",X"9F",X"00",X"00",X"99",X"9F",X"00",X"00",X"FF",X"99",X"00",
		X"00",X"FF",X"F9",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"99",X"F5",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",
		X"00",X"59",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"90",X"99",X"00",
		X"09",X"90",X"95",X"00",X"09",X"90",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9F",X"55",X"00",X"00",X"9F",X"99",X"00",X"00",X"F9",X"9F",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"99",X"9F",X"00",X"00",X"FF",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"F9",X"FF",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"9F",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"FF",X"F9",X"00",X"00",X"F9",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"99",X"00",
		X"00",X"FF",X"F9",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",
		X"00",X"59",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"90",X"99",X"00",
		X"09",X"90",X"95",X"00",X"09",X"90",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"09",X"02",X"00",X"00",X"09",X"00",X"00",X"99",X"09",X"00",X"00",X"F9",
		X"00",X"02",X"00",X"F9",X"09",X"92",X"96",X"F9",X"09",X"99",X"99",X"F9",X"09",X"99",X"90",X"FF",
		X"00",X"99",X"69",X"FF",X"00",X"99",X"99",X"F9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"19",X"00",X"00",X"49",X"99",X"00",
		X"00",X"49",X"93",X"00",X"09",X"99",X"99",X"99",X"99",X"19",X"99",X"F9",X"9F",X"19",X"79",X"FF",
		X"9F",X"90",X"97",X"F9",X"99",X"90",X"97",X"F9",X"09",X"00",X"99",X"99",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"30",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"90",X"AA",X"00",X"00",X"99",X"A3",X"99",X"99",X"A9",X"AA",X"59",X"95",X"A9",
		X"33",X"99",X"99",X"A9",X"A3",X"99",X"99",X"AA",X"AA",X"99",X"99",X"A9",X"AA",X"99",X"99",X"3A",
		X"AA",X"99",X"99",X"AA",X"33",X"99",X"99",X"33",X"AA",X"94",X"49",X"A3",X"AA",X"94",X"49",X"A3",
		X"AA",X"44",X"44",X"A3",X"A3",X"49",X"94",X"AA",X"A3",X"49",X"94",X"5A",X"AA",X"49",X"94",X"35",
		X"AA",X"49",X"94",X"33",X"A9",X"49",X"94",X"A3",X"A9",X"49",X"94",X"A3",X"A9",X"49",X"94",X"A3",
		X"A9",X"94",X"49",X"AA",X"99",X"99",X"99",X"AA",X"99",X"59",X"95",X"9A",X"90",X"95",X"59",X"99",
		X"90",X"99",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"90",X"09",X"09",X"00",X"90",X"09",X"09",
		X"00",X"99",X"09",X"00",X"00",X"A9",X"99",X"00",X"00",X"39",X"9A",X"00",X"00",X"3A",X"AA",X"00",
		X"00",X"3A",X"A3",X"00",X"00",X"A3",X"A3",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"95",X"00",
		X"00",X"9A",X"A9",X"00",X"00",X"9A",X"A9",X"00",X"00",X"9A",X"A9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"49",X"00",X"00",X"94",X"49",X"00",
		X"00",X"44",X"44",X"00",X"00",X"49",X"94",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"49",X"94",X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"94",X"00",
		X"00",X"94",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"95",X"59",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"A3",X"A3",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"9A",X"00",
		X"00",X"9A",X"A9",X"00",X"00",X"9A",X"A9",X"00",X"00",X"9A",X"A9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"49",X"00",X"00",X"94",X"49",X"00",
		X"00",X"44",X"44",X"00",X"00",X"49",X"94",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"49",X"94",X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"94",X"00",
		X"00",X"94",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"95",X"59",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"AA",X"AA",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"44",X"49",X"00",
		X"00",X"99",X"94",X"00",X"09",X"22",X"99",X"00",X"99",X"22",X"A9",X"00",X"94",X"99",X"A2",X"99",
		X"11",X"99",X"A9",X"49",X"11",X"99",X"A9",X"11",X"15",X"99",X"A1",X"19",X"55",X"11",X"11",X"EE",
		X"EE",X"11",X"11",X"E9",X"9E",X"19",X"19",X"99",X"99",X"E7",X"EE",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"44",X"49",X"00",
		X"00",X"99",X"94",X"00",X"09",X"22",X"29",X"00",X"99",X"29",X"A2",X"00",X"94",X"99",X"A2",X"99",
		X"11",X"99",X"A9",X"49",X"11",X"99",X"A9",X"11",X"17",X"99",X"A1",X"19",X"77",X"11",X"11",X"EE",
		X"EE",X"11",X"11",X"E9",X"9E",X"19",X"19",X"99",X"99",X"E5",X"EE",X"00",X"00",X"99",X"99",X"00",
		X"99",X"E0",X"E0",X"90",X"93",X"E0",X"E0",X"90",X"93",X"EE",X"99",X"90",X"93",X"99",X"F9",X"90",
		X"93",X"39",X"4F",X"90",X"93",X"9F",X"FF",X"90",X"93",X"94",X"FF",X"00",X"99",X"9F",X"99",X"00",
		X"09",X"9F",X"99",X"00",X"09",X"9F",X"FF",X"00",X"00",X"99",X"4F",X"00",X"00",X"39",X"99",X"00",
		X"00",X"33",X"33",X"00",X"00",X"99",X"93",X"00",X"00",X"99",X"33",X"00",X"50",X"9F",X"33",X"05",
		X"05",X"99",X"33",X"50",X"00",X"93",X"33",X"00",X"00",X"99",X"93",X"05",X"00",X"9B",X"99",X"55",
		X"00",X"99",X"99",X"00",X"00",X"39",X"99",X"00",X"11",X"33",X"39",X"04",X"A1",X"39",X"39",X"00",
		X"A4",X"A4",X"79",X"10",X"99",X"54",X"74",X"04",X"51",X"94",X"91",X"00",X"94",X"77",X"41",X"00",
		X"00",X"41",X"11",X"00",X"00",X"15",X"91",X"00",X"00",X"15",X"01",X"00",X"00",X"00",X"00",X"50",
		X"00",X"E0",X"E0",X"00",X"99",X"E0",X"9E",X"90",X"93",X"EE",X"EE",X"90",X"93",X"99",X"E9",X"90",
		X"93",X"33",X"99",X"90",X"93",X"39",X"AA",X"90",X"93",X"99",X"FF",X"00",X"99",X"9A",X"FF",X"00",
		X"09",X"9F",X"99",X"00",X"09",X"9F",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",X"39",X"99",X"00",
		X"00",X"33",X"33",X"00",X"00",X"39",X"39",X"00",X"00",X"99",X"33",X"00",X"00",X"B3",X"33",X"00",
		X"00",X"B3",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"93",X"00",X"00",X"93",X"99",X"00",
		X"00",X"33",X"99",X"00",X"00",X"93",X"39",X"00",X"00",X"93",X"39",X"00",X"09",X"33",X"33",X"00",
		X"09",X"33",X"93",X"00",X"09",X"99",X"99",X"00",X"09",X"33",X"09",X"00",X"00",X"33",X"99",X"00",
		X"00",X"33",X"93",X"00",X"00",X"99",X"93",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"55",X"00",X"00",X"9F",X"F5",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",
		X"00",X"59",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"90",X"99",X"00",
		X"09",X"90",X"95",X"00",X"09",X"90",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"09",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"99",X"00",
		X"99",X"9B",X"94",X"99",X"19",X"BB",X"94",X"9B",X"19",X"BB",X"99",X"BB",X"11",X"BB",X"BB",X"99",
		X"E1",X"B9",X"BB",X"99",X"EE",X"99",X"99",X"B9",X"EE",X"99",X"99",X"99",X"E1",X"B9",X"99",X"00",
		X"E1",X"BB",X"99",X"00",X"11",X"9B",X"99",X"99",X"11",X"99",X"49",X"9B",X"11",X"B9",X"99",X"BB",
		X"11",X"BB",X"BB",X"BB",X"11",X"99",X"99",X"9B",X"11",X"99",X"7B",X"9B",X"99",X"9B",X"77",X"91",
		X"9B",X"BB",X"77",X"00",X"99",X"BB",X"77",X"00",X"11",X"B9",X"BB",X"00",X"11",X"B9",X"BB",X"99",
		X"91",X"99",X"BB",X"9B",X"91",X"99",X"B9",X"BB",X"99",X"99",X"99",X"BB",X"00",X"99",X"90",X"BB",
		X"00",X"99",X"00",X"B9",X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"11",X"00",X"99",X"00",X"E1",X"99",X"99",X"00",
		X"EE",X"9B",X"94",X"99",X"EE",X"BB",X"94",X"9B",X"EE",X"BB",X"99",X"BB",X"1E",X"BB",X"BB",X"99",
		X"11",X"BB",X"BB",X"99",X"11",X"BB",X"99",X"B9",X"11",X"BB",X"99",X"99",X"11",X"BB",X"99",X"99",
		X"11",X"BB",X"49",X"9B",X"11",X"99",X"BB",X"9B",X"19",X"B9",X"99",X"BB",X"19",X"BB",X"99",X"9B",
		X"99",X"BB",X"B9",X"99",X"9B",X"BB",X"B9",X"00",X"B9",X"9B",X"7B",X"00",X"99",X"BB",X"77",X"00",
		X"00",X"BB",X"77",X"00",X"00",X"BB",X"77",X"00",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"BB",X"99",
		X"00",X"99",X"B9",X"9B",X"00",X"99",X"B9",X"BB",X"00",X"99",X"99",X"BB",X"00",X"99",X"90",X"BB",
		X"00",X"99",X"00",X"B9",X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"99",X"00",X"00",X"66",X"99",X"00",
		X"00",X"66",X"96",X"00",X"99",X"66",X"99",X"00",X"EE",X"96",X"69",X"00",X"9E",X"99",X"66",X"00",
		X"99",X"EE",X"66",X"00",X"94",X"EE",X"66",X"00",X"94",X"CE",X"66",X"00",X"99",X"9E",X"66",X"00",
		X"C9",X"9C",X"66",X"00",X"99",X"9C",X"66",X"00",X"99",X"9C",X"66",X"00",X"99",X"9C",X"66",X"00",
		X"C9",X"9C",X"66",X"00",X"CC",X"CC",X"66",X"00",X"9C",X"CC",X"69",X"00",X"99",X"CC",X"69",X"00",
		X"09",X"99",X"99",X"00",X"09",X"96",X"99",X"00",X"99",X"66",X"96",X"00",X"C9",X"99",X"66",X"00",
		X"9C",X"CC",X"66",X"00",X"9C",X"CC",X"66",X"00",X"9C",X"9C",X"66",X"00",X"99",X"9C",X"66",X"00",
		X"00",X"99",X"99",X"00",X"00",X"77",X"77",X"00",X"00",X"99",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"90",X"00",X"00",X"66",X"69",X"00",
		X"99",X"66",X"96",X"00",X"E9",X"96",X"99",X"00",X"9E",X"99",X"69",X"00",X"99",X"EE",X"66",X"00",
		X"94",X"EE",X"66",X"00",X"94",X"CE",X"66",X"00",X"99",X"99",X"66",X"00",X"C9",X"99",X"66",X"00",
		X"99",X"99",X"66",X"00",X"99",X"9C",X"66",X"00",X"99",X"99",X"66",X"00",X"C9",X"59",X"66",X"00",
		X"CC",X"99",X"66",X"00",X"9C",X"9C",X"66",X"00",X"99",X"CC",X"66",X"00",X"09",X"99",X"66",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"69",X"99",X"99",X"00",X"69",X"CC",X"97",X"00",X"99",X"CC",X"97",X"99",X"99",X"CC",X"97",
		X"97",X"90",X"99",X"97",X"97",X"90",X"09",X"97",X"99",X"90",X"00",X"77",X"00",X"00",X"00",X"99",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"99",X"00",X"90",X"99",X"E9",X"00",
		X"99",X"99",X"B9",X"00",X"EE",X"9E",X"B9",X"90",X"E9",X"EE",X"99",X"99",X"99",X"EE",X"9E",X"EE",
		X"E9",X"E9",X"9E",X"EE",X"E9",X"99",X"99",X"E9",X"99",X"97",X"99",X"99",X"9E",X"99",X"99",X"11",
		X"99",X"99",X"9E",X"11",X"E9",X"99",X"E4",X"99",X"99",X"E9",X"44",X"EE",X"09",X"EE",X"94",X"E9",
		X"00",X"91",X"99",X"99",X"00",X"91",X"9E",X"00",X"00",X"91",X"9E",X"00",X"99",X"99",X"9E",X"00",
		X"9E",X"E9",X"EE",X"00",X"9E",X"99",X"EE",X"90",X"EE",X"90",X"99",X"90",X"99",X"90",X"E9",X"99",
		X"EE",X"90",X"E9",X"99",X"99",X"00",X"EE",X"49",X"E9",X"00",X"EE",X"49",X"99",X"00",X"99",X"99",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"99",X"00",X"00",X"9A",X"E9",X"00",
		X"00",X"99",X"B9",X"00",X"00",X"9E",X"B9",X"00",X"09",X"EE",X"99",X"00",X"99",X"EE",X"9E",X"00",
		X"91",X"99",X"99",X"00",X"91",X"79",X"99",X"99",X"99",X"99",X"99",X"99",X"9E",X"99",X"99",X"9E",
		X"9E",X"99",X"99",X"9E",X"EE",X"99",X"94",X"EE",X"E9",X"99",X"44",X"11",X"90",X"EE",X"94",X"91",
		X"99",X"91",X"99",X"99",X"99",X"91",X"9E",X"EE",X"9E",X"91",X"9B",X"EE",X"9E",X"99",X"9E",X"EE",
		X"99",X"99",X"EE",X"99",X"11",X"90",X"99",X"00",X"41",X"90",X"E9",X"90",X"91",X"90",X"E9",X"99",
		X"99",X"90",X"99",X"99",X"EE",X"90",X"1E",X"19",X"9E",X"00",X"99",X"11",X"99",X"00",X"00",X"99",
		X"99",X"00",X"99",X"00",X"77",X"90",X"77",X"99",X"79",X"99",X"77",X"39",X"99",X"79",X"77",X"99",
		X"9F",X"79",X"79",X"77",X"99",X"77",X"79",X"77",X"99",X"77",X"79",X"77",X"99",X"77",X"77",X"97",
		X"97",X"77",X"77",X"99",X"99",X"77",X"99",X"00",X"99",X"77",X"77",X"90",X"97",X"77",X"77",X"99",
		X"77",X"77",X"77",X"79",X"77",X"77",X"77",X"77",X"77",X"99",X"77",X"77",X"77",X"91",X"77",X"77",
		X"74",X"99",X"77",X"77",X"74",X"11",X"79",X"77",X"97",X"11",X"79",X"77",X"9A",X"91",X"77",X"49",
		X"99",X"99",X"77",X"49",X"99",X"94",X"77",X"79",X"90",X"94",X"99",X"A9",X"00",X"94",X"49",X"99",
		X"00",X"99",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"99",X"77",X"00",X"00",X"97",X"77",X"00",X"00",X"97",X"77",X"00",X"00",X"99",X"99",
		X"99",X"00",X"99",X"00",X"97",X"90",X"77",X"99",X"79",X"99",X"77",X"39",X"99",X"79",X"79",X"39",
		X"9F",X"79",X"99",X"99",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"94",X"97",
		X"99",X"77",X"79",X"99",X"97",X"77",X"77",X"00",X"99",X"77",X"97",X"00",X"00",X"77",X"79",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"79",X"00",X"00",X"99",X"79",X"00",X"09",X"91",X"79",X"00",
		X"09",X"99",X"99",X"90",X"99",X"11",X"94",X"90",X"97",X"11",X"94",X"99",X"97",X"91",X"97",X"79",
		X"97",X"99",X"97",X"77",X"97",X"94",X"77",X"77",X"97",X"94",X"99",X"77",X"99",X"99",X"49",X"4A",
		X"09",X"90",X"99",X"49",X"09",X"00",X"99",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"00",X"99",X"90",X"99",X"90",X"99",X"99",X"92",X"90",X"09",X"29",X"92",X"00",
		X"09",X"92",X"92",X"00",X"09",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"99",X"49",X"99",X"00",
		X"99",X"94",X"92",X"00",X"99",X"99",X"99",X"00",X"22",X"99",X"99",X"00",X"29",X"99",X"99",X"00",
		X"29",X"95",X"9D",X"00",X"99",X"99",X"99",X"00",X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"29",X"00",X"99",X"99",X"29",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"00",X"09",X"92",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"99",X"00",
		X"09",X"94",X"99",X"99",X"99",X"99",X"99",X"29",X"09",X"99",X"99",X"29",X"00",X"99",X"99",X"29",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"22",X"99",X"99",X"99",X"29",X"99",X"99",X"00",X"22",X"99",X"99",X"00",
		X"29",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"92",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"39",X"2D",X"99",X"00",X"99",X"DD",X"29",X"00",X"22",X"9D",X"29",X"00",X"22",X"9D",X"22",
		X"00",X"99",X"99",X"22",X"00",X"95",X"29",X"22",X"00",X"99",X"29",X"29",X"90",X"99",X"29",X"99",
		X"99",X"99",X"99",X"9D",X"29",X"99",X"9D",X"D2",X"22",X"59",X"9D",X"DD",X"92",X"99",X"A2",X"DD",
		X"99",X"22",X"22",X"2D",X"DD",X"29",X"22",X"22",X"22",X"99",X"29",X"D9",X"DD",X"92",X"29",X"D9",
		X"DD",X"A2",X"29",X"99",X"DD",X"22",X"29",X"00",X"92",X"22",X"29",X"00",X"9D",X"2A",X"29",X"00",
		X"99",X"92",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"22",X"00",
		X"00",X"00",X"29",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"92",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"49",X"2D",X"00",X"00",X"99",X"DD",X"00",X"00",X"22",X"9D",X"00",X"00",X"22",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"95",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"95",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"22",X"DD",X"00",X"00",X"99",X"DD",X"00",
		X"00",X"DD",X"D2",X"00",X"00",X"92",X"2D",X"00",X"00",X"92",X"DD",X"00",X"00",X"92",X"DD",X"00",
		X"00",X"92",X"DD",X"00",X"00",X"99",X"D2",X"00",X"00",X"D9",X"2D",X"00",X"00",X"D9",X"DD",X"00",
		X"00",X"D9",X"DD",X"00",X"00",X"29",X"99",X"00",X"00",X"D9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"E0",X"E0",X"00",X"99",X"E0",X"9E",X"90",X"93",X"EE",X"EE",X"90",X"93",X"99",X"E9",X"90",
		X"93",X"33",X"99",X"90",X"93",X"39",X"FF",X"90",X"93",X"99",X"FF",X"00",X"99",X"9F",X"A9",X"00",
		X"09",X"99",X"99",X"00",X"09",X"39",X"99",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"39",X"93",X"00",X"00",X"33",X"33",X"00",X"00",X"B3",X"33",X"00",
		X"00",X"B3",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"93",X"00",X"00",X"9B",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"39",X"99",X"00",X"99",X"33",X"39",X"00",X"94",X"39",X"39",X"99",
		X"11",X"3B",X"39",X"49",X"11",X"B3",X"99",X"11",X"15",X"99",X"91",X"19",X"55",X"11",X"11",X"EE",
		X"EE",X"11",X"11",X"E9",X"9E",X"19",X"19",X"99",X"99",X"E7",X"EE",X"00",X"00",X"99",X"99",X"00",
		X"00",X"E0",X"9E",X"00",X"00",X"EE",X"EE",X"99",X"99",X"99",X"E9",X"39",X"33",X"33",X"99",X"99",
		X"93",X"39",X"F9",X"90",X"93",X"99",X"99",X"00",X"99",X"9A",X"99",X"00",X"09",X"99",X"99",X"00",
		X"09",X"39",X"F9",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"39",X"93",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"B3",X"33",X"00",
		X"00",X"93",X"33",X"00",X"00",X"99",X"93",X"00",X"00",X"9B",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"39",X"99",X"00",X"00",X"33",X"99",X"00",X"99",X"39",X"39",X"00",X"94",X"39",X"39",X"99",
		X"11",X"3B",X"39",X"49",X"11",X"B3",X"99",X"11",X"17",X"99",X"91",X"19",X"77",X"11",X"11",X"EE",
		X"EE",X"11",X"11",X"E9",X"9E",X"19",X"19",X"99",X"99",X"E5",X"EE",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9F",X"55",X"00",X"00",X"9F",X"99",X"00",X"00",X"F9",X"9F",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"99",X"99",X"00",X"00",X"FF",X"A9",X"00",X"00",X"9F",X"AA",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"FF",X"00",X"00",X"9A",X"9F",X"00",X"00",X"99",X"9F",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"FF",X"F9",X"00",X"00",X"F9",X"9F",X"00",X"00",X"99",X"A9",X"00",X"00",X"F9",X"99",X"00",
		X"00",X"FF",X"F9",X"00",X"00",X"99",X"F9",X"00",X"00",X"9A",X"95",X"00",X"00",X"99",X"99",X"00",
		X"00",X"59",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"90",X"99",X"00",
		X"09",X"90",X"95",X"00",X"09",X"90",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"09",X"02",X"00",X"00",X"09",X"00",X"00",X"99",X"09",X"40",X"00",X"F9",
		X"00",X"42",X"00",X"F9",X"09",X"92",X"96",X"F9",X"09",X"99",X"9A",X"F9",X"09",X"A9",X"A0",X"FF",
		X"00",X"9A",X"69",X"FF",X"00",X"4A",X"9A",X"F9",X"00",X"A9",X"4A",X"99",X"00",X"AA",X"AA",X"00",
		X"00",X"9A",X"AA",X"00",X"00",X"4A",X"9A",X"00",X"00",X"A9",X"19",X"00",X"00",X"49",X"A9",X"00",
		X"00",X"4A",X"93",X"00",X"09",X"99",X"A9",X"99",X"99",X"19",X"A9",X"F9",X"9F",X"19",X"7A",X"FF",
		X"9F",X"90",X"97",X"F9",X"99",X"90",X"97",X"F9",X"09",X"00",X"99",X"99",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"30",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"E0",X"00",X"90",X"EE",X"E0",X"00",X"90",X"9E",X"00",X"00",X"90",X"33",X"E0",X"00",
		X"99",X"99",X"90",X"00",X"39",X"9A",X"99",X"00",X"33",X"A9",X"AA",X"00",X"39",X"F9",X"FA",X"00",
		X"3B",X"FF",X"FF",X"00",X"9B",X"FF",X"F9",X"00",X"93",X"99",X"99",X"00",X"93",X"33",X"33",X"00",
		X"09",X"33",X"33",X"00",X"09",X"99",X"33",X"00",X"00",X"49",X"33",X"00",X"99",X"94",X"33",X"00",
		X"39",X"4B",X"33",X"00",X"39",X"B3",X"33",X"00",X"33",X"3B",X"33",X"00",X"93",X"3B",X"99",X"00",
		X"99",X"39",X"09",X"00",X"09",X"33",X"09",X"00",X"00",X"93",X"99",X"00",X"90",X"33",X"33",X"00",
		X"99",X"33",X"99",X"00",X"39",X"33",X"09",X"00",X"39",X"39",X"09",X"00",X"33",X"39",X"99",X"00",
		X"39",X"33",X"33",X"00",X"39",X"33",X"93",X"00",X"99",X"33",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"29",X"00",
		X"99",X"29",X"29",X"90",X"22",X"29",X"29",X"90",X"99",X"29",X"22",X"90",X"94",X"22",X"29",X"90",
		X"99",X"22",X"29",X"90",X"DD",X"29",X"22",X"90",X"22",X"99",X"92",X"90",X"99",X"59",X"92",X"90",
		X"99",X"59",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",
		X"95",X"99",X"22",X"00",X"99",X"22",X"22",X"00",X"DD",X"29",X"22",X"00",X"29",X"22",X"22",X"00",
		X"22",X"99",X"22",X"90",X"99",X"99",X"92",X"90",X"99",X"92",X"92",X"90",X"99",X"22",X"22",X"00",
		X"92",X"22",X"22",X"00",X"92",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",
		X"00",X"09",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"99",X"00",
		X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"29",X"00",X"99",X"29",X"29",X"90",
		X"22",X"29",X"29",X"90",X"99",X"29",X"22",X"90",X"99",X"22",X"29",X"90",X"99",X"22",X"29",X"90",
		X"DD",X"29",X"22",X"90",X"22",X"99",X"92",X"90",X"99",X"59",X"92",X"90",X"99",X"59",X"92",X"00",
		X"99",X"99",X"92",X"00",X"22",X"92",X"92",X"00",X"22",X"22",X"92",X"00",X"29",X"22",X"22",X"00",
		X"99",X"22",X"22",X"00",X"99",X"92",X"22",X"00",X"99",X"99",X"22",X"00",X"99",X"DD",X"22",X"90",
		X"29",X"22",X"92",X"90",X"29",X"22",X"92",X"90",X"99",X"22",X"22",X"00",X"92",X"22",X"22",X"00",
		X"92",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",
		X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"9A",X"00",
		X"99",X"22",X"99",X"00",X"9A",X"22",X"99",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"22",X"00",
		X"22",X"22",X"22",X"00",X"99",X"22",X"22",X"00",X"22",X"99",X"22",X"00",X"22",X"9D",X"22",X"00",
		X"99",X"9D",X"22",X"00",X"00",X"99",X"22",X"00",X"99",X"00",X"29",X"00",X"29",X"00",X"29",X"00",
		X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",
		X"22",X"00",X"99",X"00",X"99",X"00",X"22",X"00",X"90",X"00",X"29",X"00",X"90",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"99",X"90",
		X"00",X"09",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"92",X"22",X"90",X"00",X"99",X"99",X"90",
		X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"99",X"22",X"92",X"00",
		X"9A",X"92",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"22",X"92",X"00",X"22",X"92",X"29",X"00",
		X"99",X"92",X"99",X"00",X"29",X"22",X"92",X"90",X"99",X"22",X"92",X"99",X"92",X"22",X"92",X"29",
		X"22",X"22",X"99",X"29",X"22",X"22",X"09",X"29",X"22",X"19",X"00",X"29",X"22",X"00",X"99",X"99",
		X"22",X"00",X"22",X"90",X"22",X"00",X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",X"22",X"00",
		X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"92",X"00",X"92",X"00",X"99",X"00",X"99",X"90",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"29",
		X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"00",
		X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"90",X"00",X"09",X"BB",X"90",X"00",X"99",X"BB",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"99",X"BB",X"00",X"99",X"BB",X"BB",X"00",X"9B",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"9B",X"00",X"BB",X"99",X"99",X"00",X"BB",X"95",X"99",X"00",
		X"99",X"95",X"99",X"00",X"99",X"95",X"99",X"00",X"94",X"99",X"99",X"00",X"44",X"BB",X"99",X"00",
		X"4B",X"BB",X"BB",X"00",X"9B",X"BB",X"BB",X"00",X"BB",X"99",X"BB",X"00",X"99",X"9B",X"BB",X"00",
		X"00",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"B9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"77",X"9B",X"00",X"09",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",X"9B",X"99",X"BB",X"00",
		X"BB",X"11",X"BB",X"00",X"B9",X"77",X"BB",X"00",X"99",X"99",X"BB",X"00",X"97",X"11",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"90",X"00",X"09",X"BB",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"99",X"BB",X"90",X"00",X"99",X"BB",X"00",X"99",X"BB",X"BB",X"00",
		X"9B",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"99",X"9B",X"00",X"99",X"95",X"99",X"00",X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",
		X"44",X"99",X"99",X"00",X"B4",X"BB",X"99",X"00",X"9B",X"BB",X"BB",X"00",X"BB",X"99",X"BB",X"00",
		X"99",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"99",X"00",
		X"00",X"99",X"9B",X"00",X"00",X"77",X"BB",X"00",X"09",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",
		X"9B",X"99",X"BB",X"00",X"BB",X"11",X"BB",X"00",X"B9",X"77",X"BB",X"00",X"99",X"99",X"BB",X"00",
		X"97",X"77",X"BB",X"09",X"99",X"99",X"BB",X"9B",X"11",X"11",X"BB",X"9B",X"77",X"77",X"BB",X"9B",
		X"77",X"77",X"BB",X"BB",X"99",X"77",X"BB",X"B9",X"11",X"17",X"BB",X"B9",X"77",X"79",X"BB",X"B9",
		X"77",X"99",X"BB",X"19",X"99",X"9B",X"BB",X"B9",X"11",X"B9",X"BB",X"B9",X"77",X"B9",X"B9",X"B9",
		X"77",X"B9",X"B9",X"B9",X"77",X"BB",X"B9",X"B9",X"99",X"9B",X"BB",X"99",X"91",X"9B",X"9B",X"90",
		X"99",X"99",X"9B",X"90",X"B9",X"79",X"99",X"00",X"B9",X"79",X"BB",X"00",X"BB",X"99",X"BB",X"00",
		X"99",X"00",X"99",X"00",X"BB",X"00",X"BB",X"99",X"BB",X"00",X"B9",X"B9",X"BB",X"00",X"B9",X"B9",
		X"99",X"00",X"B9",X"B9",X"BB",X"00",X"BB",X"B9",X"BB",X"00",X"BB",X"B9",X"BB",X"00",X"BB",X"99",
		X"BB",X"00",X"99",X"90",X"BB",X"00",X"00",X"90",X"B9",X"00",X"09",X"90",X"99",X"00",X"09",X"90",
		X"97",X"11",X"BB",X"00",X"97",X"77",X"BB",X"09",X"99",X"99",X"BB",X"9B",X"1B",X"B9",X"BB",X"BB",
		X"9B",X"BB",X"BB",X"BB",X"99",X"BB",X"BB",X"BB",X"99",X"BB",X"B9",X"B9",X"11",X"BB",X"99",X"B9",
		X"77",X"B9",X"B9",X"B9",X"77",X"99",X"99",X"B9",X"99",X"9B",X"90",X"B9",X"11",X"BB",X"90",X"B9",
		X"77",X"BB",X"00",X"B9",X"77",X"BB",X"00",X"B9",X"77",X"BB",X"90",X"B9",X"99",X"9B",X"99",X"99",
		X"91",X"9B",X"BB",X"90",X"99",X"99",X"BB",X"90",X"09",X"79",X"BB",X"00",X"09",X"79",X"BB",X"00",
		X"00",X"99",X"BB",X"00",X"00",X"B9",X"99",X"00",X"00",X"B9",X"90",X"00",X"00",X"B9",X"00",X"00",
		X"00",X"B9",X"00",X"00",X"99",X"B9",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"99",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",
		X"09",X"66",X"99",X"00",X"09",X"66",X"69",X"00",X"99",X"66",X"69",X"00",X"96",X"66",X"99",X"00",
		X"66",X"66",X"66",X"00",X"69",X"99",X"66",X"00",X"99",X"E9",X"66",X"00",X"9E",X"99",X"69",X"00",
		X"9E",X"E9",X"69",X"00",X"EE",X"E9",X"99",X"00",X"EE",X"E9",X"96",X"00",X"EE",X"EE",X"96",X"00",
		X"EE",X"EE",X"96",X"00",X"EE",X"CC",X"66",X"00",X"EE",X"C9",X"66",X"00",X"99",X"99",X"66",X"00",
		X"C9",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",
		X"CC",X"99",X"66",X"00",X"99",X"99",X"66",X"00",X"99",X"9C",X"66",X"00",X"99",X"CC",X"66",X"00",
		X"99",X"C9",X"66",X"00",X"99",X"99",X"66",X"00",X"CC",X"DD",X"66",X"00",X"99",X"66",X"66",X"00",
		X"00",X"99",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",
		X"99",X"66",X"90",X"00",X"66",X"66",X"99",X"00",X"66",X"66",X"66",X"00",X"69",X"99",X"66",X"00",
		X"99",X"E9",X"66",X"00",X"9E",X"99",X"69",X"00",X"9E",X"E9",X"69",X"00",X"EE",X"E9",X"99",X"00",
		X"EE",X"E9",X"96",X"00",X"EE",X"EE",X"96",X"00",X"EE",X"EE",X"96",X"00",X"EE",X"CC",X"66",X"00",
		X"EE",X"C9",X"66",X"00",X"99",X"99",X"66",X"00",X"C9",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",
		X"CC",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",X"CC",X"9C",X"66",X"00",X"99",X"CC",X"66",X"00",
		X"99",X"CC",X"66",X"00",X"99",X"CC",X"66",X"00",X"99",X"C9",X"66",X"00",X"CC",X"99",X"66",X"00",
		X"99",X"DD",X"66",X"00",X"6D",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",
		X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"90",X"66",X"66",X"66",X"90",
		X"66",X"66",X"96",X"90",X"66",X"66",X"96",X"90",X"99",X"66",X"66",X"90",X"95",X"66",X"66",X"90",
		X"95",X"99",X"66",X"90",X"95",X"DD",X"66",X"90",X"95",X"DD",X"66",X"90",X"95",X"DD",X"66",X"90",
		X"99",X"99",X"96",X"90",X"66",X"66",X"96",X"90",X"66",X"66",X"96",X"90",X"D6",X"66",X"96",X"90",
		X"9D",X"66",X"96",X"90",X"9D",X"66",X"96",X"90",X"96",X"69",X"96",X"90",X"96",X"99",X"96",X"90",
		X"66",X"99",X"96",X"90",X"66",X"9D",X"99",X"90",X"66",X"99",X"9C",X"90",X"66",X"09",X"99",X"90",
		X"66",X"09",X"99",X"00",X"69",X"09",X"99",X"00",X"69",X"09",X"99",X"90",X"99",X"99",X"99",X"99",
		X"90",X"99",X"09",X"C9",X"90",X"97",X"09",X"99",X"90",X"77",X"09",X"C9",X"90",X"99",X"09",X"99",
		X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"96",X"00",X"66",X"66",X"96",X"00",
		X"99",X"66",X"66",X"00",X"95",X"66",X"66",X"00",X"95",X"99",X"66",X"00",X"95",X"DD",X"66",X"00",
		X"95",X"DD",X"66",X"00",X"95",X"DD",X"66",X"00",X"99",X"99",X"66",X"00",X"66",X"66",X"66",X"00",
		X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"96",X"66",X"66",X"00",X"99",X"66",X"66",X"00",
		X"D9",X"66",X"66",X"00",X"99",X"66",X"66",X"00",X"C9",X"66",X"66",X"00",X"C9",X"66",X"99",X"00",
		X"C9",X"66",X"CC",X"00",X"C9",X"66",X"CC",X"00",X"99",X"66",X"CC",X"00",X"97",X"66",X"9C",X"00",
		X"77",X"99",X"9C",X"00",X"77",X"77",X"CC",X"00",X"79",X"77",X"CC",X"00",X"99",X"77",X"CC",X"00",
		X"77",X"99",X"CC",X"00",X"77",X"00",X"CC",X"00",X"99",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",
		X"00",X"E9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9E",X"00",X"00",X"99",X"9E",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9E",X"00",X"00",X"9E",X"99",X"00",X"09",X"EE",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"E9",X"00",X"99",X"99",X"9E",X"00",X"99",X"99",X"9B",X"00",
		X"E9",X"99",X"99",X"00",X"E9",X"99",X"E9",X"00",X"E9",X"9E",X"EE",X"00",X"9E",X"E9",X"E9",X"00",
		X"99",X"99",X"E9",X"00",X"99",X"9E",X"E9",X"00",X"EE",X"9E",X"E9",X"00",X"EE",X"EE",X"9B",X"00",
		X"99",X"E9",X"9E",X"00",X"9E",X"E9",X"9B",X"00",X"9E",X"99",X"9B",X"00",X"EE",X"EE",X"E9",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"E9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"9E",X"00",X"00",X"99",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9E",X"00",
		X"00",X"9E",X"99",X"00",X"09",X"EE",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"E9",X"00",
		X"99",X"99",X"9E",X"00",X"99",X"99",X"9B",X"00",X"E9",X"99",X"99",X"00",X"E9",X"99",X"99",X"00",
		X"E9",X"99",X"9E",X"00",X"9E",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"9E",X"99",X"00",
		X"EE",X"9E",X"E9",X"00",X"EE",X"EE",X"9B",X"00",X"99",X"E9",X"9E",X"00",X"9E",X"E9",X"9B",X"00",
		X"9E",X"99",X"9B",X"00",X"EE",X"E9",X"E9",X"00",X"EE",X"EE",X"E9",X"00",X"EE",X"EE",X"E9",X"00",
		X"9E",X"99",X"E9",X"00",X"9E",X"BE",X"E9",X"00",X"99",X"9B",X"E9",X"00",X"EE",X"9B",X"EE",X"00",
		X"E9",X"99",X"E4",X"00",X"99",X"E9",X"EE",X"00",X"99",X"E9",X"9E",X"00",X"E9",X"9E",X"9E",X"00",
		X"E9",X"99",X"9E",X"00",X"9E",X"E9",X"EE",X"00",X"99",X"99",X"E9",X"00",X"99",X"99",X"99",X"00",
		X"E9",X"9E",X"9E",X"00",X"E9",X"9E",X"99",X"00",X"99",X"99",X"E9",X"00",X"9E",X"9B",X"EE",X"00",
		X"9E",X"99",X"E9",X"00",X"99",X"09",X"E9",X"00",X"E9",X"09",X"99",X"00",X"E9",X"09",X"E9",X"00",
		X"99",X"00",X"99",X"00",X"E9",X"00",X"9B",X"00",X"E9",X"00",X"9B",X"00",X"9E",X"00",X"9B",X"00",
		X"9E",X"09",X"99",X"00",X"94",X"99",X"E9",X"00",X"99",X"9E",X"99",X"00",X"E9",X"99",X"EE",X"00",
		X"EE",X"E9",X"EE",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"9E",X"E9",X"00",X"9E",X"9E",X"E9",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"BE",X"E9",X"00",
		X"99",X"9B",X"E9",X"00",X"EE",X"99",X"E9",X"00",X"E9",X"99",X"E9",X"00",X"99",X"99",X"99",X"00",
		X"99",X"EE",X"99",X"00",X"E9",X"9E",X"99",X"00",X"E9",X"99",X"9B",X"00",X"9E",X"E9",X"9E",X"00",
		X"99",X"99",X"B9",X"00",X"E9",X"99",X"99",X"00",X"E9",X"9E",X"9E",X"00",X"99",X"9E",X"9E",X"00",
		X"E9",X"99",X"99",X"00",X"EE",X"9E",X"99",X"00",X"EE",X"99",X"9E",X"00",X"E9",X"09",X"9E",X"00",
		X"99",X"00",X"99",X"00",X"E9",X"00",X"9E",X"00",X"E9",X"00",X"EE",X"00",X"E9",X"00",X"E9",X"90",
		X"B9",X"00",X"E9",X"90",X"99",X"00",X"99",X"99",X"BB",X"00",X"99",X"E9",X"9E",X"00",X"E9",X"E9",
		X"99",X"00",X"EE",X"99",X"9B",X"90",X"9E",X"90",X"9E",X"90",X"9E",X"00",X"99",X"90",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"97",X"99",
		X"99",X"09",X"77",X"97",X"99",X"49",X"99",X"97",X"94",X"49",X"99",X"99",X"44",X"49",X"99",X"90",
		X"49",X"04",X"99",X"00",X"99",X"04",X"79",X"00",X"77",X"00",X"77",X"00",X"79",X"40",X"99",X"00",
		X"79",X"90",X"E9",X"00",X"99",X"94",X"EE",X"00",X"99",X"99",X"7E",X"00",X"99",X"79",X"77",X"00",
		X"94",X"79",X"77",X"00",X"94",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"99",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"09",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"97",X"77",X"77",X"00",X"77",X"97",X"79",X"00",
		X"77",X"99",X"99",X"00",X"99",X"44",X"97",X"00",X"94",X"99",X"77",X"00",X"44",X"49",X"77",X"00",
		X"00",X"00",X"09",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"93",X"00",X"00",X"99",X"99",X"09",
		X"00",X"79",X"77",X"00",X"99",X"79",X"99",X"00",X"77",X"99",X"9F",X"00",X"97",X"09",X"99",X"00",
		X"97",X"00",X"99",X"00",X"97",X"00",X"79",X"00",X"97",X"00",X"77",X"00",X"79",X"00",X"77",X"00",
		X"99",X"00",X"99",X"00",X"99",X"40",X"E7",X"00",X"F9",X"90",X"77",X"00",X"99",X"94",X"77",X"00",
		X"97",X"99",X"77",X"00",X"77",X"79",X"77",X"00",X"77",X"79",X"77",X"00",X"99",X"79",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"97",X"97",X"79",X"00",
		X"77",X"99",X"99",X"00",X"99",X"44",X"97",X"00",X"94",X"99",X"77",X"00",X"44",X"49",X"77",X"00",
		X"44",X"49",X"77",X"00",X"99",X"99",X"77",X"00",X"11",X"91",X"77",X"00",X"91",X"99",X"77",X"00",
		X"91",X"19",X"77",X"00",X"99",X"99",X"77",X"00",X"91",X"94",X"77",X"00",X"91",X"99",X"77",X"00",
		X"99",X"19",X"77",X"00",X"94",X"99",X"97",X"00",X"94",X"91",X"97",X"00",X"94",X"99",X"97",X"00",
		X"94",X"19",X"97",X"00",X"99",X"99",X"99",X"00",X"91",X"44",X"99",X"00",X"91",X"44",X"99",X"00",
		X"91",X"99",X"99",X"00",X"99",X"11",X"09",X"00",X"91",X"19",X"00",X"00",X"91",X"99",X"00",X"09",
		X"91",X"19",X"00",X"09",X"99",X"19",X"00",X"99",X"94",X"99",X"00",X"97",X"99",X"97",X"00",X"97",
		X"79",X"97",X"00",X"77",X"79",X"97",X"99",X"77",X"79",X"99",X"77",X"77",X"79",X"19",X"77",X"77",
		X"77",X"19",X"77",X"79",X"97",X"99",X"77",X"99",X"99",X"44",X"97",X"90",X"09",X"99",X"99",X"00",
		X"44",X"49",X"77",X"00",X"99",X"99",X"77",X"00",X"11",X"91",X"77",X"00",X"91",X"99",X"77",X"00",
		X"91",X"19",X"77",X"00",X"99",X"99",X"77",X"00",X"91",X"94",X"77",X"00",X"91",X"99",X"97",X"00",
		X"99",X"19",X"97",X"00",X"94",X"99",X"97",X"90",X"94",X"91",X"99",X"90",X"94",X"99",X"E9",X"99",
		X"94",X"19",X"79",X"79",X"99",X"99",X"79",X"79",X"91",X"44",X"99",X"99",X"91",X"44",X"90",X"00",
		X"91",X"99",X"90",X"99",X"99",X"11",X"00",X"79",X"91",X"19",X"00",X"79",X"91",X"99",X"00",X"79",
		X"91",X"19",X"00",X"79",X"99",X"19",X"00",X"79",X"94",X"99",X"99",X"99",X"99",X"97",X"77",X"00",
		X"79",X"97",X"77",X"00",X"79",X"97",X"77",X"00",X"79",X"99",X"77",X"00",X"79",X"19",X"77",X"00",
		X"97",X"19",X"77",X"00",X"99",X"99",X"79",X"00",X"09",X"44",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"29",X"00",X"90",X"99",X"29",X"99",
		X"99",X"99",X"29",X"99",X"99",X"99",X"29",X"90",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"90",
		X"99",X"92",X"99",X"99",X"99",X"92",X"29",X"90",X"99",X"92",X"99",X"00",X"99",X"29",X"99",X"09",
		X"99",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"22",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",
		X"90",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"90",
		X"99",X"92",X"99",X"99",X"99",X"92",X"29",X"90",X"99",X"92",X"99",X"00",X"99",X"29",X"99",X"00",
		X"99",X"29",X"99",X"00",X"99",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"22",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"22",
		X"99",X"99",X"D9",X"22",X"99",X"99",X"D9",X"22",X"99",X"99",X"D9",X"29",X"99",X"99",X"99",X"99",
		X"99",X"99",X"9D",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"90",
		X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"92",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"92",X"9D",X"00",X"99",X"99",X"D9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"E9",X"00",X"00",X"99",X"EE",X"09",X"00",X"39",X"EE",X"99",X"00",X"39",X"99",X"93",X"00",
		X"33",X"9F",X"33",X"00",X"39",X"99",X"33",X"00",X"99",X"F9",X"39",X"00",X"99",X"F9",X"99",X"00",
		X"93",X"9F",X"99",X"00",X"39",X"9F",X"39",X"00",X"99",X"99",X"93",X"00",X"93",X"33",X"93",X"00",
		X"99",X"33",X"99",X"00",X"09",X"33",X"99",X"00",X"09",X"33",X"90",X"00",X"00",X"33",X"99",X"00",
		X"00",X"33",X"39",X"00",X"90",X"39",X"33",X"00",X"99",X"99",X"93",X"00",X"39",X"9B",X"99",X"00",
		X"33",X"33",X"93",X"00",X"99",X"33",X"33",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"99",X"00",
		X"00",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"33",X"39",X"00",X"00",X"93",X"99",X"00",X"00",
		X"93",X"99",X"90",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"39",X"00",X"09",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"00",X"99",X"00",X"D9",X"00",X"9D",X"00",X"9D",X"00",X"D9",X"00",X"9D",X"00",X"D9",X"90",
		X"99",X"00",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",
		X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"09",
		X"09",X"99",X"09",X"09",X"00",X"99",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"D9",X"99",X"9D",X"00",X"9D",X"99",X"D9",X"00",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"DD",X"99",X"99",
		X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"90",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"DD",X"99",X"99",X"00",X"DD",X"99",X"D9",X"00",X"9D",X"DD",X"D9",X"00",X"99",X"DD",X"99",X"00",
		X"99",X"DD",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"0A",X"00",X"00",X"FF",X"AF",X"00",X"00",X"AA",X"AF",X"00",X"00",X"AF",X"FF",X"00",
		X"00",X"AF",X"FF",X"00",X"00",X"FF",X"AF",X"00",X"00",X"FF",X"AF",X"00",X"AA",X"FA",X"AA",X"00",
		X"FF",X"AA",X"FA",X"00",X"FF",X"AF",X"FF",X"A0",X"FF",X"FF",X"FF",X"A0",X"FF",X"FF",X"FF",X"A0",
		X"AF",X"AA",X"AF",X"00",X"AF",X"AF",X"AF",X"00",X"AF",X"AF",X"FF",X"00",X"FF",X"FF",X"AF",X"A0",
		X"FF",X"AA",X"AF",X"A0",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FA",X"00",X"AF",X"FF",X"FF",X"00",
		X"AF",X"FA",X"FF",X"00",X"AA",X"FA",X"FF",X"00",X"AA",X"FF",X"FA",X"00",X"FA",X"FF",X"AA",X"00",
		X"FA",X"AA",X"FF",X"00",X"AA",X"FA",X"FF",X"00",X"00",X"AA",X"FA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"AA",X"00",
		X"FA",X"00",X"FF",X"A0",X"AA",X"00",X"FF",X"AA",X"A0",X"00",X"FF",X"FA",X"A0",X"00",X"FF",X"AA",
		X"00",X"00",X"FF",X"A0",X"00",X"00",X"AF",X"A0",X"00",X"AA",X"AA",X"A0",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FA",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"A0",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"FA",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"0A",X"00",
		X"FF",X"00",X"0A",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"F3",X"F0",X"33",X"00",
		X"F0",X"F0",X"00",X"00",X"FF",X"F0",X"FF",X"AA",X"F3",X"F0",X"33",X"00",X"F0",X"F0",X"00",X"00",
		X"F0",X"30",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"A0",X"A0",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"90",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"F9",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"9F",X"59",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"F9",X"F5",X"00",X"00",X"F9",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9F",X"F5",X"00",X"00",X"99",X"F5",X"00",X"00",X"F9",X"F5",X"00",
		X"00",X"99",X"F5",X"00",X"00",X"9F",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"9F",X"59",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"F9",X"F5",X"00",X"00",X"F9",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9F",X"F5",X"00",X"00",X"99",X"F5",X"00",X"00",X"F9",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"FF",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"99",X"59",X"00",X"00",X"9F",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",
		X"9F",X"09",X"00",X"00",X"9F",X"99",X"60",X"00",X"F9",X"99",X"93",X"90",X"99",X"29",X"90",X"90",
		X"00",X"99",X"93",X"90",X"00",X"99",X"A0",X"90",X"00",X"99",X"9A",X"00",X"02",X"99",X"94",X"00",
		X"00",X"99",X"9A",X"00",X"10",X"99",X"97",X"00",X"00",X"99",X"9A",X"50",X"00",X"99",X"A0",X"00",
		X"04",X"99",X"A0",X"00",X"90",X"99",X"30",X"00",X"F9",X"99",X"44",X"90",X"F9",X"9E",X"00",X"90",
		X"FF",X"0E",X"00",X"90",X"F9",X"0E",X"00",X"00",X"F9",X"0E",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"03",X"50",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"09",X"90",X"09",X"00",X"00",X"99",X"09",X"00",
		X"90",X"94",X"09",X"00",X"99",X"94",X"99",X"00",X"A9",X"94",X"95",X"00",X"AA",X"44",X"55",X"00",
		X"AA",X"94",X"59",X"90",X"3A",X"A9",X"99",X"90",X"33",X"9A",X"AA",X"99",X"AA",X"AA",X"A3",X"A9",
		X"33",X"99",X"A3",X"39",X"3A",X"99",X"AA",X"A9",X"A5",X"44",X"9A",X"A9",X"33",X"44",X"99",X"59",
		X"3A",X"99",X"49",X"A9",X"3A",X"9F",X"49",X"39",X"A9",X"9F",X"49",X"A9",X"99",X"9F",X"49",X"39",
		X"90",X"9F",X"99",X"A9",X"90",X"9A",X"99",X"A9",X"00",X"99",X"90",X"A9",X"00",X"94",X"90",X"A9",
		X"00",X"49",X"99",X"39",X"00",X"99",X"59",X"A9",X"00",X"90",X"95",X"39",X"09",X"99",X"99",X"A9",
		X"09",X"59",X"59",X"A9",X"09",X"99",X"99",X"A9",X"00",X"00",X"59",X"A9",X"00",X"00",X"99",X"99",
		X"09",X"00",X"99",X"00",X"09",X"00",X"A9",X"00",X"09",X"90",X"A9",X"00",X"00",X"99",X"39",X"00",
		X"00",X"94",X"39",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"44",X"55",X"00",
		X"00",X"94",X"59",X"00",X"00",X"A9",X"99",X"00",X"00",X"9A",X"33",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"99",X"AA",X"00",X"00",X"99",X"A3",X"00",X"00",X"44",X"9A",X"00",X"00",X"44",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"9F",X"49",X"00",X"00",X"9F",X"49",X"00",X"00",X"9F",X"49",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"94",X"9A",X"00",
		X"00",X"49",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"59",X"59",X"00",X"09",X"99",X"99",X"00",X"09",X"00",X"A9",X"00",X"09",X"00",X"9A",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"94",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"44",X"55",X"00",
		X"00",X"94",X"A9",X"00",X"00",X"A9",X"99",X"00",X"00",X"AA",X"33",X"00",X"00",X"AA",X"AA",X"00",
		X"09",X"99",X"3A",X"00",X"09",X"99",X"A3",X"00",X"09",X"44",X"9A",X"00",X"09",X"44",X"99",X"00",
		X"09",X"99",X"49",X"00",X"09",X"9F",X"49",X"00",X"09",X"9F",X"49",X"00",X"99",X"9F",X"49",X"00",
		X"9A",X"9A",X"99",X"00",X"9A",X"99",X"99",X"00",X"9A",X"99",X"9A",X"00",X"9A",X"94",X"9A",X"00",
		X"9A",X"49",X"99",X"00",X"9A",X"99",X"59",X"00",X"9A",X"90",X"95",X"00",X"99",X"99",X"59",X"00",
		X"09",X"59",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"90",X"00",
		X"99",X"99",X"49",X"00",X"94",X"22",X"44",X"00",X"44",X"99",X"94",X"00",X"44",X"99",X"99",X"00",
		X"15",X"99",X"95",X"99",X"55",X"99",X"55",X"19",X"51",X"99",X"15",X"E9",X"11",X"17",X"11",X"99",
		X"91",X"77",X"11",X"90",X"EE",X"77",X"EE",X"00",X"99",X"77",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"90",X"00",
		X"99",X"99",X"49",X"00",X"94",X"22",X"44",X"00",X"44",X"99",X"94",X"00",X"44",X"99",X"29",X"00",
		X"17",X"99",X"97",X"99",X"77",X"99",X"77",X"19",X"71",X"99",X"17",X"E9",X"11",X"15",X"11",X"99",
		X"91",X"55",X"11",X"90",X"EE",X"55",X"EE",X"00",X"99",X"55",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"90",X"E0",X"00",X"00",X"90",X"EE",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"FF",X"90",X"00",
		X"99",X"F4",X"F9",X"00",X"39",X"FF",X"4F",X"00",X"33",X"FF",X"FF",X"00",X"39",X"99",X"FF",X"00",
		X"3B",X"99",X"F4",X"00",X"9B",X"FF",X"FF",X"00",X"93",X"FF",X"99",X"00",X"93",X"99",X"33",X"00",
		X"09",X"33",X"33",X"07",X"09",X"99",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"9F",X"33",X"00",
		X"50",X"99",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"50",X"10",X"3B",X"99",X"00",
		X"11",X"39",X"99",X"00",X"A1",X"33",X"99",X"07",X"99",X"33",X"94",X"40",X"14",X"43",X"79",X"00",
		X"95",X"49",X"95",X"00",X"57",X"B5",X"54",X"50",X"71",X"45",X"11",X"45",X"49",X"17",X"A1",X"00",
		X"04",X"59",X"59",X"00",X"11",X"9A",X"55",X"00",X"05",X"0A",X"10",X"40",X"00",X"00",X"11",X"04",
		X"00",X"0E",X"E0",X"00",X"90",X"EE",X"E0",X"00",X"90",X"9E",X"00",X"00",X"90",X"33",X"E0",X"00",
		X"99",X"99",X"90",X"00",X"39",X"9A",X"99",X"00",X"33",X"AF",X"A3",X"00",X"39",X"FF",X"FF",X"00",
		X"3B",X"99",X"FF",X"00",X"9B",X"99",X"F9",X"00",X"93",X"FF",X"99",X"00",X"93",X"99",X"33",X"00",
		X"09",X"33",X"33",X"00",X"09",X"93",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"B9",X"33",X"00",
		X"00",X"3B",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"00",X"00",X"3B",X"99",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"09",X"33",X"90",X"00",X"99",X"33",X"99",X"00",
		X"33",X"33",X"39",X"00",X"39",X"93",X"99",X"00",X"99",X"93",X"93",X"00",X"09",X"19",X"33",X"00",
		X"00",X"39",X"33",X"00",X"00",X"39",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"90",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"59",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"9F",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"49",X"00",X"00",X"99",X"49",X"00",
		X"09",X"BB",X"99",X"90",X"09",X"BB",X"9B",X"90",X"99",X"BB",X"BB",X"90",X"99",X"BB",X"B9",X"90",
		X"11",X"99",X"B9",X"90",X"E1",X"99",X"BB",X"00",X"EE",X"99",X"99",X"00",X"1E",X"99",X"59",X"00",
		X"1E",X"99",X"99",X"00",X"11",X"B9",X"99",X"99",X"11",X"BB",X"9B",X"B1",X"11",X"9B",X"BB",X"99",
		X"11",X"99",X"99",X"B9",X"11",X"BB",X"90",X"91",X"99",X"BB",X"90",X"99",X"9B",X"BB",X"90",X"90",
		X"BB",X"BB",X"90",X"00",X"9B",X"BB",X"90",X"00",X"9B",X"1B",X"99",X"00",X"99",X"9B",X"99",X"19",
		X"90",X"B9",X"9B",X"B9",X"90",X"B9",X"9B",X"19",X"90",X"BB",X"9B",X"B9",X"00",X"BB",X"99",X"99",
		X"00",X"BB",X"09",X"90",X"00",X"BB",X"09",X"00",X"00",X"9B",X"09",X"00",X"00",X"99",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9E",X"00",X"99",X"00",X"99",X"00",X"39",X"00",X"19",X"99",X"39",X"00",
		X"11",X"BB",X"99",X"90",X"E1",X"BB",X"9B",X"90",X"EE",X"BB",X"BB",X"90",X"EE",X"BB",X"B9",X"90",
		X"1E",X"B9",X"B9",X"90",X"11",X"99",X"BB",X"00",X"11",X"99",X"99",X"00",X"11",X"99",X"59",X"90",
		X"11",X"B9",X"99",X"90",X"11",X"BB",X"BB",X"99",X"99",X"9B",X"99",X"B9",X"BB",X"99",X"BB",X"B9",
		X"B9",X"BB",X"BB",X"99",X"BB",X"BB",X"99",X"00",X"9B",X"BB",X"99",X"00",X"09",X"BB",X"90",X"00",
		X"00",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"1B",X"99",X"00",X"00",X"9B",X"99",X"19",
		X"00",X"B9",X"9B",X"B9",X"00",X"B9",X"9B",X"19",X"00",X"BB",X"9B",X"B9",X"00",X"BB",X"99",X"99",
		X"00",X"BB",X"09",X"90",X"00",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",
		X"00",X"66",X"99",X"00",X"99",X"66",X"69",X"00",X"99",X"66",X"99",X"00",X"EE",X"96",X"99",X"00",
		X"9E",X"99",X"96",X"00",X"49",X"E9",X"96",X"00",X"49",X"EC",X"96",X"00",X"99",X"E9",X"96",X"00",
		X"99",X"C9",X"96",X"00",X"CC",X"CC",X"96",X"00",X"CC",X"99",X"96",X"00",X"9C",X"C9",X"96",X"00",
		X"99",X"C9",X"99",X"00",X"99",X"C9",X"99",X"00",X"CC",X"C9",X"99",X"00",X"CC",X"99",X"66",X"00",
		X"9C",X"96",X"66",X"00",X"99",X"69",X"66",X"00",X"66",X"69",X"69",X"00",X"66",X"99",X"99",X"00",
		X"96",X"96",X"90",X"00",X"99",X"99",X"90",X"00",X"C9",X"CC",X"90",X"00",X"99",X"CC",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"79",X"00",X"00",X"97",X"79",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",
		X"09",X"66",X"99",X"00",X"99",X"66",X"69",X"00",X"EE",X"96",X"96",X"00",X"99",X"99",X"96",X"00",
		X"49",X"E9",X"96",X"00",X"49",X"EC",X"96",X"00",X"99",X"E9",X"96",X"00",X"99",X"C9",X"96",X"00",
		X"CC",X"CC",X"96",X"00",X"CC",X"99",X"96",X"00",X"9C",X"C9",X"96",X"00",X"99",X"C9",X"96",X"00",
		X"99",X"C9",X"96",X"00",X"99",X"C9",X"99",X"00",X"CC",X"99",X"99",X"00",X"9C",X"99",X"99",X"00",
		X"99",X"66",X"96",X"00",X"00",X"66",X"96",X"00",X"00",X"69",X"96",X"00",X"00",X"69",X"96",X"00",
		X"09",X"99",X"96",X"99",X"09",X"90",X"96",X"79",X"09",X"90",X"96",X"79",X"99",X"00",X"96",X"79",
		X"77",X"00",X"96",X"79",X"77",X"00",X"99",X"79",X"99",X"00",X"00",X"79",X"00",X"00",X"00",X"99",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"99",X"99",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"99",X"E9",X"99",X"BB",X"9E",X"EE",X"E9",
		X"BB",X"99",X"EE",X"99",X"99",X"99",X"E9",X"00",X"E9",X"99",X"99",X"90",X"E9",X"99",X"EE",X"90",
		X"E9",X"99",X"EE",X"90",X"EB",X"99",X"99",X"90",X"9B",X"99",X"9E",X"90",X"99",X"E9",X"9E",X"90",
		X"99",X"E9",X"99",X"00",X"99",X"E9",X"99",X"00",X"99",X"9E",X"90",X"00",X"9E",X"9E",X"99",X"00",
		X"9E",X"99",X"E9",X"00",X"99",X"09",X"E9",X"00",X"EE",X"09",X"EE",X"00",X"99",X"09",X"E9",X"00",
		X"E9",X"09",X"99",X"00",X"E9",X"00",X"9E",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"99",X"00",X"99",X"99",X"E9",X"00",X"E9",X"99",X"EE",X"00",X"E9",X"9E",X"99",X"00",
		X"E9",X"99",X"E9",X"00",X"E9",X"99",X"E1",X"00",X"99",X"99",X"E9",X"90",X"E9",X"99",X"99",X"90",
		X"99",X"99",X"E9",X"99",X"9E",X"99",X"99",X"E9",X"9E",X"99",X"9E",X"E9",X"99",X"E9",X"99",X"99",
		X"9B",X"E9",X"90",X"99",X"9B",X"E9",X"90",X"E9",X"9B",X"9E",X"99",X"99",X"9E",X"9E",X"E9",X"90",
		X"9E",X"99",X"99",X"90",X"99",X"00",X"9B",X"00",X"49",X"00",X"EB",X"00",X"49",X"00",X"99",X"00",
		X"99",X"00",X"E9",X"00",X"9E",X"00",X"E9",X"90",X"9B",X"00",X"99",X"90",X"99",X"00",X"09",X"90",
		X"99",X"00",X"99",X"00",X"77",X"00",X"77",X"00",X"97",X"00",X"77",X"00",X"99",X"00",X"99",X"90",
		X"99",X"99",X"9F",X"99",X"97",X"79",X"99",X"79",X"77",X"79",X"99",X"79",X"77",X"79",X"99",X"99",
		X"79",X"77",X"77",X"90",X"99",X"77",X"99",X"00",X"97",X"77",X"99",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"90",X"77",X"77",X"77",X"99",X"77",X"99",X"97",X"79",X"97",X"94",X"97",X"79",
		X"94",X"94",X"97",X"79",X"94",X"94",X"97",X"79",X"9A",X"99",X"97",X"79",X"99",X"19",X"97",X"79",
		X"90",X"99",X"99",X"49",X"00",X"91",X"77",X"49",X"00",X"99",X"77",X"A9",X"00",X"91",X"97",X"99",
		X"00",X"91",X"99",X"90",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"97",X"90",X"00",X"00",X"77",X"90",X"00",X"00",X"77",X"90",X"00",X"00",X"99",X"90",
		X"99",X"00",X"99",X"00",X"77",X"00",X"77",X"00",X"97",X"00",X"77",X"00",X"99",X"00",X"99",X"90",
		X"99",X"99",X"9F",X"99",X"99",X"79",X"99",X"79",X"99",X"79",X"99",X"79",X"49",X"79",X"49",X"99",
		X"97",X"77",X"49",X"90",X"77",X"77",X"97",X"00",X"99",X"77",X"77",X"00",X"09",X"77",X"99",X"00",
		X"99",X"77",X"77",X"00",X"97",X"77",X"77",X"00",X"97",X"99",X"77",X"00",X"97",X"94",X"77",X"00",
		X"77",X"94",X"77",X"00",X"77",X"94",X"77",X"00",X"77",X"99",X"77",X"00",X"77",X"19",X"79",X"90",
		X"77",X"99",X"49",X"90",X"77",X"91",X"49",X"90",X"77",X"99",X"79",X"99",X"77",X"91",X"79",X"99",
		X"77",X"99",X"A9",X"99",X"99",X"00",X"99",X"79",X"09",X"00",X"09",X"99",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"29",X"00",X"99",X"92",X"29",X"00",X"99",X"99",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"90",X"29",X"00",X"99",X"99",X"29",X"00",
		X"99",X"22",X"29",X"00",X"09",X"92",X"22",X"00",X"09",X"99",X"92",X"00",X"99",X"99",X"92",X"00",
		X"99",X"49",X"29",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"59",X"99",X"90",
		X"09",X"99",X"99",X"90",X"09",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"59",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"D9",X"00",X"00",X"29",X"D9",X"00",
		X"00",X"29",X"D9",X"00",X"09",X"29",X"D9",X"00",X"49",X"22",X"D9",X"99",X"92",X"22",X"D9",X"29",
		X"99",X"99",X"D9",X"29",X"09",X"95",X"99",X"99",X"00",X"99",X"99",X"90",X"99",X"99",X"22",X"90",
		X"92",X"99",X"2A",X"90",X"99",X"99",X"22",X"99",X"29",X"59",X"29",X"D9",X"A2",X"99",X"99",X"D9",
		X"99",X"22",X"9D",X"D9",X"99",X"99",X"9D",X"D9",X"DD",X"92",X"9D",X"90",X"DD",X"22",X"D2",X"00",
		X"D2",X"22",X"DD",X"00",X"2D",X"2A",X"DD",X"00",X"DD",X"22",X"D9",X"00",X"DD",X"22",X"99",X"00",
		X"9D",X"22",X"90",X"00",X"99",X"22",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"92",X"00",X"09",X"00",X"99",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"D9",X"00",X"00",X"29",X"D9",X"00",
		X"00",X"29",X"D9",X"00",X"09",X"29",X"D9",X"00",X"99",X"22",X"D9",X"00",X"92",X"22",X"D9",X"00",
		X"99",X"99",X"99",X"00",X"09",X"95",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",X"00",
		X"92",X"95",X"D9",X"00",X"99",X"99",X"D9",X"00",X"09",X"22",X"DD",X"00",X"00",X"99",X"2D",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"A2",X"DD",X"00",X"00",X"99",X"DD",X"00",X"00",X"92",X"D2",X"00",
		X"00",X"92",X"2D",X"00",X"00",X"99",X"DD",X"00",X"00",X"29",X"DD",X"00",X"00",X"D9",X"DD",X"00",
		X"00",X"99",X"DD",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"0E",X"E0",X"00",X"90",X"EE",X"E0",X"00",X"90",X"9E",X"00",X"00",X"90",X"33",X"E0",X"00",
		X"99",X"99",X"90",X"00",X"39",X"9F",X"99",X"00",X"33",X"FF",X"93",X"00",X"39",X"FF",X"93",X"00",
		X"3B",X"AF",X"93",X"00",X"9B",X"9A",X"93",X"00",X"93",X"99",X"39",X"00",X"93",X"33",X"33",X"00",
		X"09",X"33",X"33",X"00",X"09",X"99",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"33",X"00",
		X"00",X"39",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"00",X"00",X"3B",X"99",X"00",
		X"00",X"39",X"99",X"00",X"99",X"33",X"44",X"00",X"94",X"33",X"94",X"00",X"44",X"93",X"99",X"00",
		X"15",X"99",X"95",X"99",X"55",X"B9",X"55",X"19",X"51",X"99",X"15",X"E9",X"11",X"17",X"11",X"99",
		X"91",X"77",X"11",X"90",X"EE",X"77",X"EE",X"00",X"99",X"77",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"9E",X"00",X"00",X"90",X"E3",X"00",X"00",X"99",X"99",X"99",X"00",
		X"39",X"9F",X"39",X"00",X"33",X"F9",X"93",X"00",X"39",X"F9",X"93",X"00",X"3B",X"A9",X"93",X"00",
		X"9B",X"9F",X"93",X"00",X"93",X"99",X"39",X"00",X"93",X"33",X"33",X"00",X"09",X"33",X"33",X"00",
		X"09",X"99",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"99",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"99",X"00",X"00",X"39",X"00",X"00",
		X"00",X"33",X"99",X"00",X"99",X"33",X"44",X"00",X"94",X"33",X"94",X"00",X"44",X"93",X"99",X"00",
		X"17",X"99",X"97",X"99",X"77",X"B9",X"77",X"19",X"71",X"99",X"17",X"E9",X"11",X"15",X"11",X"99",
		X"91",X"55",X"11",X"90",X"EE",X"55",X"EE",X"00",X"99",X"55",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9A",X"99",X"00",X"00",X"9A",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"F9",X"95",X"00",X"00",X"F9",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"94",X"F5",X"00",X"00",X"99",X"F5",X"00",X"00",X"F9",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"F9",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"94",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",
		X"9F",X"04",X"00",X"00",X"9F",X"94",X"60",X"00",X"F9",X"94",X"A3",X"90",X"99",X"29",X"90",X"90",
		X"00",X"94",X"93",X"90",X"00",X"99",X"A0",X"90",X"00",X"4A",X"9A",X"00",X"02",X"94",X"94",X"00",
		X"00",X"94",X"9A",X"00",X"10",X"99",X"97",X"00",X"00",X"49",X"9A",X"50",X"00",X"99",X"A0",X"00",
		X"04",X"9A",X"A0",X"00",X"90",X"4A",X"30",X"00",X"F9",X"49",X"44",X"90",X"F9",X"9A",X"00",X"90",
		X"FF",X"0E",X"00",X"90",X"F9",X"0E",X"00",X"00",X"F9",X"0E",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"03",X"50",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
