library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom3 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"20",X"4C",X"45",X"53",X"20",X"50",X"49",X"45",X"43",X"45",X"D3",X"42",X"4F",X"4E",X"55",X"53",
		X"20",X"56",X"49",X"4C",X"4C",X"C5",X"42",X"4F",X"4E",X"55",X"53",X"20",X"50",X"4F",X"49",X"4E",
		X"54",X"D3",X"58",X"20",X"50",X"4F",X"49",X"4E",X"54",X"D3",X"46",X"49",X"CE",X"31",X"20",X"50",
		X"49",X"45",X"43",X"45",X"20",X"32",X"20",X"4A",X"4F",X"55",X"45",X"55",X"52",X"D3",X"31",X"20",
		X"50",X"49",X"45",X"43",X"45",X"20",X"31",X"20",X"4A",X"4F",X"55",X"45",X"55",X"D2",X"32",X"20",
		X"50",X"49",X"45",X"43",X"45",X"53",X"20",X"31",X"20",X"4A",X"4F",X"55",X"45",X"55",X"D2",X"53",
		X"50",X"4C",X"45",X"4E",X"44",X"49",X"44",X"45",X"20",X"53",X"43",X"4F",X"52",X"C5",X"53",X"56",
		X"50",X"20",X"45",X"4E",X"54",X"52",X"45",X"5A",X"20",X"56",X"4F",X"53",X"20",X"49",X"4E",X"49",
		X"54",X"49",X"41",X"4C",X"45",X"D3",X"54",X"4F",X"55",X"52",X"4E",X"45",X"5A",X"20",X"42",X"4F",
		X"55",X"4C",X"45",X"20",X"50",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",
		X"C5",X"50",X"4F",X"55",X"53",X"53",X"45",X"5A",X"20",X"46",X"45",X"55",X"20",X"51",X"55",X"41",
		X"4E",X"44",X"20",X"43",X"4F",X"52",X"52",X"45",X"43",X"54",X"C5",X"4D",X"45",X"49",X"4C",X"4C",
		X"45",X"55",X"52",X"53",X"20",X"53",X"43",X"4F",X"52",X"45",X"D3",X"44",X"45",X"46",X"45",X"4E",
		X"53",X"45",X"5A",X"20",X"20",X"20",X"20",X"20",X"56",X"49",X"4C",X"4C",X"45",X"D3",X"42",X"41",
		X"D3",X"56",X"49",X"44",X"C5",X"C1",X"53",X"50",X"49",X"45",X"4C",X"45",X"D2",X"53",X"50",X"49",
		X"45",X"4C",X"45",X"4E",X"44",X"C5",X"53",X"54",X"41",X"52",X"54",X"4B",X"4E",X"24",X"50",X"46",
		X"45",X"20",X"44",X"52",X"25",X"43",X"4B",X"45",X"CE",X"47",X"45",X"4C",X"44",X"20",X"45",X"49",
		X"4E",X"57",X"45",X"52",X"46",X"45",X"CE",X"42",X"4F",X"4E",X"55",X"53",X"53",X"54",X"41",X"44",
		X"D4",X"42",X"4F",X"4E",X"55",X"53",X"50",X"55",X"4E",X"4B",X"54",X"C5",X"58",X"20",X"50",X"55",
		X"4E",X"4B",X"54",X"C5",X"45",X"4E",X"44",X"C5",X"31",X"20",X"4D",X"25",X"4E",X"5A",X"20",X"32",
		X"20",X"53",X"50",X"49",X"45",X"4C",X"C5",X"31",X"20",X"4D",X"25",X"4E",X"5A",X"45",X"20",X"31",
		X"20",X"53",X"50",X"49",X"45",X"CC",X"32",X"20",X"4D",X"25",X"4E",X"5A",X"45",X"4E",X"20",X"31",
		X"20",X"53",X"50",X"49",X"45",X"CC",X"4B",X"52",X"45",X"44",X"49",X"54",X"45",X"BA",X"50",X"52",
		X"49",X"4D",X"41",X"20",X"45",X"52",X"47",X"45",X"42",X"4E",X"49",X"D3",X"47",X"45",X"42",X"45",
		X"4E",X"20",X"53",X"49",X"45",X"20",X"49",X"48",X"52",X"45",X"20",X"49",X"4E",X"49",X"54",X"49",
		X"41",X"4C",X"45",X"4E",X"20",X"45",X"49",X"CE",X"42",X"41",X"4C",X"4C",X"20",X"44",X"52",X"45",
		X"48",X"45",X"4E",X"20",X"46",X"25",X"52",X"20",X"41",X"4C",X"4C",X"45",X"20",X"42",X"55",X"43",
		X"48",X"53",X"54",X"41",X"42",X"45",X"CE",X"46",X"49",X"52",X"45",X"20",X"44",X"52",X"25",X"43",
		X"4B",X"45",X"4E",X"20",X"57",X"45",X"4E",X"4E",X"20",X"52",X"49",X"43",X"48",X"54",X"49",X"C7",
		X"48",X"24",X"43",X"48",X"53",X"54",X"5A",X"41",X"48",X"4C",X"45",X"CE",X"53",X"54",X"23",X"44",
		X"54",X"45",X"20",X"20",X"20",X"20",X"20",X"56",X"45",X"52",X"54",X"45",X"49",X"44",X"49",X"47",
		X"45",X"CE",X"57",X"45",X"4E",X"49",X"C7",X"4C",X"45",X"45",X"D2",X"4A",X"45",X"44",X"C5",X"4A",
		X"55",X"47",X"41",X"44",X"4F",X"D2",X"4A",X"55",X"45",X"47",X"4F",X"20",X"54",X"45",X"52",X"4D",
		X"49",X"4E",X"41",X"44",X"CF",X"50",X"55",X"4C",X"53",X"41",X"52",X"20",X"53",X"54",X"41",X"52",
		X"D4",X"49",X"4E",X"53",X"45",X"52",X"54",X"45",X"20",X"46",X"49",X"43",X"48",X"41",X"D3",X"43",
		X"49",X"55",X"44",X"41",X"44",X"20",X"45",X"58",X"54",X"52",X"C1",X"42",X"4F",X"4E",X"49",X"46",
		X"49",X"43",X"41",X"43",X"49",X"4F",X"4E",X"20",X"44",X"45",X"20",X"50",X"55",X"4E",X"54",X"4F",
		X"D3",X"58",X"20",X"50",X"55",X"4E",X"54",X"4F",X"D3",X"31",X"20",X"4D",X"4F",X"4E",X"45",X"44",
		X"41",X"20",X"32",X"20",X"4A",X"55",X"45",X"47",X"4F",X"D3",X"31",X"20",X"4D",X"4F",X"4E",X"45",
		X"44",X"41",X"20",X"31",X"20",X"4A",X"55",X"45",X"47",X"CF",X"32",X"20",X"4D",X"4F",X"4E",X"45",
		X"44",X"41",X"53",X"20",X"31",X"20",X"4A",X"55",X"45",X"47",X"CF",X"43",X"52",X"45",X"44",X"49",
		X"54",X"4F",X"53",X"BA",X"47",X"52",X"41",X"4E",X"20",X"50",X"55",X"4E",X"54",X"41",X"4A",X"C5",
		X"45",X"4E",X"54",X"52",X"45",X"20",X"53",X"55",X"53",X"20",X"49",X"4E",X"49",X"43",X"49",X"41",
		X"4C",X"45",X"D3",X"47",X"49",X"52",X"45",X"20",X"4C",X"41",X"20",X"42",X"4F",X"4C",X"41",X"20",
		X"50",X"41",X"52",X"41",X"20",X"43",X"41",X"4D",X"42",X"49",X"41",X"52",X"20",X"4C",X"45",X"54",
		X"52",X"41",X"D3",X"4F",X"50",X"52",X"49",X"4D",X"41",X"20",X"46",X"49",X"52",X"45",X"20",X"50",
		X"4F",X"52",X"20",X"4C",X"41",X"20",X"4C",X"45",X"54",X"52",X"C1",X"52",X"45",X"43",X"4F",X"52",
		X"44",X"D3",X"44",X"45",X"46",X"49",X"45",X"4E",X"44",X"41",X"20",X"20",X"20",X"20",X"20",X"43",
		X"49",X"55",X"44",X"41",X"44",X"45",X"D3",X"50",X"4F",X"43",X"CF",X"53",X"49",X"CE",X"43",X"41",
		X"44",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"C6",X"C6",X"C6",X"44",
		X"38",X"00",X"FC",X"30",X"30",X"30",X"30",X"70",X"30",X"00",X"FE",X"E0",X"78",X"3C",X"0E",X"C6",
		X"7C",X"00",X"7C",X"C6",X"06",X"3C",X"18",X"0C",X"7E",X"00",X"0C",X"0C",X"FE",X"CC",X"6C",X"3C",
		X"1C",X"00",X"7C",X"C6",X"06",X"06",X"FC",X"C0",X"FC",X"00",X"7C",X"C6",X"C6",X"FC",X"C0",X"60",
		X"3C",X"00",X"30",X"30",X"30",X"18",X"0C",X"C6",X"FE",X"00",X"7C",X"86",X"9E",X"78",X"E4",X"C4",
		X"78",X"00",X"78",X"0C",X"06",X"7E",X"C6",X"C6",X"7C",X"00",X"C6",X"C6",X"FE",X"C6",X"C6",X"6C",
		X"38",X"00",X"FC",X"C6",X"C6",X"FC",X"C6",X"C6",X"FC",X"00",X"3C",X"66",X"C0",X"C0",X"C0",X"66",
		X"3C",X"00",X"F8",X"CC",X"C6",X"C6",X"C6",X"CC",X"F8",X"00",X"FC",X"C0",X"C0",X"F8",X"C0",X"C0",
		X"FC",X"00",X"C0",X"C0",X"C0",X"FC",X"C0",X"C0",X"FE",X"00",X"3E",X"66",X"C6",X"CE",X"C0",X"60",
		X"3E",X"00",X"C6",X"C6",X"C6",X"FE",X"C6",X"C6",X"C6",X"00",X"FC",X"30",X"30",X"30",X"30",X"30",
		X"FC",X"00",X"7C",X"C6",X"06",X"06",X"06",X"06",X"06",X"00",X"CE",X"DC",X"F8",X"F0",X"D8",X"CC",
		X"C6",X"00",X"FC",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"C6",X"C6",X"D6",X"FE",X"FE",X"EE",
		X"C6",X"00",X"C6",X"CE",X"DE",X"FE",X"F6",X"E6",X"C6",X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",
		X"7C",X"00",X"C0",X"C0",X"FC",X"C6",X"C6",X"C6",X"FC",X"00",X"7A",X"CC",X"DE",X"C6",X"C6",X"C6",
		X"7C",X"00",X"CE",X"DC",X"F8",X"CE",X"C6",X"C6",X"FC",X"00",X"7C",X"C6",X"06",X"7C",X"C0",X"C6",
		X"7C",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"FC",X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",
		X"C6",X"00",X"10",X"38",X"6C",X"EE",X"C6",X"C6",X"C6",X"00",X"C6",X"EE",X"FE",X"FE",X"D6",X"C6",
		X"C6",X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"30",X"30",X"30",X"78",X"CC",X"CC",
		X"CC",X"00",X"FE",X"E0",X"70",X"38",X"1C",X"0E",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"3C",X"7E",X"FF",X"FF",X"BD",X"3C",X"3C",X"7F",X"FF",X"7F",X"7E",X"34",X"30",
		X"20",X"00",X"7C",X"37",X"25",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FE",X"FE",X"FA",X"50",
		X"10",X"10",X"3E",X"6C",X"C8",X"C0",X"80",X"00",X"00",X"00",X"1C",X"38",X"7F",X"FF",X"FF",X"7F",
		X"38",X"1C",X"38",X"1C",X"FE",X"FF",X"FF",X"FE",X"1C",X"38",X"3C",X"42",X"99",X"91",X"99",X"42",
		X"3C",X"00",X"30",X"30",X"00",X"30",X"30",X"00",X"00",X"00",X"3C",X"52",X"9D",X"95",X"9D",X"42",
		X"3C",X"00",X"C6",X"FE",X"C6",X"6C",X"38",X"10",X"44",X"00",X"7C",X"C6",X"C6",X"C6",X"7C",X"00",
		X"28",X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"00",X"28",X"00",X"A5",X"F4",X"29",X"70",X"C9",X"70",
		X"F0",X"2E",X"A9",X"1B",X"20",X"51",X"6A",X"A9",X"19",X"20",X"51",X"6A",X"A9",X"1A",X"20",X"51",
		X"6A",X"A9",X"00",X"85",X"D1",X"A5",X"F4",X"29",X"70",X"4A",X"4A",X"4A",X"AA",X"BD",X"82",X"60",
		X"85",X"D2",X"BD",X"83",X"60",X"85",X"D3",X"A2",X"90",X"A0",X"58",X"A9",X"40",X"20",X"F6",X"6A",
		X"60",X"A2",X"17",X"BD",X"F3",X"74",X"9D",X"2C",X"00",X"BD",X"0B",X"75",X"9D",X"44",X"00",X"CA",
		X"10",X"F1",X"60",X"47",X"4A",X"4C",X"44",X"45",X"57",X"4A",X"45",X"44",X"4D",X"4A",X"50",X"52",
		X"44",X"41",X"53",X"52",X"43",X"44",X"4C",X"53",X"44",X"46",X"D4",X"50",X"69",X"00",X"05",X"70",
		X"00",X"50",X"71",X"00",X"00",X"72",X"00",X"50",X"72",X"00",X"30",X"73",X"00",X"95",X"74",X"00",
		X"00",X"75",X"00",X"AD",X"59",X"00",X"85",X"D1",X"AD",X"5A",X"00",X"85",X"D2",X"AD",X"5B",X"00",
		X"85",X"D3",X"A2",X"64",X"A0",X"E2",X"A9",X"40",X"20",X"F6",X"6A",X"4C",X"E1",X"5F",X"22",X"20",
		X"E4",X"76",X"A5",X"93",X"D0",X"07",X"A0",X"1C",X"84",X"91",X"B8",X"50",X"3D",X"A2",X"01",X"86",
		X"8D",X"A0",X"15",X"B9",X"46",X"00",X"DD",X"DA",X"01",X"D0",X"0E",X"B9",X"45",X"00",X"DD",X"D8",
		X"01",X"D0",X"06",X"B9",X"44",X"00",X"DD",X"D6",X"01",X"B0",X"03",X"20",X"8B",X"75",X"88",X"88",
		X"88",X"10",X"E0",X"CA",X"10",X"DB",X"20",X"33",X"6C",X"A5",X"8D",X"10",X"09",X"20",X"21",X"69",
		X"20",X"E4",X"75",X"B8",X"50",X"04",X"A0",X"06",X"84",X"91",X"60",X"84",X"98",X"A0",X"00",X"C4",
		X"98",X"D0",X"27",X"BD",X"DA",X"01",X"99",X"46",X"00",X"BD",X"D8",X"01",X"99",X"45",X"00",X"BD",
		X"D6",X"01",X"99",X"44",X"00",X"E8",X"8A",X"CA",X"99",X"2C",X"00",X"A9",X"5B",X"99",X"2D",X"00",
		X"99",X"2E",X"00",X"A0",X"00",X"A9",X"FF",X"85",X"8D",X"60",X"B9",X"49",X"00",X"99",X"46",X"00",
		X"B9",X"48",X"00",X"99",X"45",X"00",X"B9",X"47",X"00",X"99",X"44",X"00",X"B9",X"31",X"00",X"99",
		X"2E",X"00",X"B9",X"30",X"00",X"99",X"2D",X"00",X"B9",X"2F",X"00",X"99",X"2C",X"00",X"C8",X"C8",
		X"C8",X"10",X"AC",X"60",X"A0",X"15",X"B9",X"2C",X"00",X"F0",X"40",X"C9",X"03",X"B0",X"3C",X"85",
		X"B9",X"C6",X"B9",X"84",X"16",X"20",X"80",X"69",X"20",X"2F",X"67",X"20",X"48",X"5F",X"20",X"CE",
		X"65",X"20",X"23",X"75",X"A9",X"09",X"20",X"51",X"6A",X"A9",X"12",X"20",X"51",X"6A",X"A9",X"13",
		X"20",X"51",X"6A",X"A9",X"14",X"20",X"51",X"6A",X"A9",X"FF",X"85",X"0F",X"A2",X"00",X"86",X"A5",
		X"86",X"FA",X"A9",X"02",X"85",X"0A",X"A9",X"1A",X"85",X"91",X"60",X"88",X"88",X"88",X"10",X"B6",
		X"20",X"80",X"69",X"A9",X"00",X"85",X"B9",X"A5",X"FC",X"29",X"80",X"85",X"FC",X"A9",X"1C",X"85",
		X"91",X"60",X"82",X"78",X"6E",X"A5",X"F1",X"49",X"FF",X"29",X"18",X"D0",X"E3",X"A5",X"CA",X"29",
		X"0F",X"D0",X"07",X"C6",X"0F",X"D0",X"03",X"4C",X"30",X"76",X"A2",X"00",X"A5",X"94",X"86",X"94",
		X"18",X"65",X"95",X"86",X"95",X"0A",X"0A",X"10",X"02",X"C6",X"A5",X"18",X"65",X"A3",X"85",X"A3",
		X"A9",X"00",X"65",X"A5",X"10",X"05",X"A9",X"1A",X"B8",X"50",X"06",X"C9",X"1B",X"90",X"02",X"A9",
		X"00",X"85",X"A5",X"A4",X"0A",X"B9",X"42",X"76",X"85",X"1D",X"A9",X"B0",X"85",X"1E",X"A5",X"A5",
		X"18",X"69",X"41",X"20",X"BA",X"76",X"A5",X"FA",X"29",X"07",X"F0",X"1D",X"A5",X"A5",X"18",X"69",
		X"41",X"A4",X"16",X"99",X"2C",X"00",X"E6",X"16",X"A9",X"84",X"85",X"0F",X"A2",X"00",X"86",X"FA",
		X"86",X"A5",X"C6",X"0A",X"10",X"03",X"20",X"E4",X"75",X"60",X"84",X"24",X"86",X"23",X"20",X"9D",
		X"69",X"A5",X"1D",X"85",X"00",X"A5",X"1E",X"85",X"01",X"A9",X"00",X"85",X"08",X"A9",X"40",X"85",
		X"0B",X"A9",X"00",X"85",X"0C",X"20",X"27",X"66",X"A5",X"1D",X"18",X"69",X"0A",X"85",X"1D",X"A6",
		X"23",X"A4",X"24",X"60",X"A0",X"15",X"B9",X"2C",X"00",X"F0",X"0F",X"C9",X"03",X"B0",X"0B",X"A9",
		X"5B",X"99",X"2C",X"00",X"99",X"2D",X"00",X"99",X"2E",X"00",X"88",X"88",X"88",X"10",X"E7",X"60",
		X"20",X"80",X"69",X"A9",X"00",X"85",X"B9",X"85",X"93",X"85",X"AE",X"A5",X"FC",X"29",X"80",X"85",
		X"FC",X"20",X"23",X"75",X"A9",X"01",X"20",X"51",X"6A",X"A9",X"C0",X"85",X"20",X"20",X"21",X"69",
		X"20",X"E4",X"76",X"A0",X"15",X"B9",X"46",X"00",X"19",X"45",X"00",X"19",X"44",X"00",X"D0",X"04",
		X"A8",X"B8",X"50",X"3D",X"B9",X"46",X"00",X"85",X"D3",X"B9",X"45",X"00",X"85",X"D2",X"B9",X"44",
		X"00",X"85",X"D1",X"98",X"48",X"A9",X"40",X"A2",X"80",X"A4",X"20",X"20",X"F6",X"6A",X"68",X"A8",
		X"A9",X"50",X"85",X"1D",X"A5",X"20",X"85",X"1E",X"B9",X"2C",X"00",X"20",X"BA",X"76",X"B9",X"2D",
		X"00",X"20",X"BA",X"76",X"B9",X"2E",X"00",X"20",X"BA",X"76",X"A5",X"20",X"38",X"E9",X"0A",X"85",
		X"20",X"88",X"88",X"88",X"10",X"AF",X"20",X"AA",X"74",X"A9",X"14",X"85",X"92",X"A9",X"22",X"85",
		X"91",X"A9",X"FF",X"85",X"AF",X"60",X"20",X"33",X"6C",X"20",X"2F",X"67",X"20",X"86",X"69",X"A9",
		X"01",X"85",X"A7",X"20",X"21",X"69",X"A9",X"0C",X"20",X"51",X"6A",X"A9",X"20",X"85",X"91",X"A5",
		X"66",X"F0",X"04",X"A9",X"14",X"85",X"91",X"60",X"A9",X"FF",X"D0",X"02",X"A9",X"00",X"85",X"98",
		X"A0",X"0C",X"A6",X"97",X"BD",X"5D",X"01",X"18",X"79",X"E2",X"77",X"49",X"FF",X"85",X"07",X"BD",
		X"28",X"01",X"18",X"79",X"D5",X"77",X"85",X"06",X"B9",X"EF",X"77",X"A2",X"00",X"25",X"98",X"81",
		X"06",X"88",X"10",X"DE",X"60",X"00",X"FF",X"00",X"01",X"FE",X"FF",X"00",X"01",X"02",X"FF",X"00",
		X"01",X"00",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FE",X"40",
		X"40",X"80",X"40",X"40",X"80",X"00",X"80",X"40",X"40",X"80",X"40",X"40",X"A2",X"02",X"AD",X"ED",
		X"00",X"E0",X"01",X"F0",X"03",X"B0",X"02",X"0A",X"0A",X"0A",X"B5",X"5C",X"29",X"1F",X"B0",X"37",
		X"F0",X"10",X"C9",X"1B",X"B0",X"0A",X"A8",X"A5",X"FB",X"29",X"07",X"C9",X"07",X"98",X"90",X"02",
		X"E9",X"01",X"95",X"5C",X"AD",X"EE",X"00",X"29",X"20",X"D0",X"04",X"A9",X"F0",X"85",X"5F",X"A5",
		X"5F",X"F0",X"08",X"C6",X"5F",X"A9",X"00",X"95",X"5C",X"95",X"60",X"18",X"B5",X"60",X"F0",X"23",
		X"D6",X"60",X"D0",X"1F",X"38",X"B0",X"1C",X"C9",X"1B",X"B0",X"09",X"B5",X"5C",X"69",X"20",X"90",
		X"D1",X"F0",X"01",X"18",X"A9",X"1F",X"B0",X"CA",X"95",X"5C",X"B5",X"60",X"F0",X"01",X"38",X"A9",
		X"78",X"95",X"60",X"B0",X"03",X"4C",X"A3",X"78",X"A9",X"00",X"E0",X"01",X"90",X"16",X"F0",X"0C",
		X"A5",X"F3",X"29",X"0C",X"4A",X"4A",X"F0",X"0C",X"69",X"02",X"D0",X"08",X"A5",X"F3",X"29",X"10",
		X"F0",X"02",X"A9",X"01",X"38",X"A8",X"65",X"67",X"85",X"67",X"A5",X"F4",X"29",X"04",X"F0",X"11",
		X"98",X"38",X"65",X"68",X"C9",X"04",X"90",X"07",X"38",X"E9",X"04",X"E6",X"66",X"D0",X"F5",X"85",
		X"68",X"F6",X"63",X"CA",X"30",X"03",X"4C",X"FE",X"77",X"A5",X"F3",X"29",X"03",X"A8",X"F0",X"12",
		X"4A",X"69",X"00",X"49",X"FF",X"38",X"65",X"67",X"90",X"0A",X"C0",X"02",X"B0",X"02",X"E6",X"66",
		X"E6",X"66",X"85",X"67",X"A5",X"FB",X"4A",X"B0",X"27",X"A0",X"00",X"A2",X"02",X"B5",X"63",X"F0",
		X"09",X"C9",X"10",X"90",X"05",X"69",X"EF",X"C8",X"95",X"63",X"CA",X"10",X"F0",X"98",X"D0",X"10",
		X"A2",X"02",X"B5",X"63",X"F0",X"07",X"18",X"69",X"EF",X"95",X"63",X"30",X"03",X"CA",X"10",X"F2",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"7D",X"83",X"01",X"07",X"0D",X"13",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"19",X"33",X"00",X"00",X"41",X"47",X"00",X"00",X"00",X"00",X"00",
		X"00",X"5D",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"97",X"9D",X"A3",X"00",X"00",X"00",
		X"00",X"4D",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",
		X"B3",X"00",X"A0",X"10",X"04",X"10",X"00",X"00",X"86",X"40",X"FE",X"04",X"00",X"00",X"C0",X"10",
		X"04",X"10",X"00",X"00",X"86",X"40",X"FE",X"04",X"00",X"00",X"60",X"10",X"00",X"01",X"50",X"10",
		X"F8",X"01",X"48",X"10",X"18",X"01",X"60",X"18",X"F0",X"01",X"60",X"10",X"F8",X"01",X"60",X"10",
		X"08",X"10",X"00",X"00",X"82",X"20",X"02",X"01",X"84",X"10",X"00",X"04",X"84",X"38",X"FF",X"04",
		X"00",X"00",X"10",X"04",X"00",X"01",X"00",X"00",X"2F",X"04",X"0F",X"01",X"00",X"00",X"18",X"18",
		X"00",X"18",X"00",X"00",X"A4",X"18",X"00",X"18",X"A0",X"10",X"00",X"02",X"00",X"00",X"10",X"02",
		X"01",X"20",X"10",X"02",X"01",X"20",X"10",X"02",X"01",X"20",X"10",X"02",X"01",X"20",X"10",X"02",
		X"01",X"20",X"10",X"02",X"01",X"20",X"00",X"00",X"A4",X"02",X"00",X"C0",X"00",X"00",X"20",X"80",
		X"00",X"03",X"00",X"00",X"A3",X"40",X"FD",X"02",X"A3",X"40",X"FD",X"02",X"A3",X"40",X"FD",X"02",
		X"00",X"00",X"40",X"FF",X"02",X"08",X"00",X"00",X"88",X"FF",X"FF",X"08",X"00",X"00",X"C0",X"FF",
		X"02",X"08",X"00",X"00",X"88",X"FF",X"FF",X"08",X"00",X"00",X"18",X"02",X"FF",X"10",X"08",X"20",
		X"00",X"01",X"00",X"00",X"A4",X"10",X"FF",X"04",X"00",X"00",X"A9",X"02",X"2C",X"93",X"00",X"10",
		X"3A",X"8D",X"02",X"00",X"85",X"69",X"8E",X"98",X"00",X"8C",X"99",X"00",X"AA",X"F0",X"08",X"A2",
		X"08",X"0E",X"02",X"00",X"CA",X"90",X"FA",X"8A",X"0A",X"0A",X"0A",X"69",X"07",X"A8",X"C0",X"47",
		X"B0",X"13",X"A2",X"07",X"B9",X"F1",X"78",X"F0",X"08",X"95",X"6A",X"A9",X"01",X"95",X"7A",X"95",
		X"82",X"88",X"CA",X"10",X"EF",X"AE",X"98",X"00",X"AC",X"99",X"00",X"60",X"A9",X"18",X"A0",X"AF",
		X"8D",X"00",X"40",X"8C",X"01",X"40",X"60",X"AD",X"E0",X"00",X"D0",X"F0",X"A2",X"07",X"D6",X"7A",
		X"D0",X"56",X"B4",X"6A",X"F0",X"52",X"D6",X"82",X"D0",X"30",X"B9",X"31",X"79",X"95",X"72",X"B9",
		X"32",X"79",X"95",X"7A",X"D0",X"15",X"95",X"6A",X"8A",X"D0",X"3D",X"A9",X"00",X"95",X"72",X"9D",
		X"00",X"40",X"A9",X"00",X"95",X"6A",X"CA",X"10",X"D5",X"30",X"35",X"B9",X"34",X"79",X"95",X"82",
		X"B5",X"6A",X"18",X"69",X"04",X"95",X"6A",X"4C",X"98",X"7A",X"B9",X"2E",X"79",X"95",X"7A",X"B5",
		X"72",X"18",X"79",X"2F",X"79",X"24",X"69",X"50",X"0D",X"E0",X"01",X"F0",X"09",X"AD",X"0A",X"40",
		X"29",X"1E",X"D0",X"02",X"A9",X"1E",X"95",X"72",X"B5",X"72",X"9D",X"00",X"40",X"CA",X"10",X"9E",
		X"A5",X"70",X"D0",X"26",X"A5",X"8A",X"F0",X"22",X"2A",X"2A",X"2A",X"29",X"03",X"AA",X"A5",X"8B",
		X"DD",X"CA",X"7A",X"D0",X"06",X"BD",X"CD",X"7A",X"B8",X"50",X"03",X"38",X"E9",X"02",X"8D",X"06",
		X"40",X"85",X"8B",X"A9",X"A4",X"8D",X"07",X"40",X"85",X"79",X"60",X"30",X"00",X"00",X"70",X"30",
		X"30",X"A9",X"30",X"85",X"8B",X"A5",X"8A",X"09",X"80",X"85",X"8A",X"60",X"A5",X"8A",X"09",X"40",
		X"85",X"8A",X"30",X"04",X"A9",X"70",X"85",X"8B",X"60",X"AD",X"DA",X"00",X"D0",X"1D",X"A5",X"8A",
		X"29",X"7F",X"85",X"8A",X"24",X"8A",X"70",X"E4",X"A5",X"8A",X"29",X"BF",X"85",X"8A",X"AD",X"DA",
		X"00",X"D0",X"08",X"85",X"8A",X"8D",X"06",X"40",X"8D",X"07",X"40",X"60",X"A9",X"00",X"8D",X"0F",
		X"40",X"A9",X"03",X"8D",X"0F",X"40",X"A2",X"07",X"A9",X"00",X"9D",X"00",X"40",X"95",X"6A",X"95",
		X"72",X"CA",X"10",X"F6",X"A9",X"20",X"8D",X"08",X"40",X"60",X"48",X"8A",X"48",X"98",X"48",X"D8",
		X"BA",X"E0",X"E0",X"90",X"16",X"BD",X"04",X"01",X"29",X"10",X"D0",X"0F",X"BD",X"06",X"01",X"C9",
		X"50",X"90",X"08",X"C9",X"80",X"B0",X"04",X"A5",X"9F",X"10",X"1F",X"A2",X"FF",X"9A",X"D8",X"E8",
		X"8A",X"78",X"95",X"00",X"9D",X"00",X"01",X"CA",X"D0",X"F8",X"A9",X"40",X"8D",X"00",X"48",X"2C",
		X"00",X"49",X"50",X"03",X"4C",X"01",X"50",X"4C",X"82",X"7C",X"8D",X"00",X"4C",X"E6",X"FB",X"AD",
		X"00",X"49",X"10",X"34",X"E6",X"9F",X"A5",X"D8",X"F0",X"02",X"C6",X"D8",X"A5",X"EC",X"85",X"F3",
		X"A2",X"07",X"06",X"F3",X"90",X"02",X"F6",X"E4",X"B5",X"E4",X"9D",X"00",X"4B",X"CA",X"10",X"F2",
		X"AD",X"00",X"4A",X"49",X"02",X"85",X"F3",X"A5",X"F5",X"29",X"BF",X"A8",X"A5",X"FC",X"29",X"3E",
		X"D0",X"04",X"98",X"09",X"40",X"A8",X"84",X"F5",X"AE",X"00",X"49",X"86",X"EE",X"A5",X"F5",X"29",
		X"FE",X"A8",X"AE",X"00",X"48",X"86",X"F6",X"8C",X"00",X"48",X"AE",X"00",X"48",X"86",X"ED",X"09",
		X"01",X"8D",X"00",X"48",X"AE",X"00",X"48",X"86",X"F8",X"A5",X"F6",X"38",X"E5",X"F7",X"29",X"0F",
		X"C9",X"08",X"90",X"02",X"09",X"F0",X"18",X"65",X"94",X"85",X"94",X"A5",X"F6",X"38",X"09",X"0F",
		X"E5",X"F7",X"4A",X"4A",X"4A",X"4A",X"C9",X"08",X"90",X"02",X"09",X"F0",X"18",X"65",X"95",X"85",
		X"95",X"A5",X"F8",X"85",X"F7",X"A9",X"07",X"8D",X"0F",X"40",X"8D",X"0B",X"40",X"AD",X"08",X"40",
		X"49",X"7F",X"85",X"F4",X"24",X"F2",X"50",X"06",X"20",X"37",X"7A",X"20",X"FC",X"77",X"A2",X"01",
		X"B4",X"ED",X"B5",X"EF",X"94",X"EF",X"A8",X"35",X"EF",X"15",X"F1",X"95",X"F1",X"98",X"15",X"EF",
		X"35",X"F1",X"95",X"F1",X"CA",X"10",X"E9",X"A4",X"F2",X"A5",X"FC",X"29",X"3E",X"F0",X"02",X"A4",
		X"F1",X"98",X"49",X"FF",X"25",X"F9",X"45",X"FA",X"85",X"FA",X"84",X"F9",X"A5",X"F5",X"29",X"40",
		X"09",X"06",X"A6",X"AE",X"E8",X"A4",X"93",X"D0",X"10",X"A2",X"00",X"A4",X"FB",X"C0",X"40",X"90",
		X"08",X"A6",X"66",X"E0",X"02",X"90",X"02",X"A2",X"03",X"3D",X"7E",X"7C",X"A4",X"63",X"10",X"02",
		X"09",X"20",X"A4",X"64",X"10",X"02",X"09",X"10",X"A4",X"65",X"10",X"02",X"09",X"08",X"85",X"F5",
		X"2C",X"00",X"49",X"30",X"FB",X"8D",X"00",X"4D",X"68",X"A8",X"68",X"AA",X"68",X"40",X"FF",X"FD",
		X"FB",X"F9",X"A9",X"00",X"8D",X"0F",X"40",X"8D",X"05",X"40",X"8D",X"07",X"40",X"8D",X"08",X"40",
		X"A9",X"03",X"8D",X"0F",X"40",X"A9",X"08",X"8D",X"03",X"40",X"A9",X"C0",X"8D",X"02",X"40",X"A9",
		X"44",X"8D",X"00",X"48",X"A0",X"60",X"2C",X"00",X"49",X"30",X"FB",X"2C",X"00",X"49",X"10",X"FB",
		X"8D",X"00",X"4C",X"88",X"10",X"F0",X"A9",X"A2",X"8D",X"03",X"40",X"A0",X"00",X"A2",X"00",X"94",
		X"00",X"C8",X"98",X"9D",X"00",X"01",X"E8",X"D0",X"F6",X"8D",X"00",X"4C",X"98",X"55",X"00",X"95",
		X"00",X"D0",X"1D",X"C8",X"98",X"5D",X"00",X"01",X"9D",X"00",X"01",X"D0",X"13",X"E8",X"D0",X"EC",
		X"C8",X"D0",X"DA",X"A9",X"40",X"8D",X"02",X"40",X"A9",X"42",X"8D",X"00",X"48",X"4C",X"39",X"7D",
		X"A2",X"07",X"A0",X"00",X"8C",X"03",X"40",X"9A",X"BA",X"2A",X"A0",X"A0",X"90",X"02",X"A0",X"10",
		X"8C",X"00",X"40",X"A0",X"A8",X"8C",X"01",X"40",X"A0",X"20",X"2C",X"00",X"49",X"30",X"FB",X"2C",
		X"00",X"49",X"10",X"FB",X"8D",X"00",X"4C",X"88",X"10",X"F0",X"A0",X"00",X"8C",X"01",X"40",X"A0",
		X"14",X"2C",X"00",X"49",X"30",X"FB",X"2C",X"00",X"49",X"10",X"FB",X"8D",X"00",X"4C",X"88",X"10",
		X"F0",X"BA",X"CA",X"9A",X"10",X"C2",X"4C",X"4B",X"7B",X"A2",X"00",X"86",X"06",X"86",X"8D",X"9A",
		X"A9",X"50",X"85",X"07",X"A2",X"2F",X"A9",X"12",X"85",X"99",X"A0",X"00",X"8E",X"00",X"4C",X"51",
		X"06",X"C8",X"D0",X"FB",X"A8",X"8A",X"29",X"07",X"C9",X"01",X"98",X"B0",X"18",X"F0",X"10",X"48",
		X"8A",X"48",X"4A",X"4A",X"4A",X"AA",X"BD",X"F9",X"60",X"05",X"8D",X"85",X"8D",X"68",X"AA",X"A5",
		X"99",X"69",X"22",X"85",X"99",X"E6",X"07",X"CA",X"10",X"D0",X"58",X"20",X"86",X"69",X"20",X"2F",
		X"67",X"A9",X"00",X"85",X"EA",X"A9",X"0E",X"85",X"E4",X"85",X"93",X"A9",X"22",X"BA",X"D0",X"02",
		X"A9",X"20",X"A2",X"FF",X"9A",X"20",X"3B",X"7F",X"A9",X"80",X"85",X"00",X"85",X"01",X"A2",X"00",
		X"A9",X"C0",X"81",X"00",X"A0",X"24",X"AD",X"20",X"20",X"29",X"11",X"C9",X"11",X"F0",X"02",X"A0",
		X"23",X"98",X"20",X"51",X"6A",X"AD",X"0A",X"40",X"85",X"FD",X"A0",X"10",X"AD",X"0A",X"40",X"C5",
		X"FD",X"D0",X"0A",X"85",X"FD",X"88",X"10",X"F4",X"A9",X"27",X"20",X"51",X"6A",X"A9",X"1F",X"20",
		X"51",X"6A",X"A9",X"02",X"85",X"AE",X"A9",X"00",X"85",X"B9",X"20",X"5C",X"65",X"A5",X"F3",X"49",
		X"FF",X"85",X"FD",X"A9",X"01",X"85",X"FF",X"8D",X"08",X"40",X"46",X"9F",X"90",X"FC",X"A5",X"F2",
		X"29",X"24",X"D0",X"05",X"85",X"FF",X"20",X"7F",X"7F",X"A5",X"F2",X"29",X"21",X"D0",X"05",X"85",
		X"FF",X"20",X"62",X"7F",X"A9",X"00",X"8D",X"01",X"40",X"8D",X"03",X"40",X"A5",X"F2",X"29",X"22",
		X"D0",X"05",X"85",X"FF",X"20",X"EB",X"7E",X"20",X"32",X"51",X"A5",X"F1",X"49",X"FF",X"8D",X"00",
		X"40",X"F0",X"07",X"A9",X"A8",X"8D",X"01",X"40",X"E6",X"E4",X"A5",X"F2",X"49",X"FF",X"29",X"27",
		X"8D",X"02",X"40",X"F0",X"07",X"A9",X"A8",X"8D",X"03",X"40",X"E6",X"E4",X"A5",X"FA",X"29",X"07",
		X"F0",X"17",X"A5",X"B9",X"49",X"01",X"85",X"B9",X"A9",X"00",X"85",X"FA",X"20",X"86",X"69",X"A5",
		X"FD",X"49",X"FF",X"85",X"FD",X"A9",X"01",X"85",X"FF",X"20",X"6B",X"7E",X"24",X"F2",X"50",X"8A",
		X"4C",X"4B",X"7B",X"11",X"14",X"15",X"16",X"21",X"24",X"25",X"26",X"A5",X"FF",X"F0",X"7B",X"A5",
		X"F3",X"C5",X"FD",X"85",X"FD",X"D0",X"06",X"A5",X"F4",X"C5",X"FE",X"85",X"FE",X"F0",X"6B",X"A9",
		X"25",X"20",X"49",X"6A",X"A9",X"1B",X"20",X"49",X"6A",X"20",X"2F",X"67",X"A5",X"F3",X"29",X"03",
		X"AA",X"BD",X"2F",X"6C",X"20",X"51",X"6A",X"A5",X"F3",X"29",X"1C",X"4A",X"4A",X"AA",X"BD",X"63",
		X"7E",X"48",X"4A",X"4A",X"4A",X"4A",X"A2",X"40",X"A0",X"28",X"20",X"9D",X"6A",X"68",X"29",X"07",
		X"A2",X"50",X"20",X"9D",X"6A",X"A9",X"70",X"85",X"1D",X"A9",X"28",X"85",X"1E",X"A5",X"F4",X"29",
		X"08",X"F0",X"02",X"A9",X"46",X"20",X"BA",X"76",X"A5",X"F4",X"29",X"04",X"F0",X"02",X"A9",X"58",
		X"20",X"BA",X"76",X"A5",X"F4",X"29",X"03",X"AA",X"BD",X"08",X"5B",X"A2",X"40",X"A0",X"34",X"20",
		X"9D",X"6A",X"A9",X"26",X"20",X"51",X"6A",X"20",X"AA",X"74",X"60",X"20",X"62",X"7F",X"20",X"86",
		X"69",X"78",X"A9",X"00",X"85",X"8D",X"A9",X"1F",X"85",X"99",X"A9",X"02",X"85",X"07",X"A9",X"AA",
		X"91",X"06",X"C8",X"B1",X"06",X"F0",X"03",X"20",X"32",X"7F",X"C8",X"D0",X"F6",X"B1",X"06",X"C9",
		X"AA",X"F0",X"03",X"20",X"30",X"7F",X"A9",X"00",X"91",X"06",X"85",X"9F",X"8D",X"00",X"4C",X"E6",
		X"06",X"D0",X"DB",X"E6",X"07",X"A5",X"07",X"C9",X"3F",X"D0",X"D3",X"A5",X"99",X"4C",X"3B",X"7F",
		X"49",X"AA",X"05",X"8D",X"85",X"8D",X"A9",X"21",X"85",X"99",X"60",X"58",X"20",X"51",X"6A",X"A5",
		X"8D",X"A2",X"08",X"0A",X"90",X"18",X"48",X"86",X"C5",X"A9",X"E0",X"85",X"0B",X"8A",X"0A",X"0A",
		X"0A",X"18",X"69",X"88",X"A8",X"8A",X"A2",X"A0",X"20",X"9D",X"6A",X"A6",X"C5",X"68",X"CA",X"D0",
		X"E2",X"60",X"A2",X"07",X"8A",X"0A",X"95",X"E4",X"CA",X"10",X"F9",X"E8",X"86",X"06",X"A0",X"18",
		X"84",X"07",X"A5",X"06",X"81",X"06",X"E6",X"07",X"D0",X"F8",X"E6",X"06",X"D0",X"F0",X"60",X"A9",
		X"0E",X"A2",X"07",X"95",X"E4",X"CA",X"10",X"FB",X"A9",X"00",X"85",X"E6",X"20",X"86",X"69",X"A2",
		X"00",X"A0",X"05",X"A9",X"19",X"85",X"07",X"B9",X"E2",X"7F",X"85",X"06",X"A9",X"40",X"81",X"06",
		X"E6",X"07",X"D0",X"FA",X"88",X"10",X"EC",X"A0",X"05",X"B9",X"E8",X"7F",X"85",X"07",X"86",X"06",
		X"A9",X"40",X"81",X"06",X"E6",X"06",X"D0",X"FA",X"88",X"10",X"EE",X"A0",X"04",X"B9",X"E2",X"7F",
		X"18",X"79",X"E3",X"7F",X"6A",X"85",X"06",X"84",X"98",X"A0",X"04",X"B9",X"E8",X"7F",X"18",X"79",
		X"E9",X"7F",X"6A",X"85",X"07",X"A9",X"40",X"81",X"06",X"88",X"10",X"EF",X"A4",X"98",X"88",X"10",
		X"DC",X"60",X"00",X"33",X"66",X"99",X"CC",X"FF",X"19",X"46",X"74",X"A2",X"D0",X"FF",X"D8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"7B",X"4B",X"7B",X"2A",X"7B");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
