library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(3 downto 0)
);
end entity;

architecture prom of snd is
	type rom is array(0 to  1023) of std_logic_vector(3 downto 0);
	signal rom_data: rom := (
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",X"F",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",
		X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",
		X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",
		X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",
		X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",
		X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"2",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",
		X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3",X"3");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
