library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity k3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of k3 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"EE",X"EE",X"EE",X"0E",X"EE",X"EE",
		X"EE",X"E0",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"0E",X"EE",X"EE",
		X"0E",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"22",X"3B",X"1F",X"09",X"1E",X"00",X"00",X"08",X"50",X"70",X"E0",X"78",X"30",
		X"06",X"0D",X"1F",X"32",X"04",X"00",X"00",X"00",X"60",X"F0",X"B8",X"E8",X"44",X"00",X"00",X"00",
		X"40",X"70",X"3B",X"1F",X"1D",X"0B",X"0E",X"7C",X"00",X"02",X"4E",X"FC",X"C8",X"7C",X"38",X"30",
		X"0E",X"1F",X"1D",X"0B",X"1F",X"32",X"60",X"00",X"78",X"38",X"EC",X"F8",X"6C",X"66",X"02",X"00",
		X"8E",X"64",X"79",X"3F",X"97",X"9D",X"38",X"75",X"53",X"86",X"8C",X"DD",X"FD",X"69",X"10",X"BF",
		X"FC",X"19",X"DF",X"BB",X"7F",X"64",X"C0",X"9C",X"B8",X"3C",X"5E",X"F0",X"F9",X"DC",X"B6",X"B3",
		X"00",X"00",X"04",X"04",X"08",X"10",X"A0",X"C0",X"00",X"00",X"00",X"08",X"02",X"78",X"FE",X"D6",
		X"00",X"00",X"28",X"38",X"24",X"00",X"1C",X"7F",X"00",X"00",X"20",X"30",X"18",X"09",X"0D",X"03",
		X"00",X"08",X"E4",X"F0",X"B0",X"60",X"E0",X"C0",X"AB",X"FD",X"FE",X"7F",X"77",X"2F",X"4F",X"E3",
		X"67",X"DB",X"FE",X"FE",X"FD",X"6D",X"F1",X"D7",X"04",X"04",X"09",X"11",X"01",X"07",X"0F",X"1B",
		X"B0",X"F4",X"66",X"B4",X"B6",X"61",X"C0",X"80",X"CF",X"AF",X"17",X"A7",X"F3",X"DF",X"FF",X"E7",
		X"7B",X"F6",X"E8",X"E6",X"FE",X"B6",X"6D",X"FF",X"1D",X"1B",X"0D",X"1E",X"1D",X"0F",X"03",X"00",
		X"30",X"40",X"A0",X"90",X"48",X"04",X"00",X"00",X"FA",X"BC",X"7C",X"F8",X"E2",X"04",X"00",X"00",
		X"6F",X"36",X"39",X"1F",X"4E",X"20",X"20",X"00",X"04",X"02",X"0D",X"09",X"10",X"20",X"20",X"00",
		X"00",X"02",X"0C",X"98",X"C8",X"C0",X"58",X"FC",X"00",X"1E",X"7F",X"73",X"6D",X"FE",X"FF",X"FF",
		X"00",X"00",X"0F",X"DE",X"F7",X"DF",X"FF",X"FF",X"80",X"C4",X"62",X"30",X"19",X"13",X"03",X"0F",
		X"FE",X"EE",X"F6",X"F7",X"EF",X"DE",X"F8",X"FF",X"FF",X"EF",X"CB",X"17",X"2F",X"5D",X"8B",X"EF",
		X"BF",X"7D",X"DC",X"C5",X"D3",X"ED",X"E1",X"83",X"0F",X"06",X"19",X"3F",X"3D",X"1B",X"1B",X"5D",
		X"FF",X"7F",X"EF",X"F7",X"FA",X"F7",X"FB",X"F7",X"87",X"D8",X"2F",X"0F",X"67",X"FB",X"FF",X"B7",
		X"E7",X"AD",X"61",X"C1",X"9C",X"FD",X"FF",X"BF",X"7F",X"EF",X"FF",X"FB",X"FF",X"6F",X"07",X"0D",
		X"EF",X"DE",X"3C",X"F0",X"84",X"94",X"0A",X"01",X"CF",X"FE",X"FF",X"7F",X"B5",X"CB",X"FF",X"74",
		X"3F",X"FF",X"DE",X"9F",X"83",X"3D",X"48",X"50",X"0E",X"0F",X"0F",X"27",X"13",X"28",X"48",X"80",
		X"00",X"03",X"03",X"01",X"01",X"01",X"73",X"77",X"00",X"80",X"80",X"00",X"00",X"00",X"9C",X"DC",
		X"7F",X"7F",X"7F",X"7F",X"77",X"70",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"DC",X"1C",X"00",X"00",
		X"00",X"70",X"77",X"7F",X"7F",X"7F",X"7F",X"77",X"00",X"1C",X"DC",X"FC",X"FC",X"FC",X"FC",X"DC",
		X"73",X"01",X"01",X"01",X"03",X"03",X"00",X"00",X"9C",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"7F",X"7F",X"7F",X"1E",X"3F",X"3F",X"3F",X"00",X"80",X"80",X"80",X"00",X"00",X"8C",X"FC",
		X"3F",X"3F",X"1E",X"7F",X"7F",X"7F",X"00",X"00",X"8C",X"00",X"00",X"80",X"80",X"80",X"00",X"00",
		X"00",X"03",X"03",X"03",X"00",X"01",X"63",X"7F",X"00",X"FC",X"FC",X"FC",X"F0",X"F8",X"F8",X"F8",
		X"63",X"01",X"00",X"03",X"03",X"03",X"00",X"00",X"F8",X"F8",X"F0",X"FC",X"FC",X"FC",X"00",X"00",
		X"00",X"03",X"03",X"01",X"71",X"77",X"7C",X"78",X"00",X"80",X"80",X"00",X"1C",X"DC",X"7C",X"3C",
		X"78",X"7C",X"76",X"73",X"71",X"70",X"00",X"00",X"3C",X"7C",X"DC",X"9C",X"1C",X"1C",X"00",X"00",
		X"00",X"70",X"71",X"73",X"76",X"7C",X"78",X"78",X"00",X"1C",X"1C",X"9C",X"DC",X"7C",X"3C",X"3C",
		X"7C",X"77",X"71",X"01",X"03",X"03",X"00",X"00",X"7C",X"DC",X"1C",X"00",X"80",X"80",X"00",X"00",
		X"00",X"7F",X"7F",X"7F",X"07",X"0C",X"18",X"30",X"00",X"E0",X"E0",X"E0",X"80",X"C0",X"4C",X"7C",
		X"18",X"0C",X"07",X"7F",X"7F",X"7F",X"00",X"00",X"4C",X"C0",X"80",X"E0",X"E0",X"E0",X"00",X"00",
		X"00",X"0F",X"0F",X"0F",X"03",X"06",X"64",X"7C",X"00",X"FC",X"FC",X"FC",X"C0",X"60",X"30",X"18",
		X"64",X"06",X"03",X"0F",X"0F",X"0F",X"00",X"00",X"30",X"60",X"C0",X"FC",X"FC",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"7C",X"82",X"82",X"82",X"7C",X"00",X"8C",X"D2",X"A2",X"82",X"84",X"00",X"00",
		X"00",X"00",X"00",X"7C",X"82",X"82",X"82",X"7C",X"00",X"0C",X"92",X"92",X"52",X"3C",X"00",X"00",
		X"00",X"7C",X"82",X"82",X"7C",X"00",X"9C",X"A2",X"A2",X"A2",X"E4",X"00",X"02",X"FE",X"42",X"00",
		X"00",X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"8C",X"D2",X"A2",X"82",X"84",
		X"00",X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"6C",X"92",X"92",X"92",X"6C",
		X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"9C",X"92",X"92",X"7C",X"00",X"FE",
		X"00",X"00",X"01",X"03",X"03",X"03",X"07",X"0F",X"00",X"60",X"F8",X"80",X"E0",X"C0",X"C0",X"E0",
		X"1F",X"0F",X"37",X"19",X"06",X"03",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"20",X"80",X"FF",X"00",
		X"00",X"00",X"21",X"41",X"45",X"4B",X"31",X"00",X"3E",X"41",X"41",X"41",X"3E",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"4A",X"49",X"49",X"30",X"00",X"3E",X"41",X"41",X"41",X"3E",X"00",X"00",X"00",
		X"00",X"42",X"7F",X"40",X"00",X"27",X"45",X"45",X"45",X"39",X"00",X"3E",X"41",X"41",X"3E",X"00",
		X"21",X"41",X"45",X"4B",X"31",X"00",X"3E",X"41",X"41",X"3E",X"00",X"3E",X"41",X"41",X"3E",X"00",
		X"36",X"49",X"49",X"49",X"36",X"00",X"3E",X"41",X"41",X"3E",X"00",X"3E",X"41",X"41",X"3E",X"00",
		X"7F",X"00",X"3E",X"49",X"49",X"39",X"00",X"3E",X"41",X"41",X"3E",X"00",X"3E",X"41",X"41",X"3E",
		X"00",X"FF",X"01",X"04",X"07",X"0F",X"0F",X"1F",X"00",X"00",X"C0",X"60",X"98",X"EC",X"F0",X"F8",
		X"07",X"03",X"03",X"07",X"01",X"1F",X"06",X"00",X"F0",X"E0",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"54",X"7D",X"3F",X"1D",X"06",X"07",X"13",X"2F",X"00",X"00",X"C0",X"E0",X"E6",X"E6",X"4C",X"FE",
		X"3F",X"23",X"07",X"06",X"1D",X"3F",X"7D",X"54",X"FE",X"4C",X"E6",X"E6",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",
		X"31",X"21",X"2C",X"2E",X"6E",X"60",X"60",X"7F",X"B0",X"30",X"30",X"70",X"F8",X"38",X"38",X"F8",
		X"00",X"00",X"03",X"07",X"67",X"67",X"32",X"7F",X"2A",X"BE",X"FC",X"B8",X"60",X"E0",X"C4",X"FC",
		X"7F",X"32",X"67",X"67",X"07",X"03",X"00",X"00",X"F4",X"C8",X"E0",X"60",X"B8",X"FC",X"BE",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",
		X"1F",X"1C",X"1C",X"1F",X"0E",X"0C",X"0C",X"0C",X"FE",X"06",X"06",X"76",X"74",X"34",X"84",X"8C",
		X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"60",X"F0",X"DA",X"CA",X"CA",X"E0",X"60",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"00",X"00",
		X"DB",X"DB",X"DF",X"1F",X"00",X"00",X"7F",X"FF",X"FF",X"00",X"00",X"7F",X"FF",X"FF",X"DB",X"DB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"E0",X"FA",X"FA",X"00",X"00",X"00",
		X"60",X"F0",X"9A",X"8A",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"1F",X"4A",X"7A",X"4A",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",X"00",X"00",X"40",X"42",X"7F",X"7F",X"40",X"40",
		X"00",X"62",X"73",X"79",X"59",X"5D",X"4F",X"46",X"00",X"20",X"61",X"49",X"4D",X"4F",X"7B",X"31",
		X"00",X"18",X"1C",X"16",X"13",X"7F",X"7F",X"10",X"00",X"27",X"67",X"45",X"45",X"45",X"7D",X"38",
		X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",X"00",X"03",X"03",X"71",X"79",X"0D",X"07",X"03",
		X"00",X"36",X"4F",X"4D",X"59",X"59",X"76",X"30",X"00",X"06",X"4F",X"49",X"49",X"69",X"3F",X"1E",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"FF",X"C3",X"C3",X"C3",X"FF",X"7E",X"00",X"00",X"7F",
		X"C3",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"C3",X"00",X"00",X"7E",X"FF",X"C3",X"C3",X"C3",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7E",X"13",X"11",X"13",X"7E",X"7C",
		X"00",X"7F",X"7F",X"49",X"49",X"49",X"7F",X"36",X"00",X"1C",X"3E",X"63",X"41",X"41",X"63",X"22",
		X"00",X"7F",X"7F",X"41",X"41",X"63",X"3E",X"1C",X"00",X"00",X"7F",X"7F",X"49",X"49",X"49",X"41",
		X"00",X"7F",X"7F",X"09",X"09",X"09",X"09",X"01",X"00",X"1C",X"3E",X"63",X"41",X"49",X"79",X"79",
		X"00",X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"41",X"7F",X"7F",X"41",X"41",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"00",X"00",X"7F",X"7F",X"40",X"40",X"40",X"40",X"00",X"7F",X"7F",X"0E",X"1C",X"0E",X"7F",X"7F",
		X"00",X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",
		X"00",X"7F",X"7F",X"11",X"11",X"11",X"1F",X"0E",X"00",X"3E",X"7F",X"41",X"51",X"71",X"3F",X"5E",
		X"00",X"7F",X"7F",X"11",X"31",X"79",X"6F",X"4E",X"00",X"26",X"6F",X"49",X"49",X"4B",X"7A",X"30",
		X"00",X"00",X"01",X"01",X"7F",X"7F",X"01",X"01",X"00",X"3F",X"7F",X"40",X"40",X"40",X"7F",X"3F",
		X"00",X"0F",X"1F",X"38",X"70",X"38",X"1F",X"0F",X"00",X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",
		X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"00",X"07",X"0F",X"78",X"78",X"0F",X"07",
		X"00",X"61",X"71",X"79",X"5D",X"4F",X"47",X"43",X"00",X"00",X"00",X"5F",X"5F",X"07",X"00",X"00",
		X"00",X"00",X"02",X"03",X"51",X"59",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"52",X"5E",X"52",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
