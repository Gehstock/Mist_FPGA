library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"70",X"F8",X"8D",X"85",X"C0",X"60",X"00",
		X"8E",X"4A",X"2E",X"10",X"E8",X"A4",X"E2",X"00",X"18",X"3C",X"7E",X"FF",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"06",X"06",X"06",X"0E",X"0C",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"BF",X"C3",X"C3",X"BF",X"81",X"81",X"FC",X"C6",X"81",X"81",X"81",X"81",X"C6",X"FC",
		X"81",X"81",X"9D",X"BD",X"BD",X"9D",X"81",X"81",X"18",X"60",X"80",X"03",X"0C",X"10",X"0C",X"03",
		X"06",X"00",X"18",X"00",X"18",X"00",X"03",X"07",X"60",X"00",X"18",X"00",X"18",X"00",X"C0",X"E0",
		X"07",X"07",X"03",X"18",X"00",X"18",X"00",X"00",X"E0",X"E0",X"C0",X"18",X"00",X"18",X"00",X"00",
		X"06",X"00",X"00",X"18",X"00",X"00",X"03",X"07",X"70",X"00",X"00",X"18",X"00",X"00",X"C0",X"E0",
		X"07",X"07",X"03",X"00",X"18",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"14",X"40",X"41",X"01",X"00",X"00",X"00",X"0A",X"0A",X"E0",X"F0",X"F0",
		X"01",X"41",X"40",X"14",X"14",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"0A",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"40",X"41",X"01",X"00",X"00",X"00",X"04",X"04",X"E0",X"F0",X"F0",
		X"01",X"41",X"40",X"08",X"08",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"04",X"04",X"00",X"00",X"00",
		X"22",X"2E",X"2C",X"2F",X"20",X"20",X"20",X"20",X"60",X"7F",X"00",X"F8",X"0F",X"0F",X"0E",X"0E",
		X"20",X"20",X"20",X"20",X"30",X"1F",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"00",X"FF",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"FC",X"00",X"00",X"02",X"FE",X"FE",X"86",X"86",X"FE",X"FE",X"02",
		X"00",X"1F",X"20",X"20",X"27",X"27",X"27",X"27",X"00",X"FF",X"00",X"00",X"00",X"42",X"7E",X"3C",
		X"00",X"FC",X"02",X"FA",X"8A",X"8A",X"FA",X"02",X"00",X"7E",X"7E",X"06",X"04",X"04",X"04",X"00",
		X"20",X"26",X"26",X"20",X"20",X"1F",X"00",X"00",X"3E",X"3E",X"3E",X"30",X"00",X"FF",X"00",X"00",
		X"00",X"24",X"66",X"FF",X"FF",X"66",X"24",X"00",X"18",X"3C",X"7E",X"18",X"18",X"7E",X"3C",X"18",
		X"1F",X"3F",X"60",X"C0",X"C0",X"60",X"3F",X"1F",X"8C",X"92",X"FF",X"92",X"92",X"FF",X"92",X"62",
		X"20",X"22",X"22",X"2E",X"2E",X"22",X"22",X"20",X"00",X"1F",X"20",X"20",X"27",X"26",X"26",X"24",
		X"00",X"FF",X"00",X"00",X"3C",X"3C",X"3C",X"00",X"F2",X"F2",X"C2",X"02",X"02",X"FC",X"00",X"00",
		X"02",X"FA",X"8A",X"02",X"02",X"FA",X"FA",X"02",X"00",X"FC",X"02",X"02",X"F2",X"72",X"72",X"32",
		X"26",X"3F",X"3F",X"26",X"26",X"1F",X"00",X"00",X"20",X"27",X"27",X"27",X"27",X"27",X"27",X"20",
		X"00",X"1F",X"20",X"20",X"26",X"26",X"26",X"20",X"7F",X"41",X"7F",X"7F",X"00",X"FF",X"00",X"00",
		X"00",X"7F",X"7F",X"41",X"67",X"67",X"7F",X"00",X"00",X"FF",X"00",X"7F",X"41",X"41",X"41",X"7F",
		X"02",X"52",X"52",X"02",X"02",X"FC",X"00",X"00",X"02",X"62",X"62",X"62",X"7A",X"5A",X"7A",X"02",
		X"00",X"FC",X"02",X"C2",X"82",X"82",X"8A",X"9A",X"2C",X"2C",X"34",X"34",X"2C",X"2C",X"34",X"34",
		X"04",X"3F",X"11",X"0F",X"04",X"03",X"01",X"00",X"04",X"3F",X"11",X"3F",X"04",X"3F",X"22",X"3F",
		X"00",X"01",X"03",X"07",X"0C",X"1F",X"31",X"3F",X"DD",X"55",X"77",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"7D",X"47",X"45",X"C5",X"45",X"7F",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"77",X"55",
		X"DD",X"55",X"00",X"FF",X"FF",X"00",X"77",X"55",X"DC",X"54",X"76",X"14",X"0C",X"04",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"52",X"52",X"52",X"7E",X"7E",X"00",X"00",X"00",
		X"44",X"24",X"1E",X"0E",X"00",X"00",X"2C",X"52",X"30",X"7E",X"7E",X"00",X"00",X"0E",X"1E",X"24",
		X"7E",X"7E",X"00",X"00",X"7E",X"7E",X"0C",X"18",X"00",X"00",X"00",X"02",X"46",X"6C",X"38",X"18",
		X"00",X"00",X"04",X"0E",X"16",X"54",X"74",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"3C",X"18",X"7E",X"7E",X"00",X"00",X"00",X"18",X"30",X"7E",X"7E",X"00",X"00",X"42",X"66",
		X"42",X"3C",X"18",X"00",X"00",X"7E",X"7E",X"0C",X"66",X"42",X"00",X"00",X"18",X"3C",X"42",X"42",
		X"00",X"00",X"00",X"42",X"66",X"3C",X"18",X"3C",X"C3",X"C3",X"C3",X"C3",X"FC",X"FC",X"FC",X"FC",
		X"C3",X"C3",X"C3",X"C3",X"3F",X"3F",X"FF",X"FF",X"C3",X"C3",X"C3",X"C3",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"80",
		X"01",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"03",X"07",X"0F",X"1C",X"3C",X"7F",X"FF",X"C3",X"C3",X"C3",X"C3",X"3C",X"3C",X"FF",X"FF",
		X"C3",X"C3",X"C3",X"C3",X"FC",X"FC",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"F8",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",X"F8",X"FC",X"FC",X"FC",X"FC",X"7C",X"3C",
		X"00",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"14",X"14",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"14",X"14",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"14",X"14",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"14",X"14",X"00",X"00",
		X"0F",X"3F",X"0F",X"3F",X"0F",X"0F",X"0F",X"0F",X"F0",X"FC",X"F0",X"FC",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"3F",X"0F",X"3F",X"0F",X"0F",X"00",X"00",X"F0",X"FC",X"F0",X"FC",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"0A",X"0A",X"3F",X"E2",X"F6",X"F6",X"00",X"00",X"0A",X"0A",X"FF",X"D1",X"DB",X"5B",
		X"F6",X"F6",X"F6",X"3F",X"0A",X"0A",X"00",X"00",X"1B",X"9B",X"DB",X"FF",X"0A",X"0A",X"00",X"00",
		X"0F",X"0B",X"38",X"0B",X"3F",X"08",X"0F",X"0E",X"F0",X"F0",X"1C",X"F0",X"FC",X"10",X"70",X"F0",
		X"08",X"0F",X"3B",X"08",X"3B",X"0F",X"07",X"07",X"10",X"F0",X"FC",X"10",X"FC",X"F0",X"E0",X"E0",
		X"00",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"1F",X"20",X"2F",X"2F",X"3F",X"1F",X"00",X"0F",X"F8",X"04",X"F4",X"F4",X"FC",X"F8",X"00",X"F0",
		X"00",X"30",X"30",X"00",X"30",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"0C",X"00",X"00",X"00",
		X"1F",X"20",X"2F",X"2F",X"3F",X"10",X"0F",X"0F",X"F8",X"04",X"F4",X"F4",X"FC",X"08",X"F0",X"F0",
		X"00",X"30",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"0C",X"00",X"00",X"00",
		X"1F",X"20",X"2F",X"2F",X"30",X"1F",X"0F",X"0F",X"F8",X"04",X"F4",X"F4",X"0C",X"F8",X"F0",X"F0",
		X"00",X"01",X"31",X"30",X"30",X"00",X"00",X"00",X"00",X"80",X"8C",X"0C",X"0C",X"00",X"00",X"00",
		X"1F",X"20",X"2F",X"20",X"3F",X"1F",X"0F",X"0F",X"F8",X"04",X"F4",X"04",X"FC",X"F8",X"F0",X"F0",
		X"03",X"05",X"09",X"11",X"21",X"0F",X"08",X"08",X"80",X"80",X"FC",X"80",X"80",X"F0",X"10",X"10",
		X"08",X"0F",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"10",X"F0",X"F0",X"F0",X"70",X"60",X"40",X"00",
		X"09",X"09",X"09",X"09",X"09",X"0F",X"08",X"08",X"C0",X"A0",X"90",X"88",X"84",X"F0",X"10",X"10",
		X"08",X"0F",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"10",X"F0",X"F0",X"F0",X"70",X"60",X"40",X"00",
		X"1F",X"3F",X"2F",X"1F",X"3F",X"1F",X"1F",X"1F",X"F8",X"FC",X"F4",X"F8",X"FC",X"F8",X"F8",X"F8",
		X"1B",X"1B",X"3B",X"18",X"2C",X"3F",X"11",X"01",X"D8",X"D8",X"DC",X"18",X"34",X"FC",X"88",X"80",
		X"1F",X"3E",X"1E",X"28",X"38",X"18",X"1E",X"1E",X"F8",X"7C",X"78",X"14",X"1C",X"18",X"78",X"78",
		X"1B",X"1B",X"3B",X"28",X"1C",X"3F",X"1F",X"0F",X"D8",X"D8",X"DC",X"14",X"38",X"FC",X"F8",X"F0",
		X"21",X"11",X"09",X"05",X"03",X"0F",X"08",X"08",X"90",X"90",X"90",X"90",X"90",X"F0",X"10",X"10",
		X"08",X"0F",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"10",X"F0",X"F0",X"F0",X"70",X"60",X"40",X"00",
		X"01",X"01",X"3F",X"01",X"01",X"0F",X"08",X"08",X"84",X"88",X"90",X"A0",X"C0",X"F0",X"10",X"10",
		X"08",X"0F",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"10",X"F0",X"F0",X"F0",X"70",X"60",X"40",X"00",
		X"80",X"C0",X"E0",X"F0",X"38",X"3C",X"FE",X"FF",X"3E",X"7F",X"C3",X"C3",X"C3",X"C3",X"7F",X"3E",
		X"00",X"00",X"00",X"FF",X"81",X"FF",X"00",X"00",X"00",X"FC",X"02",X"82",X"82",X"82",X"C2",X"7A",
		X"0D",X"3D",X"7D",X"7D",X"7D",X"3D",X"0D",X"07",X"02",X"02",X"02",X"02",X"02",X"FC",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"4C",X"52",X"52",X"20",X"20",X"2F",X"2F",X"20",X"1F",X"3C",X"3C",
		X"22",X"00",X"3E",X"48",X"48",X"3E",X"00",X"4E",X"FC",X"FC",X"3C",X"FC",X"FC",X"3C",X"FC",X"FC",
		X"4A",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"3C",X"1F",X"20",X"20",X"21",X"23",X"23",X"2F",
		X"18",X"3C",X"7E",X"FF",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"FF",X"7E",X"3C",X"18",
		X"10",X"30",X"7F",X"FF",X"FF",X"7F",X"30",X"10",X"08",X"0C",X"FE",X"FF",X"FF",X"FE",X"0C",X"08",
		X"00",X"00",X"00",X"00",X"10",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",
		X"00",X"08",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"84",X"10",X"00",X"00",X"40",X"04",X"00",X"00",X"50",X"00",X"22",
		X"8A",X"00",X"00",X"00",X"04",X"00",X"20",X"04",X"00",X"80",X"10",X"00",X"14",X"80",X"20",X"00",
		X"00",X"00",X"08",X"04",X"00",X"01",X"23",X"01",X"00",X"00",X"41",X"02",X"08",X"C0",X"B2",X"68",
		X"86",X"13",X"20",X"07",X"03",X"00",X"10",X"00",X"48",X"D4",X"B0",X"64",X"C0",X"08",X"01",X"10",
		X"00",X"00",X"00",X"2C",X"EF",X"3D",X"30",X"F0",X"00",X"00",X"00",X"16",X"F7",X"FF",X"01",X"FE",
		X"F0",X"30",X"3D",X"EF",X"2C",X"00",X"00",X"00",X"FE",X"01",X"FF",X"F7",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"34",X"F7",X"FC",X"F0",X"F0",X"00",X"00",X"00",X"1A",X"FB",X"FF",X"00",X"FE",
		X"F0",X"F0",X"FC",X"F7",X"34",X"00",X"00",X"00",X"FE",X"00",X"FF",X"FB",X"1A",X"00",X"00",X"00",
		X"0F",X"0F",X"1F",X"1F",X"04",X"1C",X"08",X"08",X"F0",X"F0",X"F8",X"F8",X"20",X"38",X"10",X"10",
		X"0D",X"0D",X"0D",X"1D",X"1D",X"05",X"1D",X"0C",X"B0",X"B0",X"B0",X"B8",X"B8",X"A0",X"B8",X"30",
		X"09",X"09",X"1F",X"07",X"1C",X"1C",X"08",X"0C",X"90",X"90",X"F8",X"E0",X"38",X"38",X"10",X"30",
		X"0D",X"0D",X"0D",X"1D",X"05",X"1D",X"1D",X"0E",X"B0",X"B0",X"B0",X"B8",X"A0",X"B8",X"B8",X"70",
		X"80",X"C0",X"E0",X"F0",X"38",X"3C",X"3E",X"3F",X"01",X"03",X"07",X"0F",X"1C",X"3C",X"7C",X"FC",
		X"C3",X"C3",X"C3",X"C3",X"3C",X"3C",X"3C",X"3C",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
