library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity d1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of d1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"34",X"00",X"36",X"00",X"36",X"00",X"0E",X"00",
		X"0F",X"00",X"6F",X"00",X"2F",X"00",X"31",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"FC",X"00",X"F0",X"01",X"E0",X"03",
		X"40",X"00",X"78",X"00",X"18",X"00",X"B0",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"80",X"0F",X"90",X"0F",
		X"B0",X"07",X"20",X"07",X"00",X"03",X"40",X"01",X"C0",X"01",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"1F",X"00",X"07",X"80",X"07",X"80",X"07",
		X"C0",X"12",X"C0",X"12",X"80",X"37",X"00",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"40",X"48",X"41",X"08",X"42",X"C8",X"42",X"03",X"C0",X"00",X"07",X"E0",X"00",X"0D",X"B0",
		X"00",X"19",X"98",X"00",X"11",X"88",X"00",X"91",X"89",X"00",X"D5",X"AB",X"00",X"FD",X"BF",X"00",
		X"FD",X"BF",X"00",X"D5",X"AB",X"00",X"91",X"89",X"00",X"11",X"88",X"00",X"19",X"98",X"00",X"0D",
		X"B0",X"00",X"07",X"E0",X"00",X"03",X"C0",X"00",X"0C",X"00",X"03",X"1C",X"80",X"03",X"34",X"C0",
		X"02",X"64",X"60",X"02",X"44",X"20",X"02",X"44",X"26",X"02",X"54",X"AF",X"02",X"F4",X"FF",X"02",
		X"F4",X"FF",X"02",X"54",X"AF",X"02",X"44",X"26",X"02",X"44",X"20",X"02",X"64",X"60",X"02",X"34",
		X"C0",X"02",X"1C",X"80",X"03",X"0C",X"00",X"03",X"30",X"00",X"0C",X"70",X"00",X"0E",X"D0",X"00",
		X"0B",X"90",X"81",X"09",X"10",X"81",X"08",X"10",X"99",X"08",X"50",X"BD",X"0A",X"D0",X"FF",X"0B",
		X"D0",X"FF",X"0B",X"50",X"BD",X"0A",X"10",X"99",X"08",X"10",X"81",X"08",X"90",X"81",X"09",X"D0",
		X"00",X"0B",X"70",X"00",X"0E",X"30",X"00",X"0C",X"C0",X"00",X"30",X"C0",X"01",X"38",X"40",X"03",
		X"2C",X"40",X"06",X"26",X"40",X"04",X"22",X"40",X"64",X"22",X"40",X"F5",X"2A",X"40",X"FF",X"2F",
		X"40",X"FF",X"2F",X"40",X"F5",X"2A",X"40",X"64",X"22",X"40",X"04",X"22",X"40",X"06",X"26",X"40",
		X"03",X"2C",X"C0",X"01",X"38",X"C0",X"00",X"30",X"F8",X"00",X"00",X"8C",X"00",X"00",X"CE",X"00",
		X"00",X"7F",X"00",X"00",X"39",X"00",X"00",X"F9",X"01",X"00",X"ED",X"03",X"00",X"E7",X"07",X"00",
		X"E0",X"E7",X"00",X"C0",X"B7",X"00",X"80",X"9F",X"00",X"00",X"9C",X"00",X"00",X"FE",X"00",X"00",
		X"73",X"00",X"00",X"31",X"00",X"00",X"1F",X"00",X"E0",X"03",X"00",X"30",X"02",X"00",X"38",X"03",
		X"00",X"FC",X"01",X"00",X"E4",X"00",X"00",X"E4",X"07",X"00",X"B4",X"0F",X"00",X"9C",X"1F",X"00",
		X"80",X"9F",X"03",X"00",X"DF",X"02",X"00",X"7E",X"02",X"00",X"70",X"02",X"00",X"F8",X"03",X"00",
		X"CC",X"01",X"00",X"C4",X"00",X"00",X"7C",X"00",X"80",X"0F",X"00",X"C0",X"08",X"00",X"E0",X"0C",
		X"00",X"F0",X"07",X"00",X"90",X"03",X"00",X"90",X"1F",X"00",X"D0",X"3E",X"00",X"70",X"7E",X"00",
		X"00",X"7E",X"0E",X"00",X"7C",X"0B",X"00",X"F8",X"09",X"00",X"C0",X"09",X"00",X"E0",X"0F",X"00",
		X"30",X"07",X"00",X"10",X"03",X"00",X"F0",X"01",X"00",X"3E",X"00",X"00",X"23",X"00",X"80",X"33",
		X"00",X"C0",X"1F",X"00",X"40",X"0E",X"00",X"40",X"7E",X"00",X"40",X"FB",X"00",X"C0",X"F9",X"01",
		X"00",X"F8",X"39",X"00",X"F0",X"2D",X"00",X"E0",X"27",X"00",X"00",X"27",X"00",X"80",X"3F",X"00",
		X"C0",X"1C",X"00",X"40",X"0C",X"00",X"C0",X"07",X"FF",X"FF",X"00",X"03",X"C0",X"00",X"C6",X"63",
		X"00",X"8C",X"31",X"00",X"F8",X"1F",X"00",X"80",X"01",X"00",X"C0",X"03",X"00",X"E0",X"07",X"00",
		X"E0",X"07",X"00",X"C0",X"03",X"00",X"80",X"01",X"00",X"F8",X"1F",X"00",X"8C",X"31",X"00",X"C6",
		X"63",X"00",X"03",X"C0",X"00",X"FF",X"FF",X"00",X"FC",X"FF",X"03",X"0C",X"00",X"03",X"18",X"8F",
		X"01",X"30",X"C6",X"00",X"E0",X"7F",X"00",X"00",X"06",X"00",X"00",X"0F",X"00",X"80",X"1F",X"00",
		X"80",X"1F",X"00",X"00",X"0F",X"00",X"00",X"06",X"00",X"E0",X"7F",X"00",X"30",X"C6",X"00",X"18",
		X"8F",X"01",X"0C",X"00",X"03",X"FC",X"FF",X"03",X"F0",X"FF",X"0F",X"30",X"00",X"0C",X"60",X"3C",
		X"06",X"C0",X"18",X"03",X"80",X"FF",X"01",X"00",X"18",X"00",X"00",X"3C",X"00",X"00",X"7E",X"00",
		X"00",X"7E",X"00",X"00",X"3C",X"00",X"00",X"18",X"00",X"80",X"FF",X"01",X"C0",X"18",X"03",X"60",
		X"3C",X"06",X"30",X"00",X"0C",X"F0",X"FF",X"0F",X"C0",X"FF",X"3F",X"C0",X"00",X"30",X"80",X"F1",
		X"18",X"00",X"63",X"0C",X"00",X"FE",X"07",X"00",X"60",X"00",X"00",X"F0",X"00",X"00",X"F8",X"01",
		X"00",X"F8",X"01",X"00",X"F0",X"00",X"00",X"60",X"00",X"00",X"FE",X"07",X"00",X"63",X"0C",X"80",
		X"F1",X"18",X"C0",X"00",X"30",X"C0",X"FF",X"3F",X"00",X"1F",X"00",X"00",X"31",X"00",X"00",X"73",
		X"00",X"00",X"FE",X"00",X"00",X"9C",X"00",X"80",X"9F",X"00",X"C0",X"B7",X"00",X"E0",X"E7",X"00",
		X"E7",X"07",X"00",X"ED",X"03",X"00",X"F9",X"01",X"00",X"39",X"00",X"00",X"7F",X"00",X"00",X"CE",
		X"00",X"00",X"8C",X"00",X"00",X"F8",X"00",X"00",X"00",X"7C",X"00",X"00",X"C4",X"00",X"00",X"CC",
		X"01",X"00",X"F8",X"03",X"00",X"70",X"02",X"00",X"7E",X"02",X"00",X"DF",X"02",X"80",X"9F",X"03",
		X"9C",X"1F",X"00",X"B4",X"0F",X"00",X"E4",X"07",X"00",X"E4",X"00",X"00",X"FC",X"01",X"00",X"38",
		X"03",X"00",X"30",X"02",X"00",X"E0",X"03",X"00",X"00",X"F0",X"01",X"00",X"10",X"03",X"00",X"30",
		X"07",X"00",X"E0",X"0F",X"00",X"C0",X"09",X"00",X"F8",X"09",X"00",X"7C",X"0B",X"00",X"7E",X"0E",
		X"70",X"7E",X"00",X"D0",X"3E",X"00",X"90",X"1F",X"00",X"90",X"03",X"00",X"F0",X"07",X"00",X"E0",
		X"0C",X"00",X"C0",X"08",X"00",X"80",X"0F",X"00",X"00",X"C0",X"07",X"00",X"40",X"0C",X"00",X"C0",
		X"1C",X"00",X"80",X"3F",X"00",X"00",X"27",X"00",X"E0",X"27",X"00",X"F0",X"2D",X"00",X"F8",X"39",
		X"C0",X"F9",X"01",X"40",X"FB",X"00",X"40",X"7E",X"00",X"40",X"0E",X"00",X"C0",X"1F",X"00",X"80",
		X"33",X"00",X"00",X"23",X"00",X"00",X"3E",X"00",X"08",X"00",X"36",X"00",X"41",X"00",X"22",X"00",
		X"41",X"00",X"36",X"00",X"08",X"00",X"00",X"00",X"20",X"00",X"D8",X"00",X"04",X"01",X"88",X"00",
		X"04",X"01",X"D8",X"00",X"20",X"00",X"00",X"00",X"80",X"00",X"60",X"03",X"10",X"04",X"20",X"02",
		X"10",X"04",X"60",X"03",X"80",X"00",X"00",X"00",X"00",X"02",X"80",X"0D",X"40",X"10",X"80",X"08",
		X"40",X"10",X"80",X"0D",X"00",X"02",X"00",X"00",X"41",X"63",X"6B",X"7F",X"6B",X"63",X"41",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"F0",X"44",X"CD",X"0D",X"44",X"C9",X"C3",X"0F",X"45",X"C3",X"72",X"44",X"3A",X"D9",X"20",
		X"B7",X"C8",X"3A",X"E2",X"21",X"B7",X"C2",X"28",X"44",X"AF",X"21",X"10",X"22",X"BE",X"CA",X"38",
		X"44",X"21",X"30",X"22",X"BE",X"CA",X"38",X"44",X"AF",X"21",X"50",X"22",X"BE",X"CA",X"38",X"44",
		X"21",X"70",X"22",X"BE",X"CA",X"38",X"44",X"C9",X"3A",X"19",X"23",X"B7",X"CA",X"A8",X"44",X"3D",
		X"32",X"19",X"23",X"7D",X"D6",X"10",X"6F",X"EB",X"2A",X"1A",X"23",X"22",X"20",X"23",X"22",X"22",
		X"23",X"7D",X"D6",X"0C",X"6F",X"22",X"1A",X"23",X"21",X"20",X"23",X"06",X"20",X"FF",X"7B",X"D6",
		X"16",X"5F",X"3A",X"56",X"23",X"C6",X"02",X"E6",X"07",X"32",X"56",X"23",X"47",X"1A",X"90",X"12",
		X"C9",X"C9",X"21",X"03",X"22",X"11",X"0D",X"00",X"01",X"13",X"00",X"7E",X"19",X"FE",X"2F",X"D2",
		X"85",X"44",X"7E",X"B7",X"C0",X"09",X"7E",X"19",X"FE",X"2F",X"D2",X"90",X"44",X"7E",X"B7",X"C0",
		X"09",X"7E",X"19",X"FE",X"2F",X"D2",X"9B",X"44",X"7E",X"B7",X"C0",X"09",X"7E",X"19",X"FE",X"2F",
		X"D2",X"A6",X"44",X"7E",X"B7",X"C0",X"AF",X"C9",X"CD",X"0A",X"44",X"C0",X"21",X"03",X"23",X"7E",
		X"34",X"FE",X"04",X"DA",X"BA",X"44",X"3E",X"02",X"36",X"03",X"00",X"00",X"00",X"E6",X"03",X"07",
		X"07",X"07",X"47",X"07",X"07",X"80",X"21",X"6C",X"06",X"85",X"D2",X"CE",X"44",X"24",X"6F",X"11",
		X"18",X"23",X"06",X"28",X"FF",X"21",X"7E",X"47",X"F7",X"3A",X"03",X"23",X"3D",X"85",X"D2",X"E2",
		X"44",X"24",X"6F",X"7E",X"32",X"18",X"23",X"CD",X"2A",X"50",X"C3",X"F0",X"44",X"00",X"00",X"00",
		X"21",X"18",X"23",X"7E",X"B7",X"C8",X"35",X"23",X"34",X"2A",X"1E",X"23",X"44",X"4D",X"21",X"1C",
		X"23",X"CD",X"3F",X"14",X"2A",X"1C",X"23",X"7D",X"D6",X"0C",X"6F",X"22",X"1C",X"23",X"C9",X"01",
		X"E3",X"21",X"0A",X"FE",X"02",X"D4",X"AF",X"47",X"07",X"E6",X"0E",X"21",X"2B",X"45",X"85",X"D2",
		X"23",X"45",X"24",X"6F",X"5E",X"23",X"56",X"EB",X"50",X"59",X"E9",X"3B",X"45",X"85",X"45",X"CD",
		X"45",X"E7",X"45",X"39",X"46",X"FD",X"46",X"17",X"47",X"34",X"47",X"21",X"E0",X"21",X"CD",X"6B",
		X"47",X"C0",X"3A",X"22",X"20",X"B7",X"C8",X"3A",X"90",X"21",X"B7",X"C0",X"21",X"E8",X"21",X"7E",
		X"07",X"E6",X"06",X"34",X"01",X"73",X"45",X"81",X"D2",X"5C",X"45",X"04",X"4F",X"0A",X"6F",X"03",
		X"0A",X"67",X"22",X"E0",X"21",X"EB",X"34",X"2B",X"36",X"FF",X"21",X"EB",X"21",X"36",X"1E",X"23",
		X"36",X"00",X"C9",X"00",X"04",X"00",X"08",X"00",X"02",X"00",X"01",X"EB",X"36",X"00",X"21",X"B4",
		X"00",X"22",X"E0",X"21",X"C9",X"3A",X"22",X"20",X"B7",X"CA",X"7B",X"45",X"3A",X"10",X"22",X"21",
		X"30",X"22",X"B6",X"C0",X"E5",X"21",X"EB",X"21",X"EF",X"23",X"36",X"FF",X"E1",X"C0",X"EB",X"34",
		X"11",X"80",X"22",X"21",X"00",X"58",X"06",X"40",X"FF",X"CD",X"8C",X"5A",X"3A",X"0A",X"20",X"3D",
		X"32",X"97",X"22",X"32",X"B7",X"22",X"21",X"F1",X"22",X"36",X"00",X"21",X"00",X"00",X"22",X"D2",
		X"22",X"21",X"F3",X"22",X"36",X"FF",X"21",X"D9",X"22",X"7E",X"07",X"77",X"C9",X"3A",X"91",X"22",
		X"21",X"B1",X"22",X"B6",X"CA",X"DC",X"45",X"EB",X"34",X"C3",X"0E",X"46",X"3A",X"90",X"22",X"21",
		X"B0",X"22",X"B6",X"C0",X"C3",X"37",X"47",X"21",X"E6",X"21",X"EF",X"C0",X"3E",X"52",X"32",X"4B",
		X"22",X"32",X"6B",X"22",X"36",X"03",X"21",X"E5",X"21",X"34",X"4E",X"7E",X"FE",X"11",X"D2",X"0B",
		X"46",X"CD",X"15",X"46",X"21",X"D0",X"58",X"CD",X"29",X"46",X"C9",X"EB",X"34",X"C9",X"21",X"AA",
		X"0A",X"22",X"54",X"23",X"C9",X"3A",X"0A",X"20",X"C6",X"11",X"91",X"26",X"00",X"6F",X"29",X"29",
		X"29",X"29",X"29",X"11",X"0B",X"24",X"19",X"EB",X"C9",X"06",X"09",X"FF",X"7B",X"C6",X"17",X"D2",
		X"33",X"46",X"14",X"5F",X"0D",X"C2",X"29",X"46",X"C9",X"3A",X"54",X"23",X"FE",X"83",X"D2",X"6A",
		X"46",X"21",X"E5",X"21",X"35",X"4E",X"7E",X"FE",X"00",X"CA",X"37",X"47",X"CD",X"15",X"46",X"21",
		X"40",X"58",X"06",X"09",X"3E",X"00",X"12",X"13",X"05",X"C2",X"56",X"46",X"7B",X"C6",X"17",X"D2",
		X"63",X"46",X"14",X"5F",X"0D",X"C8",X"CD",X"29",X"46",X"C9",X"21",X"EA",X"21",X"EF",X"C0",X"36",
		X"07",X"CD",X"D5",X"46",X"CD",X"96",X"47",X"21",X"90",X"22",X"7E",X"2F",X"23",X"B6",X"C8",X"21",
		X"B0",X"22",X"7E",X"2F",X"23",X"B6",X"C8",X"11",X"AC",X"2C",X"2A",X"54",X"23",X"E5",X"06",X"08",
		X"1A",X"E6",X"E0",X"4F",X"7E",X"B1",X"12",X"23",X"7B",X"C6",X"20",X"D2",X"9F",X"46",X"14",X"5F",
		X"05",X"C2",X"90",X"46",X"E1",X"E5",X"11",X"B0",X"2C",X"06",X"08",X"1A",X"E6",X"3F",X"4F",X"7E",
		X"0F",X"0F",X"E6",X"C0",X"B1",X"12",X"13",X"1A",X"E6",X"F8",X"4F",X"7E",X"0F",X"0F",X"E6",X"07",
		X"B1",X"12",X"23",X"7B",X"C6",X"1F",X"D2",X"CA",X"46",X"14",X"5F",X"05",X"C2",X"AB",X"46",X"E1",
		X"2B",X"22",X"54",X"23",X"C9",X"3A",X"E5",X"21",X"3D",X"C8",X"4F",X"CD",X"15",X"46",X"21",X"D0",
		X"58",X"CD",X"E5",X"46",X"C9",X"06",X"09",X"1A",X"B6",X"12",X"13",X"23",X"05",X"C2",X"E7",X"46",
		X"7B",X"C6",X"17",X"D2",X"F7",X"46",X"14",X"5F",X"0D",X"C2",X"E5",X"46",X"C9",X"CD",X"18",X"47",
		X"21",X"43",X"20",X"7E",X"E6",X"F3",X"77",X"21",X"E6",X"21",X"EF",X"C0",X"21",X"43",X"20",X"7E",
		X"F6",X"0C",X"77",X"EB",X"34",X"34",X"C9",X"C9",X"0E",X"10",X"21",X"2B",X"2C",X"3E",X"00",X"06",
		X"09",X"77",X"23",X"05",X"C2",X"21",X"47",X"7D",X"C6",X"17",X"D2",X"2E",X"47",X"24",X"6F",X"0D",
		X"C2",X"1D",X"47",X"C9",X"CD",X"18",X"47",X"21",X"E2",X"21",X"3E",X"00",X"77",X"23",X"77",X"23",
		X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"3E",X"38",X"32",X"4B",X"22",X"32",X"6B",X"22",X"21",
		X"43",X"20",X"7E",X"F6",X"0C",X"77",X"21",X"F3",X"22",X"AF",X"BE",X"CA",X"69",X"47",X"77",X"21",
		X"D9",X"22",X"7E",X"07",X"1F",X"1F",X"E6",X"7F",X"77",X"00",X"C9",X"7E",X"23",X"B6",X"2B",X"C8",
		X"D5",X"5E",X"23",X"56",X"1B",X"72",X"2B",X"73",X"7A",X"B3",X"D1",X"C0",X"37",X"C9",X"86",X"47",
		X"8A",X"47",X"8E",X"47",X"92",X"47",X"04",X"06",X"08",X"08",X"04",X"06",X"08",X"0A",X"06",X"08",
		X"0A",X"0C",X"06",X"0A",X"0C",X"0E",X"21",X"8E",X"21",X"EF",X"C0",X"36",X"02",X"23",X"AF",X"BE",
		X"2F",X"77",X"C8",X"11",X"D0",X"43",X"21",X"AF",X"2C",X"06",X"07",X"CD",X"0A",X"0E",X"C9",X"C5",
		X"F5",X"D5",X"21",X"90",X"22",X"7E",X"2F",X"23",X"B6",X"C2",X"D2",X"47",X"EB",X"21",X"83",X"22",
		X"3A",X"6B",X"20",X"C6",X"0A",X"BE",X"DA",X"D2",X"47",X"EB",X"2B",X"CD",X"80",X"5A",X"D1",X"F1",
		X"C1",X"C9",X"21",X"B0",X"22",X"7E",X"2F",X"23",X"B6",X"C2",X"CE",X"47",X"EB",X"21",X"A3",X"22",
		X"3A",X"6B",X"20",X"C6",X"0A",X"BE",X"DA",X"CE",X"47",X"C3",X"C9",X"47",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
