library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4C",X"54",X"A0",X"4C",X"09",X"A0",X"85",X"EF",X"EA",X"78",X"D8",X"AD",X"03",X"40",X"29",X"20",
		X"D0",X"06",X"4C",X"03",X"90",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"00",X"A2",X"FF",X"9A",X"A9",
		X"00",X"8D",X"00",X"40",X"8D",X"02",X"40",X"8D",X"03",X"40",X"8D",X"04",X"40",X"8D",X"05",X"40",
		X"8D",X"00",X"08",X"20",X"80",X"A4",X"A2",X"00",X"20",X"D7",X"A4",X"20",X"FA",X"A4",X"20",X"6E",
		X"A4",X"20",X"91",X"CE",X"AD",X"10",X"07",X"85",X"16",X"AD",X"11",X"07",X"85",X"15",X"4C",X"B0",
		X"A1",X"85",X"EF",X"EA",X"48",X"8A",X"48",X"98",X"48",X"AD",X"03",X"40",X"29",X"20",X"D0",X"06",
		X"4C",X"00",X"90",X"85",X"EF",X"EA",X"A5",X"00",X"F0",X"06",X"4C",X"00",X"90",X"85",X"EF",X"EA",
		X"A9",X"00",X"85",X"00",X"D8",X"A5",X"0B",X"F0",X"73",X"AD",X"04",X"40",X"49",X"FF",X"29",X"E0",
		X"85",X"0D",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"20",X"50",X"A1",X"AD",X"02",X"40",X"29",X"C0",
		X"F0",X"5A",X"85",X"0C",X"20",X"50",X"A1",X"AD",X"02",X"40",X"25",X"0C",X"F0",X"4E",X"20",X"50",
		X"A1",X"AD",X"02",X"40",X"25",X"0C",X"F0",X"44",X"20",X"50",X"A1",X"AD",X"02",X"40",X"25",X"0C",
		X"F0",X"3A",X"E6",X"0F",X"A9",X"10",X"8D",X"03",X"40",X"A5",X"0D",X"C9",X"80",X"F0",X"39",X"A2",
		X"00",X"AD",X"03",X"40",X"49",X"FF",X"29",X"0F",X"06",X"0C",X"90",X"05",X"4A",X"4A",X"85",X"EF",
		X"EA",X"29",X"03",X"F0",X"51",X"E8",X"C9",X"01",X"F0",X"4C",X"E8",X"C9",X"02",X"F0",X"3C",X"E8",
		X"85",X"EF",X"EA",X"A5",X"0F",X"C9",X"02",X"B0",X"2A",X"85",X"EF",X"EA",X"8D",X"00",X"40",X"68",
		X"A8",X"68",X"AA",X"68",X"40",X"85",X"EF",X"EA",X"A2",X"05",X"A5",X"0C",X"C9",X"40",X"F0",X"26",
		X"E8",X"C9",X"80",X"F0",X"21",X"E8",X"C9",X"C0",X"F0",X"D9",X"4C",X"EC",X"A0",X"85",X"EF",X"6E",
		X"85",X"EF",X"EA",X"C6",X"0F",X"A4",X"26",X"A1",X"85",X"EF",X"EA",X"A5",X"0D",X"C9",X"60",X"D0",
		X"05",X"A2",X"04",X"85",X"EF",X"6E",X"A5",X"0E",X"F8",X"18",X"7D",X"5F",X"A1",X"D9",X"67",X"A1",
		X"90",X"06",X"B9",X"67",X"A1",X"85",X"EF",X"6E",X"85",X"0E",X"D8",X"C6",X"0F",X"C9",X"10",X"D0",
		X"AB",X"8D",X"00",X"40",X"4D",X"01",X"85",X"10",X"A2",X"FF",X"9A",X"4C",X"72",X"A1",X"85",X"EF",
		X"EA",X"A2",X"E7",X"85",X"EF",X"6E",X"A5",X"FF",X"A5",X"FF",X"EA",X"CA",X"D0",X"F8",X"60",X"01",
		X"02",X"03",X"01",X"06",X"08",X"03",X"01",X"09",X"09",X"16",X"16",X"16",X"09",X"09",X"09",X"85",
		X"EF",X"EA",X"20",X"B8",X"A5",X"20",X"A0",X"A4",X"20",X"19",X"C9",X"20",X"E6",X"DA",X"85",X"EF",
		X"EA",X"20",X"98",X"D3",X"20",X"14",X"DB",X"A9",X"00",X"85",X"11",X"AD",X"02",X"40",X"49",X"FF",
		X"29",X"03",X"F0",X"ED",X"C9",X"01",X"F0",X"12",X"C9",X"02",X"D0",X"E5",X"A5",X"0E",X"C9",X"02",
		X"90",X"DF",X"20",X"2A",X"A6",X"E6",X"11",X"C1",X"EF",X"EA",X"20",X"2A",X"A6",X"85",X"EF",X"6E",
		X"E6",X"11",X"85",X"EF",X"6E",X"A2",X"1D",X"20",X"73",X"A4",X"A2",X"01",X"20",X"D7",X"A4",X"A9",
		X"00",X"8D",X"04",X"40",X"08",X"80",X"A4",X"20",X"08",X"C9",X"20",X"AD",X"CE",X"20",X"C4",X"CE",
		X"20",X"E0",X"CE",X"20",X"E4",X"D3",X"85",X"EF",X"EA",X"20",X"37",X"A6",X"20",X"29",X"D4",X"20",
		X"BA",X"D4",X"20",X"29",X"D0",X"A9",X"01",X"85",X"0B",X"A9",X"00",X"85",X"12",X"08",X"A0",X"A4",
		X"A9",X"FF",X"85",X"20",X"C1",X"30",X"4D",X"00",X"85",X"21",X"85",X"31",X"4D",X"80",X"85",X"1E",
		X"85",X"2E",X"A5",X"10",X"D0",X"0C",X"20",X"B8",X"A5",X"20",X"7B",X"D8",X"20",X"18",X"D9",X"85",
		X"EF",X"EA",X"C6",X"1F",X"C6",X"2F",X"85",X"EF",X"EA",X"20",X"C1",X"A5",X"A2",X"80",X"20",X"C9",
		X"CE",X"20",X"75",X"D4",X"20",X"70",X"C1",X"A9",X"00",X"8D",X"04",X"40",X"A5",X"12",X"8D",X"02",
		X"40",X"A9",X"A2",X"48",X"A9",X"46",X"48",X"A5",X"3E",X"10",X"06",X"4C",X"46",X"A3",X"85",X"EF",
		X"EA",X"4C",X"86",X"A3",X"85",X"EF",X"EA",X"20",X"FB",X"D3",X"20",X"F1",X"A5",X"20",X"29",X"D4",
		X"20",X"59",X"DB",X"20",X"5A",X"A5",X"20",X"D5",X"A6",X"A9",X"20",X"20",X"74",X"A6",X"20",X"A0",
		X"A4",X"20",X"45",X"CD",X"85",X"EF",X"EA",X"20",X"4F",X"A4",X"20",X"F8",X"A6",X"20",X"22",X"A7",
		X"20",X"97",X"C6",X"20",X"25",X"C4",X"20",X"9D",X"CE",X"20",X"E9",X"A7",X"20",X"B1",X"AE",X"20",
		X"FF",X"AD",X"20",X"97",X"B2",X"20",X"8D",X"BE",X"20",X"65",X"B3",X"20",X"20",X"AF",X"20",X"B7",
		X"B2",X"20",X"66",X"AC",X"20",X"F8",X"CE",X"20",X"35",X"CF",X"20",X"22",X"CA",X"20",X"17",X"D3",
		X"20",X"45",X"D3",X"20",X"6D",X"D3",X"20",X"5E",X"CD",X"A5",X"10",X"F0",X"09",X"20",X"33",X"D0",
		X"20",X"29",X"D0",X"85",X"EF",X"EA",X"33",X"1D",X"10",X"AD",X"A9",X"00",X"20",X"86",X"D3",X"20",
		X"A0",X"A4",X"20",X"B8",X"A5",X"24",X"1D",X"70",X"05",X"C6",X"3F",X"85",X"EF",X"EA",X"20",X"D8",
		X"A5",X"20",X"04",X"A6",X"24",X"1D",X"50",X"06",X"4C",X"19",X"A2",X"85",X"EF",X"EA",X"A5",X"10",
		X"F0",X"46",X"A5",X"3F",X"30",X"1A",X"A5",X"11",X"C9",X"02",X"B0",X"06",X"4C",X"19",X"A2",X"85",
		X"EF",X"EA",X"E6",X"12",X"A5",X"12",X"29",X"01",X"85",X"12",X"4C",X"19",X"A2",X"85",X"EF",X"EA",
		X"20",X"12",X"D4",X"A9",X"FF",X"20",X"74",X"A6",X"20",X"6D",X"DB",X"C6",X"11",X"70",X"E3",X"A9",
		X"00",X"8D",X"02",X"40",X"C1",X"12",X"C9",X"0E",X"D0",X"08",X"85",X"10",X"A4",X"B0",X"A1",X"85",
		X"EF",X"EA",X"4C",X"72",X"A1",X"85",X"EF",X"6E",X"E6",X"1C",X"A5",X"1C",X"C9",X"04",X"90",X"0A",
		X"A9",X"00",X"85",X"1C",X"A4",X"00",X"A3",X"85",X"EF",X"EA",X"A9",X"80",X"85",X"1E",X"EA",X"1F",
		X"4C",X"19",X"A2",X"85",X"EF",X"6E",X"E6",X"40",X"F8",X"A5",X"41",X"38",X"69",X"00",X"85",X"41",
		X"D8",X"A2",X"4F",X"20",X"73",X"A4",X"20",X"81",X"C1",X"A9",X"00",X"85",X"59",X"C1",X"5A",X"C9",
		X"3E",X"29",X"20",X"09",X"01",X"85",X"3E",X"4D",X"80",X"85",X"C7",X"A9",X"00",X"85",X"1D",X"C1",
		X"EF",X"EA",X"A9",X"00",X"85",X"4C",X"4D",X"10",X"85",X"49",X"A9",X"0F",X"85",X"4A",X"4D",X"03",
		X"85",X"4B",X"60",X"85",X"EF",X"6E",X"A2",X"4F",X"20",X"73",X"A4",X"20",X"A0",X"A4",X"A9",X"42",
		X"20",X"86",X"D3",X"A5",X"3E",X"29",X"20",X"85",X"3E",X"A9",X"00",X"85",X"1D",X"C1",X"C7",X"C1",
		X"59",X"85",X"5A",X"20",X"C5",X"A7",X"A9",X"80",X"85",X"9D",X"85",X"D7",X"C9",X"46",X"38",X"E9",
		X"98",X"85",X"48",X"F0",X"07",X"90",X"24",X"B0",X"54",X"85",X"EF",X"EA",X"A5",X"45",X"85",X"7E",
		X"85",X"80",X"A5",X"46",X"85",X"7F",X"C1",X"81",X"A5",X"47",X"85",X"7C",X"C1",X"EF",X"6E",X"A9",
		X"80",X"85",X"7B",X"A9",X"00",X"85",X"48",X"28",X"85",X"EF",X"EA",X"A5",X"48",X"49",X"FF",X"38",
		X"69",X"00",X"85",X"48",X"C9",X"49",X"38",X"E5",X"48",X"85",X"49",X"B0",X"05",X"E6",X"4C",X"C1",
		X"EF",X"EA",X"A5",X"46",X"18",X"65",X"48",X"85",X"46",X"A5",X"4A",X"38",X"E5",X"48",X"85",X"4A",
		X"B0",X"05",X"C6",X"4B",X"85",X"EF",X"EA",X"4C",X"BC",X"A3",X"85",X"EF",X"EA",X"A5",X"4A",X"18",
		X"65",X"48",X"85",X"02",X"A5",X"4B",X"69",X"00",X"85",X"03",X"C9",X"03",X"90",X"0F",X"A5",X"02",
		X"C9",X"0F",X"90",X"09",X"20",X"9E",X"A7",X"4C",X"72",X"A3",X"85",X"EF",X"EA",X"A5",X"46",X"38",
		X"E5",X"48",X"85",X"46",X"A5",X"49",X"18",X"65",X"48",X"85",X"49",X"90",X"05",X"C6",X"4C",X"85",
		X"EF",X"EA",X"A5",X"02",X"85",X"4A",X"A5",X"03",X"85",X"4B",X"4C",X"BC",X"A3",X"85",X"EF",X"EA",
		X"AD",X"03",X"40",X"10",X"FB",X"20",X"88",X"A5",X"20",X"91",X"A6",X"20",X"43",X"CE",X"58",X"EA",
		X"EA",X"EA",X"78",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"30",X"FB",X"60",X"85",X"EF",X"EA",X"A2",
		X"01",X"85",X"EF",X"EA",X"A9",X"00",X"95",X"00",X"E8",X"E0",X"EE",X"90",X"F7",X"60",X"85",X"EF",
		X"EA",X"A9",X"10",X"85",X"02",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"01",X"A8",X"85",X"EF",X"EA",
		X"91",X"01",X"C8",X"D0",X"FB",X"E6",X"02",X"A5",X"02",X"C9",X"18",X"90",X"EB",X"60",X"85",X"EF",
		X"EA",X"A9",X"10",X"85",X"02",X"85",X"EF",X"EA",X"A0",X"E1",X"85",X"EF",X"EA",X"A9",X"00",X"85",
		X"01",X"85",X"EF",X"EA",X"91",X"01",X"C8",X"D0",X"05",X"E6",X"02",X"85",X"EF",X"EA",X"C0",X"A0",
		X"D0",X"F2",X"A5",X"02",X"C9",X"17",X"F0",X"0C",X"C9",X"13",X"D0",X"E1",X"E6",X"02",X"4C",X"A8",
		X"A4",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A9",X"02",X"85",X"02",X"85",X"EF",X"EA",X"A9",
		X"00",X"85",X"01",X"A8",X"85",X"EF",X"EA",X"91",X"01",X"C8",X"D0",X"FB",X"E6",X"02",X"A5",X"02",
		X"DD",X"F6",X"A4",X"90",X"EA",X"60",X"08",X"07",X"85",X"EF",X"EA",X"A2",X"07",X"85",X"EF",X"EA",
		X"BD",X"10",X"A5",X"9D",X"00",X"0C",X"DD",X"18",X"A5",X"9D",X"08",X"0C",X"66",X"10",X"F1",X"60",
		X"FF",X"38",X"C0",X"3F",X"00",X"F8",X"FF",X"07",X"F8",X"C0",X"88",X"FF",X"3F",X"75",X"F8",X"88",
		X"D0",X"C7",X"38",X"FF",X"3F",X"75",X"D0",X"38",X"CF",X"00",X"C0",X"FF",X"3F",X"75",X"CF",X"C0",
		X"78",X"F8",X"F8",X"FF",X"3F",X"75",X"78",X"F8",X"3F",X"C0",X"88",X"FF",X"38",X"72",X"3F",X"88",
		X"D0",X"C7",X"3F",X"FF",X"38",X"72",X"D0",X"3F",X"CF",X"00",X"C0",X"FF",X"38",X"72",X"CF",X"C0",
		X"F8",X"F8",X"C0",X"FF",X"38",X"72",X"F8",X"C0",X"85",X"EF",X"EA",X"A5",X"40",X"38",X"85",X"EF",
		X"EA",X"E9",X"08",X"B0",X"FC",X"69",X"08",X"AA",X"A9",X"F8",X"85",X"EF",X"6E",X"18",X"69",X"08",
		X"CA",X"10",X"FA",X"AA",X"A0",X"00",X"85",X"EF",X"EA",X"BD",X"18",X"A5",X"99",X"08",X"0C",X"6C",
		X"C8",X"C0",X"08",X"90",X"F4",X"60",X"85",X"EF",X"EA",X"A5",X"C7",X"30",X"1E",X"F0",X"1C",X"A6",
		X"B4",X"A5",X"40",X"85",X"EF",X"6E",X"38",X"E9",X"04",X"B0",X"FB",X"7D",X"B4",X"A5",X"AA",X"85",
		X"EF",X"EA",X"BD",X"AC",X"A5",X"8D",X"01",X"0C",X"85",X"EF",X"EA",X"60",X"C0",X"C7",X"F8",X"C7",
		X"00",X"F8",X"88",X"07",X"04",X"08",X"85",X"EF",X"EA",X"A9",X"FF",X"8D",X"08",X"0C",X"28",X"85",
		X"EF",X"EA",X"A4",X"12",X"BE",X"ED",X"A5",X"A0",X"0F",X"85",X"EF",X"EA",X"B5",X"00",X"99",X"3E",
		X"00",X"CA",X"88",X"10",X"F7",X"60",X"85",X"EF",X"EA",X"A4",X"12",X"BE",X"ED",X"A5",X"A0",X"0F",
		X"85",X"EF",X"EA",X"B9",X"3E",X"00",X"95",X"00",X"CA",X"88",X"10",X"F7",X"60",X"2D",X"3D",X"85",
		X"EF",X"EA",X"20",X"17",X"A6",X"85",X"EF",X"6E",X"B1",X"01",X"9D",X"00",X"03",X"64",X"E8",X"D0",
		X"F7",X"60",X"85",X"EF",X"EA",X"20",X"17",X"A6",X"85",X"EF",X"EA",X"BD",X"00",X"03",X"91",X"01",
		X"E8",X"C8",X"D0",X"F7",X"60",X"85",X"EF",X"EA",X"A6",X"12",X"BD",X"26",X"A6",X"85",X"02",X"A9",
		X"00",X"85",X"01",X"AA",X"A8",X"60",X"05",X"06",X"85",X"EF",X"EA",X"F8",X"38",X"A5",X"0E",X"E9",
		X"01",X"85",X"0E",X"D8",X"60",X"85",X"EF",X"EA",X"AD",X"04",X"40",X"49",X"FF",X"48",X"29",X"01",
		X"AA",X"BD",X"60",X"A6",X"85",X"1F",X"85",X"2F",X"68",X"4A",X"29",X"03",X"A8",X"BE",X"62",X"A6",
		X"BD",X"66",X"A6",X"85",X"17",X"BD",X"67",X"A6",X"85",X"18",X"BD",X"68",X"A6",X"85",X"19",X"60",
		X"03",X"05",X"00",X"03",X"06",X"09",X"00",X"50",X"01",X"00",X"00",X"02",X"00",X"50",X"02",X"00",
		X"00",X"03",X"85",X"EF",X"EA",X"AA",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"10",X"FB",X"58",X"EA",
		X"EA",X"EA",X"78",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"30",X"FB",X"CA",X"D0",X"EB",X"60",X"85",
		X"EF",X"EA",X"A5",X"D0",X"D0",X"40",X"A5",X"3E",X"29",X"DF",X"D0",X"3A",X"A5",X"49",X"38",X"E9",
		X"01",X"85",X"49",X"B0",X"05",X"E6",X"4C",X"85",X"EF",X"EA",X"E6",X"7F",X"E6",X"91",X"EE",X"04",
		X"02",X"EE",X"24",X"02",X"EE",X"44",X"02",X"EE",X"64",X"02",X"EE",X"84",X"02",X"E6",X"EA",X"A5",
		X"4A",X"38",X"E9",X"01",X"85",X"4A",X"A5",X"4B",X"E9",X"00",X"85",X"4B",X"E6",X"48",X"A9",X"00",
		X"20",X"DE",X"D2",X"85",X"EF",X"EA",X"A5",X"49",X"8D",X"05",X"40",X"A6",X"4C",X"BD",X"E6",X"A6",
		X"8D",X"04",X"40",X"85",X"4D",X"60",X"13",X"12",X"11",X"10",X"17",X"16",X"15",X"14",X"1B",X"1A",
		X"19",X"18",X"1F",X"1E",X"1D",X"1C",X"85",X"EF",X"EA",X"A2",X"00",X"85",X"EF",X"EA",X"BD",X"18",
		X"A7",X"38",X"E5",X"4A",X"BD",X"19",X"A7",X"E5",X"4B",X"90",X"08",X"E8",X"E8",X"4C",X"FE",X"A6",
		X"85",X"EF",X"EA",X"8A",X"4A",X"85",X"4E",X"28",X"38",X"02",X"98",X"01",X"20",X"01",X"00",X"00",
		X"85",X"EF",X"EA",X"C6",X"D0",X"10",X"0A",X"A6",X"4E",X"BD",X"98",X"A7",X"85",X"D0",X"C1",X"EF",
		X"EA",X"C6",X"D1",X"10",X"07",X"A9",X"01",X"85",X"D1",X"85",X"EF",X"EA",X"C6",X"D7",X"10",X"07",
		X"A9",X"01",X"85",X"D7",X"C1",X"EF",X"6E",X"C6",X"D6",X"10",X"07",X"A9",X"20",X"85",X"D6",X"C1",
		X"EF",X"EA",X"C6",X"D4",X"10",X"07",X"A9",X"00",X"85",X"D4",X"85",X"EF",X"6E",X"C6",X"D5",X"10",
		X"07",X"A9",X"03",X"85",X"D5",X"C1",X"EF",X"6E",X"C6",X"D8",X"10",X"07",X"A9",X"04",X"85",X"D8",
		X"85",X"EF",X"EA",X"C6",X"D9",X"10",X"07",X"A9",X"04",X"85",X"D9",X"85",X"EF",X"6E",X"A5",X"DA",
		X"38",X"E9",X"01",X"B0",X"05",X"A9",X"00",X"85",X"EF",X"EA",X"85",X"DA",X"E2",X"ED",X"10",X"07",
		X"A9",X"01",X"85",X"ED",X"C1",X"EF",X"6E",X"60",X"06",X"05",X"04",X"03",X"85",X"EF",X"6E",X"A9",
		X"80",X"85",X"7B",X"85",X"83",X"C9",X"40",X"29",X"FC",X"08",X"A5",X"40",X"29",X"03",X"28",X"F0",
		X"06",X"18",X"69",X"04",X"85",X"EF",X"6E",X"0A",X"A8",X"B9",X"D1",X"A7",X"85",X"7E",X"5D",X"D2",
		X"A7",X"85",X"7F",X"85",X"EF",X"6E",X"A9",X"08",X"85",X"A9",X"A9",X"FF",X"85",X"B9",X"C1",X"BB",
		X"60",X"60",X"B0",X"B0",X"C0",X"40",X"D0",X"80",X"D0",X"A0",X"D0",X"A0",X"D0",X"20",X"D0",X"80",
		X"D0",X"85",X"EF",X"EA",X"4C",X"90",X"A8",X"85",X"EF",X"EA",X"A5",X"9D",X"F0",X"F6",X"A5",X"D1",
		X"D0",X"F2",X"A5",X"7B",X"29",X"08",X"F0",X"06",X"4C",X"C7",X"AB",X"85",X"EF",X"6E",X"A5",X"7B",
		X"29",X"04",X"F0",X"06",X"4C",X"B3",X"A8",X"85",X"EF",X"EA",X"A5",X"7B",X"29",X"BF",X"85",X"7B",
		X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"7B",X"95",X"5B",X"CA",X"10",X"F9",X"A5",X"8A",X"D0",X"06",
		X"20",X"90",X"AA",X"85",X"EF",X"EA",X"A5",X"5B",X"10",X"66",X"20",X"BA",X"B1",X"20",X"E1",X"CA",
		X"20",X"07",X"B3",X"20",X"B0",X"AF",X"20",X"3D",X"CC",X"20",X"E4",X"AD",X"85",X"EF",X"EA",X"A5",
		X"61",X"C9",X"46",X"90",X"4B",X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"5B",X"95",X"7B",X"CA",X"10",
		X"F9",X"A5",X"7B",X"29",X"04",X"F0",X"09",X"A5",X"7B",X"09",X"40",X"85",X"7B",X"85",X"EF",X"EA",
		X"20",X"E0",X"AC",X"A5",X"10",X"F0",X"07",X"A5",X"8A",X"D0",X"10",X"85",X"EF",X"EA",X"A5",X"81",
		X"C9",X"F0",X"B0",X"2A",X"C9",X"46",X"90",X"1C",X"85",X"EF",X"EA",X"A5",X"80",X"C9",X"10",X"90",
		X"13",X"C9",X"F0",X"B0",X"0F",X"A5",X"81",X"85",X"7F",X"A5",X"80",X"85",X"7E",X"85",X"EF",X"EA",
		X"60",X"85",X"EF",X"EA",X"A5",X"7B",X"29",X"F8",X"85",X"7B",X"60",X"85",X"EF",X"EA",X"A5",X"7B",
		X"29",X"7F",X"09",X"10",X"85",X"7B",X"20",X"10",X"AF",X"A5",X"3E",X"09",X"40",X"85",X"3E",X"60",
		X"85",X"EF",X"EA",X"A9",X"00",X"85",X"D1",X"A5",X"8B",X"29",X"82",X"85",X"8B",X"A9",X"00",X"85",
		X"8C",X"A5",X"B6",X"D0",X"5C",X"A9",X"00",X"8D",X"3C",X"07",X"A9",X"04",X"85",X"A0",X"A9",X"04",
		X"85",X"A4",X"85",X"A1",X"A9",X"05",X"85",X"B6",X"A9",X"02",X"20",X"86",X"D3",X"A0",X"7E",X"20",
		X"E9",X"A8",X"A5",X"BA",X"85",X"B8",X"60",X"85",X"EF",X"EA",X"A9",X"30",X"85",X"09",X"A9",X"F8",
		X"85",X"0A",X"98",X"48",X"20",X"AA",X"D0",X"68",X"A8",X"A6",X"CC",X"85",X"EF",X"EA",X"CA",X"CA",
		X"CA",X"CA",X"30",X"19",X"BD",X"01",X"04",X"D9",X"00",X"00",X"D0",X"F2",X"BD",X"02",X"04",X"D9",
		X"01",X"00",X"D0",X"EA",X"BD",X"00",X"04",X"85",X"BA",X"60",X"85",X"EF",X"6E",X"00",X"C1",X"EF",
		X"EA",X"C9",X"05",X"D0",X"1F",X"A5",X"A3",X"C9",X"03",X"D0",X"15",X"A5",X"A2",X"C9",X"01",X"30",
		X"0F",X"C6",X"B6",X"A5",X"9F",X"29",X"FE",X"85",X"9F",X"A9",X"00",X"85",X"B7",X"C1",X"EF",X"6E",
		X"60",X"85",X"EF",X"EA",X"C9",X"04",X"D0",X"09",X"C6",X"B6",X"85",X"EF",X"6E",X"60",X"85",X"EF",
		X"EA",X"C9",X"03",X"F0",X"06",X"4C",X"19",X"AA",X"85",X"EF",X"EA",X"A5",X"B8",X"85",X"BA",X"E1",
		X"B9",X"D0",X"03",X"4C",X"F1",X"A9",X"A9",X"FF",X"85",X"08",X"A9",X"48",X"85",X"09",X"4D",X"D8",
		X"85",X"0A",X"20",X"AA",X"D0",X"A6",X"CC",X"F0",X"78",X"20",X"9D",X"CE",X"A5",X"1A",X"65",X"7F",
		X"29",X"0F",X"A8",X"B9",X"7E",X"AA",X"85",X"57",X"85",X"EF",X"EA",X"18",X"65",X"BA",X"85",X"B8",
		X"85",X"EF",X"EA",X"A4",X"CC",X"85",X"EF",X"6E",X"88",X"88",X"88",X"88",X"30",X"29",X"B9",X"00",
		X"04",X"C5",X"B8",X"D0",X"F3",X"85",X"EF",X"6E",X"85",X"B9",X"B9",X"01",X"04",X"85",X"7E",X"C1",
		X"E9",X"B9",X"02",X"04",X"85",X"7F",X"C1",X"EA",X"B9",X"03",X"04",X"85",X"7D",X"81",X"E8",X"85",
		X"E8",X"C6",X"B6",X"60",X"85",X"EF",X"6E",X"86",X"07",X"A6",X"08",X"30",X"16",X"E6",X"08",X"DD",
		X"DB",X"A9",X"08",X"A6",X"07",X"28",X"F0",X"19",X"4C",X"8B",X"A9",X"FF",X"03",X"04",X"05",X"00",
		X"85",X"EF",X"EA",X"A5",X"57",X"49",X"03",X"E6",X"08",X"A6",X"07",X"4C",X"8B",X"A9",X"85",X"EF",
		X"EA",X"A9",X"00",X"85",X"09",X"4D",X"FF",X"85",X"0A",X"20",X"AA",X"D0",X"A4",X"CC",X"85",X"EF",
		X"EA",X"88",X"88",X"88",X"88",X"10",X"06",X"4C",X"1D",X"A9",X"85",X"EF",X"EA",X"B9",X"00",X"04",
		X"C5",X"BA",X"D0",X"ED",X"F0",X"92",X"85",X"EF",X"EA",X"C9",X"02",X"D0",X"27",X"A9",X"08",X"85",
		X"A0",X"A9",X"04",X"85",X"A4",X"A5",X"7D",X"C9",X"01",X"F0",X"07",X"A9",X"01",X"10",X"08",X"85",
		X"EF",X"EA",X"A9",X"03",X"85",X"EF",X"EA",X"85",X"9F",X"C6",X"B6",X"A9",X"03",X"20",X"86",X"D3",
		X"60",X"85",X"EF",X"EA",X"C9",X"01",X"D0",X"35",X"A5",X"A3",X"C9",X"03",X"30",X"2B",X"A5",X"A2",
		X"C9",X"01",X"30",X"25",X"A9",X"02",X"85",X"A0",X"A9",X"03",X"85",X"8A",X"A5",X"7B",X"29",X"FB",
		X"85",X"7B",X"A9",X"80",X"05",X"E8",X"85",X"E8",X"C6",X"B6",X"A9",X"30",X"85",X"D7",X"A9",X"40",
		X"85",X"D0",X"A9",X"30",X"85",X"ED",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"00",X"01",X"02",
		X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"01",X"85",X"EF",
		X"EA",X"A5",X"10",X"F0",X"53",X"A6",X"12",X"AD",X"03",X"40",X"29",X"40",X"D0",X"05",X"A2",X"00",
		X"85",X"EF",X"EA",X"BD",X"00",X"40",X"49",X"FF",X"29",X"0F",X"AA",X"BD",X"D5",X"AA",X"48",X"30",
		X"20",X"A6",X"63",X"30",X"0D",X"C5",X"5C",X"F0",X"18",X"49",X"02",X"C5",X"5C",X"F0",X"12",X"85",
		X"EF",X"EA",X"A5",X"5B",X"09",X"01",X"85",X"5B",X"A5",X"63",X"29",X"7F",X"85",X"63",X"85",X"EF",
		X"EA",X"68",X"85",X"5D",X"60",X"FF",X"00",X"02",X"FF",X"03",X"00",X"03",X"FF",X"01",X"01",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"85",X"EF",X"EA",X"A5",X"6A",X"D0",X"3D",X"A5",X"40",X"29",X"03",
		X"0A",X"AA",X"BD",X"2A",X"AB",X"85",X"01",X"BD",X"2B",X"AB",X"85",X"02",X"A4",X"E7",X"B1",X"01",
		X"48",X"C9",X"FF",X"F0",X"16",X"10",X"0B",X"A2",X"A9",X"86",X"8B",X"68",X"29",X"03",X"48",X"C1",
		X"EF",X"EA",X"A5",X"5B",X"09",X"01",X"85",X"5B",X"85",X"EF",X"EA",X"68",X"85",X"5D",X"64",X"B1",
		X"01",X"C8",X"85",X"6A",X"C0",X"E7",X"C1",X"EF",X"EA",X"60",X"32",X"AB",X"64",X"AB",X"86",X"AB",
		X"A6",X"AB",X"00",X"0E",X"03",X"07",X"02",X"07",X"03",X"07",X"02",X"07",X"03",X"0E",X"00",X"07",
		X"01",X"07",X"00",X"16",X"82",X"07",X"03",X"07",X"00",X"07",X"01",X"04",X"02",X"0E",X"03",X"0E",
		X"00",X"07",X"01",X"0E",X"02",X"07",X"01",X"07",X"02",X"07",X"01",X"07",X"02",X"07",X"03",X"0E",
		X"83",X"00",X"FF",X"7F",X"00",X"07",X"02",X"07",X"03",X"16",X"02",X"01",X"82",X"07",X"03",X"0E",
		X"81",X"04",X"02",X"07",X"03",X"07",X"02",X"07",X"03",X"07",X"02",X"07",X"03",X"16",X"02",X"0E",
		X"01",X"14",X"00",X"07",X"FF",X"7F",X"00",X"07",X"01",X"07",X"03",X"07",X"00",X"07",X"01",X"07",
		X"00",X"07",X"01",X"07",X"00",X"07",X"01",X"07",X"00",X"07",X"01",X"07",X"00",X"07",X"03",X"07",
		X"00",X"07",X"01",X"07",X"FF",X"7F",X"00",X"07",X"03",X"07",X"FF",X"7F",X"05",X"05",X"05",X"FF",
		X"05",X"05",X"05",X"FF",X"02",X"FE",X"02",X"00",X"02",X"02",X"00",X"03",X"FE",X"FE",X"FE",X"00",
		X"FE",X"02",X"00",X"03",X"85",X"EF",X"6E",X"A5",X"C7",X"30",X"08",X"A9",X"40",X"85",X"C7",X"28",
		X"85",X"EF",X"EA",X"AD",X"D0",X"02",X"F0",X"0C",X"A9",X"10",X"0D",X"D0",X"02",X"8D",X"D0",X"02",
		X"60",X"85",X"EF",X"EA",X"A5",X"BB",X"10",X"32",X"A9",X"0E",X"20",X"86",X"D3",X"A5",X"7E",X"30",
		X"0D",X"A9",X"00",X"85",X"BB",X"4D",X"04",X"85",X"BC",X"10",X"0E",X"85",X"EF",X"6E",X"A9",X"04",
		X"85",X"BB",X"A9",X"08",X"85",X"BC",X"85",X"EF",X"EA",X"A0",X"07",X"85",X"EF",X"EA",X"B9",X"AC",
		X"AB",X"99",X"BD",X"00",X"88",X"10",X"F7",X"85",X"EF",X"EA",X"A5",X"BB",X"AA",X"D6",X"BD",X"D0",
		X"0B",X"E6",X"BB",X"A5",X"BB",X"C5",X"BC",X"F0",X"3A",X"85",X"EF",X"EA",X"A9",X"81",X"85",X"9F",
		X"8A",X"0A",X"AA",X"A9",X"0C",X"85",X"A0",X"A9",X"02",X"85",X"A4",X"A5",X"7E",X"18",X"7D",X"B4",
		X"AB",X"85",X"7E",X"A5",X"7F",X"18",X"7D",X"B5",X"AB",X"85",X"7F",X"C9",X"F0",X"90",X"10",X"A9",
		X"00",X"85",X"7B",X"A9",X"01",X"85",X"B2",X"A9",X"0D",X"20",X"86",X"D3",X"85",X"EF",X"EA",X"60",
		X"85",X"EF",X"EA",X"00",X"85",X"EF",X"EA",X"A0",X"0C",X"85",X"EF",X"EA",X"B9",X"A0",X"02",X"10",
		X"4E",X"48",X"C9",X"B8",X"D0",X"23",X"98",X"48",X"B9",X"A1",X"02",X"85",X"01",X"B9",X"A2",X"02",
		X"85",X"02",X"B9",X"A3",X"02",X"0A",X"AA",X"BD",X"C6",X"AC",X"A0",X"00",X"91",X"01",X"BD",X"C7",
		X"AC",X"C8",X"91",X"01",X"68",X"A8",X"85",X"EF",X"EA",X"68",X"C9",X"80",X"D0",X"19",X"B9",X"A1",
		X"02",X"85",X"01",X"B9",X"A2",X"02",X"85",X"02",X"98",X"48",X"A0",X"00",X"98",X"91",X"01",X"C8",
		X"91",X"01",X"68",X"A8",X"85",X"EF",X"EA",X"98",X"AA",X"DE",X"A0",X"02",X"85",X"EF",X"EA",X"88",
		X"88",X"88",X"88",X"10",X"A7",X"60",X"C4",X"C1",X"C7",X"C1",X"C5",X"C1",X"C9",X"C1",X"C6",X"C1",
		X"CB",X"C1",X"85",X"EF",X"EA",X"4C",X"A1",X"AD",X"85",X"EF",X"EA",X"4C",X"AD",X"AD",X"85",X"EF",
		X"EA",X"A5",X"7E",X"85",X"01",X"A5",X"7F",X"85",X"02",X"20",X"C8",X"C5",X"A0",X"00",X"B1",X"01",
		X"C9",X"40",X"90",X"E7",X"C9",X"C0",X"B0",X"E3",X"A4",X"59",X"85",X"EF",X"EA",X"B9",X"00",X"03",
		X"29",X"C0",X"D0",X"D1",X"B9",X"04",X"03",X"18",X"69",X"03",X"38",X"E5",X"7F",X"B0",X"07",X"49",
		X"FF",X"69",X"01",X"85",X"EF",X"6E",X"C9",X"03",X"B0",X"BB",X"B9",X"01",X"03",X"18",X"69",X"08",
		X"38",X"E5",X"7E",X"B0",X"07",X"49",X"FF",X"69",X"01",X"85",X"EF",X"EA",X"C9",X"06",X"B0",X"71",
		X"B9",X"00",X"03",X"09",X"40",X"99",X"00",X"03",X"29",X"07",X"48",X"B9",X"01",X"03",X"85",X"01",
		X"B9",X"04",X"03",X"85",X"02",X"08",X"C8",X"C5",X"A2",X"0C",X"85",X"EF",X"6E",X"BD",X"A0",X"02",
		X"10",X"0B",X"CA",X"CA",X"CA",X"CA",X"10",X"F5",X"68",X"60",X"85",X"EF",X"6E",X"68",X"85",X"0A",
		X"C9",X"04",X"D0",X"05",X"A9",X"02",X"85",X"EF",X"EA",X"C9",X"03",X"F0",X"4A",X"48",X"4D",X"01",
		X"20",X"86",X"D3",X"68",X"86",X"04",X"06",X"A6",X"7C",X"1D",X"D2",X"AD",X"48",X"4E",X"BD",X"DC",
		X"AD",X"20",X"DE",X"D2",X"68",X"AA",X"BD",X"D6",X"AD",X"A6",X"04",X"9D",X"A3",X"02",X"4D",X"C0",
		X"9D",X"A0",X"02",X"A5",X"01",X"9D",X"A1",X"02",X"A5",X"02",X"9D",X"A2",X"02",X"28",X"85",X"EF",
		X"EA",X"C8",X"C8",X"C8",X"C8",X"C8",X"C4",X"5A",X"D0",X"07",X"85",X"EF",X"6E",X"60",X"85",X"EF",
		X"EA",X"4C",X"FD",X"AC",X"85",X"EF",X"6E",X"A5",X"7B",X"09",X"08",X"85",X"7B",X"08",X"10",X"AF",
		X"A9",X"40",X"05",X"3E",X"85",X"3E",X"C9",X"E8",X"09",X"40",X"85",X"E8",X"4D",X"0C",X"20",X"86",
		X"D3",X"60",X"01",X"00",X"00",X"01",X"01",X"00",X"03",X"02",X"05",X"04",X"05",X"03",X"06",X"07",
		X"09",X"04",X"85",X"EF",X"6E",X"A5",X"5B",X"29",X"02",X"F0",X"11",X"A5",X"5F",X"85",X"E5",X"C9",
		X"3E",X"09",X"82",X"85",X"3E",X"4D",X"80",X"85",X"C7",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",
		X"A5",X"B2",X"F0",X"45",X"29",X"04",X"D0",X"52",X"A5",X"B2",X"29",X"01",X"D0",X"3F",X"A5",X"7E",
		X"18",X"69",X"08",X"49",X"FF",X"8D",X"3A",X"07",X"38",X"E9",X"10",X"8D",X"3E",X"07",X"18",X"69",
		X"20",X"8D",X"36",X"07",X"A9",X"04",X"85",X"BD",X"85",X"BE",X"85",X"BF",X"A9",X"20",X"85",X"C0",
		X"A9",X"00",X"85",X"C4",X"85",X"DF",X"A9",X"D8",X"8D",X"3B",X"07",X"8D",X"37",X"07",X"8D",X"3F",
		X"07",X"85",X"EF",X"EA",X"06",X"B2",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"20",X"45",X"CD",
		X"A9",X"00",X"85",X"9F",X"4C",X"44",X"AE",X"85",X"EF",X"EA",X"A6",X"C4",X"D6",X"BD",X"D0",X"0F",
		X"E8",X"86",X"C4",X"E0",X"04",X"D0",X"08",X"A9",X"80",X"85",X"1D",X"60",X"85",X"EF",X"EA",X"8A",
		X"0A",X"A8",X"B9",X"97",X"AE",X"8D",X"35",X"07",X"B9",X"98",X"AE",X"8D",X"34",X"07",X"B9",X"9F",
		X"AE",X"8D",X"39",X"07",X"B9",X"A0",X"AE",X"8D",X"38",X"07",X"B9",X"A7",X"AE",X"8D",X"3D",X"07",
		X"B9",X"A8",X"AE",X"8D",X"3C",X"07",X"60",X"17",X"01",X"18",X"01",X"19",X"01",X"00",X"00",X"14",
		X"01",X"15",X"01",X"16",X"01",X"00",X"00",X"17",X"03",X"18",X"03",X"19",X"03",X"00",X"00",X"85",
		X"EF",X"EA",X"A5",X"7B",X"29",X"10",X"F0",X"28",X"A5",X"B1",X"D0",X"28",X"A9",X"0D",X"20",X"86",
		X"D3",X"A9",X"40",X"85",X"C7",X"20",X"10",X"AF",X"A9",X"05",X"85",X"9F",X"A9",X"0C",X"85",X"A0",
		X"A9",X"02",X"85",X"A4",X"A9",X"10",X"85",X"A1",X"20",X"08",X"C9",X"E6",X"B1",X"85",X"EF",X"EA",
		X"60",X"85",X"EF",X"EA",X"A6",X"A3",X"BD",X"0C",X"AF",X"85",X"7F",X"A5",X"B1",X"C9",X"20",X"90",
		X"0C",X"E6",X"7E",X"A5",X"7E",X"C9",X"FC",X"B0",X"0A",X"60",X"85",X"EF",X"EA",X"E6",X"B1",X"60",
		X"85",X"EF",X"EA",X"A9",X"80",X"85",X"1D",X"4D",X"00",X"85",X"DF",X"60",X"F0",X"F4",X"85",X"EF",
		X"EA",X"A5",X"7E",X"85",X"45",X"C9",X"7F",X"85",X"46",X"A5",X"7C",X"85",X"47",X"28",X"85",X"EF",
		X"EA",X"A5",X"9F",X"D0",X"08",X"8D",X"20",X"07",X"F0",X"4A",X"85",X"EF",X"6E",X"A5",X"A5",X"C5",
		X"A0",X"D0",X"09",X"A5",X"A6",X"C5",X"9F",X"F0",X"0E",X"85",X"EF",X"EA",X"A5",X"A1",X"85",X"A2",
		X"A9",X"00",X"85",X"A3",X"C1",X"EF",X"6E",X"C6",X"A2",X"D0",X"13",X"A5",X"A1",X"85",X"A2",X"EA",
		X"A3",X"A5",X"A3",X"C5",X"A4",X"D0",X"07",X"A9",X"00",X"85",X"A3",X"85",X"EF",X"6E",X"A5",X"A3",
		X"18",X"65",X"A0",X"8D",X"21",X"07",X"C9",X"9F",X"8D",X"20",X"07",X"85",X"A6",X"C9",X"A0",X"85",
		X"A5",X"85",X"EF",X"EA",X"A2",X"00",X"A5",X"7C",X"29",X"01",X"F0",X"04",X"E8",X"85",X"EF",X"6E",
		X"AD",X"03",X"40",X"29",X"40",X"F0",X"09",X"A5",X"12",X"F0",X"05",X"E8",X"E8",X"85",X"EF",X"6E",
		X"A5",X"7E",X"18",X"7D",X"AA",X"AF",X"18",X"69",X"08",X"49",X"FF",X"8D",X"22",X"07",X"C9",X"7F",
		X"38",X"E9",X"0E",X"8D",X"23",X"07",X"C1",X"EF",X"EA",X"60",X"00",X"02",X"FE",X"00",X"85",X"EF",
		X"EA",X"A5",X"8B",X"29",X"01",X"F0",X"07",X"A9",X"02",X"85",X"67",X"85",X"EF",X"6E",X"60",X"85",
		X"EF",X"EA",X"A5",X"8B",X"29",X"02",X"D0",X"08",X"A9",X"00",X"85",X"A7",X"28",X"85",X"EF",X"6E",
		X"A9",X"01",X"85",X"A7",X"28",X"85",X"EF",X"6E",X"A5",X"8B",X"29",X"20",X"F0",X"7A",X"A9",X"80",
		X"85",X"8D",X"A5",X"7C",X"4A",X"90",X"07",X"A9",X"01",X"10",X"08",X"85",X"EF",X"6E",X"A9",X"02",
		X"85",X"EF",X"EA",X"85",X"8F",X"C9",X"7E",X"85",X"90",X"85",X"92",X"A5",X"7F",X"85",X"91",X"C1",
		X"4C",X"54",X"A0",X"4C",X"09",X"A0",X"85",X"EF",X"EA",X"78",X"D8",X"AD",X"03",X"40",X"29",X"20",
		X"D0",X"06",X"4C",X"03",X"90",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"00",X"A2",X"FF",X"9A",X"A9",
		X"00",X"8D",X"00",X"40",X"8D",X"02",X"40",X"8D",X"03",X"40",X"8D",X"04",X"40",X"8D",X"05",X"40",
		X"8D",X"00",X"08",X"20",X"80",X"A4",X"A2",X"00",X"20",X"D7",X"A4",X"20",X"FA",X"A4",X"20",X"6E",
		X"A4",X"20",X"91",X"CE",X"AD",X"10",X"07",X"85",X"16",X"AD",X"11",X"07",X"85",X"15",X"4C",X"B0",
		X"A1",X"85",X"EF",X"EA",X"48",X"8A",X"48",X"98",X"48",X"AD",X"03",X"40",X"29",X"20",X"D0",X"06",
		X"4C",X"00",X"90",X"85",X"EF",X"EA",X"A5",X"00",X"F0",X"06",X"4C",X"00",X"90",X"85",X"EF",X"EA",
		X"A9",X"00",X"85",X"00",X"D8",X"A5",X"0B",X"F0",X"73",X"AD",X"04",X"40",X"49",X"FF",X"29",X"E0",
		X"85",X"0D",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"20",X"50",X"A1",X"AD",X"02",X"40",X"29",X"C0",
		X"F0",X"5A",X"85",X"0C",X"20",X"50",X"A1",X"AD",X"02",X"40",X"25",X"0C",X"F0",X"4E",X"20",X"50",
		X"A1",X"AD",X"02",X"40",X"25",X"0C",X"F0",X"44",X"20",X"50",X"A1",X"AD",X"02",X"40",X"25",X"0C",
		X"F0",X"3A",X"E6",X"0F",X"A9",X"10",X"8D",X"03",X"40",X"A5",X"0D",X"C9",X"80",X"F0",X"39",X"A2",
		X"00",X"AD",X"03",X"40",X"49",X"FF",X"29",X"0F",X"06",X"0C",X"90",X"05",X"4A",X"4A",X"85",X"EF",
		X"EA",X"29",X"03",X"F0",X"51",X"E8",X"C9",X"01",X"F0",X"4C",X"E8",X"C9",X"02",X"F0",X"3C",X"E8",
		X"85",X"EF",X"EA",X"A5",X"0F",X"C9",X"02",X"B0",X"2A",X"85",X"EF",X"EA",X"8D",X"00",X"40",X"68",
		X"A8",X"68",X"AA",X"68",X"40",X"85",X"EF",X"EA",X"A2",X"05",X"A5",X"0C",X"C9",X"40",X"F0",X"26",
		X"E8",X"C9",X"80",X"F0",X"21",X"E8",X"C9",X"C0",X"F0",X"D9",X"4C",X"EC",X"A0",X"85",X"EF",X"6E",
		X"85",X"EF",X"EA",X"C6",X"0F",X"A4",X"26",X"A1",X"85",X"EF",X"EA",X"A5",X"0D",X"C9",X"60",X"D0",
		X"05",X"A2",X"04",X"85",X"EF",X"6E",X"A5",X"0E",X"F8",X"18",X"7D",X"5F",X"A1",X"D9",X"67",X"A1",
		X"90",X"06",X"B9",X"67",X"A1",X"85",X"EF",X"6E",X"85",X"0E",X"D8",X"C6",X"0F",X"C9",X"10",X"D0",
		X"AB",X"8D",X"00",X"40",X"4D",X"01",X"85",X"10",X"A2",X"FF",X"9A",X"4C",X"72",X"A1",X"85",X"EF",
		X"EA",X"A2",X"E7",X"85",X"EF",X"6E",X"A5",X"FF",X"A5",X"FF",X"EA",X"CA",X"D0",X"F8",X"60",X"01",
		X"02",X"03",X"01",X"06",X"08",X"03",X"01",X"09",X"09",X"16",X"16",X"16",X"09",X"09",X"09",X"85",
		X"EF",X"EA",X"20",X"B8",X"A5",X"20",X"A0",X"A4",X"20",X"19",X"C9",X"20",X"E6",X"DA",X"85",X"EF",
		X"EA",X"20",X"98",X"D3",X"20",X"14",X"DB",X"A9",X"00",X"85",X"11",X"AD",X"02",X"40",X"49",X"FF",
		X"29",X"03",X"F0",X"ED",X"C9",X"01",X"F0",X"12",X"C9",X"02",X"D0",X"E5",X"A5",X"0E",X"C9",X"02",
		X"90",X"DF",X"20",X"2A",X"A6",X"E6",X"11",X"C1",X"EF",X"EA",X"20",X"2A",X"A6",X"85",X"EF",X"6E",
		X"E6",X"11",X"85",X"EF",X"6E",X"A2",X"1D",X"20",X"73",X"A4",X"A2",X"01",X"20",X"D7",X"A4",X"A9",
		X"00",X"8D",X"04",X"40",X"08",X"80",X"A4",X"20",X"08",X"C9",X"20",X"AD",X"CE",X"20",X"C4",X"CE",
		X"20",X"E0",X"CE",X"20",X"E4",X"D3",X"85",X"EF",X"EA",X"20",X"37",X"A6",X"20",X"29",X"D4",X"20",
		X"BA",X"D4",X"20",X"29",X"D0",X"A9",X"01",X"85",X"0B",X"A9",X"00",X"85",X"12",X"08",X"A0",X"A4",
		X"A9",X"FF",X"85",X"20",X"C1",X"30",X"4D",X"00",X"85",X"21",X"85",X"31",X"4D",X"80",X"85",X"1E",
		X"85",X"2E",X"A5",X"10",X"D0",X"0C",X"20",X"B8",X"A5",X"20",X"7B",X"D8",X"20",X"18",X"D9",X"85",
		X"EF",X"EA",X"C6",X"1F",X"C6",X"2F",X"85",X"EF",X"EA",X"20",X"C1",X"A5",X"A2",X"80",X"20",X"C9",
		X"CE",X"20",X"75",X"D4",X"20",X"70",X"C1",X"A9",X"00",X"8D",X"04",X"40",X"A5",X"12",X"8D",X"02",
		X"40",X"A9",X"A2",X"48",X"A9",X"46",X"48",X"A5",X"3E",X"10",X"06",X"4C",X"46",X"A3",X"85",X"EF",
		X"EA",X"4C",X"86",X"A3",X"85",X"EF",X"EA",X"20",X"FB",X"D3",X"20",X"F1",X"A5",X"20",X"29",X"D4",
		X"20",X"59",X"DB",X"20",X"5A",X"A5",X"20",X"D5",X"A6",X"A9",X"20",X"20",X"74",X"A6",X"20",X"A0",
		X"A4",X"20",X"45",X"CD",X"85",X"EF",X"EA",X"20",X"4F",X"A4",X"20",X"F8",X"A6",X"20",X"22",X"A7",
		X"20",X"97",X"C6",X"20",X"25",X"C4",X"20",X"9D",X"CE",X"20",X"E9",X"A7",X"20",X"B1",X"AE",X"20",
		X"FF",X"AD",X"20",X"97",X"B2",X"20",X"8D",X"BE",X"20",X"65",X"B3",X"20",X"20",X"AF",X"20",X"B7",
		X"B2",X"20",X"66",X"AC",X"20",X"F8",X"CE",X"20",X"35",X"CF",X"20",X"22",X"CA",X"20",X"17",X"D3",
		X"20",X"45",X"D3",X"20",X"6D",X"D3",X"20",X"5E",X"CD",X"A5",X"10",X"F0",X"09",X"20",X"33",X"D0",
		X"20",X"29",X"D0",X"85",X"EF",X"EA",X"33",X"1D",X"10",X"AD",X"A9",X"00",X"20",X"86",X"D3",X"20",
		X"A0",X"A4",X"20",X"B8",X"A5",X"24",X"1D",X"70",X"05",X"C6",X"3F",X"85",X"EF",X"EA",X"20",X"D8",
		X"A5",X"20",X"04",X"A6",X"24",X"1D",X"50",X"06",X"4C",X"19",X"A2",X"85",X"EF",X"EA",X"A5",X"10",
		X"F0",X"46",X"A5",X"3F",X"30",X"1A",X"A5",X"11",X"C9",X"02",X"B0",X"06",X"4C",X"19",X"A2",X"85",
		X"EF",X"EA",X"E6",X"12",X"A5",X"12",X"29",X"01",X"85",X"12",X"4C",X"19",X"A2",X"85",X"EF",X"EA",
		X"20",X"12",X"D4",X"A9",X"FF",X"20",X"74",X"A6",X"20",X"6D",X"DB",X"C6",X"11",X"70",X"E3",X"A9",
		X"00",X"8D",X"02",X"40",X"C1",X"12",X"C9",X"0E",X"D0",X"08",X"85",X"10",X"A4",X"B0",X"A1",X"85",
		X"EF",X"EA",X"4C",X"72",X"A1",X"85",X"EF",X"6E",X"E6",X"1C",X"A5",X"1C",X"C9",X"04",X"90",X"0A",
		X"A9",X"00",X"85",X"1C",X"A4",X"00",X"A3",X"85",X"EF",X"EA",X"A9",X"80",X"85",X"1E",X"EA",X"1F",
		X"4C",X"19",X"A2",X"85",X"EF",X"6E",X"E6",X"40",X"F8",X"A5",X"41",X"38",X"69",X"00",X"85",X"41",
		X"D8",X"A2",X"4F",X"20",X"73",X"A4",X"20",X"81",X"C1",X"A9",X"00",X"85",X"59",X"C1",X"5A",X"C9",
		X"3E",X"29",X"20",X"09",X"01",X"85",X"3E",X"4D",X"80",X"85",X"C7",X"A9",X"00",X"85",X"1D",X"C1",
		X"EF",X"EA",X"A9",X"00",X"85",X"4C",X"4D",X"10",X"85",X"49",X"A9",X"0F",X"85",X"4A",X"4D",X"03",
		X"85",X"4B",X"60",X"85",X"EF",X"6E",X"A2",X"4F",X"20",X"73",X"A4",X"20",X"A0",X"A4",X"A9",X"42",
		X"20",X"86",X"D3",X"A5",X"3E",X"29",X"20",X"85",X"3E",X"A9",X"00",X"85",X"1D",X"C1",X"C7",X"C1",
		X"59",X"85",X"5A",X"20",X"C5",X"A7",X"A9",X"80",X"85",X"9D",X"85",X"D7",X"C9",X"46",X"38",X"E9",
		X"98",X"85",X"48",X"F0",X"07",X"90",X"24",X"B0",X"54",X"85",X"EF",X"EA",X"A5",X"45",X"85",X"7E",
		X"85",X"80",X"A5",X"46",X"85",X"7F",X"C1",X"81",X"A5",X"47",X"85",X"7C",X"C1",X"EF",X"6E",X"A9",
		X"80",X"85",X"7B",X"A9",X"00",X"85",X"48",X"28",X"85",X"EF",X"EA",X"A5",X"48",X"49",X"FF",X"38",
		X"69",X"00",X"85",X"48",X"C9",X"49",X"38",X"E5",X"48",X"85",X"49",X"B0",X"05",X"E6",X"4C",X"C1",
		X"EF",X"EA",X"A5",X"46",X"18",X"65",X"48",X"85",X"46",X"A5",X"4A",X"38",X"E5",X"48",X"85",X"4A",
		X"B0",X"05",X"C6",X"4B",X"85",X"EF",X"EA",X"4C",X"BC",X"A3",X"85",X"EF",X"EA",X"A5",X"4A",X"18",
		X"65",X"48",X"85",X"02",X"A5",X"4B",X"69",X"00",X"85",X"03",X"C9",X"03",X"90",X"0F",X"A5",X"02",
		X"C9",X"0F",X"90",X"09",X"20",X"9E",X"A7",X"4C",X"72",X"A3",X"85",X"EF",X"EA",X"A5",X"46",X"38",
		X"E5",X"48",X"85",X"46",X"A5",X"49",X"18",X"65",X"48",X"85",X"49",X"90",X"05",X"C6",X"4C",X"85",
		X"EF",X"EA",X"A5",X"02",X"85",X"4A",X"A5",X"03",X"85",X"4B",X"4C",X"BC",X"A3",X"85",X"EF",X"EA",
		X"AD",X"03",X"40",X"10",X"FB",X"20",X"88",X"A5",X"20",X"91",X"A6",X"20",X"43",X"CE",X"58",X"EA",
		X"EA",X"EA",X"78",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"30",X"FB",X"60",X"85",X"EF",X"EA",X"A2",
		X"01",X"85",X"EF",X"EA",X"A9",X"00",X"95",X"00",X"E8",X"E0",X"EE",X"90",X"F7",X"60",X"85",X"EF",
		X"EA",X"A9",X"10",X"85",X"02",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"01",X"A8",X"85",X"EF",X"EA",
		X"91",X"01",X"C8",X"D0",X"FB",X"E6",X"02",X"A5",X"02",X"C9",X"18",X"90",X"EB",X"60",X"85",X"EF",
		X"EA",X"A9",X"10",X"85",X"02",X"85",X"EF",X"EA",X"A0",X"E1",X"85",X"EF",X"EA",X"A9",X"00",X"85",
		X"01",X"85",X"EF",X"EA",X"91",X"01",X"C8",X"D0",X"05",X"E6",X"02",X"85",X"EF",X"EA",X"C0",X"A0",
		X"D0",X"F2",X"A5",X"02",X"C9",X"17",X"F0",X"0C",X"C9",X"13",X"D0",X"E1",X"E6",X"02",X"4C",X"A8",
		X"A4",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A9",X"02",X"85",X"02",X"85",X"EF",X"EA",X"A9",
		X"00",X"85",X"01",X"A8",X"85",X"EF",X"EA",X"91",X"01",X"C8",X"D0",X"FB",X"E6",X"02",X"A5",X"02",
		X"DD",X"F6",X"A4",X"90",X"EA",X"60",X"08",X"07",X"85",X"EF",X"EA",X"A2",X"07",X"85",X"EF",X"EA",
		X"BD",X"10",X"A5",X"9D",X"00",X"0C",X"DD",X"18",X"A5",X"9D",X"08",X"0C",X"66",X"10",X"F1",X"60",
		X"FF",X"38",X"C0",X"3F",X"00",X"F8",X"FF",X"07",X"F8",X"C0",X"88",X"FF",X"3F",X"75",X"F8",X"88",
		X"D0",X"C7",X"38",X"FF",X"3F",X"75",X"D0",X"38",X"CF",X"00",X"C0",X"FF",X"3F",X"75",X"CF",X"C0",
		X"78",X"F8",X"F8",X"FF",X"3F",X"75",X"78",X"F8",X"3F",X"C0",X"88",X"FF",X"38",X"72",X"3F",X"88",
		X"D0",X"C7",X"3F",X"FF",X"38",X"72",X"D0",X"3F",X"CF",X"00",X"C0",X"FF",X"38",X"72",X"CF",X"C0",
		X"F8",X"F8",X"C0",X"FF",X"38",X"72",X"F8",X"C0",X"85",X"EF",X"EA",X"A5",X"40",X"38",X"85",X"EF",
		X"EA",X"E9",X"08",X"B0",X"FC",X"69",X"08",X"AA",X"A9",X"F8",X"85",X"EF",X"6E",X"18",X"69",X"08",
		X"CA",X"10",X"FA",X"AA",X"A0",X"00",X"85",X"EF",X"EA",X"BD",X"18",X"A5",X"99",X"08",X"0C",X"6C",
		X"C8",X"C0",X"08",X"90",X"F4",X"60",X"85",X"EF",X"EA",X"A5",X"C7",X"30",X"1E",X"F0",X"1C",X"A6",
		X"B4",X"A5",X"40",X"85",X"EF",X"6E",X"38",X"E9",X"04",X"B0",X"FB",X"7D",X"B4",X"A5",X"AA",X"85",
		X"EF",X"EA",X"BD",X"AC",X"A5",X"8D",X"01",X"0C",X"85",X"EF",X"EA",X"60",X"C0",X"C7",X"F8",X"C7",
		X"00",X"F8",X"88",X"07",X"04",X"08",X"85",X"EF",X"EA",X"A9",X"FF",X"8D",X"08",X"0C",X"28",X"85",
		X"EF",X"EA",X"A4",X"12",X"BE",X"ED",X"A5",X"A0",X"0F",X"85",X"EF",X"EA",X"B5",X"00",X"99",X"3E",
		X"00",X"CA",X"88",X"10",X"F7",X"60",X"85",X"EF",X"EA",X"A4",X"12",X"BE",X"ED",X"A5",X"A0",X"0F",
		X"85",X"EF",X"EA",X"B9",X"3E",X"00",X"95",X"00",X"CA",X"88",X"10",X"F7",X"60",X"2D",X"3D",X"85",
		X"EF",X"EA",X"20",X"17",X"A6",X"85",X"EF",X"6E",X"B1",X"01",X"9D",X"00",X"03",X"64",X"E8",X"D0",
		X"F7",X"60",X"85",X"EF",X"EA",X"20",X"17",X"A6",X"85",X"EF",X"EA",X"BD",X"00",X"03",X"91",X"01",
		X"E8",X"C8",X"D0",X"F7",X"60",X"85",X"EF",X"EA",X"A6",X"12",X"BD",X"26",X"A6",X"85",X"02",X"A9",
		X"00",X"85",X"01",X"AA",X"A8",X"60",X"05",X"06",X"85",X"EF",X"EA",X"F8",X"38",X"A5",X"0E",X"E9",
		X"01",X"85",X"0E",X"D8",X"60",X"85",X"EF",X"EA",X"AD",X"04",X"40",X"49",X"FF",X"48",X"29",X"01",
		X"AA",X"BD",X"60",X"A6",X"85",X"1F",X"85",X"2F",X"68",X"4A",X"29",X"03",X"A8",X"BE",X"62",X"A6",
		X"BD",X"66",X"A6",X"85",X"17",X"BD",X"67",X"A6",X"85",X"18",X"BD",X"68",X"A6",X"85",X"19",X"60",
		X"03",X"05",X"00",X"03",X"06",X"09",X"00",X"50",X"01",X"00",X"00",X"02",X"00",X"50",X"02",X"00",
		X"00",X"03",X"85",X"EF",X"EA",X"AA",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"10",X"FB",X"58",X"EA",
		X"EA",X"EA",X"78",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"30",X"FB",X"CA",X"D0",X"EB",X"60",X"85",
		X"EF",X"EA",X"A5",X"D0",X"D0",X"40",X"A5",X"3E",X"29",X"DF",X"D0",X"3A",X"A5",X"49",X"38",X"E9",
		X"01",X"85",X"49",X"B0",X"05",X"E6",X"4C",X"85",X"EF",X"EA",X"E6",X"7F",X"E6",X"91",X"EE",X"04",
		X"02",X"EE",X"24",X"02",X"EE",X"44",X"02",X"EE",X"64",X"02",X"EE",X"84",X"02",X"E6",X"EA",X"A5",
		X"4A",X"38",X"E9",X"01",X"85",X"4A",X"A5",X"4B",X"E9",X"00",X"85",X"4B",X"E6",X"48",X"A9",X"00",
		X"20",X"DE",X"D2",X"85",X"EF",X"EA",X"A5",X"49",X"8D",X"05",X"40",X"A6",X"4C",X"BD",X"E6",X"A6",
		X"8D",X"04",X"40",X"85",X"4D",X"60",X"13",X"12",X"11",X"10",X"17",X"16",X"15",X"14",X"1B",X"1A",
		X"19",X"18",X"1F",X"1E",X"1D",X"1C",X"85",X"EF",X"EA",X"A2",X"00",X"85",X"EF",X"EA",X"BD",X"18",
		X"A7",X"38",X"E5",X"4A",X"BD",X"19",X"A7",X"E5",X"4B",X"90",X"08",X"E8",X"E8",X"4C",X"FE",X"A6",
		X"85",X"EF",X"EA",X"8A",X"4A",X"85",X"4E",X"28",X"38",X"02",X"98",X"01",X"20",X"01",X"00",X"00",
		X"85",X"EF",X"EA",X"C6",X"D0",X"10",X"0A",X"A6",X"4E",X"BD",X"98",X"A7",X"85",X"D0",X"C1",X"EF",
		X"EA",X"C6",X"D1",X"10",X"07",X"A9",X"01",X"85",X"D1",X"85",X"EF",X"EA",X"C6",X"D7",X"10",X"07",
		X"A9",X"01",X"85",X"D7",X"C1",X"EF",X"6E",X"C6",X"D6",X"10",X"07",X"A9",X"20",X"85",X"D6",X"C1",
		X"EF",X"EA",X"C6",X"D4",X"10",X"07",X"A9",X"00",X"85",X"D4",X"85",X"EF",X"6E",X"C6",X"D5",X"10",
		X"07",X"A9",X"03",X"85",X"D5",X"C1",X"EF",X"6E",X"C6",X"D8",X"10",X"07",X"A9",X"04",X"85",X"D8",
		X"85",X"EF",X"EA",X"C6",X"D9",X"10",X"07",X"A9",X"04",X"85",X"D9",X"85",X"EF",X"6E",X"A5",X"DA",
		X"38",X"E9",X"01",X"B0",X"05",X"A9",X"00",X"85",X"EF",X"EA",X"85",X"DA",X"E2",X"ED",X"10",X"07",
		X"A9",X"01",X"85",X"ED",X"C1",X"EF",X"6E",X"60",X"06",X"05",X"04",X"03",X"85",X"EF",X"6E",X"A9",
		X"80",X"85",X"7B",X"85",X"83",X"C9",X"40",X"29",X"FC",X"08",X"A5",X"40",X"29",X"03",X"28",X"F0",
		X"06",X"18",X"69",X"04",X"85",X"EF",X"6E",X"0A",X"A8",X"B9",X"D1",X"A7",X"85",X"7E",X"5D",X"D2",
		X"A7",X"85",X"7F",X"85",X"EF",X"6E",X"A9",X"08",X"85",X"A9",X"A9",X"FF",X"85",X"B9",X"C1",X"BB",
		X"60",X"60",X"B0",X"B0",X"C0",X"40",X"D0",X"80",X"D0",X"A0",X"D0",X"A0",X"D0",X"20",X"D0",X"80",
		X"D0",X"85",X"EF",X"EA",X"4C",X"90",X"A8",X"85",X"EF",X"EA",X"A5",X"9D",X"F0",X"F6",X"A5",X"D1",
		X"D0",X"F2",X"A5",X"7B",X"29",X"08",X"F0",X"06",X"4C",X"C7",X"AB",X"85",X"EF",X"6E",X"A5",X"7B",
		X"29",X"04",X"F0",X"06",X"4C",X"B3",X"A8",X"85",X"EF",X"EA",X"A5",X"7B",X"29",X"BF",X"85",X"7B",
		X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"7B",X"95",X"5B",X"CA",X"10",X"F9",X"A5",X"8A",X"D0",X"06",
		X"20",X"90",X"AA",X"85",X"EF",X"EA",X"A5",X"5B",X"10",X"66",X"20",X"BA",X"B1",X"20",X"E1",X"CA",
		X"20",X"07",X"B3",X"20",X"B0",X"AF",X"20",X"3D",X"CC",X"20",X"E4",X"AD",X"85",X"EF",X"EA",X"A5",
		X"61",X"C9",X"46",X"90",X"4B",X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"5B",X"95",X"7B",X"CA",X"10",
		X"F9",X"A5",X"7B",X"29",X"04",X"F0",X"09",X"A5",X"7B",X"09",X"40",X"85",X"7B",X"85",X"EF",X"EA",
		X"20",X"E0",X"AC",X"A5",X"10",X"F0",X"07",X"A5",X"8A",X"D0",X"10",X"85",X"EF",X"EA",X"A5",X"81",
		X"C9",X"F0",X"B0",X"2A",X"C9",X"46",X"90",X"1C",X"85",X"EF",X"EA",X"A5",X"80",X"C9",X"10",X"90",
		X"13",X"C9",X"F0",X"B0",X"0F",X"A5",X"81",X"85",X"7F",X"A5",X"80",X"85",X"7E",X"85",X"EF",X"EA",
		X"60",X"85",X"EF",X"EA",X"A5",X"7B",X"29",X"F8",X"85",X"7B",X"60",X"85",X"EF",X"EA",X"A5",X"7B",
		X"29",X"7F",X"09",X"10",X"85",X"7B",X"20",X"10",X"AF",X"A5",X"3E",X"09",X"40",X"85",X"3E",X"60",
		X"85",X"EF",X"EA",X"A9",X"00",X"85",X"D1",X"A5",X"8B",X"29",X"82",X"85",X"8B",X"A9",X"00",X"85",
		X"8C",X"A5",X"B6",X"D0",X"5C",X"A9",X"00",X"8D",X"3C",X"07",X"A9",X"04",X"85",X"A0",X"A9",X"04",
		X"85",X"A4",X"85",X"A1",X"A9",X"05",X"85",X"B6",X"A9",X"02",X"20",X"86",X"D3",X"A0",X"7E",X"20",
		X"E9",X"A8",X"A5",X"BA",X"85",X"B8",X"60",X"85",X"EF",X"EA",X"A9",X"30",X"85",X"09",X"A9",X"F8",
		X"85",X"0A",X"98",X"48",X"20",X"AA",X"D0",X"68",X"A8",X"A6",X"CC",X"85",X"EF",X"EA",X"CA",X"CA",
		X"CA",X"CA",X"30",X"19",X"BD",X"01",X"04",X"D9",X"00",X"00",X"D0",X"F2",X"BD",X"02",X"04",X"D9",
		X"01",X"00",X"D0",X"EA",X"BD",X"00",X"04",X"85",X"BA",X"60",X"85",X"EF",X"6E",X"00",X"C1",X"EF",
		X"EA",X"C9",X"05",X"D0",X"1F",X"A5",X"A3",X"C9",X"03",X"D0",X"15",X"A5",X"A2",X"C9",X"01",X"30",
		X"0F",X"C6",X"B6",X"A5",X"9F",X"29",X"FE",X"85",X"9F",X"A9",X"00",X"85",X"B7",X"C1",X"EF",X"6E",
		X"60",X"85",X"EF",X"EA",X"C9",X"04",X"D0",X"09",X"C6",X"B6",X"85",X"EF",X"6E",X"60",X"85",X"EF",
		X"EA",X"C9",X"03",X"F0",X"06",X"4C",X"19",X"AA",X"85",X"EF",X"EA",X"A5",X"B8",X"85",X"BA",X"E1",
		X"B9",X"D0",X"03",X"4C",X"F1",X"A9",X"A9",X"FF",X"85",X"08",X"A9",X"48",X"85",X"09",X"4D",X"D8",
		X"85",X"0A",X"20",X"AA",X"D0",X"A6",X"CC",X"F0",X"78",X"20",X"9D",X"CE",X"A5",X"1A",X"65",X"7F",
		X"29",X"0F",X"A8",X"B9",X"7E",X"AA",X"85",X"57",X"85",X"EF",X"EA",X"18",X"65",X"BA",X"85",X"B8",
		X"85",X"EF",X"EA",X"A4",X"CC",X"85",X"EF",X"6E",X"88",X"88",X"88",X"88",X"30",X"29",X"B9",X"00",
		X"04",X"C5",X"B8",X"D0",X"F3",X"85",X"EF",X"6E",X"85",X"B9",X"B9",X"01",X"04",X"85",X"7E",X"C1",
		X"E9",X"B9",X"02",X"04",X"85",X"7F",X"C1",X"EA",X"B9",X"03",X"04",X"85",X"7D",X"81",X"E8",X"85",
		X"E8",X"C6",X"B6",X"60",X"85",X"EF",X"6E",X"86",X"07",X"A6",X"08",X"30",X"16",X"E6",X"08",X"DD",
		X"DB",X"A9",X"08",X"A6",X"07",X"28",X"F0",X"19",X"4C",X"8B",X"A9",X"FF",X"03",X"04",X"05",X"00",
		X"85",X"EF",X"EA",X"A5",X"57",X"49",X"03",X"E6",X"08",X"A6",X"07",X"4C",X"8B",X"A9",X"85",X"EF",
		X"EA",X"A9",X"00",X"85",X"09",X"4D",X"FF",X"85",X"0A",X"20",X"AA",X"D0",X"A4",X"CC",X"85",X"EF",
		X"EA",X"88",X"88",X"88",X"88",X"10",X"06",X"4C",X"1D",X"A9",X"85",X"EF",X"EA",X"B9",X"00",X"04",
		X"C5",X"BA",X"D0",X"ED",X"F0",X"92",X"85",X"EF",X"EA",X"C9",X"02",X"D0",X"27",X"A9",X"08",X"85",
		X"A0",X"A9",X"04",X"85",X"A4",X"A5",X"7D",X"C9",X"01",X"F0",X"07",X"A9",X"01",X"10",X"08",X"85",
		X"EF",X"EA",X"A9",X"03",X"85",X"EF",X"EA",X"85",X"9F",X"C6",X"B6",X"A9",X"03",X"20",X"86",X"D3",
		X"60",X"85",X"EF",X"EA",X"C9",X"01",X"D0",X"35",X"A5",X"A3",X"C9",X"03",X"30",X"2B",X"A5",X"A2",
		X"C9",X"01",X"30",X"25",X"A9",X"02",X"85",X"A0",X"A9",X"03",X"85",X"8A",X"A5",X"7B",X"29",X"FB",
		X"85",X"7B",X"A9",X"80",X"05",X"E8",X"85",X"E8",X"C6",X"B6",X"A9",X"30",X"85",X"D7",X"A9",X"40",
		X"85",X"D0",X"A9",X"30",X"85",X"ED",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"00",X"01",X"02",
		X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"01",X"85",X"EF",
		X"EA",X"A5",X"10",X"F0",X"53",X"A6",X"12",X"AD",X"03",X"40",X"29",X"40",X"D0",X"05",X"A2",X"00",
		X"85",X"EF",X"EA",X"BD",X"00",X"40",X"49",X"FF",X"29",X"0F",X"AA",X"BD",X"D5",X"AA",X"48",X"30",
		X"20",X"A6",X"63",X"30",X"0D",X"C5",X"5C",X"F0",X"18",X"49",X"02",X"C5",X"5C",X"F0",X"12",X"85",
		X"EF",X"EA",X"A5",X"5B",X"09",X"01",X"85",X"5B",X"A5",X"63",X"29",X"7F",X"85",X"63",X"85",X"EF",
		X"EA",X"68",X"85",X"5D",X"60",X"FF",X"00",X"02",X"FF",X"03",X"00",X"03",X"FF",X"01",X"01",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"85",X"EF",X"EA",X"A5",X"6A",X"D0",X"3D",X"A5",X"40",X"29",X"03",
		X"0A",X"AA",X"BD",X"2A",X"AB",X"85",X"01",X"BD",X"2B",X"AB",X"85",X"02",X"A4",X"E7",X"B1",X"01",
		X"48",X"C9",X"FF",X"F0",X"16",X"10",X"0B",X"A2",X"A9",X"86",X"8B",X"68",X"29",X"03",X"48",X"C1",
		X"EF",X"EA",X"A5",X"5B",X"09",X"01",X"85",X"5B",X"85",X"EF",X"EA",X"68",X"85",X"5D",X"64",X"B1",
		X"01",X"C8",X"85",X"6A",X"C0",X"E7",X"C1",X"EF",X"EA",X"60",X"32",X"AB",X"64",X"AB",X"86",X"AB",
		X"A6",X"AB",X"00",X"0E",X"03",X"07",X"02",X"07",X"03",X"07",X"02",X"07",X"03",X"0E",X"00",X"07",
		X"01",X"07",X"00",X"16",X"82",X"07",X"03",X"07",X"00",X"07",X"01",X"04",X"02",X"0E",X"03",X"0E",
		X"00",X"07",X"01",X"0E",X"02",X"07",X"01",X"07",X"02",X"07",X"01",X"07",X"02",X"07",X"03",X"0E",
		X"83",X"00",X"FF",X"7F",X"00",X"07",X"02",X"07",X"03",X"16",X"02",X"01",X"82",X"07",X"03",X"0E",
		X"81",X"04",X"02",X"07",X"03",X"07",X"02",X"07",X"03",X"07",X"02",X"07",X"03",X"16",X"02",X"0E",
		X"01",X"14",X"00",X"07",X"FF",X"7F",X"00",X"07",X"01",X"07",X"03",X"07",X"00",X"07",X"01",X"07",
		X"00",X"07",X"01",X"07",X"00",X"07",X"01",X"07",X"00",X"07",X"01",X"07",X"00",X"07",X"03",X"07",
		X"00",X"07",X"01",X"07",X"FF",X"7F",X"00",X"07",X"03",X"07",X"FF",X"7F",X"05",X"05",X"05",X"FF",
		X"05",X"05",X"05",X"FF",X"02",X"FE",X"02",X"00",X"02",X"02",X"00",X"03",X"FE",X"FE",X"FE",X"00",
		X"FE",X"02",X"00",X"03",X"85",X"EF",X"6E",X"A5",X"C7",X"30",X"08",X"A9",X"40",X"85",X"C7",X"28",
		X"85",X"EF",X"EA",X"AD",X"D0",X"02",X"F0",X"0C",X"A9",X"10",X"0D",X"D0",X"02",X"8D",X"D0",X"02",
		X"60",X"85",X"EF",X"EA",X"A5",X"BB",X"10",X"32",X"A9",X"0E",X"20",X"86",X"D3",X"A5",X"7E",X"30",
		X"0D",X"A9",X"00",X"85",X"BB",X"4D",X"04",X"85",X"BC",X"10",X"0E",X"85",X"EF",X"6E",X"A9",X"04",
		X"85",X"BB",X"A9",X"08",X"85",X"BC",X"85",X"EF",X"EA",X"A0",X"07",X"85",X"EF",X"EA",X"B9",X"AC",
		X"AB",X"99",X"BD",X"00",X"88",X"10",X"F7",X"85",X"EF",X"EA",X"A5",X"BB",X"AA",X"D6",X"BD",X"D0",
		X"0B",X"E6",X"BB",X"A5",X"BB",X"C5",X"BC",X"F0",X"3A",X"85",X"EF",X"EA",X"A9",X"81",X"85",X"9F",
		X"8A",X"0A",X"AA",X"A9",X"0C",X"85",X"A0",X"A9",X"02",X"85",X"A4",X"A5",X"7E",X"18",X"7D",X"B4",
		X"AB",X"85",X"7E",X"A5",X"7F",X"18",X"7D",X"B5",X"AB",X"85",X"7F",X"C9",X"F0",X"90",X"10",X"A9",
		X"00",X"85",X"7B",X"A9",X"01",X"85",X"B2",X"A9",X"0D",X"20",X"86",X"D3",X"85",X"EF",X"EA",X"60",
		X"85",X"EF",X"EA",X"00",X"85",X"EF",X"EA",X"A0",X"0C",X"85",X"EF",X"EA",X"B9",X"A0",X"02",X"10",
		X"4E",X"48",X"C9",X"B8",X"D0",X"23",X"98",X"48",X"B9",X"A1",X"02",X"85",X"01",X"B9",X"A2",X"02",
		X"85",X"02",X"B9",X"A3",X"02",X"0A",X"AA",X"BD",X"C6",X"AC",X"A0",X"00",X"91",X"01",X"BD",X"C7",
		X"AC",X"C8",X"91",X"01",X"68",X"A8",X"85",X"EF",X"EA",X"68",X"C9",X"80",X"D0",X"19",X"B9",X"A1",
		X"02",X"85",X"01",X"B9",X"A2",X"02",X"85",X"02",X"98",X"48",X"A0",X"00",X"98",X"91",X"01",X"C8",
		X"91",X"01",X"68",X"A8",X"85",X"EF",X"EA",X"98",X"AA",X"DE",X"A0",X"02",X"85",X"EF",X"EA",X"88",
		X"88",X"88",X"88",X"10",X"A7",X"60",X"C4",X"C1",X"C7",X"C1",X"C5",X"C1",X"C9",X"C1",X"C6",X"C1",
		X"CB",X"C1",X"85",X"EF",X"EA",X"4C",X"A1",X"AD",X"85",X"EF",X"EA",X"4C",X"AD",X"AD",X"85",X"EF",
		X"EA",X"A5",X"7E",X"85",X"01",X"A5",X"7F",X"85",X"02",X"20",X"C8",X"C5",X"A0",X"00",X"B1",X"01",
		X"C9",X"40",X"90",X"E7",X"C9",X"C0",X"B0",X"E3",X"A4",X"59",X"85",X"EF",X"EA",X"B9",X"00",X"03",
		X"29",X"C0",X"D0",X"D1",X"B9",X"04",X"03",X"18",X"69",X"03",X"38",X"E5",X"7F",X"B0",X"07",X"49",
		X"FF",X"69",X"01",X"85",X"EF",X"6E",X"C9",X"03",X"B0",X"BB",X"B9",X"01",X"03",X"18",X"69",X"08",
		X"38",X"E5",X"7E",X"B0",X"07",X"49",X"FF",X"69",X"01",X"85",X"EF",X"EA",X"C9",X"06",X"B0",X"71",
		X"B9",X"00",X"03",X"09",X"40",X"99",X"00",X"03",X"29",X"07",X"48",X"B9",X"01",X"03",X"85",X"01",
		X"B9",X"04",X"03",X"85",X"02",X"08",X"C8",X"C5",X"A2",X"0C",X"85",X"EF",X"6E",X"BD",X"A0",X"02",
		X"10",X"0B",X"CA",X"CA",X"CA",X"CA",X"10",X"F5",X"68",X"60",X"85",X"EF",X"6E",X"68",X"85",X"0A",
		X"C9",X"04",X"D0",X"05",X"A9",X"02",X"85",X"EF",X"EA",X"C9",X"03",X"F0",X"4A",X"48",X"4D",X"01",
		X"20",X"86",X"D3",X"68",X"86",X"04",X"06",X"A6",X"7C",X"1D",X"D2",X"AD",X"48",X"4E",X"BD",X"DC",
		X"AD",X"20",X"DE",X"D2",X"68",X"AA",X"BD",X"D6",X"AD",X"A6",X"04",X"9D",X"A3",X"02",X"4D",X"C0",
		X"9D",X"A0",X"02",X"A5",X"01",X"9D",X"A1",X"02",X"A5",X"02",X"9D",X"A2",X"02",X"28",X"85",X"EF",
		X"EA",X"C8",X"C8",X"C8",X"C8",X"C8",X"C4",X"5A",X"D0",X"07",X"85",X"EF",X"6E",X"60",X"85",X"EF",
		X"EA",X"4C",X"FD",X"AC",X"85",X"EF",X"6E",X"A5",X"7B",X"09",X"08",X"85",X"7B",X"08",X"10",X"AF",
		X"A9",X"40",X"05",X"3E",X"85",X"3E",X"C9",X"E8",X"09",X"40",X"85",X"E8",X"4D",X"0C",X"20",X"86",
		X"D3",X"60",X"01",X"00",X"00",X"01",X"01",X"00",X"03",X"02",X"05",X"04",X"05",X"03",X"06",X"07",
		X"09",X"04",X"85",X"EF",X"6E",X"A5",X"5B",X"29",X"02",X"F0",X"11",X"A5",X"5F",X"85",X"E5",X"C9",
		X"3E",X"09",X"82",X"85",X"3E",X"4D",X"80",X"85",X"C7",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",
		X"A5",X"B2",X"F0",X"45",X"29",X"04",X"D0",X"52",X"A5",X"B2",X"29",X"01",X"D0",X"3F",X"A5",X"7E",
		X"18",X"69",X"08",X"49",X"FF",X"8D",X"3A",X"07",X"38",X"E9",X"10",X"8D",X"3E",X"07",X"18",X"69",
		X"20",X"8D",X"36",X"07",X"A9",X"04",X"85",X"BD",X"85",X"BE",X"85",X"BF",X"A9",X"20",X"85",X"C0",
		X"A9",X"00",X"85",X"C4",X"85",X"DF",X"A9",X"D8",X"8D",X"3B",X"07",X"8D",X"37",X"07",X"8D",X"3F",
		X"07",X"85",X"EF",X"EA",X"06",X"B2",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"20",X"45",X"CD",
		X"A9",X"00",X"85",X"9F",X"4C",X"44",X"AE",X"85",X"EF",X"EA",X"A6",X"C4",X"D6",X"BD",X"D0",X"0F",
		X"E8",X"86",X"C4",X"E0",X"04",X"D0",X"08",X"A9",X"80",X"85",X"1D",X"60",X"85",X"EF",X"EA",X"8A",
		X"0A",X"A8",X"B9",X"97",X"AE",X"8D",X"35",X"07",X"B9",X"98",X"AE",X"8D",X"34",X"07",X"B9",X"9F",
		X"AE",X"8D",X"39",X"07",X"B9",X"A0",X"AE",X"8D",X"38",X"07",X"B9",X"A7",X"AE",X"8D",X"3D",X"07",
		X"B9",X"A8",X"AE",X"8D",X"3C",X"07",X"60",X"17",X"01",X"18",X"01",X"19",X"01",X"00",X"00",X"14",
		X"01",X"15",X"01",X"16",X"01",X"00",X"00",X"17",X"03",X"18",X"03",X"19",X"03",X"00",X"00",X"85",
		X"EF",X"EA",X"A5",X"7B",X"29",X"10",X"F0",X"28",X"A5",X"B1",X"D0",X"28",X"A9",X"0D",X"20",X"86",
		X"D3",X"A9",X"40",X"85",X"C7",X"20",X"10",X"AF",X"A9",X"05",X"85",X"9F",X"A9",X"0C",X"85",X"A0",
		X"A9",X"02",X"85",X"A4",X"A9",X"10",X"85",X"A1",X"20",X"08",X"C9",X"E6",X"B1",X"85",X"EF",X"EA",
		X"60",X"85",X"EF",X"EA",X"A6",X"A3",X"BD",X"0C",X"AF",X"85",X"7F",X"A5",X"B1",X"C9",X"20",X"90",
		X"0C",X"E6",X"7E",X"A5",X"7E",X"C9",X"FC",X"B0",X"0A",X"60",X"85",X"EF",X"EA",X"E6",X"B1",X"60",
		X"85",X"EF",X"EA",X"A9",X"80",X"85",X"1D",X"4D",X"00",X"85",X"DF",X"60",X"F0",X"F4",X"85",X"EF",
		X"EA",X"A5",X"7E",X"85",X"45",X"C9",X"7F",X"85",X"46",X"A5",X"7C",X"85",X"47",X"28",X"85",X"EF",
		X"EA",X"A5",X"9F",X"D0",X"08",X"8D",X"20",X"07",X"F0",X"4A",X"85",X"EF",X"6E",X"A5",X"A5",X"C5",
		X"A0",X"D0",X"09",X"A5",X"A6",X"C5",X"9F",X"F0",X"0E",X"85",X"EF",X"EA",X"A5",X"A1",X"85",X"A2",
		X"A9",X"00",X"85",X"A3",X"C1",X"EF",X"6E",X"C6",X"A2",X"D0",X"13",X"A5",X"A1",X"85",X"A2",X"EA",
		X"A3",X"A5",X"A3",X"C5",X"A4",X"D0",X"07",X"A9",X"00",X"85",X"A3",X"85",X"EF",X"6E",X"A5",X"A3",
		X"18",X"65",X"A0",X"8D",X"21",X"07",X"C9",X"9F",X"8D",X"20",X"07",X"85",X"A6",X"C9",X"A0",X"85",
		X"A5",X"85",X"EF",X"EA",X"A2",X"00",X"A5",X"7C",X"29",X"01",X"F0",X"04",X"E8",X"85",X"EF",X"6E",
		X"AD",X"03",X"40",X"29",X"40",X"F0",X"09",X"A5",X"12",X"F0",X"05",X"E8",X"E8",X"85",X"EF",X"6E",
		X"A5",X"7E",X"18",X"7D",X"AA",X"AF",X"18",X"69",X"08",X"49",X"FF",X"8D",X"22",X"07",X"C9",X"7F",
		X"38",X"E9",X"0E",X"8D",X"23",X"07",X"C1",X"EF",X"EA",X"60",X"00",X"02",X"FE",X"00",X"85",X"EF",
		X"EA",X"A5",X"8B",X"29",X"01",X"F0",X"07",X"A9",X"02",X"85",X"67",X"85",X"EF",X"6E",X"60",X"85",
		X"EF",X"EA",X"A5",X"8B",X"29",X"02",X"D0",X"08",X"A9",X"00",X"85",X"A7",X"28",X"85",X"EF",X"6E",
		X"A9",X"01",X"85",X"A7",X"28",X"85",X"EF",X"6E",X"A5",X"8B",X"29",X"20",X"F0",X"7A",X"A9",X"80",
		X"85",X"8D",X"A5",X"7C",X"4A",X"90",X"07",X"A9",X"01",X"10",X"08",X"85",X"EF",X"6E",X"A9",X"02",
		X"85",X"EF",X"EA",X"85",X"8F",X"C9",X"7E",X"85",X"90",X"85",X"92",X"A5",X"7F",X"85",X"91",X"C1",
		X"93",X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"8D",X"95",X"5B",X"CA",X"10",X"F9",X"20",X"E1",X"CA",
		X"A5",X"67",X"C9",X"03",X"D0",X"0E",X"A5",X"8B",X"29",X"10",X"85",X"8B",X"A9",X"00",X"85",X"8D",
		X"60",X"85",X"EF",X"EA",X"A5",X"8F",X"49",X"02",X"09",X"01",X"85",X"9F",X"85",X"A7",X"A9",X"0E",
		X"85",X"A8",X"A9",X"0F",X"85",X"A0",X"A5",X"91",X"38",X"E9",X"10",X"85",X"91",X"85",X"93",X"A9",
		X"01",X"85",X"A4",X"85",X"AC",X"A5",X"8B",X"29",X"D7",X"09",X"40",X"85",X"8B",X"A9",X"0A",X"85",
		X"8C",X"A9",X"FF",X"85",X"B3",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"8B",X"29",X"04",
		X"F0",X"26",X"A5",X"8B",X"29",X"F9",X"09",X"02",X"85",X"8B",X"A9",X"10",X"85",X"9C",X"A5",X"7F",
		X"85",X"91",X"85",X"93",X"A9",X"13",X"85",X"A8",X"A9",X"00",X"85",X"87",X"85",X"9E",X"A9",X"01",
		X"85",X"AA",X"20",X"07",X"B3",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"8B",X"29",X"02",
		X"D0",X"04",X"60",X"85",X"EF",X"EA",X"A5",X"8B",X"29",X"FE",X"85",X"8B",X"85",X"EF",X"EA",X"A5",
		X"D4",X"D0",X"53",X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"8D",X"95",X"5B",X"CA",X"10",X"F9",X"85",
		X"EF",X"EA",X"20",X"E1",X"CA",X"A5",X"67",X"C9",X"02",X"B0",X"3F",X"A9",X"00",X"85",X"AF",X"20",
		X"3D",X"CC",X"85",X"EF",X"EA",X"A2",X"0F",X"85",X"EF",X"EA",X"B5",X"5B",X"95",X"8D",X"CA",X"10",
		X"F9",X"A5",X"92",X"85",X"90",X"A5",X"93",X"85",X"91",X"C9",X"E8",X"B0",X"2E",X"A5",X"8B",X"29",
		X"02",X"D0",X"09",X"A9",X"00",X"85",X"A7",X"F0",X"0A",X"85",X"EF",X"EA",X"A9",X"01",X"85",X"A7",
		X"85",X"EF",X"EA",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"8B",X"29",X"F8",X"85",X"8B",
		X"A9",X"80",X"85",X"B0",X"C1",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"8B",X"29",X"F8",X"85",
		X"8B",X"A9",X"18",X"85",X"D3",X"4D",X"01",X"85",X"A7",X"A9",X"14",X"85",X"A8",X"4D",X"04",X"20",
		X"86",X"D3",X"60",X"85",X"EF",X"6E",X"A5",X"B0",X"10",X"1D",X"A5",X"91",X"18",X"69",X"03",X"85",
		X"91",X"C9",X"E8",X"90",X"12",X"06",X"B0",X"4D",X"18",X"85",X"D3",X"A9",X"14",X"85",X"A8",X"4D",
		X"04",X"20",X"86",X"D3",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"D3",X"F0",X"3B",X"C6",
		X"D3",X"08",X"C9",X"10",X"D0",X"05",X"E6",X"A8",X"85",X"EF",X"EA",X"C9",X"08",X"D0",X"05",X"E6",
		X"A8",X"85",X"EF",X"EA",X"28",X"D0",X"23",X"A5",X"B3",X"C9",X"01",X"30",X"0B",X"A5",X"B4",X"C9",
		X"01",X"F0",X"05",X"E6",X"B4",X"C1",X"EF",X"6E",X"A5",X"8B",X"29",X"78",X"85",X"8B",X"4D",X"00",
		X"85",X"A7",X"85",X"8D",X"C5",X"24",X"07",X"C1",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A5",X"8C",
		X"F0",X"25",X"A5",X"8C",X"C9",X"05",X"D0",X"10",X"A9",X"10",X"85",X"A8",X"4D",X"11",X"85",X"A0",
		X"A9",X"09",X"20",X"86",X"D3",X"85",X"EF",X"6E",X"C6",X"8C",X"D0",X"0B",X"A5",X"8B",X"29",X"BF",
		X"09",X"04",X"85",X"8B",X"C1",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"10",X"F0",X"3F",X"A6",
		X"12",X"AD",X"03",X"40",X"29",X"40",X"D0",X"05",X"A2",X"00",X"85",X"EF",X"6E",X"BD",X"00",X"40",
		X"49",X"FF",X"29",X"10",X"48",X"78",X"13",X"45",X"8B",X"29",X"10",X"F0",X"10",X"A9",X"A9",X"85",
		X"8B",X"A9",X"00",X"85",X"D3",X"C1",X"B0",X"C1",X"EF",X"EA",X"85",X"EF",X"6E",X"85",X"EF",X"6E",
		X"A5",X"8B",X"29",X"EF",X"85",X"8B",X"2C",X"05",X"8B",X"85",X"8B",X"85",X"EF",X"6E",X"60",X"85",
		X"EF",X"EA",X"A5",X"8B",X"29",X"02",X"D0",X"08",X"A5",X"B0",X"30",X"04",X"60",X"85",X"EF",X"EA",
		X"A2",X"00",X"A5",X"96",X"F0",X"06",X"E8",X"C6",X"96",X"85",X"EF",X"EA",X"A5",X"91",X"38",X"FD",
		X"93",X"B2",X"85",X"03",X"A2",X"09",X"85",X"EF",X"EA",X"BD",X"9E",X"B4",X"85",X"02",X"CA",X"BD",
		X"9E",X"B4",X"85",X"01",X"A0",X"00",X"B1",X"01",X"10",X"52",X"29",X"0C",X"D0",X"4E",X"A0",X"04",
		X"B1",X"01",X"38",X"E5",X"03",X"B0",X"07",X"49",X"FF",X"69",X"01",X"85",X"EF",X"EA",X"C9",X"08",
		X"B0",X"3A",X"88",X"B1",X"01",X"38",X"F9",X"8D",X"00",X"B0",X"07",X"49",X"FF",X"69",X"01",X"85",
		X"EF",X"EA",X"C9",X"08",X"B0",X"26",X"A9",X"0A",X"20",X"86",X"D3",X"A0",X"00",X"B1",X"01",X"09",
		X"08",X"91",X"01",X"29",X"40",X"F0",X"0A",X"A9",X"0B",X"20",X"86",X"D3",X"E6",X"B3",X"85",X"EF",
		X"EA",X"A0",X"1A",X"B1",X"01",X"09",X"20",X"91",X"01",X"85",X"EF",X"EA",X"CA",X"10",X"9A",X"85",
		X"EF",X"EA",X"60",X"00",X"08",X"85",X"EF",X"EA",X"A5",X"8B",X"10",X"18",X"20",X"25",X"B1",X"20",
		X"01",X"B2",X"20",X"8D",X"B1",X"20",X"8B",X"B0",X"20",X"D7",X"AF",X"20",X"5B",X"B0",X"20",X"4A",
		X"B1",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"8B",X"10",X"48",X"A5",X"8B",X"29",X"02",
		X"F0",X"23",X"C6",X"AA",X"D0",X"1F",X"A5",X"A9",X"85",X"AA",X"A5",X"A7",X"49",X"04",X"85",X"A7",
		X"29",X"02",X"D0",X"05",X"E6",X"AC",X"85",X"EF",X"EA",X"A5",X"AC",X"29",X"01",X"18",X"69",X"12",
		X"85",X"A8",X"85",X"EF",X"EA",X"A5",X"A7",X"8D",X"24",X"07",X"A5",X"A8",X"8D",X"25",X"07",X"A5",
		X"90",X"18",X"69",X"08",X"49",X"FF",X"8D",X"26",X"07",X"A5",X"91",X"38",X"E9",X"0E",X"8D",X"27",
		X"07",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A9",X"06",X"85",X"A1",X"C9",X"87",X"C9",X"02",
		X"D0",X"08",X"A9",X"06",X"85",X"A2",X"28",X"85",X"EF",X"EA",X"A9",X"02",X"85",X"A4",X"C9",X"7C",
		X"C9",X"03",X"48",X"D0",X"0B",X"A9",X"01",X"85",X"9F",X"A9",X"00",X"85",X"A0",X"C1",X"EF",X"6E",
		X"68",X"C9",X"02",X"48",X"70",X"0B",X"A9",X"01",X"85",X"9F",X"A9",X"02",X"85",X"A0",X"C1",X"EF",
		X"EA",X"68",X"C9",X"01",X"48",X"70",X"0B",X"A9",X"03",X"85",X"9F",X"A9",X"02",X"85",X"A0",X"C1",
		X"EF",X"EA",X"68",X"48",X"70",X"0B",X"A9",X"03",X"85",X"9F",X"A9",X"00",X"85",X"A0",X"C1",X"EF",
		X"EA",X"68",X"60",X"85",X"EF",X"6E",X"24",X"C7",X"30",X"0B",X"70",X"3E",X"A5",X"D7",X"D0",X"05",
		X"F0",X"07",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A2",X"00",X"85",X"EF",X"6E",X"BD",X"9D",
		X"B3",X"38",X"E5",X"4A",X"BD",X"9E",X"B3",X"E5",X"4B",X"90",X"08",X"E8",X"E8",X"4C",X"7E",X"B3",
		X"85",X"EF",X"EA",X"8A",X"4A",X"AA",X"E8",X"86",X"C7",X"20",X"CE",X"B3",X"60",X"98",X"02",X"28",
		X"02",X"98",X"01",X"28",X"01",X"00",X"00",X"85",X"EF",X"EA",X"20",X"B2",X"B3",X"06",X"C7",X"28",
		X"85",X"EF",X"EA",X"A9",X"00",X"A2",X"18",X"85",X"EF",X"EA",X"9D",X"28",X"07",X"66",X"10",X"FA",
		X"A2",X"A1",X"85",X"EF",X"6E",X"9D",X"FF",X"01",X"CA",X"D0",X"FA",X"60",X"85",X"EF",X"6E",X"A9",
		X"00",X"85",X"C5",X"85",X"EF",X"6E",X"A9",X"00",X"20",X"71",X"B4",X"A5",X"5B",X"30",X"03",X"4C",
		X"69",X"B4",X"29",X"0C",X"D0",X"77",X"20",X"00",X"B5",X"20",X"B6",X"B4",X"20",X"57",X"B5",X"20",
		X"07",X"B7",X"20",X"78",X"B7",X"20",X"3D",X"CC",X"20",X"67",X"B7",X"85",X"EF",X"6E",X"20",X"AA",
		X"B4",X"85",X"EF",X"EA",X"20",X"B4",X"B7",X"85",X"EF",X"EA",X"20",X"37",X"B8",X"20",X"A0",X"B8",
		X"85",X"EF",X"EA",X"A9",X"01",X"20",X"71",X"B4",X"E6",X"C6",X"A5",X"40",X"29",X"02",X"4A",X"AA",
		X"A5",X"C6",X"DD",X"58",X"B4",X"90",X"07",X"A9",X"00",X"85",X"C6",X"85",X"EF",X"EA",X"E6",X"C5",
		X"A2",X"07",X"AD",X"04",X"40",X"29",X"10",X"F0",X"0F",X"A5",X"40",X"C9",X"08",X"90",X"05",X"A9",
		X"07",X"85",X"EF",X"EA",X"AA",X"85",X"EF",X"EA",X"A5",X"C5",X"DD",X"50",X"B4",X"90",X"87",X"60",
		X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"05",X"04",X"85",X"EF",X"EA",X"20",X"8F",X"B9",
		X"20",X"FA",X"BA",X"4C",X"04",X"B4",X"85",X"EF",X"EA",X"20",X"5C",X"BD",X"4C",X"13",X"B4",X"85",
		X"EF",X"EA",X"48",X"A5",X"C6",X"0A",X"AA",X"BD",X"9E",X"B4",X"85",X"01",X"BD",X"9F",X"B4",X"85",
		X"02",X"A0",X"1F",X"68",X"D0",X"0F",X"85",X"EF",X"EA",X"B1",X"01",X"99",X"5B",X"00",X"88",X"10",
		X"F8",X"60",X"85",X"EF",X"EA",X"B9",X"5B",X"00",X"91",X"01",X"88",X"10",X"F8",X"60",X"00",X"02",
		X"20",X"02",X"40",X"02",X"60",X"02",X"80",X"02",X"85",X"EF",X"EA",X"A5",X"60",X"85",X"5E",X"A5",
		X"61",X"85",X"5F",X"60",X"85",X"EF",X"EA",X"23",X"5B",X"50",X"3A",X"A5",X"6A",X"D0",X"36",X"A5",
		X"D6",X"D0",X"05",X"C6",X"6C",X"85",X"EF",X"EA",X"A5",X"6C",X"D0",X"1C",X"A4",X"6D",X"B9",X"F6",
		X"B4",X"85",X"6B",X"C8",X"B9",X"F6",X"B4",X"85",X"6C",X"C8",X"C0",X"08",X"90",X"05",X"A0",X"00",
		X"85",X"EF",X"EA",X"84",X"6D",X"85",X"EF",X"EA",X"A5",X"61",X"C5",X"7F",X"90",X"07",X"A9",X"00",
		X"85",X"6B",X"85",X"EF",X"EA",X"60",X"00",X"0C",X"01",X"09",X"00",X"06",X"01",X"04",X"85",X"EF",
		X"EA",X"A5",X"5B",X"29",X"1C",X"C9",X"10",X"D0",X"19",X"20",X"6D",X"B9",X"A0",X"01",X"B1",X"01",
		X"C9",X"41",X"B0",X"12",X"C9",X"40",X"F0",X"29",X"85",X"EF",X"EA",X"A9",X"02",X"85",X"67",X"C1",
		X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A9",X"3F",X"85",X"6E",X"A5",X"6F",X"29",X"F0",X"09",X"02",
		X"85",X"6F",X"A9",X"04",X"85",X"70",X"C1",X"72",X"A9",X"00",X"85",X"71",X"78",X"DD",X"85",X"EF",
		X"EA",X"A5",X"72",X"C9",X"01",X"D0",X"0B",X"A5",X"5B",X"29",X"88",X"09",X"40",X"85",X"5B",X"C1",
		X"EF",X"EA",X"4C",X"1B",X"B5",X"85",X"EF",X"6E",X"A5",X"6A",X"D0",X"39",X"A5",X"5B",X"29",X"10",
		X"D0",X"33",X"A9",X"1F",X"85",X"03",X"4D",X"CD",X"85",X"04",X"A9",X"21",X"85",X"05",X"4D",X"CD",
		X"85",X"06",X"A2",X"01",X"20",X"D3",X"CC",X"90",X"1C",X"A5",X"5B",X"09",X"01",X"85",X"5B",X"4D",
		X"04",X"85",X"6A",X"85",X"EF",X"6E",X"73",X"5B",X"50",X"3C",X"A5",X"6B",X"29",X"01",X"F0",X"09",
		X"D0",X"27",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"85",X"EF",X"EA",X"A5",X"7E",X"85",X"01",
		X"A5",X"7F",X"85",X"02",X"C1",X"EF",X"6E",X"A5",X"5E",X"85",X"03",X"A5",X"5F",X"85",X"04",X"08",
		X"F8",X"B5",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"20",X"9D",X"CE",X"A5",X"1A",X"29",X"03",
		X"85",X"5D",X"60",X"85",X"EF",X"6E",X"A5",X"5B",X"29",X"20",X"F0",X"18",X"C6",X"78",X"10",X"14",
		X"A5",X"61",X"C9",X"56",X"90",X"0E",X"A5",X"5B",X"09",X"10",X"85",X"5B",X"4D",X"02",X"85",X"67",
		X"60",X"85",X"EF",X"EA",X"20",X"9D",X"CE",X"A5",X"1A",X"65",X"7F",X"29",X"01",X"AA",X"BD",X"F4",
		X"B5",X"85",X"5D",X"60",X"01",X"02",X"85",X"EF",X"EA",X"A5",X"01",X"38",X"E5",X"03",X"26",X"05",
		X"A5",X"02",X"38",X"E5",X"04",X"26",X"05",X"A5",X"05",X"29",X"03",X"AA",X"BD",X"12",X"B6",X"85",
		X"5D",X"60",X"03",X"02",X"00",X"01",X"85",X"EF",X"EA",X"A5",X"7F",X"85",X"0A",X"A9",X"00",X"85",
		X"09",X"85",X"EF",X"EA",X"20",X"AA",X"D0",X"A6",X"CC",X"D0",X"0A",X"A9",X"D8",X"85",X"0A",X"4C",
		X"24",X"B6",X"85",X"EF",X"EA",X"A6",X"CB",X"E4",X"CC",X"90",X"05",X"A2",X"00",X"85",X"EF",X"EA",
		X"A0",X"00",X"85",X"EF",X"EA",X"BD",X"01",X"04",X"99",X"CD",X"00",X"E8",X"C8",X"C0",X"03",X"90",
		X"F4",X"E8",X"86",X"CB",X"BD",X"FC",X"03",X"C5",X"B9",X"D0",X"06",X"20",X"44",X"BD",X"85",X"EF",
		X"EA",X"60",X"85",X"EF",X"EA",X"A9",X"46",X"85",X"09",X"A9",X"D8",X"85",X"0A",X"20",X"AA",X"D0",
		X"A9",X"FF",X"85",X"04",X"85",X"08",X"A2",X"00",X"85",X"EF",X"EA",X"BD",X"00",X"04",X"30",X"50",
		X"BD",X"02",X"04",X"38",X"E5",X"7F",X"B0",X"21",X"49",X"FF",X"C5",X"04",X"B0",X"38",X"85",X"04",
		X"BD",X"00",X"04",X"85",X"09",X"BD",X"01",X"04",X"85",X"01",X"BD",X"02",X"04",X"85",X"02",X"BD",
		X"03",X"04",X"85",X"03",X"10",X"20",X"85",X"EF",X"EA",X"C5",X"08",X"B0",X"19",X"85",X"08",X"BD",
		X"00",X"04",X"85",X"0A",X"BD",X"01",X"04",X"85",X"05",X"BD",X"02",X"04",X"85",X"06",X"BD",X"03",
		X"04",X"85",X"07",X"85",X"EF",X"EA",X"E8",X"E8",X"E8",X"E8",X"4C",X"7B",X"B6",X"85",X"EF",X"EA",
		X"A2",X"00",X"A5",X"04",X"30",X"09",X"A5",X"09",X"C5",X"B9",X"D0",X"1C",X"85",X"EF",X"EA",X"A5",
		X"08",X"30",X"09",X"A5",X"0A",X"C5",X"B9",X"D0",X"0A",X"85",X"EF",X"EA",X"20",X"44",X"BD",X"60",
		X"85",X"EF",X"EA",X"A2",X"04",X"85",X"EF",X"EA",X"B5",X"01",X"85",X"CD",X"B5",X"02",X"85",X"CE",
		X"B5",X"03",X"85",X"CF",X"28",X"85",X"EF",X"6E",X"A5",X"5B",X"29",X"1C",X"D0",X"50",X"A9",X"00",
		X"85",X"C8",X"A5",X"5C",X"49",X"02",X"C5",X"5D",X"D0",X"07",X"A5",X"5C",X"85",X"5D",X"C1",X"EF",
		X"EA",X"20",X"E1",X"CA",X"A5",X"67",X"C9",X"02",X"D0",X"34",X"A5",X"5B",X"09",X"01",X"85",X"5B",
		X"A9",X"04",X"85",X"6A",X"EA",X"C8",X"08",X"EC",X"BA",X"A5",X"C8",X"DD",X"5F",X"B7",X"B0",X"0F",
		X"A6",X"C8",X"A5",X"5D",X"5D",X"61",X"B7",X"85",X"5D",X"4C",X"21",X"B7",X"85",X"EF",X"6E",X"A5",
		X"5B",X"09",X"08",X"85",X"5B",X"4D",X"40",X"05",X"75",X"85",X"75",X"85",X"EF",X"6E",X"60",X"02",
		X"04",X"00",X"03",X"02",X"03",X"85",X"EF",X"6E",X"A5",X"62",X"10",X"09",X"A5",X"5B",X"09",X"08",
		X"85",X"5B",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"61",X"C9",X"48",X"90",X"08",X"C9",
		X"E8",X"B0",X"20",X"60",X"85",X"EF",X"6E",X"E3",X"5B",X"50",X"14",X"A5",X"5D",X"49",X"02",X"85",
		X"5D",X"A9",X"00",X"85",X"6C",X"4D",X"04",X"85",X"6A",X"20",X"E1",X"CA",X"85",X"EF",X"6E",X"60",
		X"85",X"EF",X"EA",X"A5",X"5B",X"29",X"F0",X"09",X"08",X"85",X"5B",X"A5",X"75",X"09",X"40",X"85",
		X"75",X"60",X"85",X"EF",X"6E",X"A0",X"00",X"A5",X"5B",X"10",X"6E",X"29",X"04",X"D0",X"6A",X"A5",
		X"5B",X"29",X"08",X"F0",X"0D",X"24",X"5B",X"70",X"60",X"A5",X"75",X"29",X"20",X"D0",X"5A",X"85",
		X"EF",X"EA",X"A5",X"7B",X"10",X"53",X"29",X"0C",X"D0",X"4F",X"A5",X"7E",X"38",X"E5",X"5E",X"B0",
		X"08",X"49",X"FF",X"AA",X"E8",X"8A",X"85",X"EF",X"EA",X"D9",X"2E",X"B8",X"B0",X"3B",X"A6",X"64",
		X"A5",X"5F",X"18",X"7D",X"32",X"B8",X"85",X"01",X"A5",X"7F",X"38",X"E5",X"01",X"B0",X"08",X"49",
		X"FF",X"AA",X"E8",X"8A",X"85",X"EF",X"EA",X"D9",X"30",X"B8",X"B0",X"1D",X"A5",X"7B",X"09",X"08",
		X"85",X"7B",X"20",X"10",X"AF",X"A9",X"40",X"05",X"3E",X"85",X"3E",X"A5",X"E8",X"09",X"40",X"85",
		X"E8",X"A9",X"0C",X"20",X"86",X"D3",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"64",X"60",X"06",X"06",
		X"03",X"06",X"00",X"08",X"F8",X"85",X"EF",X"EA",X"A5",X"5B",X"10",X"57",X"29",X"1C",X"D0",X"53",
		X"A5",X"5C",X"29",X"02",X"49",X"02",X"0A",X"0A",X"0A",X"09",X"01",X"85",X"02",X"24",X"5B",X"70",
		X"08",X"A2",X"08",X"4C",X"60",X"B8",X"85",X"EF",X"EA",X"A5",X"5C",X"0A",X"AA",X"85",X"EF",X"EA",
		X"BD",X"94",X"B8",X"85",X"01",X"BD",X"95",X"B8",X"85",X"03",X"A5",X"01",X"C5",X"6E",X"D0",X"09",
		X"A5",X"02",X"C5",X"6F",X"F0",X"0E",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"71",X"A5",X"03",X"85",
		X"72",X"85",X"EF",X"EA",X"A5",X"01",X"85",X"6E",X"A5",X"02",X"85",X"6F",X"A5",X"03",X"85",X"70",
		X"85",X"EF",X"EA",X"60",X"30",X"03",X"32",X"03",X"32",X"03",X"30",X"03",X"41",X"03",X"85",X"EF",
		X"EA",X"20",X"6D",X"B9",X"A5",X"5B",X"0A",X"26",X"03",X"A2",X"00",X"A5",X"61",X"C9",X"37",X"90",
		X"04",X"E8",X"85",X"EF",X"EA",X"A5",X"03",X"3D",X"3F",X"B9",X"85",X"03",X"A5",X"6F",X"48",X"10",
		X"09",X"A9",X"80",X"05",X"03",X"85",X"03",X"85",X"EF",X"EA",X"68",X"29",X"7F",X"4A",X"4A",X"4A",
		X"05",X"03",X"A0",X"00",X"91",X"01",X"C8",X"C6",X"72",X"D0",X"15",X"A5",X"70",X"85",X"72",X"E6",
		X"71",X"A5",X"6F",X"29",X"0F",X"C5",X"71",X"B0",X"07",X"A9",X"00",X"85",X"71",X"85",X"EF",X"EA",
		X"A5",X"6E",X"18",X"65",X"71",X"91",X"01",X"C8",X"20",X"43",X"B9",X"85",X"EF",X"EA",X"A5",X"60",
		X"18",X"7D",X"3B",X"B9",X"49",X"FF",X"91",X"01",X"C8",X"A5",X"61",X"48",X"1C",X"E9",X"0E",X"91",
		X"01",X"68",X"C9",X"36",X"90",X"0B",X"C9",X"46",X"B0",X"07",X"24",X"5B",X"50",X"07",X"85",X"EF",
		X"EA",X"60",X"85",X"EF",X"6E",X"49",X"FF",X"38",X"E9",X"09",X"29",X"0F",X"18",X"69",X"B0",X"A0",
		X"01",X"91",X"01",X"88",X"B1",X"01",X"29",X"FB",X"91",X"01",X"60",X"08",X"0A",X"06",X"08",X"00",
		X"01",X"85",X"EF",X"EA",X"A2",X"00",X"A5",X"5B",X"29",X"04",X"F0",X"1E",X"A5",X"5C",X"29",X"01",
		X"F0",X"08",X"A5",X"73",X"30",X"04",X"E8",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"29",X"40",X"F0",
		X"09",X"A5",X"12",X"F0",X"05",X"E8",X"E8",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A5",X"C6",
		X"0A",X"AA",X"BD",X"81",X"B9",X"85",X"01",X"DD",X"82",X"B9",X"85",X"02",X"28",X"20",X"07",X"24",
		X"07",X"28",X"07",X"2C",X"07",X"30",X"07",X"34",X"07",X"38",X"07",X"3C",X"07",X"85",X"EF",X"6E",
		X"A5",X"5B",X"29",X"04",X"F0",X"12",X"20",X"AB",X"B9",X"20",X"D8",X"B9",X"20",X"15",X"BA",X"20",
		X"7D",X"BA",X"20",X"C6",X"BA",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"73",X"D0",X"25",
		X"A9",X"36",X"85",X"6E",X"C9",X"5C",X"29",X"02",X"49",X"02",X"0A",X"0A",X"0A",X"09",X"03",X"85",
		X"6F",X"A9",X"02",X"85",X"70",X"C1",X"72",X"4D",X"00",X"85",X"71",X"A9",X"10",X"85",X"73",X"08",
		X"8D",X"CC",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"73",X"29",X"10",X"F0",X"33",X"20",
		X"6D",X"B9",X"A0",X"01",X"B1",X"01",X"C9",X"39",X"D0",X"22",X"A5",X"72",X"C9",X"01",X"D0",X"1C",
		X"A9",X"FF",X"85",X"6E",X"4D",X"00",X"85",X"6F",X"85",X"71",X"06",X"73",X"08",X"9D",X"CE",X"A5",
		X"1A",X"65",X"7F",X"29",X"0F",X"05",X"73",X"85",X"73",X"85",X"EF",X"EA",X"20",X"8D",X"CC",X"85",
		X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"73",X"29",X"20",X"F0",X"0B",X"A5",X"73",X"29",X"0F",
		X"F0",X"09",X"C6",X"73",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"24",X"5B",X"70",X"09",X"20",
		X"18",X"B6",X"4C",X"3E",X"BA",X"85",X"EF",X"EA",X"20",X"64",X"B6",X"85",X"EF",X"EA",X"A5",X"CD",
		X"85",X"5E",X"A5",X"CE",X"85",X"5F",X"A5",X"CF",X"85",X"5C",X"85",X"5D",X"20",X"EC",X"BA",X"BD",
		X"79",X"BA",X"85",X"6E",X"A5",X"5C",X"29",X"02",X"49",X"02",X"0A",X"0A",X"0A",X"09",X"03",X"85",
		X"6F",X"A9",X"02",X"85",X"70",X"85",X"72",X"A9",X"00",X"85",X"71",X"20",X"8D",X"CC",X"A5",X"73",
		X"29",X"F0",X"0A",X"85",X"73",X"85",X"EF",X"EA",X"60",X"43",X"3A",X"85",X"EF",X"EA",X"A5",X"73",
		X"29",X"40",X"F0",X"3B",X"20",X"6D",X"B9",X"20",X"EC",X"BA",X"A0",X"01",X"B1",X"01",X"DD",X"C0",
		X"BA",X"D0",X"26",X"A5",X"72",X"C9",X"01",X"D0",X"20",X"BD",X"C2",X"BA",X"85",X"6E",X"A5",X"6F",
		X"29",X"F0",X"09",X"01",X"85",X"6F",X"A9",X"04",X"85",X"70",X"85",X"72",X"A9",X"00",X"85",X"71",
		X"06",X"73",X"A9",X"02",X"85",X"6A",X"85",X"EF",X"EA",X"20",X"8D",X"CC",X"85",X"EF",X"EA",X"60",
		X"46",X"3D",X"41",X"32",X"85",X"EF",X"EA",X"A5",X"73",X"10",X"1E",X"A5",X"D2",X"D0",X"1A",X"20",
		X"E1",X"CA",X"20",X"3D",X"CC",X"20",X"AA",X"B4",X"A5",X"6A",X"D0",X"0D",X"A9",X"00",X"85",X"73",
		X"A5",X"5B",X"29",X"FB",X"85",X"5B",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A2",X"00",X"24",
		X"5B",X"50",X"04",X"E8",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"5B",X"29",X"08",X"F0",
		X"32",X"24",X"5B",X"70",X"16",X"24",X"75",X"50",X"2E",X"A5",X"74",X"C9",X"02",X"B0",X"06",X"20",
		X"8A",X"BB",X"85",X"EF",X"6E",X"4C",X"24",X"BB",X"85",X"EF",X"EA",X"20",X"9E",X"BB",X"20",X"E1",
		X"BB",X"85",X"EF",X"EA",X"20",X"5F",X"BC",X"20",X"99",X"BC",X"20",X"B9",X"BC",X"20",X"2F",X"BD",
		X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A5",X"6E",X"C9",X"30",X"90",X"12",X"C9",X"43",X"90",
		X"1E",X"20",X"6D",X"B9",X"A0",X"01",X"B1",X"01",X"C9",X"4B",X"F0",X"2C",X"85",X"EF",X"6E",X"20",
		X"B9",X"BC",X"20",X"2F",X"BD",X"20",X"8D",X"CC",X"20",X"AA",X"B4",X"60",X"85",X"EF",X"6E",X"A9",
		X"49",X"85",X"6E",X"A9",X"05",X"85",X"70",X"C1",X"72",X"A5",X"6F",X"09",X"02",X"85",X"6F",X"4D",
		X"00",X"85",X"71",X"F0",X"DA",X"85",X"EF",X"6E",X"A5",X"72",X"C9",X"01",X"D0",X"07",X"A9",X"08",
		X"85",X"74",X"85",X"EF",X"6E",X"4C",X"4F",X"BB",X"85",X"EF",X"EA",X"A9",X"47",X"85",X"6E",X"C9",
		X"70",X"85",X"72",X"A9",X"00",X"85",X"71",X"4D",X"02",X"85",X"74",X"60",X"85",X"EF",X"6E",X"A5",
		X"74",X"D0",X"3B",X"A5",X"B4",X"85",X"B5",X"4A",X"00",X"A5",X"5E",X"C9",X"80",X"B0",X"05",X"A2",
		X"01",X"85",X"EF",X"EA",X"8A",X"18",X"65",X"B3",X"6A",X"6A",X"29",X"80",X"48",X"81",X"75",X"85",
		X"75",X"68",X"4A",X"4A",X"4A",X"09",X"81",X"85",X"6F",X"A9",X"01",X"85",X"74",X"4D",X"34",X"85",
		X"6E",X"A9",X"03",X"85",X"70",X"C1",X"72",X"4D",X"00",X"85",X"71",X"85",X"EF",X"6E",X"60",X"85",
		X"EF",X"EA",X"A5",X"74",X"29",X"01",X"F0",X"27",X"C6",X"77",X"30",X"27",X"A5",X"76",X"0A",X"AA",
		X"BD",X"4D",X"BC",X"18",X"65",X"60",X"85",X"60",X"BD",X"4E",X"BC",X"18",X"65",X"61",X"C9",X"46",
		X"B0",X"05",X"A9",X"46",X"85",X"EF",X"EA",X"85",X"61",X"20",X"AA",X"B4",X"85",X"EF",X"EA",X"60",
		X"85",X"EF",X"EA",X"A5",X"75",X"48",X"29",X"0F",X"0A",X"AA",X"BD",X"3D",X"BC",X"30",X"1A",X"85",
		X"76",X"BD",X"3E",X"BC",X"85",X"77",X"68",X"10",X"0A",X"A6",X"76",X"BD",X"45",X"BC",X"85",X"76",
		X"85",X"EF",X"EA",X"E6",X"75",X"60",X"85",X"EF",X"EA",X"68",X"06",X"74",X"60",X"07",X"08",X"06",
		X"08",X"05",X"08",X"FF",X"FF",X"00",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"FE",X"02",
		X"FE",X"02",X"00",X"02",X"02",X"00",X"02",X"FE",X"02",X"FE",X"00",X"FE",X"FE",X"85",X"EF",X"EA",
		X"A5",X"74",X"29",X"02",X"F0",X"30",X"A5",X"61",X"18",X"69",X"07",X"85",X"61",X"20",X"AA",X"B4",
		X"A5",X"61",X"C9",X"EE",X"90",X"20",X"A9",X"E6",X"85",X"61",X"A9",X"14",X"85",X"6E",X"A9",X"02",
		X"85",X"6F",X"A9",X"04",X"85",X"70",X"85",X"72",X"A9",X"00",X"85",X"71",X"06",X"74",X"A9",X"04",
		X"20",X"86",X"D3",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"74",X"29",X"04",X"F0",X"16",
		X"20",X"6D",X"B9",X"A0",X"01",X"B1",X"01",X"C9",X"16",X"D0",X"0B",X"A5",X"72",X"C9",X"01",X"D0",
		X"05",X"06",X"74",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"74",X"29",X"08",X"F0",X"54",
		X"A5",X"75",X"29",X"20",X"F0",X"49",X"A9",X"00",X"24",X"5B",X"50",X"06",X"38",X"65",X"B5",X"85",
		X"EF",X"EA",X"85",X"01",X"A5",X"40",X"38",X"85",X"EF",X"EA",X"E9",X"04",X"B0",X"FC",X"69",X"04",
		X"A8",X"A9",X"FD",X"85",X"EF",X"EA",X"18",X"69",X"03",X"88",X"10",X"FA",X"18",X"65",X"01",X"48",
		X"AA",X"BD",X"15",X"BD",X"20",X"DE",X"D2",X"68",X"AA",X"BD",X"21",X"BD",X"85",X"6E",X"A9",X"80",
		X"85",X"6F",X"A9",X"28",X"85",X"70",X"C1",X"72",X"A9",X"00",X"85",X"71",X"C1",X"EF",X"6E",X"06",
		X"74",X"85",X"EF",X"EA",X"60",X"01",X"02",X"07",X"01",X"07",X"05",X"01",X"07",X"06",X"01",X"05",
		X"06",X"23",X"24",X"25",X"23",X"25",X"26",X"23",X"25",X"27",X"23",X"26",X"27",X"85",X"EF",X"6E",
		X"A5",X"74",X"29",X"10",X"F0",X"23",X"A5",X"75",X"29",X"20",X"F0",X"09",X"A5",X"72",X"C9",X"01",
		X"D0",X"17",X"85",X"EF",X"6E",X"C6",X"C9",X"C9",X"5B",X"29",X"60",X"F0",X"05",X"C6",X"CA",X"C1",
		X"EF",X"EA",X"A9",X"00",X"85",X"5B",X"C1",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A2",X"1F",X"A9",
		X"00",X"85",X"EF",X"EA",X"95",X"5B",X"66",X"10",X"FB",X"A5",X"40",X"C9",X"07",X"90",X"07",X"29",
		X"07",X"09",X"04",X"85",X"EF",X"6E",X"A8",X"A9",X"FA",X"85",X"EF",X"EA",X"18",X"69",X"06",X"88",
		X"10",X"FA",X"18",X"65",X"C7",X"AA",X"AD",X"04",X"40",X"29",X"08",X"D0",X"08",X"8A",X"18",X"69",
		X"30",X"AA",X"85",X"EF",X"6E",X"A5",X"C9",X"DD",X"CB",X"BD",X"B0",X"2E",X"A5",X"CA",X"DD",X"2B",
		X"BE",X"B0",X"18",X"A5",X"5B",X"09",X"20",X"85",X"5B",X"20",X"9D",X"CE",X"A5",X"1A",X"65",X"7F",
		X"09",X"01",X"29",X"03",X"85",X"78",X"EA",X"CA",X"85",X"EF",X"EA",X"E6",X"C9",X"4D",X"84",X"05",
		X"5B",X"85",X"5B",X"A9",X"20",X"85",X"73",X"C1",X"EF",X"EA",X"60",X"00",X"01",X"01",X"01",X"01",
		X"00",X"00",X"02",X"02",X"03",X"03",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"03",X"03",
		X"04",X"04",X"00",X"00",X"03",X"04",X"05",X"05",X"00",X"00",X"04",X"04",X"05",X"05",X"00",X"00",
		X"04",X"04",X"04",X"04",X"00",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"02",X"03",X"03",X"04",
		X"00",X"00",X"03",X"03",X"04",X"04",X"00",X"00",X"02",X"02",X"02",X"03",X"00",X"00",X"03",X"03",
		X"04",X"04",X"00",X"00",X"03",X"04",X"05",X"05",X"00",X"00",X"04",X"04",X"05",X"05",X"00",X"00",
		X"04",X"04",X"04",X"04",X"00",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"00",X"01",X"01",X"02",X"00",X"00",X"03",X"03",
		X"04",X"04",X"00",X"00",X"03",X"03",X"03",X"04",X"00",X"00",X"03",X"03",X"03",X"03",X"00",X"00",
		X"03",X"03",X"03",X"04",X"00",X"00",X"03",X"03",X"04",X"04",X"00",X"00",X"02",X"03",X"03",X"04",
		X"00",X"00",X"03",X"03",X"04",X"04",X"00",X"00",X"02",X"02",X"02",X"03",X"00",X"00",X"03",X"03",
		X"04",X"04",X"00",X"00",X"03",X"03",X"03",X"04",X"00",X"00",X"03",X"03",X"03",X"03",X"00",X"00",
		X"03",X"03",X"03",X"04",X"00",X"00",X"03",X"03",X"04",X"04",X"00",X"85",X"EF",X"EA",X"20",X"97",
		X"BE",X"20",X"F0",X"BE",X"60",X"85",X"EF",X"EA",X"A5",X"3E",X"29",X"03",X"D0",X"3F",X"A5",X"40",
		X"29",X"02",X"F0",X"39",X"A5",X"7B",X"29",X"18",X"D0",X"33",X"AD",X"D0",X"02",X"29",X"C0",X"D0",
		X"2C",X"A5",X"D6",X"D0",X"28",X"C6",X"EB",X"10",X"24",X"A5",X"7B",X"29",X"04",X"D0",X"1E",X"A9",
		X"80",X"8D",X"D0",X"02",X"E6",X"EC",X"A5",X"EC",X"C9",X"10",X"90",X"07",X"A9",X"0F",X"85",X"EC",
		X"85",X"EF",X"EA",X"A6",X"EC",X"BD",X"DE",X"BE",X"85",X"EB",X"85",X"EF",X"EA",X"60",X"07",X"07",
		X"06",X"06",X"05",X"05",X"04",X"04",X"03",X"03",X"02",X"02",X"01",X"01",X"00",X"00",X"85",X"EF",
		X"EA",X"A5",X"ED",X"D0",X"1B",X"AD",X"D0",X"02",X"F0",X"16",X"C9",X"80",X"D0",X"09",X"20",X"13",
		X"BF",X"20",X"38",X"BF",X"85",X"EF",X"6E",X"20",X"B3",X"BF",X"20",X"53",X"C1",X"85",X"EF",X"6E",
		X"60",X"85",X"EF",X"EA",X"A5",X"7E",X"C9",X"80",X"2A",X"29",X"01",X"85",X"01",X"C9",X"7F",X"C9",
		X"90",X"2A",X"29",X"01",X"0A",X"18",X"65",X"01",X"8D",X"D9",X"02",X"A5",X"40",X"29",X"01",X"8D",
		X"D7",X"02",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A5",X"7E",X"85",X"01",X"C9",X"7F",X"85",
		X"02",X"AD",X"D9",X"02",X"4A",X"48",X"50",X"09",X"A5",X"01",X"49",X"FF",X"85",X"01",X"C1",X"EF",
		X"EA",X"68",X"4A",X"90",X"0C",X"A5",X"02",X"49",X"FF",X"18",X"69",X"20",X"85",X"02",X"C1",X"EF",
		X"EA",X"A5",X"02",X"4A",X"4A",X"4A",X"4A",X"38",X"E9",X"04",X"AA",X"A9",X"F8",X"85",X"EF",X"6E",
		X"18",X"69",X"08",X"CA",X"10",X"FA",X"85",X"02",X"A5",X"01",X"4A",X"4A",X"4A",X"4A",X"18",X"65",
		X"02",X"AA",X"BD",X"89",X"BF",X"8D",X"D8",X"02",X"60",X"03",X"03",X"02",X"02",X"02",X"01",X"00",
		X"00",X"03",X"03",X"03",X"02",X"02",X"01",X"01",X"00",X"04",X"03",X"03",X"03",X"02",X"02",X"01",
		X"00",X"04",X"04",X"04",X"03",X"03",X"02",X"02",X"01",X"04",X"04",X"04",X"04",X"04",X"03",X"02",
		X"02",X"85",X"EF",X"EA",X"2C",X"D0",X"02",X"30",X"06",X"70",X"43",X"60",X"85",X"EF",X"6E",X"AD",
		X"D0",X"02",X"49",X"C0",X"8D",X"D0",X"02",X"CD",X"D9",X"02",X"0A",X"0A",X"0D",X"D9",X"02",X"AA",
		X"A0",X"00",X"85",X"EF",X"6E",X"BD",X"13",X"C1",X"99",X"D1",X"02",X"E8",X"C8",X"C0",X"05",X"D0",
		X"F4",X"A9",X"00",X"8D",X"D6",X"02",X"CD",X"D9",X"02",X"29",X"01",X"AA",X"BD",X"FF",X"C0",X"8D",
		X"38",X"07",X"AE",X"D7",X"02",X"BD",X"FD",X"C0",X"8D",X"D7",X"02",X"85",X"EF",X"6E",X"AD",X"D0",
		X"02",X"29",X"10",X"D0",X"3B",X"AD",X"D8",X"02",X"4A",X"90",X"09",X"AD",X"D6",X"02",X"4A",X"90",
		X"1F",X"85",X"EF",X"EA",X"AD",X"D3",X"02",X"18",X"6D",X"D1",X"02",X"8D",X"D3",X"02",X"AD",X"D4",
		X"02",X"18",X"6D",X"D2",X"02",X"8D",X"D4",X"02",X"CE",X"D5",X"02",X"F0",X"09",X"85",X"EF",X"EA",
		X"4C",X"D2",X"C0",X"85",X"EF",X"EA",X"AD",X"D0",X"02",X"29",X"20",X"F0",X"09",X"85",X"EF",X"EA",
		X"4C",X"C7",X"C0",X"85",X"EF",X"EA",X"AD",X"D8",X"02",X"0A",X"AA",X"BD",X"27",X"C1",X"85",X"01",
		X"BD",X"28",X"C1",X"85",X"02",X"AD",X"D0",X"02",X"29",X"01",X"AA",X"BC",X"01",X"C1",X"B1",X"01",
		X"8D",X"D1",X"02",X"C8",X"B1",X"01",X"8D",X"D2",X"02",X"C8",X"B1",X"01",X"8D",X"D5",X"02",X"C8",
		X"B1",X"01",X"F0",X"0B",X"AD",X"D0",X"02",X"09",X"20",X"8D",X"D0",X"02",X"85",X"EF",X"EA",X"AD",
		X"D0",X"02",X"09",X"01",X"8D",X"D0",X"02",X"85",X"EF",X"EA",X"AD",X"D9",X"02",X"F0",X"43",X"C9",
		X"01",X"D0",X"11",X"CE",X"D1",X"02",X"AD",X"D1",X"02",X"49",X"FF",X"8D",X"D1",X"02",X"4C",X"D2",
		X"C0",X"85",X"EF",X"EA",X"C9",X"02",X"F0",X"0E",X"CE",X"D1",X"02",X"AD",X"D1",X"02",X"49",X"FF",
		X"8D",X"D1",X"02",X"85",X"EF",X"EA",X"CE",X"D2",X"02",X"AD",X"D2",X"02",X"49",X"FF",X"8D",X"D2",
		X"02",X"4C",X"D2",X"C0",X"85",X"EF",X"EA",X"A9",X"00",X"8D",X"D0",X"02",X"8D",X"38",X"07",X"85",
		X"EF",X"EA",X"AD",X"D6",X"02",X"29",X"38",X"4A",X"4A",X"4A",X"18",X"6D",X"D7",X"02",X"AA",X"BD",
		X"03",X"C1",X"8D",X"39",X"07",X"EE",X"D6",X"02",X"AD",X"D3",X"02",X"18",X"69",X"08",X"49",X"FF",
		X"8D",X"3A",X"07",X"AD",X"D4",X"02",X"38",X"E9",X"08",X"8D",X"3B",X"07",X"60",X"00",X"08",X"81",
		X"83",X"00",X"04",X"2C",X"2D",X"2E",X"2F",X"2F",X"2E",X"2D",X"2C",X"2C",X"2D",X"2E",X"2F",X"2F",
		X"2E",X"2D",X"2C",X"FC",X"00",X"00",X"D8",X"0E",X"04",X"00",X"00",X"D8",X"0E",X"FC",X"00",X"00",
		X"40",X"0C",X"04",X"00",X"00",X"40",X"0C",X"31",X"C1",X"39",X"C1",X"41",X"C1",X"49",X"C1",X"4D",
		X"C1",X"FC",X"FA",X"19",X"00",X"FC",X"00",X"19",X"FF",X"FC",X"FB",X"1E",X"00",X"FC",X"00",X"14",
		X"FF",X"FC",X"FC",X"26",X"00",X"FC",X"00",X"0C",X"FF",X"FC",X"FD",X"32",X"FF",X"FC",X"FE",X"32",
		X"FF",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"64",X"AD",X"D3",X"02",X"85",X"5E",X"CD",X"D4",X"02",
		X"18",X"69",X"06",X"85",X"5F",X"48",X"01",X"20",X"D1",X"B7",X"85",X"EF",X"6E",X"60",X"85",X"EF",
		X"EA",X"A2",X"09",X"85",X"EF",X"6E",X"A9",X"00",X"9D",X"D0",X"02",X"CA",X"10",X"F8",X"60",X"85",
		X"EF",X"EA",X"20",X"8B",X"C1",X"20",X"04",X"A6",X"60",X"85",X"EF",X"EA",X"A5",X"40",X"29",X"FC",
		X"08",X"A5",X"40",X"29",X"03",X"28",X"F0",X"06",X"18",X"69",X"04",X"85",X"EF",X"6E",X"0A",X"AA",
		X"BD",X"CF",X"C1",X"85",X"01",X"DD",X"D0",X"C1",X"85",X"02",X"A0",X"00",X"A2",X"00",X"85",X"EF",
		X"EA",X"A9",X"03",X"85",X"03",X"C1",X"EF",X"6E",X"B1",X"01",X"9D",X"00",X"03",X"64",X"E8",X"C6",
		X"03",X"10",X"F5",X"A9",X"00",X"9D",X"00",X"03",X"E8",X"BD",X"FE",X"02",X"10",X"E3",X"60",X"DF",
		X"C1",X"0B",X"C2",X"47",X"C2",X"8B",X"C2",X"D7",X"C2",X"2B",X"C3",X"7F",X"C3",X"D7",X"C3",X"00",
		X"D8",X"9C",X"02",X"01",X"18",X"7C",X"02",X"00",X"68",X"4C",X"02",X"01",X"38",X"1C",X"02",X"00",
		X"C8",X"EC",X"01",X"00",X"48",X"8C",X"01",X"01",X"C8",X"6C",X"01",X"00",X"38",X"3C",X"01",X"00",
		X"48",X"EC",X"00",X"01",X"98",X"DC",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"B8",X"BC",X"02",X"01",
		X"B8",X"9C",X"02",X"00",X"A8",X"6C",X"02",X"01",X"48",X"6C",X"02",X"01",X"A8",X"0C",X"02",X"03",
		X"78",X"DC",X"01",X"01",X"38",X"DC",X"01",X"01",X"38",X"BC",X"01",X"00",X"B8",X"9C",X"01",X"00",
		X"58",X"5C",X"01",X"03",X"58",X"1C",X"01",X"00",X"C8",X"0C",X"01",X"01",X"B8",X"DC",X"00",X"01",
		X"48",X"CC",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"58",X"DC",X"02",X"02",X"18",X"BC",X"02",X"03",
		X"D8",X"9C",X"02",X"01",X"C8",X"94",X"02",X"01",X"18",X"7C",X"02",X"01",X"D8",X"1C",X"02",X"01",
		X"28",X"F4",X"01",X"02",X"98",X"DC",X"01",X"01",X"D8",X"9C",X"01",X"01",X"58",X"9C",X"01",X"02",
		X"A8",X"6C",X"01",X"03",X"58",X"5C",X"01",X"00",X"D8",X"1C",X"01",X"03",X"28",X"F4",X"00",X"01",
		X"B8",X"DC",X"00",X"02",X"58",X"DC",X"00",X"FF",X"FF",X"FF",X"FF",X"03",X"A8",X"CC",X"02",X"02",
		X"B8",X"BC",X"02",X"00",X"58",X"BC",X"02",X"01",X"18",X"7C",X"02",X"01",X"98",X"5C",X"02",X"02",
		X"78",X"3C",X"02",X"03",X"88",X"2C",X"02",X"02",X"28",X"EC",X"01",X"02",X"B8",X"DC",X"01",X"01",
		X"78",X"BC",X"01",X"01",X"D8",X"9C",X"01",X"00",X"68",X"8C",X"01",X"03",X"48",X"6C",X"01",X"02",
		X"48",X"4C",X"01",X"01",X"98",X"3C",X"01",X"03",X"D8",X"FC",X"00",X"02",X"B8",X"DC",X"00",X"02",
		X"28",X"CC",X"00",X"FF",X"FF",X"FF",X"FF",X"03",X"48",X"CC",X"02",X"02",X"58",X"BC",X"02",X"00",
		X"A8",X"AC",X"02",X"02",X"D8",X"7C",X"02",X"02",X"18",X"7C",X"02",X"03",X"78",X"64",X"02",X"02",
		X"58",X"3C",X"02",X"02",X"48",X"0C",X"02",X"01",X"98",X"FC",X"01",X"03",X"48",X"EC",X"01",X"00",
		X"B8",X"BC",X"01",X"03",X"78",X"A4",X"01",X"01",X"48",X"8C",X"01",X"03",X"C8",X"6C",X"01",X"02",
		X"38",X"64",X"01",X"02",X"A8",X"4C",X"01",X"03",X"B8",X"3C",X"01",X"01",X"88",X"0C",X"01",X"01",
		X"48",X"EC",X"00",X"02",X"98",X"DC",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"D8",X"DC",X"02",X"03",
		X"48",X"CC",X"02",X"02",X"B8",X"9C",X"02",X"03",X"38",X"9C",X"02",X"02",X"38",X"64",X"02",X"02",
		X"38",X"3C",X"02",X"03",X"C8",X"2C",X"02",X"02",X"A8",X"0C",X"02",X"03",X"78",X"DC",X"01",X"02",
		X"38",X"DC",X"01",X"03",X"A8",X"AC",X"01",X"03",X"58",X"9C",X"01",X"01",X"C8",X"8C",X"01",X"02",
		X"88",X"4C",X"01",X"03",X"B8",X"1C",X"01",X"02",X"58",X"04",X"01",X"03",X"38",X"FC",X"00",X"01",
		X"68",X"EC",X"00",X"02",X"B8",X"DC",X"00",X"02",X"48",X"CC",X"00",X"FF",X"FF",X"FF",X"FF",X"03",
		X"A8",X"CC",X"02",X"02",X"18",X"BC",X"02",X"02",X"48",X"B4",X"02",X"02",X"D8",X"9C",X"02",X"03",
		X"C8",X"94",X"02",X"02",X"A8",X"6C",X"02",X"02",X"48",X"4C",X"02",X"03",X"D8",X"1C",X"02",X"02",
		X"28",X"0C",X"02",X"03",X"28",X"F4",X"01",X"01",X"58",X"DC",X"01",X"02",X"48",X"CC",X"01",X"02",
		X"B8",X"BC",X"01",X"03",X"D8",X"9C",X"01",X"01",X"A8",X"6C",X"01",X"02",X"78",X"5C",X"01",X"02",
		X"58",X"3C",X"01",X"03",X"D8",X"1C",X"01",X"02",X"C8",X"14",X"01",X"03",X"38",X"FC",X"00",X"02",
		X"58",X"DC",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"B8",X"DC",X"02",X"02",X"58",X"DC",X"02",X"02",
		X"78",X"BC",X"02",X"03",X"B8",X"9C",X"02",X"02",X"A8",X"8C",X"02",X"03",X"38",X"7C",X"02",X"02",
		X"78",X"3C",X"02",X"03",X"A8",X"2C",X"02",X"03",X"48",X"2C",X"02",X"03",X"88",X"0C",X"02",X"02",
		X"28",X"EC",X"01",X"02",X"28",X"AC",X"01",X"02",X"68",X"8C",X"01",X"02",X"98",X"3C",X"01",X"02",
		X"98",X"1C",X"01",X"03",X"D8",X"FC",X"01",X"02",X"B8",X"DC",X"00",X"02",X"28",X"CC",X"00",X"FF",
		X"FF",X"FF",X"FF",X"85",X"EF",X"EA",X"A5",X"3E",X"29",X"02",X"D0",X"17",X"A5",X"D0",X"D0",X"13",
		X"20",X"46",X"C4",X"20",X"83",X"C4",X"20",X"DE",X"C4",X"20",X"14",X"C5",X"A9",X"00",X"85",X"48",
		X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A6",X"59",X"85",X"EF",X"EA",X"E4",X"5A",X"90",X"04",
		X"60",X"85",X"EF",X"EA",X"BD",X"04",X"03",X"18",X"65",X"48",X"9D",X"04",X"03",X"08",X"A5",X"48",
		X"30",X"16",X"28",X"08",X"B0",X"07",X"C9",X"E8",X"90",X"0E",X"85",X"EF",X"EA",X"BD",X"00",X"03",
		X"09",X"40",X"9D",X"00",X"03",X"85",X"EF",X"EA",X"E8",X"E8",X"E8",X"E8",X"E8",X"28",X"4C",X"4C",
		X"C4",X"85",X"EF",X"EA",X"A6",X"5A",X"85",X"EF",X"EA",X"BD",X"00",X"03",X"A8",X"C9",X"FF",X"F0",
		X"43",X"98",X"30",X"35",X"A5",X"4A",X"38",X"FD",X"02",X"03",X"85",X"01",X"A5",X"4B",X"FD",X"03",
		X"03",X"10",X"0B",X"A9",X"80",X"9D",X"00",X"03",X"4C",X"C9",X"C4",X"85",X"EF",X"EA",X"D0",X"24",
		X"A5",X"01",X"49",X"FF",X"38",X"69",X"00",X"C9",X"34",X"90",X"19",X"9D",X"04",X"03",X"BD",X"00",
		X"03",X"09",X"20",X"9D",X"00",X"03",X"85",X"EF",X"EA",X"E8",X"E8",X"E8",X"E8",X"E8",X"4C",X"89",
		X"C4",X"85",X"EF",X"EA",X"86",X"5A",X"A9",X"00",X"9D",X"04",X"03",X"60",X"85",X"EF",X"EA",X"A6",
		X"59",X"85",X"EF",X"EA",X"BD",X"00",X"03",X"A8",X"C9",X"FF",X"F0",X"23",X"98",X"30",X"12",X"BD",
		X"04",X"03",X"C9",X"E8",X"90",X"19",X"BD",X"00",X"03",X"09",X"40",X"9D",X"00",X"03",X"85",X"EF",
		X"EA",X"98",X"10",X"0B",X"E8",X"E8",X"E8",X"E8",X"E8",X"4C",X"E4",X"C4",X"85",X"EF",X"6E",X"86",
		X"59",X"60",X"85",X"EF",X"6E",X"A6",X"59",X"85",X"EF",X"EA",X"BD",X"00",X"03",X"30",X"30",X"A8",
		X"29",X"60",X"F0",X"2B",X"A9",X"01",X"85",X"0A",X"98",X"29",X"40",X"D0",X"10",X"C6",X"0A",X"DD",
		X"04",X"03",X"C9",X"3C",X"90",X"13",X"29",X"03",X"D0",X"0F",X"85",X"EF",X"6E",X"20",X"5B",X"C5",
		X"C6",X"0A",X"10",X"0B",X"30",X"03",X"85",X"EF",X"EA",X"20",X"E5",X"C5",X"85",X"EF",X"6E",X"E8",
		X"E8",X"E8",X"E8",X"E8",X"E4",X"5A",X"90",X"C2",X"60",X"85",X"EF",X"EA",X"20",X"56",X"C6",X"A5",
		X"0A",X"F0",X"0A",X"BD",X"04",X"03",X"29",X"03",X"D0",X"17",X"85",X"EF",X"6E",X"A5",X"01",X"38",
		X"E9",X"20",X"85",X"01",X"58",X"05",X"C6",X"02",X"85",X"EF",X"EA",X"4C",X"87",X"C5",X"85",X"EF",
		X"EA",X"1E",X"00",X"03",X"C1",X"EF",X"6E",X"A9",X"00",X"A0",X"00",X"20",X"7B",X"C6",X"90",X"05",
		X"91",X"01",X"85",X"EF",X"6E",X"C8",X"20",X"7B",X"C6",X"90",X"05",X"91",X"01",X"C1",X"EF",X"6E",
		X"A5",X"01",X"18",X"69",X"20",X"85",X"01",X"50",X"05",X"E6",X"02",X"85",X"EF",X"6E",X"A9",X"00",
		X"20",X"7B",X"C6",X"90",X"05",X"91",X"01",X"C1",X"EF",X"EA",X"88",X"20",X"7B",X"C6",X"90",X"05",
		X"91",X"01",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"46",X"02",X"46",X"02",X"A2",X"02",X"A2",
		X"02",X"66",X"01",X"46",X"02",X"AA",X"01",X"A2",X"02",X"66",X"01",X"A5",X"02",X"18",X"69",X"10",
		X"85",X"02",X"60",X"85",X"EF",X"6E",X"20",X"56",X"C6",X"BD",X"04",X"03",X"18",X"69",X"04",X"29",
		X"07",X"A8",X"A9",X"FC",X"85",X"EF",X"6E",X"18",X"69",X"04",X"88",X"10",X"FA",X"48",X"DD",X"00",
		X"03",X"29",X"07",X"A8",X"68",X"18",X"79",X"4F",X"C6",X"A0",X"00",X"20",X"7B",X"C6",X"90",X"05",
		X"91",X"01",X"85",X"EF",X"EA",X"18",X"69",X"01",X"C8",X"20",X"7B",X"C6",X"90",X"05",X"91",X"01",
		X"85",X"EF",X"EA",X"48",X"A5",X"01",X"18",X"69",X"20",X"85",X"01",X"90",X"05",X"E6",X"02",X"85",
		X"EF",X"EA",X"68",X"18",X"69",X"02",X"20",X"7B",X"C6",X"90",X"05",X"91",X"01",X"85",X"EF",X"EA",
		X"88",X"38",X"E9",X"01",X"20",X"7B",X"C6",X"90",X"05",X"91",X"01",X"85",X"EF",X"EA",X"60",X"40",
		X"60",X"80",X"A0",X"80",X"85",X"EF",X"EA",X"BD",X"01",X"03",X"85",X"01",X"BD",X"04",X"03",X"85",
		X"02",X"48",X"20",X"C8",X"C5",X"68",X"29",X"04",X"D0",X"0E",X"A5",X"01",X"38",X"E9",X"20",X"85",
		X"01",X"B0",X"05",X"C6",X"02",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"48",X"B1",X"01",X"F0",
		X"0B",X"C9",X"40",X"90",X"0D",X"C9",X"C0",X"B0",X"09",X"85",X"EF",X"EA",X"38",X"68",X"60",X"85",
		X"EF",X"EA",X"18",X"68",X"60",X"85",X"EF",X"EA",X"A5",X"3E",X"29",X"03",X"AA",X"F0",X"65",X"A5",
		X"DF",X"29",X"0F",X"D0",X"15",X"A9",X"80",X"85",X"DF",X"E0",X"01",X"D0",X"08",X"A5",X"40",X"D0",
		X"04",X"AA",X"85",X"EF",X"EA",X"86",X"E1",X"85",X"EF",X"EA",X"A5",X"E1",X"0A",X"AA",X"BD",X"13",
		X"C7",X"85",X"01",X"BD",X"14",X"C7",X"85",X"02",X"A9",X"C6",X"48",X"A9",X"D5",X"48",X"6C",X"01",
		X"00",X"EA",X"EA",X"85",X"EF",X"EA",X"A5",X"DF",X"30",X"2A",X"A5",X"3E",X"29",X"02",X"F0",X"28",
		X"A9",X"00",X"8D",X"20",X"07",X"8D",X"00",X"18",X"85",X"9F",X"A9",X"38",X"8D",X"01",X"0C",X"A9",
		X"C0",X"85",X"1D",X"85",X"EF",X"EA",X"A5",X"3E",X"29",X"FC",X"85",X"3E",X"A9",X"42",X"20",X"86",
		X"D3",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A9",X"00",X"85",X"C7",X"4D",X"80",X"85",X"D7",
		X"4C",X"F6",X"C6",X"BD",X"C7",X"F4",X"C9",X"F7",X"C9",X"85",X"EF",X"EA",X"C6",X"DD",X"10",X"0E",
		X"AD",X"44",X"C7",X"85",X"DD",X"C9",X"DF",X"49",X"20",X"85",X"DF",X"85",X"EF",X"6E",X"A5",X"DF",
		X"29",X"20",X"4A",X"4A",X"4A",X"4A",X"4A",X"AA",X"A5",X"DB",X"18",X"7D",X"45",X"C7",X"85",X"DB",
		X"85",X"EF",X"EA",X"60",X"05",X"FF",X"01",X"85",X"EF",X"EA",X"A5",X"DC",X"18",X"69",X"10",X"49",
		X"FF",X"85",X"01",X"A2",X"03",X"85",X"EF",X"6E",X"8A",X"0A",X"0A",X"A8",X"A5",X"01",X"38",X"FD",
		X"72",X"C7",X"99",X"26",X"07",X"C9",X"DB",X"38",X"FD",X"76",X"C7",X"99",X"27",X"07",X"66",X"10",
		X"E7",X"60",X"10",X"20",X"10",X"00",X"04",X"00",X"00",X"00",X"85",X"EF",X"6E",X"C6",X"DE",X"10",
		X"2F",X"AD",X"B1",X"C7",X"85",X"DE",X"C9",X"DF",X"49",X"40",X"85",X"DF",X"0D",X"40",X"4A",X"4A",
		X"4A",X"4A",X"4A",X"4A",X"AA",X"BD",X"B2",X"C7",X"8D",X"31",X"07",X"BD",X"B4",X"C7",X"8D",X"2D",
		X"07",X"BD",X"B6",X"C7",X"8D",X"29",X"07",X"DD",X"B8",X"C7",X"8D",X"25",X"07",X"C1",X"EF",X"6E",
		X"60",X"04",X"1A",X"1B",X"1C",X"1D",X"1A",X"1B",X"00",X"00",X"85",X"EF",X"6E",X"A5",X"D9",X"D0",
		X"24",X"A5",X"DF",X"10",X"20",X"29",X"0F",X"0A",X"AA",X"BD",X"E6",X"C7",X"85",X"01",X"DD",X"E7",
		X"C7",X"85",X"02",X"A9",X"C7",X"48",X"4D",X"DE",X"48",X"6C",X"01",X"00",X"85",X"EF",X"6E",X"20",
		X"B3",X"C8",X"85",X"EF",X"6E",X"60",X"DF",X"C8",X"F3",X"C7",X"24",X"C8",X"75",X"C8",X"92",X"C8",
		X"85",X"EF",X"EA",X"A2",X"06",X"85",X"EF",X"6E",X"8A",X"0A",X"0A",X"A8",X"BD",X"1A",X"C8",X"99",
		X"25",X"07",X"CA",X"10",X"F3",X"A9",X"81",X"8D",X"24",X"07",X"A9",X"85",X"8D",X"30",X"07",X"A9",
		X"30",X"85",X"DB",X"A9",X"F8",X"85",X"DC",X"E6",X"DF",X"60",X"1E",X"1F",X"1E",X"1E",X"1F",X"1E",
		X"20",X"85",X"EF",X"EA",X"A5",X"DB",X"18",X"6D",X"71",X"C8",X"85",X"DB",X"A5",X"DC",X"38",X"ED",
		X"70",X"C8",X"85",X"DC",X"C9",X"E8",X"B0",X"37",X"A9",X"81",X"8D",X"28",X"07",X"A9",X"81",X"8D",
		X"34",X"07",X"A9",X"81",X"8D",X"3C",X"07",X"A9",X"21",X"8D",X"35",X"07",X"A9",X"22",X"8D",X"3D",
		X"07",X"8A",X"49",X"FF",X"2D",X"20",X"07",X"8D",X"20",X"07",X"A5",X"DC",X"C9",X"D8",X"B0",X"0F",
		X"A9",X"83",X"8D",X"2C",X"07",X"A9",X"87",X"8D",X"38",X"07",X"E6",X"DF",X"85",X"EF",X"EA",X"60",
		X"04",X"02",X"85",X"EF",X"EA",X"A5",X"DB",X"18",X"6D",X"71",X"C8",X"85",X"DB",X"A5",X"DC",X"38",
		X"ED",X"70",X"C8",X"85",X"DC",X"C9",X"58",X"B0",X"05",X"E6",X"DF",X"85",X"EF",X"EA",X"60",X"85",
		X"EF",X"EA",X"A0",X"80",X"84",X"9D",X"20",X"9E",X"A7",X"20",X"08",X"C9",X"A9",X"00",X"85",X"E0",
		X"85",X"DF",X"60",X"00",X"F0",X"E0",X"00",X"F0",X"E0",X"F0",X"00",X"00",X"00",X"10",X"10",X"10",
		X"20",X"85",X"EF",X"EA",X"A5",X"DC",X"18",X"69",X"10",X"49",X"FF",X"85",X"01",X"A2",X"06",X"85",
		X"EF",X"EA",X"8A",X"0A",X"0A",X"A8",X"BD",X"A3",X"C8",X"18",X"65",X"01",X"99",X"26",X"07",X"BD",
		X"AA",X"C8",X"18",X"65",X"DB",X"99",X"27",X"07",X"CA",X"10",X"E7",X"60",X"85",X"EF",X"EA",X"A9",
		X"C1",X"20",X"86",X"D3",X"20",X"08",X"C9",X"20",X"A0",X"A4",X"20",X"B2",X"B3",X"A9",X"F8",X"8D",
		X"01",X"0C",X"A2",X"46",X"A5",X"3E",X"29",X"01",X"F0",X"05",X"A2",X"41",X"85",X"EF",X"EA",X"8A",
		X"20",X"86",X"D3",X"E6",X"DF",X"28",X"85",X"EF",X"EA",X"A2",X"1F",X"A9",X"00",X"85",X"EF",X"6E",
		X"9D",X"20",X"07",X"CA",X"10",X"FA",X"60",X"85",X"EF",X"EA",X"A2",X"00",X"85",X"EF",X"6E",X"A9",
		X"00",X"9D",X"00",X"18",X"6C",X"E0",X"20",X"D0",X"F6",X"60",X"85",X"EF",X"6E",X"A5",X"3E",X"29",
		X"02",X"F0",X"45",X"A5",X"E4",X"D0",X"10",X"20",X"B8",X"A5",X"A9",X"00",X"85",X"9D",X"C1",X"A3",
		X"A9",X"01",X"85",X"A4",X"C1",X"EF",X"6E",X"A5",X"DA",X"D0",X"32",X"A9",X"10",X"85",X"DA",X"08",
		X"08",X"C9",X"20",X"A0",X"A4",X"A5",X"E3",X"F0",X"06",X"20",X"80",X"C9",X"85",X"EF",X"6E",X"A5",
		X"E3",X"49",X"01",X"85",X"E3",X"EA",X"E4",X"C9",X"E4",X"C9",X"0F",X"90",X"10",X"A5",X"0A",X"18",
		X"69",X"09",X"20",X"DE",X"D2",X"85",X"EF",X"6E",X"E6",X"DF",X"85",X"EF",X"6E",X"60",X"85",X"EF",
		X"EA",X"A5",X"E5",X"C9",X"C0",X"90",X"06",X"38",X"E9",X"08",X"85",X"EF",X"6E",X"85",X"02",X"4D",
		X"40",X"85",X"01",X"20",X"C8",X"C5",X"A0",X"04",X"85",X"EF",X"EA",X"B9",X"D8",X"C9",X"91",X"01",
		X"88",X"10",X"F8",X"A2",X"00",X"A5",X"E5",X"85",X"EF",X"EA",X"DD",X"D3",X"C9",X"B0",X"06",X"E8",
		X"10",X"F8",X"85",X"EF",X"6E",X"86",X"0A",X"46",X"0A",X"0A",X"AA",X"A5",X"01",X"18",X"69",X"0C",
		X"85",X"01",X"A0",X"00",X"85",X"EF",X"6E",X"BD",X"DD",X"C9",X"91",X"01",X"6C",X"C8",X"C0",X"04",
		X"90",X"F5",X"60",X"A8",X"78",X"58",X"48",X"00",X"0C",X"19",X"18",X"1F",X"1D",X"02",X"01",X"01",
		X"01",X"02",X"06",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"06",X"01",X"01",X"04",X"01",X"01",
		X"01",X"85",X"EF",X"EA",X"85",X"EF",X"6E",X"A5",X"DF",X"10",X"0A",X"29",X"0F",X"D0",X"0A",X"20",
		X"DE",X"C8",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"C9",X"01",X"D0",X"07",X"20",X"2C",X"C9",
		X"60",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"DF",X"A9",X"80",X"85",X"9D",X"20",X"9E",X"A7",X"60",
		X"85",X"EF",X"EA",X"A5",X"7B",X"29",X"18",X"F0",X"14",X"A9",X"00",X"85",X"E8",X"8D",X"3C",X"07",
		X"8D",X"3D",X"07",X"8D",X"3E",X"07",X"8D",X"3F",X"07",X"60",X"85",X"EF",X"EA",X"A5",X"B2",X"F0",
		X"01",X"60",X"A5",X"3E",X"29",X"03",X"F0",X"01",X"60",X"24",X"E8",X"50",X"01",X"60",X"10",X"64",
		X"A2",X"08",X"85",X"EF",X"EA",X"BD",X"9E",X"B4",X"85",X"01",X"BD",X"9F",X"B4",X"85",X"02",X"A0",
		X"00",X"B1",X"01",X"29",X"04",X"F0",X"12",X"A0",X"03",X"B1",X"01",X"45",X"E9",X"D0",X"0A",X"C8",
		X"B1",X"01",X"45",X"EA",X"F0",X"60",X"85",X"EF",X"EA",X"CA",X"CA",X"10",X"D8",X"85",X"EF",X"EA",
		X"A2",X"00",X"A5",X"E8",X"29",X"01",X"F0",X"04",X"E8",X"85",X"EF",X"EA",X"AD",X"03",X"40",X"F0",
		X"09",X"A5",X"12",X"F0",X"05",X"E8",X"E8",X"85",X"EF",X"EA",X"BD",X"D7",X"CA",X"8D",X"3C",X"07",
		X"A5",X"E9",X"18",X"7D",X"DB",X"CA",X"49",X"FF",X"8D",X"3E",X"07",X"A5",X"E8",X"29",X"F0",X"85",
		X"E8",X"85",X"EF",X"EA",X"A9",X"28",X"8D",X"3D",X"07",X"A5",X"EA",X"38",X"E9",X"0F",X"8D",X"3F",
		X"07",X"A5",X"E8",X"29",X"0F",X"85",X"E8",X"AD",X"3F",X"07",X"C9",X"E0",X"90",X"08",X"A9",X"00",
		X"8D",X"3C",X"07",X"85",X"EF",X"EA",X"60",X"01",X"03",X"01",X"03",X"08",X"0A",X"06",X"08",X"85",
		X"EF",X"EA",X"20",X"05",X"CB",X"85",X"EF",X"EA",X"20",X"2A",X"CB",X"20",X"2A",X"CC",X"A5",X"5B",
		X"29",X"01",X"F0",X"0E",X"20",X"BE",X"CC",X"90",X"09",X"20",X"25",X"CD",X"4C",X"E8",X"CA",X"85",
		X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A5",X"5D",X"AA",X"E8",X"BD",X"1E",X"CB",X"18",X"65",X"5E",
		X"85",X"60",X"BD",X"23",X"CB",X"18",X"65",X"5F",X"85",X"61",X"85",X"EF",X"6E",X"60",X"00",X"02",
		X"02",X"FE",X"FE",X"00",X"FF",X"01",X"01",X"FF",X"85",X"EF",X"EA",X"A5",X"61",X"49",X"FF",X"85",
		X"01",X"A5",X"4A",X"38",X"E5",X"01",X"48",X"0D",X"F0",X"85",X"4F",X"A5",X"4B",X"E9",X"00",X"85",
		X"50",X"E6",X"50",X"68",X"29",X"0F",X"85",X"02",X"A5",X"60",X"4A",X"4A",X"4A",X"4A",X"05",X"4F",
		X"A8",X"A5",X"4C",X"29",X"0C",X"05",X"50",X"0A",X"AA",X"BD",X"CB",X"CB",X"85",X"4F",X"DD",X"CC",
		X"CB",X"85",X"50",X"B1",X"4F",X"85",X"58",X"65",X"01",X"D0",X"09",X"A5",X"5B",X"09",X"02",X"85",
		X"5B",X"85",X"EF",X"EA",X"A9",X"20",X"85",X"57",X"20",X"FD",X"CB",X"A9",X"00",X"85",X"05",X"4A",
		X"02",X"85",X"EF",X"EA",X"A5",X"55",X"85",X"51",X"A5",X"56",X"18",X"7D",X"EB",X"CB",X"85",X"52",
		X"A0",X"00",X"A5",X"02",X"C9",X"08",X"90",X"04",X"C8",X"85",X"EF",X"EA",X"29",X"07",X"85",X"03",
		X"A5",X"60",X"29",X"0F",X"19",X"EE",X"CB",X"85",X"04",X"A4",X"03",X"B9",X"F0",X"CB",X"85",X"03",
		X"A4",X"04",X"B1",X"51",X"25",X"03",X"F0",X"0B",X"A5",X"05",X"18",X"7D",X"F8",X"CB",X"85",X"05",
		X"85",X"EF",X"EA",X"CA",X"10",X"BE",X"A5",X"05",X"85",X"66",X"60",X"00",X"E6",X"00",X"E7",X"00",
		X"E8",X"00",X"E9",X"00",X"EA",X"00",X"EB",X"00",X"EC",X"00",X"ED",X"00",X"EE",X"00",X"EF",X"00",
		X"F0",X"00",X"F1",X"00",X"F2",X"00",X"F3",X"00",X"F4",X"00",X"F5",X"E0",X"E2",X"E4",X"00",X"10",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"01",X"02",X"04",X"85",X"EF",X"6E",X"A9",X"08",
		X"85",X"06",X"A9",X"00",X"85",X"55",X"85",X"56",X"85",X"EF",X"EA",X"06",X"55",X"26",X"56",X"06",
		X"58",X"90",X"10",X"18",X"A5",X"57",X"65",X"55",X"85",X"55",X"A5",X"56",X"69",X"00",X"85",X"56",
		X"85",X"EF",X"EA",X"C6",X"06",X"D0",X"E4",X"60",X"85",X"EF",X"EA",X"A6",X"66",X"BD",X"33",X"CC",
		X"85",X"67",X"60",X"02",X"02",X"01",X"02",X"02",X"01",X"03",X"00",X"85",X"EF",X"EA",X"A5",X"67",
		X"F0",X"15",X"C9",X"01",X"F0",X"29",X"C9",X"02",X"F0",X"44",X"C9",X"03",X"F0",X"50",X"D0",X"3E",
		X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"C6",X"6A",X"10",X"07",X"A9",X"00",X"85",X"6A",X"85",
		X"EF",X"EA",X"A5",X"5D",X"30",X"05",X"85",X"5C",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A0",
		X"00",X"A6",X"5D",X"E8",X"8A",X"29",X"02",X"F0",X"04",X"C8",X"85",X"EF",X"EA",X"A5",X"61",X"18",
		X"79",X"89",X"CC",X"85",X"61",X"C8",X"84",X"64",X"60",X"F8",X"08",X"85",X"EF",X"EA",X"A5",X"5E",
		X"85",X"60",X"A5",X"5F",X"85",X"61",X"A9",X"02",X"85",X"67",X"60",X"85",X"EF",X"EA",X"A0",X"60",
		X"20",X"E9",X"A8",X"A5",X"BA",X"C5",X"B9",X"F0",X"0A",X"A9",X"04",X"05",X"5B",X"85",X"5B",X"60",
		X"85",X"EF",X"EA",X"A5",X"62",X"09",X"80",X"85",X"62",X"4C",X"8E",X"CC",X"85",X"EF",X"EA",X"A9",
		X"0F",X"85",X"03",X"A9",X"CD",X"85",X"04",X"A9",X"17",X"85",X"05",X"A9",X"CD",X"85",X"06",X"A2",
		X"07",X"85",X"EF",X"EA",X"A5",X"5B",X"29",X"FE",X"85",X"5B",X"8A",X"A8",X"85",X"EF",X"EA",X"A5",
		X"5E",X"18",X"71",X"03",X"85",X"01",X"29",X"0F",X"F0",X"08",X"88",X"10",X"F2",X"18",X"60",X"85",
		X"EF",X"EA",X"8A",X"A8",X"85",X"EF",X"EA",X"A5",X"5F",X"18",X"71",X"05",X"85",X"02",X"18",X"65",
		X"49",X"29",X"07",X"F0",X"08",X"88",X"10",X"EF",X"18",X"60",X"85",X"EF",X"6E",X"38",X"60",X"FA",
		X"FC",X"FE",X"00",X"02",X"04",X"06",X"08",X"FD",X"FE",X"FF",X"00",X"01",X"02",X"03",X"04",X"00",
		X"02",X"00",X"01",X"85",X"EF",X"6E",X"A5",X"5D",X"0A",X"AA",X"A5",X"01",X"38",X"FD",X"3B",X"CD",
		X"85",X"60",X"A5",X"02",X"38",X"FD",X"3C",X"CD",X"85",X"61",X"60",X"00",X"01",X"00",X"00",X"02",
		X"00",X"02",X"01",X"85",X"EF",X"6E",X"A2",X"1C",X"A0",X"07",X"85",X"EF",X"6E",X"98",X"0A",X"0A",
		X"0A",X"9D",X"B0",X"02",X"44",X"CA",X"CA",X"CA",X"CA",X"10",X"F2",X"60",X"85",X"EF",X"6E",X"A0",
		X"1C",X"85",X"EF",X"EA",X"B9",X"B0",X"02",X"29",X"38",X"48",X"29",X"7F",X"4A",X"AA",X"68",X"1D",
		X"20",X"07",X"99",X"B0",X"02",X"DD",X"21",X"07",X"99",X"B1",X"02",X"BD",X"22",X"07",X"99",X"B2",
		X"02",X"BD",X"23",X"07",X"99",X"B3",X"02",X"44",X"88",X"88",X"88",X"10",X"D7",X"85",X"EF",X"6E",
		X"A9",X"00",X"85",X"01",X"4A",X"1C",X"85",X"EF",X"EA",X"BD",X"B0",X"02",X"5D",X"AC",X"02",X"30",
		X"2E",X"A0",X"00",X"BD",X"B0",X"02",X"29",X"03",X"F0",X"07",X"98",X"09",X"04",X"A8",X"85",X"EF",
		X"EA",X"BD",X"AC",X"02",X"29",X"03",X"F0",X"07",X"98",X"09",X"02",X"A8",X"85",X"EF",X"6E",X"B9",
		X"39",X"CE",X"85",X"03",X"5D",X"3A",X"CE",X"85",X"04",X"6C",X"03",X"00",X"85",X"EF",X"6E",X"BD",
		X"B0",X"02",X"30",X"4E",X"10",X"0E",X"85",X"EF",X"EA",X"BD",X"B3",X"02",X"DD",X"AF",X"02",X"B0",
		X"41",X"85",X"EF",X"EA",X"BD",X"B0",X"02",X"48",X"BD",X"AC",X"02",X"9D",X"B0",X"02",X"2C",X"9D",
		X"AC",X"02",X"BD",X"B1",X"02",X"48",X"DD",X"AD",X"02",X"9D",X"B1",X"02",X"2C",X"9D",X"AD",X"02",
		X"BD",X"B2",X"02",X"48",X"BD",X"AE",X"02",X"9D",X"B2",X"02",X"68",X"9D",X"AE",X"02",X"BD",X"B3",
		X"02",X"48",X"BD",X"AF",X"02",X"9D",X"B3",X"02",X"68",X"9D",X"AF",X"02",X"38",X"66",X"01",X"85",
		X"EF",X"EA",X"CA",X"CA",X"CA",X"CA",X"D0",X"0E",X"A5",X"01",X"10",X"06",X"4C",X"90",X"CD",X"85",
		X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"4C",X"99",X"CD",X"22",X"CE",X"22",X"CE",X"E4",X"CD",X"D9",
		X"CD",X"85",X"EF",X"EA",X"A5",X"40",X"29",X"03",X"0A",X"85",X"01",X"A2",X"1F",X"85",X"EF",X"EA",
		X"A9",X"00",X"85",X"02",X"8A",X"29",X"03",X"C9",X"01",X"D0",X"1D",X"A4",X"01",X"BD",X"B0",X"02",
		X"C9",X"30",X"90",X"14",X"C9",X"B0",X"90",X"08",X"C9",X"FF",X"F0",X"0C",X"C8",X"85",X"EF",X"EA",
		X"B9",X"85",X"CE",X"85",X"02",X"85",X"EF",X"EA",X"BD",X"B0",X"02",X"18",X"65",X"02",X"9D",X"00",
		X"18",X"CA",X"10",X"CC",X"60",X"00",X"00",X"20",X"10",X"40",X"20",X"60",X"30",X"80",X"40",X"85",
		X"EF",X"EA",X"A9",X"FC",X"85",X"1A",X"A9",X"38",X"85",X"1B",X"60",X"85",X"EF",X"EA",X"A5",X"1A",
		X"38",X"65",X"1B",X"85",X"1A",X"38",X"65",X"1B",X"85",X"1B",X"60",X"85",X"EF",X"EA",X"A2",X"3F",
		X"A9",X"3B",X"85",X"EF",X"EA",X"9D",X"C0",X"13",X"CA",X"10",X"FA",X"20",X"EB",X"CF",X"20",X"19",
		X"C9",X"60",X"85",X"EF",X"EA",X"A2",X"01",X"85",X"EF",X"EA",X"A9",X"2F",X"85",X"EF",X"EA",X"9D",
		X"00",X"10",X"E8",X"E0",X"E0",X"D0",X"F8",X"20",X"EB",X"CF",X"20",X"19",X"C9",X"60",X"85",X"EF",
		X"EA",X"A2",X"1F",X"85",X"EF",X"EA",X"8A",X"29",X"01",X"A8",X"B9",X"F4",X"CE",X"9D",X"A0",X"13",
		X"CA",X"D0",X"F3",X"60",X"37",X"39",X"85",X"EF",X"EA",X"A5",X"D5",X"D0",X"35",X"AE",X"BF",X"13",
		X"E8",X"E0",X"3B",X"D0",X"05",X"A2",X"37",X"85",X"EF",X"EA",X"8E",X"BF",X"13",X"CE",X"BE",X"13",
		X"E8",X"E0",X"3B",X"D0",X"05",X"A2",X"37",X"85",X"EF",X"EA",X"8E",X"BE",X"13",X"4A",X"1F",X"85",
		X"EF",X"EA",X"8A",X"29",X"01",X"A8",X"B9",X"BE",X"13",X"9D",X"A0",X"13",X"66",X"D0",X"F3",X"85",
		X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A5",X"7B",X"F0",X"0F",X"29",X"18",X"D0",X"0B",X"A5",X"3E",
		X"4A",X"B0",X"06",X"20",X"4C",X"CF",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A9",X"00",X"85",
		X"03",X"A5",X"3E",X"29",X"82",X"D0",X"39",X"A9",X"FF",X"38",X"E5",X"7F",X"85",X"01",X"C9",X"4A",
		X"38",X"E5",X"01",X"85",X"01",X"C9",X"4B",X"E9",X"00",X"85",X"02",X"A5",X"01",X"38",X"E9",X"C0",
		X"48",X"A5",X"02",X"E9",X"00",X"AA",X"68",X"4A",X"4A",X"4A",X"1D",X"A8",X"CF",X"85",X"02",X"4D",
		X"00",X"85",X"03",X"A2",X"FF",X"85",X"EF",X"6E",X"E8",X"E0",X"08",X"D0",X"0A",X"85",X"EF",X"6E",
		X"20",X"B5",X"CF",X"60",X"85",X"EF",X"6E",X"46",X"02",X"90",X"ED",X"F8",X"A5",X"03",X"18",X"7D",
		X"AC",X"CF",X"85",X"03",X"74",X"4C",X"88",X"CF",X"00",X"20",X"40",X"60",X"01",X"02",X"04",X"08",
		X"16",X"32",X"64",X"85",X"EF",X"6E",X"A9",X"99",X"85",X"04",X"A9",X"10",X"85",X"05",X"C9",X"03",
		X"48",X"4A",X"4A",X"4A",X"4A",X"48",X"48",X"00",X"85",X"EF",X"EA",X"68",X"29",X"0F",X"D0",X"06",
		X"B9",X"E6",X"CF",X"85",X"EF",X"6E",X"18",X"69",X"01",X"91",X"04",X"C8",X"C0",X"02",X"D0",X"EB",
		X"B9",X"E6",X"CF",X"91",X"04",X"28",X"2E",X"00",X"01",X"85",X"EF",X"EA",X"A9",X"78",X"85",X"01",
		X"A9",X"10",X"85",X"02",X"4A",X"00",X"85",X"EF",X"EA",X"A0",X"00",X"85",X"EF",X"6E",X"BD",X"15",
		X"D0",X"91",X"01",X"E8",X"C8",X"C0",X"06",X"D0",X"F5",X"A5",X"01",X"18",X"69",X"20",X"85",X"01",
		X"C9",X"D8",X"D0",X"E5",X"60",X"28",X"2C",X"2C",X"2C",X"2C",X"29",X"2D",X"2F",X"2F",X"2F",X"2E",
		X"2D",X"2A",X"2C",X"2C",X"2C",X"2C",X"2B",X"85",X"EF",X"EA",X"A2",X"16",X"A0",X"02",X"4C",X"3B",
		X"D0",X"85",X"EF",X"EA",X"A2",X"44",X"A4",X"12",X"85",X"EF",X"EA",X"B9",X"63",X"D0",X"85",X"01",
		X"A9",X"10",X"85",X"02",X"A9",X"03",X"85",X"03",X"A9",X"05",X"85",X"04",X"85",X"EF",X"EA",X"B5",
		X"00",X"48",X"4A",X"4A",X"4A",X"4A",X"20",X"68",X"D0",X"68",X"20",X"68",X"D0",X"CA",X"C6",X"03",
		X"D0",X"ED",X"60",X"42",X"58",X"4D",X"85",X"EF",X"EA",X"29",X"0F",X"D0",X"17",X"A4",X"04",X"F0",
		X"1A",X"C6",X"04",X"D0",X"1C",X"85",X"EF",X"EA",X"48",X"A0",X"00",X"84",X"04",X"68",X"4C",X"8B",
		X"D0",X"85",X"EF",X"EA",X"A4",X"04",X"D0",X"F0",X"85",X"EF",X"EA",X"18",X"69",X"01",X"85",X"EF",
		X"EA",X"A0",X"00",X"48",X"68",X"D0",X"05",X"A9",X"2F",X"85",X"EF",X"EA",X"91",X"01",X"E6",X"01",
		X"D0",X"05",X"E6",X"02",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"40",X"29",X"03",X"0A",
		X"AA",X"BD",X"30",X"D1",X"85",X"01",X"BD",X"31",X"D1",X"85",X"02",X"A9",X"00",X"AA",X"85",X"06",
		X"85",X"EF",X"EA",X"A0",X"01",X"B1",X"01",X"85",X"03",X"C8",X"B1",X"01",X"30",X"51",X"85",X"04",
		X"A5",X"4A",X"38",X"E5",X"03",X"85",X"05",X"A5",X"4B",X"E5",X"04",X"30",X"2D",X"29",X"03",X"D0",
		X"3E",X"A5",X"05",X"49",X"FF",X"C5",X"09",X"90",X"21",X"C5",X"0A",X"B0",X"1D",X"9D",X"02",X"04",
		X"A0",X"00",X"B1",X"01",X"9D",X"01",X"04",X"A0",X"03",X"B1",X"01",X"9D",X"03",X"04",X"A5",X"06",
		X"9D",X"00",X"04",X"E8",X"E8",X"E8",X"E8",X"85",X"EF",X"EA",X"A5",X"01",X"18",X"69",X"04",X"85",
		X"01",X"A5",X"02",X"69",X"00",X"85",X"02",X"EA",X"06",X"4C",X"C3",X"D0",X"85",X"EF",X"6E",X"86",
		X"CC",X"A9",X"FF",X"9D",X"00",X"04",X"D5",X"01",X"04",X"9D",X"02",X"04",X"D5",X"03",X"04",X"28",
		X"38",X"D1",X"A4",X"D1",X"0C",X"D2",X"74",X"D2",X"B6",X"C3",X"02",X"01",X"48",X"C3",X"02",X"02",
		X"28",X"A3",X"02",X"02",X"A6",X"93",X"02",X"01",X"58",X"93",X"02",X"02",X"A6",X"73",X"02",X"01",
		X"58",X"53",X"02",X"02",X"B6",X"43",X"02",X"01",X"88",X"43",X"02",X"02",X"68",X"23",X"02",X"02",
		X"86",X"F3",X"01",X"01",X"B6",X"E3",X"01",X"01",X"76",X"C3",X"01",X"01",X"48",X"C3",X"01",X"02",
		X"A6",X"B3",X"01",X"01",X"68",X"A3",X"01",X"02",X"96",X"83",X"01",X"01",X"A8",X"63",X"01",X"02",
		X"56",X"63",X"01",X"01",X"A6",X"33",X"01",X"01",X"86",X"33",X"01",X"01",X"78",X"13",X"01",X"02",
		X"A6",X"F3",X"00",X"01",X"86",X"F3",X"00",X"01",X"78",X"F3",X"00",X"02",X"78",X"D3",X"00",X"02",
		X"FF",X"FF",X"FF",X"FF",X"86",X"D3",X"02",X"01",X"56",X"C3",X"02",X"01",X"28",X"C3",X"02",X"02",
		X"68",X"A3",X"02",X"02",X"56",X"A3",X"02",X"01",X"B6",X"83",X"02",X"01",X"48",X"83",X"02",X"02",
		X"B8",X"53",X"02",X"02",X"66",X"33",X"02",X"01",X"46",X"33",X"02",X"01",X"B6",X"23",X"02",X"01",
		X"58",X"13",X"02",X"02",X"58",X"F3",X"01",X"02",X"C8",X"C3",X"01",X"02",X"A8",X"C3",X"01",X"02",
		X"58",X"93",X"01",X"02",X"38",X"73",X"01",X"02",X"96",X"63",X"01",X"01",X"C8",X"43",X"01",X"02",
		X"88",X"23",X"01",X"02",X"48",X"23",X"01",X"02",X"56",X"03",X"01",X"01",X"B8",X"F3",X"00",X"02",
		X"48",X"E3",X"00",X"02",X"78",X"D3",X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"C6",X"D3",X"02",X"01",
		X"58",X"D3",X"02",X"02",X"98",X"B3",X"02",X"02",X"46",X"B3",X"02",X"01",X"86",X"93",X"02",X"01",
		X"66",X"93",X"02",X"01",X"98",X"73",X"02",X"02",X"66",X"73",X"02",X"01",X"86",X"53",X"02",X"01",
		X"A6",X"33",X"02",X"01",X"78",X"33",X"02",X"02",X"A6",X"13",X"02",X"01",X"86",X"13",X"02",X"01",
		X"78",X"F3",X"01",X"02",X"66",X"D3",X"01",X"01",X"86",X"B3",X"01",X"01",X"98",X"73",X"01",X"02",
		X"66",X"73",X"01",X"01",X"78",X"53",X"01",X"02",X"86",X"33",X"01",X"01",X"A6",X"13",X"01",X"01",
		X"78",X"13",X"01",X"02",X"B8",X"F3",X"00",X"02",X"86",X"F3",X"00",X"01",X"86",X"D3",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"D6",X"C3",X"02",X"01",X"96",X"C3",X"02",X"01",X"28",X"C3",X"02",X"02",
		X"66",X"B3",X"02",X"01",X"A8",X"A3",X"02",X"02",X"48",X"A3",X"02",X"02",X"56",X"83",X"02",X"01",
		X"C6",X"73",X"02",X"01",X"38",X"53",X"02",X"02",X"88",X"23",X"02",X"02",X"76",X"23",X"02",X"01",
		X"36",X"23",X"02",X"01",X"B8",X"13",X"02",X"02",X"36",X"C3",X"01",X"01",X"C8",X"A3",X"01",X"02",
		X"C8",X"63",X"01",X"02",X"B6",X"63",X"01",X"01",X"56",X"63",X"01",X"01",X"48",X"63",X"01",X"02",
		X"B8",X"33",X"01",X"02",X"38",X"33",X"01",X"02",X"86",X"13",X"01",X"01",X"36",X"03",X"01",X"01",
		X"C6",X"F3",X"00",X"01",X"78",X"D3",X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"85",X"EF",X"EA",X"0A",
		X"AA",X"F8",X"BD",X"F9",X"D2",X"18",X"65",X"42",X"85",X"42",X"BD",X"FA",X"D2",X"65",X"43",X"85",
		X"43",X"A5",X"44",X"69",X"00",X"85",X"44",X"D8",X"60",X"04",X"00",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"05",X"00",X"06",X"00",X"08",X"00",X"04",X"00",X"12",X"00",X"10",X"00",X"15",X"00",
		X"20",X"00",X"25",X"00",X"30",X"85",X"EF",X"6E",X"A5",X"3E",X"29",X"20",X"D0",X"24",X"F8",X"A5",
		X"42",X"38",X"E5",X"17",X"A5",X"43",X"E5",X"18",X"A5",X"44",X"E5",X"19",X"D8",X"90",X"13",X"E6",
		X"3F",X"20",X"75",X"D4",X"A9",X"20",X"05",X"3E",X"85",X"3E",X"A9",X"0F",X"20",X"86",X"D3",X"85",
		X"EF",X"EA",X"60",X"85",X"EF",X"6E",X"A5",X"10",X"F0",X"1F",X"A5",X"14",X"F8",X"38",X"E5",X"42",
		X"A5",X"15",X"E5",X"43",X"A5",X"16",X"E5",X"44",X"B0",X"0F",X"A2",X"02",X"85",X"EF",X"6E",X"B5",
		X"42",X"95",X"14",X"CA",X"10",X"F9",X"85",X"EF",X"EA",X"D8",X"60",X"85",X"EF",X"6E",X"A6",X"4E",
		X"BD",X"80",X"D3",X"C5",X"E6",X"F0",X"08",X"85",X"E6",X"20",X"86",X"D3",X"85",X"EF",X"6E",X"60",
		X"42",X"43",X"44",X"45",X"85",X"EF",X"6E",X"48",X"A5",X"10",X"F0",X"08",X"68",X"48",X"C5",X"03",
		X"40",X"85",X"EF",X"EA",X"68",X"60",X"85",X"EF",X"EA",X"A2",X"0E",X"20",X"C4",X"D4",X"A2",X"10",
		X"A5",X"0E",X"C9",X"02",X"90",X"05",X"A2",X"12",X"85",X"EF",X"EA",X"20",X"C4",X"D4",X"A2",X"14",
		X"20",X"C4",X"D4",X"A2",X"01",X"85",X"EF",X"6E",X"A5",X"0E",X"E0",X"01",X"F0",X"07",X"4A",X"4A",
		X"4A",X"4A",X"85",X"EF",X"6E",X"29",X"0F",X"D0",X"07",X"E0",X"00",X"F0",X"14",X"85",X"EF",X"6E",
		X"18",X"69",X"51",X"9D",X"14",X"12",X"4D",X"01",X"9D",X"14",X"16",X"CA",X"10",X"DA",X"85",X"EF",
		X"EA",X"60",X"85",X"EF",X"6E",X"A2",X"00",X"20",X"C4",X"D4",X"A5",X"11",X"C9",X"02",X"90",X"08",
		X"A2",X"02",X"20",X"C4",X"D4",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A2",X"0A",X"20",X"C4",
		X"D4",X"A2",X"06",X"A5",X"12",X"F0",X"05",X"A2",X"08",X"85",X"EF",X"EA",X"20",X"C4",X"D4",X"60",
		X"85",X"EF",X"EA",X"A2",X"0C",X"20",X"C4",X"D4",X"A2",X"06",X"A5",X"12",X"F0",X"05",X"A2",X"08",
		X"85",X"EF",X"EA",X"20",X"C4",X"D4",X"60",X"85",X"EF",X"EA",X"A2",X"04",X"20",X"C4",X"D4",X"A5",
		X"41",X"48",X"29",X"F0",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"01",X"8D",X"95",X"10",X"68",X"29",
		X"0F",X"18",X"69",X"01",X"8D",X"96",X"10",X"A9",X"AD",X"85",X"01",X"A9",X"10",X"85",X"02",X"A0",
		X"00",X"A5",X"41",X"29",X"0F",X"D0",X"07",X"A5",X"41",X"29",X"10",X"85",X"EF",X"EA",X"AA",X"F0",
		X"11",X"A9",X"31",X"91",X"01",X"C8",X"F8",X"8A",X"38",X"E9",X"01",X"D8",X"4C",X"5E",X"D4",X"85",
		X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A6",X"3F",X"86",X"03",X"85",X"EF",X"EA",X"A6",X"03",X"F0",
		X"36",X"A9",X"80",X"85",X"EF",X"EA",X"18",X"69",X"02",X"CA",X"D0",X"FA",X"85",X"01",X"A9",X"10",
		X"85",X"02",X"A2",X"32",X"A0",X"00",X"8A",X"91",X"01",X"C8",X"E8",X"8A",X"91",X"01",X"A5",X"01",
		X"18",X"69",X"20",X"85",X"01",X"88",X"E8",X"8A",X"91",X"01",X"C8",X"E8",X"8A",X"91",X"01",X"C6",
		X"03",X"4C",X"7D",X"D4",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"1F",X"85",X"03",X"4C",
		X"7D",X"D4",X"85",X"EF",X"EA",X"BD",X"3C",X"D5",X"85",X"01",X"BD",X"3D",X"D5",X"85",X"02",X"A2",
		X"00",X"A0",X"00",X"B1",X"01",X"85",X"07",X"C8",X"85",X"EF",X"EA",X"B1",X"01",X"85",X"03",X"85",
		X"05",X"C8",X"B1",X"01",X"85",X"04",X"18",X"69",X"04",X"85",X"06",X"C8",X"85",X"EF",X"EA",X"B1",
		X"01",X"C8",X"C9",X"FE",X"F0",X"E5",X"C9",X"FF",X"F0",X"41",X"C9",X"FD",X"D0",X"0B",X"B1",X"01",
		X"C8",X"85",X"07",X"4C",X"EF",X"D4",X"85",X"EF",X"EA",X"C9",X"FC",X"D0",X"10",X"B1",X"01",X"C8",
		X"84",X"0A",X"20",X"74",X"A6",X"A4",X"0A",X"4C",X"EF",X"D4",X"85",X"EF",X"6E",X"81",X"03",X"C9",
		X"07",X"81",X"05",X"E6",X"03",X"70",X"05",X"E6",X"04",X"85",X"EF",X"EA",X"E6",X"05",X"70",X"05",
		X"E6",X"06",X"85",X"EF",X"6E",X"4C",X"EF",X"D4",X"85",X"EF",X"EA",X"60",X"68",X"D5",X"7A",X"D5",
		X"81",X"D5",X"8C",X"D5",X"98",X"D5",X"A4",X"D5",X"B2",X"D5",X"C0",X"D5",X"C8",X"D5",X"E0",X"D5",
		X"F8",X"D5",X"02",X"D6",X"0B",X"D6",X"20",X"D6",X"40",X"D6",X"B7",X"D6",X"9A",X"D7",X"2F",X"D6",
		X"8B",X"D6",X"A4",X"D6",X"AD",X"D6",X"B2",X"D6",X"00",X"23",X"10",X"02",X"1F",X"1A",X"FE",X"2C",
		X"10",X"12",X"13",X"27",X"1D",X"0D",X"19",X"1C",X"0F",X"FF",X"00",X"39",X"10",X"03",X"1F",X"1A",
		X"FF",X"00",X"8D",X"10",X"1A",X"0B",X"1E",X"1E",X"0F",X"1C",X"18",X"FF",X"01",X"2C",X"12",X"42",
		X"3E",X"33",X"4B",X"37",X"44",X"28",X"2A",X"FF",X"01",X"2C",X"12",X"42",X"3E",X"33",X"4B",X"37",
		X"44",X"28",X"2B",X"FF",X"01",X"6B",X"12",X"61",X"5B",X"67",X"5F",X"50",X"6D",X"6E",X"5B",X"6C",
		X"6E",X"FF",X"01",X"6B",X"12",X"61",X"5B",X"67",X"5F",X"50",X"69",X"70",X"5F",X"6C",X"76",X"FF",
		X"01",X"6E",X"11",X"42",X"47",X"45",X"3A",X"FF",X"01",X"A6",X"11",X"19",X"18",X"16",X"23",X"00",
		X"02",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"00",X"00",X"0C",X"1F",X"1E",X"1E",X"19",X"18",X"FF",
		X"01",X"A6",X"11",X"02",X"00",X"19",X"1C",X"00",X"03",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"1D",
		X"00",X"0C",X"1F",X"1E",X"1E",X"19",X"18",X"FF",X"01",X"0D",X"12",X"5D",X"6C",X"5F",X"5E",X"63",
		X"6E",X"FF",X"01",X"4A",X"12",X"0C",X"19",X"18",X"1F",X"1D",X"FF",X"01",X"A7",X"12",X"5C",X"5F",
		X"6D",X"6E",X"50",X"60",X"63",X"70",X"5F",X"50",X"6A",X"66",X"5B",X"73",X"5F",X"6C",X"6D",X"FF",
		X"01",X"EA",X"12",X"40",X"33",X"3F",X"37",X"28",X"28",X"45",X"35",X"41",X"44",X"37",X"FF",X"01",
		X"D4",X"13",X"78",X"79",X"7A",X"7B",X"7C",X"28",X"2A",X"32",X"31",X"2B",X"FF",X"85",X"EF",X"EA",
		X"00",X"23",X"11",X"40",X"41",X"00",X"FC",X"20",X"FD",X"01",X"54",X"51",X"51",X"4F",X"FC",X"20",
		X"57",X"51",X"51",X"7D",X"7E",X"FC",X"40",X"FD",X"00",X"FE",X"31",X"11",X"60",X"61",X"00",X"FC",
		X"20",X"FD",X"01",X"55",X"51",X"51",X"4F",X"FC",X"20",X"59",X"51",X"51",X"7D",X"7E",X"FC",X"40",
		X"FD",X"00",X"FE",X"6A",X"11",X"80",X"81",X"00",X"FC",X"20",X"FD",X"01",X"56",X"51",X"51",X"4F",
		X"FC",X"20",X"52",X"51",X"51",X"51",X"7D",X"7E",X"FC",X"40",X"FF",X"01",X"05",X"12",X"52",X"51",
		X"51",X"7D",X"7E",X"FE",X"0E",X"12",X"53",X"51",X"51",X"7D",X"7E",X"FE",X"16",X"12",X"55",X"51",
		X"51",X"7D",X"7E",X"FF",X"01",X"0E",X"12",X"55",X"FE",X"16",X"12",X"57",X"FF",X"01",X"16",X"12",
		X"59",X"FF",X"01",X"0E",X"12",X"57",X"FF",X"00",X"6F",X"11",X"E2",X"CC",X"CC",X"CC",X"E3",X"FE",
		X"8C",X"11",X"E2",X"CC",X"CC",X"D5",X"CC",X"E1",X"CC",X"E1",X"FE",X"AC",X"11",X"E1",X"CC",X"D6",
		X"D5",X"CC",X"CE",X"E1",X"E1",X"FE",X"C9",X"11",X"E2",X"CC",X"CC",X"D5",X"CC",X"D6",X"D5",X"CF",
		X"CC",X"CE",X"D6",X"D5",X"CC",X"E3",X"FE",X"E9",X"11",X"E1",X"CC",X"E1",X"E1",X"CC",X"CC",X"D5",
		X"E1",X"CF",X"CC",X"D6",X"D5",X"CC",X"E1",X"FE",X"06",X"12",X"E2",X"CC",X"D7",X"D5",X"CC",X"CC",
		X"D5",X"CC",X"D6",X"D5",X"CC",X"E1",X"CC",X"D6",X"D5",X"CC",X"D6",X"D9",X"DA",X"E3",X"FE",X"26",
		X"12",X"E1",X"CC",X"D8",X"D5",X"CC",X"E1",X"E1",X"CC",X"D6",X"D5",X"CC",X"CC",X"CC",X"D6",X"D5",
		X"CC",X"D6",X"DB",X"DC",X"E1",X"FE",X"43",X"12",X"E2",X"CC",X"CC",X"DD",X"CC",X"CF",X"CE",X"CC",
		X"CC",X"D5",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"D6",X"CC",X"CC",X"D6",X"DE",X"DF",X"E0",X"D9",
		X"D7",X"E3",X"FE",X"63",X"12",X"E1",X"E1",X"CC",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"E1",X"CD",X"CC",X"CE",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"D6",X"D9",X"D7",X"E1",X"FE",
		X"83",X"12",X"E1",X"E1",X"CC",X"E1",X"CD",X"CC",X"CC",X"CE",X"E1",X"CC",X"E1",X"E1",X"E1",X"CC",
		X"E1",X"CC",X"E1",X"CC",X"D1",X"E1",X"CC",X"E1",X"D6",X"DB",X"D8",X"E1",X"FE",X"A3",X"12",X"E1",
		X"E1",X"E1",X"E1",X"CC",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",
		X"CC",X"D2",X"E1",X"CC",X"E1",X"E1",X"E1",X"E1",X"E1",X"FF",X"00",X"C2",X"12",X"E2",X"CC",X"CC",
		X"CC",X"E1",X"CC",X"E1",X"E1",X"E1",X"E1",X"CC",X"E1",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",X"CC",
		X"CC",X"D1",X"CC",X"E1",X"CC",X"CC",X"CC",X"CE",X"E3",X"00",X"FE",X"E2",X"12",X"E1",X"E1",X"CC",
		X"E1",X"E1",X"CF",X"CC",X"CC",X"CE",X"E1",X"CC",X"E1",X"E1",X"E1",X"CC",X"CC",X"CC",X"E1",X"CC",
		X"D4",X"D2",X"CC",X"E1",X"CC",X"E1",X"CF",X"CC",X"E1",X"FE",X"02",X"13",X"E1",X"E1",X"CC",X"E1",
		X"E1",X"E1",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",X"CC",X"D3",
		X"CC",X"CC",X"E1",X"CC",X"E1",X"E1",X"CC",X"E1",X"FE",X"22",X"13",X"E1",X"E1",X"CC",X"E1",X"E1",
		X"CC",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",X"E1",X"E1",X"CC",X"E1",X"CC",X"E1",X"CC",X"E1",X"D4",
		X"CC",X"E1",X"CC",X"E1",X"CD",X"CC",X"E1",X"FE",X"42",X"13",X"E1",X"CC",X"CC",X"CC",X"E1",X"CF",
		X"CC",X"CC",X"D0",X"E1",X"CC",X"CC",X"CC",X"E1",X"CC",X"E1",X"CC",X"E1",X"CC",X"E1",X"D3",X"CC",
		X"E1",X"CC",X"CC",X"CC",X"D0",X"E1",X"FE",X"61",X"13",X"E2",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E3",X"00",X"E2",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E3",X"FF",X"85",X"EF",X"EA",X"20",X"A0",X"A4",X"A9",
		X"00",X"85",X"0A",X"A9",X"E1",X"8D",X"01",X"0C",X"A2",X"22",X"20",X"C4",X"D4",X"85",X"EF",X"EA",
		X"A2",X"01",X"20",X"78",X"A6",X"20",X"22",X"A7",X"20",X"F8",X"CE",X"A5",X"0A",X"D0",X"14",X"A2",
		X"1E",X"20",X"C4",X"D4",X"A2",X"20",X"20",X"C4",X"D4",X"A9",X"20",X"20",X"74",X"A6",X"E6",X"0A",
		X"85",X"EF",X"EA",X"20",X"C7",X"D8",X"A5",X"0A",X"C9",X"17",X"90",X"D4",X"20",X"A0",X"A4",X"A9",
		X"38",X"8D",X"01",X"0C",X"60",X"85",X"EF",X"EA",X"A5",X"0A",X"F0",X"45",X"A5",X"D6",X"D0",X"41",
		X"A0",X"03",X"85",X"EF",X"EA",X"B9",X"12",X"D9",X"99",X"01",X"00",X"88",X"10",X"F7",X"85",X"EF",
		X"EA",X"A0",X"1F",X"85",X"EF",X"EA",X"B1",X"03",X"91",X"01",X"88",X"10",X"F9",X"A5",X"01",X"38",
		X"E9",X"20",X"85",X"01",X"B0",X"05",X"C6",X"02",X"85",X"EF",X"EA",X"A5",X"03",X"38",X"E9",X"20",
		X"85",X"03",X"B0",X"DD",X"C6",X"04",X"C9",X"04",X"C9",X"10",X"D0",X"D5",X"E6",X"0A",X"C1",X"EF",
		X"EA",X"60",X"80",X"13",X"60",X"13",X"85",X"EF",X"EA",X"A2",X"1C",X"20",X"C4",X"D4",X"20",X"48",
		X"D9",X"20",X"B5",X"D9",X"A2",X"18",X"20",X"C4",X"D4",X"A2",X"1A",X"20",X"C4",X"D4",X"20",X"B2",
		X"DA",X"20",X"88",X"DA",X"20",X"EE",X"D9",X"20",X"38",X"DA",X"A9",X"A0",X"20",X"74",X"A6",X"20",
		X"C3",X"DA",X"20",X"A0",X"A4",X"60",X"85",X"EF",X"EA",X"A9",X"00",X"85",X"5B",X"C1",X"0A",X"C1",
		X"EF",X"EA",X"A4",X"5B",X"BE",X"A6",X"D9",X"20",X"C4",X"D4",X"A9",X"00",X"85",X"5C",X"C1",X"EF",
		X"EA",X"A4",X"5C",X"BE",X"AA",X"D9",X"A5",X"5B",X"20",X"95",X"A5",X"A6",X"0A",X"A9",X"01",X"8D",
		X"00",X"18",X"B9",X"AD",X"D9",X"18",X"7D",X"85",X"CE",X"8D",X"01",X"18",X"4D",X"70",X"8D",X"03",
		X"18",X"B9",X"B0",X"D9",X"8D",X"02",X"18",X"4D",X"40",X"20",X"74",X"A6",X"E6",X"5C",X"C9",X"5C",
		X"C9",X"03",X"90",X"CD",X"E6",X"0A",X"EA",X"0A",X"A9",X"00",X"8D",X"00",X"18",X"EA",X"5B",X"C9",
		X"5B",X"C9",X"04",X"90",X"AD",X"60",X"24",X"26",X"28",X"2A",X"00",X"00",X"01",X"41",X"32",X"32",
		X"C0",X"78",X"38",X"85",X"EF",X"6E",X"A2",X"16",X"20",X"C4",X"D4",X"A5",X"19",X"29",X"0F",X"18",
		X"69",X"01",X"8D",X"50",X"12",X"C9",X"18",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"01",X"8D",X"51",
		X"12",X"A2",X"02",X"A9",X"01",X"85",X"EF",X"6E",X"9D",X"52",X"12",X"CA",X"10",X"FA",X"A2",X"04",
		X"A9",X"02",X"85",X"EF",X"6E",X"9D",X"50",X"16",X"CA",X"10",X"FA",X"60",X"85",X"EF",X"6E",X"A9",
		X"0B",X"85",X"01",X"85",X"03",X"4D",X"13",X"85",X"02",X"A9",X"17",X"85",X"04",X"4A",X"00",X"85",
		X"EF",X"EA",X"A0",X"00",X"85",X"EF",X"EA",X"BD",X"00",X"07",X"91",X"01",X"A9",X"01",X"91",X"03",
		X"E8",X"E0",X"0F",X"90",X"04",X"60",X"85",X"EF",X"EA",X"C8",X"C0",X"03",X"90",X"E9",X"20",X"26",
		X"DA",X"4C",X"02",X"DA",X"85",X"EF",X"EA",X"A5",X"01",X"18",X"69",X"20",X"85",X"01",X"A5",X"03",
		X"18",X"69",X"20",X"85",X"03",X"60",X"85",X"EF",X"EA",X"A9",X"10",X"85",X"01",X"85",X"03",X"A9",
		X"13",X"85",X"02",X"A9",X"17",X"85",X"04",X"A2",X"00",X"85",X"EF",X"EA",X"A0",X"00",X"85",X"EF",
		X"EA",X"BD",X"10",X"07",X"48",X"29",X"F0",X"4A",X"4A",X"4A",X"4A",X"20",X"7B",X"DA",X"C8",X"68",
		X"29",X"0F",X"20",X"7B",X"DA",X"E8",X"E0",X"0F",X"90",X"04",X"60",X"85",X"EF",X"EA",X"C8",X"C0",
		X"06",X"90",X"DE",X"20",X"26",X"DA",X"4C",X"4C",X"DA",X"85",X"EF",X"EA",X"18",X"69",X"51",X"91",
		X"01",X"A9",X"01",X"91",X"03",X"60",X"85",X"EF",X"EA",X"A9",X"38",X"85",X"01",X"85",X"03",X"A9",
		X"19",X"85",X"02",X"A9",X"1D",X"85",X"04",X"A9",X"2A",X"85",X"05",X"A0",X"00",X"85",X"EF",X"EA",
		X"A5",X"05",X"91",X"01",X"A9",X"01",X"91",X"03",X"E6",X"05",X"C8",X"C0",X"05",X"90",X"F1",X"60",
		X"85",X"EF",X"EA",X"A2",X"1F",X"A9",X"36",X"85",X"EF",X"EA",X"9D",X"80",X"12",X"CA",X"10",X"FA",
		X"60",X"85",X"EF",X"EA",X"A2",X"09",X"85",X"EF",X"EA",X"BD",X"D4",X"13",X"5D",X"DA",X"DA",X"F0",
		X"05",X"EA",X"EA",X"85",X"EF",X"EA",X"CA",X"10",X"F0",X"60",X"78",X"79",X"7A",X"7B",X"7C",X"28",
		X"2A",X"32",X"31",X"2A",X"85",X"EF",X"EA",X"20",X"08",X"C9",X"20",X"45",X"CD",X"A9",X"68",X"85",
		X"DC",X"A9",X"E0",X"85",X"DB",X"A9",X"00",X"85",X"DF",X"8D",X"04",X"40",X"8D",X"20",X"07",X"85",
		X"E2",X"A9",X"03",X"8D",X"24",X"07",X"C5",X"28",X"07",X"A9",X"01",X"8D",X"2C",X"07",X"C5",X"30",
		X"07",X"60",X"85",X"EF",X"6E",X"A9",X"01",X"20",X"74",X"A6",X"20",X"22",X"A7",X"A5",X"D8",X"D0",
		X"30",X"A6",X"E2",X"A5",X"DC",X"18",X"7D",X"55",X"DB",X"85",X"DC",X"C9",X"A0",X"B0",X"07",X"C9",
		X"30",X"B0",X"0C",X"85",X"EF",X"6E",X"A5",X"E2",X"49",X"01",X"85",X"E2",X"C1",X"EF",X"6E",X"20",
		X"1B",X"C7",X"20",X"49",X"C7",X"20",X"7C",X"C7",X"20",X"5E",X"CD",X"20",X"43",X"CE",X"85",X"EF",
		X"EA",X"20",X"F8",X"CE",X"60",X"02",X"FE",X"85",X"EF",X"EA",X"A5",X"40",X"29",X"03",X"0A",X"0A",
		X"85",X"01",X"A5",X"4C",X"29",X"F3",X"05",X"01",X"85",X"4C",X"60",X"85",X"EF",X"6E",X"A5",X"10",
		X"F0",X"55",X"20",X"CA",X"DB",X"90",X"04",X"60",X"85",X"EF",X"EA",X"20",X"F1",X"DB",X"20",X"A0",
		X"A4",X"A9",X"00",X"8D",X"04",X"40",X"4A",X"18",X"20",X"C4",X"D4",X"A2",X"1A",X"20",X"C4",X"D4",
		X"20",X"B2",X"DA",X"20",X"38",X"DA",X"20",X"EE",X"D9",X"A9",X"00",X"85",X"5C",X"C1",X"5E",X"C1",
		X"5F",X"20",X"2B",X"DD",X"A9",X"30",X"85",X"5B",X"85",X"EF",X"EA",X"A9",X"01",X"20",X"74",X"A6",
		X"20",X"22",X"A7",X"20",X"F8",X"CE",X"20",X"6F",X"DC",X"20",X"C3",X"DC",X"20",X"FB",X"DC",X"90",
		X"EA",X"20",X"A0",X"A4",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"A2",X"00",X"85",X"EF",X"6E",
		X"BD",X"12",X"07",X"38",X"E5",X"42",X"BD",X"11",X"07",X"E5",X"43",X"BD",X"10",X"07",X"E5",X"44",
		X"90",X"0A",X"E8",X"E8",X"E8",X"E0",X"0F",X"90",X"E7",X"85",X"EF",X"EA",X"86",X"60",X"28",X"85",
		X"EF",X"EA",X"A9",X"01",X"85",X"0A",X"C1",X"EF",X"EA",X"A9",X"00",X"85",X"01",X"4D",X"07",X"85",
		X"02",X"A9",X"00",X"A2",X"02",X"85",X"EF",X"EA",X"95",X"03",X"CA",X"10",X"FB",X"A5",X"0A",X"F0",
		X"17",X"A9",X"10",X"85",X"01",X"A9",X"07",X"85",X"02",X"A5",X"44",X"85",X"03",X"A5",X"43",X"85",
		X"04",X"A5",X"42",X"85",X"05",X"85",X"EF",X"EA",X"A6",X"60",X"85",X"EF",X"EA",X"8A",X"A8",X"A9",
		X"02",X"85",X"06",X"85",X"EF",X"EA",X"B1",X"01",X"48",X"C8",X"C6",X"06",X"10",X"F8",X"8A",X"48",
		X"A8",X"A2",X"00",X"85",X"EF",X"EA",X"B5",X"03",X"91",X"01",X"C8",X"E8",X"E0",X"03",X"90",X"F6",
		X"68",X"AA",X"A0",X"02",X"85",X"EF",X"EA",X"68",X"99",X"03",X"00",X"88",X"10",X"F9",X"E8",X"E8",
		X"E8",X"E0",X"0F",X"90",X"C8",X"85",X"EF",X"EA",X"C6",X"0A",X"10",X"8D",X"60",X"85",X"EF",X"EA",
		X"A5",X"DA",X"D0",X"4A",X"A9",X"0F",X"85",X"DA",X"A6",X"12",X"AD",X"03",X"40",X"29",X"40",X"D0",
		X"05",X"A2",X"00",X"85",X"EF",X"EA",X"BD",X"00",X"40",X"49",X"FF",X"29",X"0F",X"F0",X"2F",X"A2",
		X"00",X"C9",X"08",X"B0",X"07",X"29",X"05",X"D0",X"07",X"85",X"EF",X"EA",X"E8",X"85",X"EF",X"EA",
		X"A5",X"5C",X"18",X"7D",X"BF",X"DC",X"10",X"05",X"A9",X"1A",X"85",X"EF",X"EA",X"C9",X"1B",X"90",
		X"05",X"A9",X"00",X"85",X"EF",X"EA",X"85",X"5C",X"20",X"2B",X"DD",X"85",X"EF",X"EA",X"60",X"01",
		X"FF",X"85",X"EF",X"EA",X"A6",X"12",X"AD",X"03",X"40",X"29",X"40",X"D0",X"05",X"A2",X"00",X"85",
		X"EF",X"EA",X"BD",X"00",X"40",X"49",X"FF",X"29",X"10",X"C5",X"5F",X"F0",X"1B",X"85",X"5F",X"AA",
		X"F0",X"16",X"AD",X"AF",X"11",X"48",X"A5",X"60",X"18",X"65",X"5E",X"AA",X"68",X"9D",X"00",X"07",
		X"E6",X"5E",X"20",X"EE",X"D9",X"85",X"EF",X"EA",X"60",X"85",X"EF",X"EA",X"A5",X"D6",X"D0",X"07",
		X"C6",X"5B",X"30",X"20",X"85",X"EF",X"6E",X"AD",X"02",X"40",X"49",X"FF",X"29",X"03",X"D0",X"14",
		X"85",X"EF",X"EA",X"A5",X"5E",X"C9",X"03",X"90",X"0F",X"85",X"EF",X"EA",X"A9",X"40",X"20",X"74",
		X"A6",X"85",X"EF",X"EA",X"38",X"85",X"EF",X"6E",X"60",X"85",X"EF",X"EA",X"20",X"38",X"DD",X"20",
		X"75",X"DD",X"20",X"AE",X"DD",X"60",X"85",X"EF",X"EA",X"A9",X"01",X"85",X"5D",X"C9",X"5C",X"85",
		X"0A",X"85",X"EF",X"EA",X"20",X"BE",X"DD",X"A5",X"0A",X"18",X"69",X"33",X"A0",X"00",X"91",X"01",
		X"A5",X"02",X"18",X"69",X"04",X"85",X"02",X"4D",X"01",X"91",X"01",X"E6",X"0A",X"C9",X"0A",X"C9",
		X"1B",X"90",X"07",X"A9",X"00",X"85",X"0A",X"C1",X"EF",X"EA",X"E6",X"5D",X"C9",X"5D",X"C9",X"1E",
		X"90",X"D2",X"60",X"85",X"EF",X"6E",X"A9",X"00",X"85",X"5D",X"85",X"EF",X"6E",X"20",X"BE",X"DD",
		X"A0",X"00",X"B1",X"01",X"48",X"C9",X"01",X"29",X"F0",X"09",X"0F",X"85",X"03",X"1C",X"E5",X"01",
		X"18",X"65",X"03",X"85",X"01",X"2C",X"91",X"01",X"A5",X"02",X"18",X"69",X"04",X"85",X"02",X"4D",
		X"01",X"91",X"01",X"E6",X"5D",X"C9",X"5D",X"C9",X"1F",X"90",X"D2",X"60",X"85",X"EF",X"6E",X"AD",
		X"AF",X"11",X"38",X"E9",X"33",X"18",X"69",X"0B",X"8D",X"AF",X"11",X"60",X"85",X"EF",X"6E",X"A5",
		X"5D",X"C9",X"15",X"B0",X"5E",X"C9",X"10",X"B0",X"34",X"C9",X"0B",X"B0",X"11",X"90",X"03",X"85",
		X"EF",X"EA",X"A5",X"5D",X"85",X"01",X"4D",X"11",X"85",X"02",X"60",X"85",X"EF",X"6E",X"A5",X"5D",
		X"38",X"E9",X"0A",X"AA",X"A9",X"0A",X"85",X"01",X"A9",X"11",X"85",X"02",X"C1",X"EF",X"6E",X"A9",
		X"21",X"18",X"65",X"01",X"85",X"01",X"66",X"D0",X"F6",X"60",X"85",X"EF",X"6E",X"A5",X"5D",X"38",
		X"E9",X"0F",X"AA",X"A9",X"AF",X"85",X"01",X"A9",X"11",X"85",X"02",X"85",X"EF",X"EA",X"A9",X"1F",
		X"18",X"65",X"01",X"85",X"01",X"90",X"05",X"E6",X"02",X"85",X"EF",X"EA",X"CA",X"D0",X"EF",X"60",
		X"85",X"EF",X"EA",X"A9",X"5E",X"85",X"01",X"A9",X"12",X"85",X"02",X"A5",X"01",X"38",X"E5",X"5D",
		X"85",X"01",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"80",X"80",X"81",X"81",X"80",X"80",X"00",X"00",X"08",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"FB",X"FD",X"FB",X"F7",X"F7",X"FF",X"0F",X"1F",X"FF",X"BF",X"BF",X"BF",X"3F",X"7F",X"FF",
		X"FF",X"FE",X"FC",X"FE",X"FD",X"FD",X"FF",X"F8",X"F0",X"FF",X"EF",X"EF",X"EF",X"9F",X"7E",X"00",
		X"FF",X"3F",X"BF",X"7F",X"BF",X"BF",X"FF",X"1F",X"0F",X"FF",X"F7",X"F7",X"F7",X"FB",X"7B",X"00",
		X"00",X"7F",X"9F",X"EF",X"EF",X"EF",X"FF",X"F0",X"F8",X"FF",X"FD",X"FD",X"FE",X"FC",X"FF",X"FF",
		X"00",X"FD",X"FD",X"FB",X"F7",X"EF",X"EF",X"F7",X"F7",X"CF",X"BF",X"BF",X"7F",X"7F",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FD",X"FD",X"FD",X"FB",X"E7",X"F7",X"CF",X"BF",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"3F",X"DF",X"DF",X"EF",X"EF",X"F7",X"FB",X"FD",X"00",
		X"00",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"80",X"BF",X"BF",X"DF",X"DF",X"EF",X"DF",X"EF",X"F7",X"F7",X"FB",X"FB",X"F9",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",
		X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F0",X"F0",X"F8",X"F8",X"FC",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FE",X"FC",X"F8",X"F8",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"80",X"00",X"01",X"01",X"00",X"80",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"01",X"03",X"07",X"07",X"0F",X"FF",X"FF",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"FF",
		X"FF",X"FE",X"FC",X"FE",X"FC",X"FC",X"F8",X"FF",X"FF",X"F0",X"E0",X"E0",X"E0",X"80",X"00",X"00",
		X"FF",X"3F",X"3F",X"7F",X"3F",X"3F",X"1F",X"FF",X"FF",X"0F",X"07",X"07",X"07",X"03",X"03",X"00",
		X"00",X"00",X"80",X"E0",X"E0",X"E0",X"F0",X"FF",X"FF",X"F8",X"FC",X"FC",X"FE",X"FC",X"FF",X"FF",
		X"00",X"01",X"01",X"03",X"07",X"0F",X"0F",X"07",X"07",X"0F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"E0",X"F0",X"C0",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"E0",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",
		X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F0",X"F0",X"F8",X"F8",X"FC",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FE",X"FC",X"F8",X"F8",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"F1",X"F9",X"FC",X"FC",X"FC",X"FC",X"FD",X"F9",X"FB",X"F3",X"F7",X"E7",X"8F",X"3F",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",
		X"FE",X"FE",X"FD",X"FD",X"FB",X"FB",X"F7",X"F7",X"EF",X"EF",X"DF",X"DF",X"BF",X"BF",X"7F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"8F",X"E7",X"F7",X"F3",X"FB",X"F9",X"FD",X"FC",X"FC",X"FC",X"FC",X"F9",X"F1",X"00",
		X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"7F",X"BF",X"BF",X"DF",X"DF",X"EF",X"EF",X"F7",X"F7",X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"C0",X"00",X"70",X"7C",X"7E",X"7E",X"7C",X"70",X"00",X"C0",X"F0",X"C0",X"00",
		X"E3",X"CF",X"03",X"6F",X"03",X"00",X"00",X"3B",X"3B",X"00",X"00",X"03",X"6F",X"03",X"CF",X"E3",
		X"FF",X"FC",X"FE",X"FC",X"F8",X"F8",X"F0",X"00",X"08",X"E8",X"C4",X"C4",X"C2",X"C2",X"81",X"01",
		X"80",X"81",X"43",X"41",X"23",X"23",X"17",X"10",X"00",X"0F",X"1F",X"1F",X"1F",X"7F",X"FF",X"FF",
		X"01",X"C1",X"C2",X"82",X"C4",X"C4",X"E8",X"08",X"00",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FF",
		X"FF",X"FF",X"7F",X"1F",X"1F",X"1F",X"0F",X"00",X"10",X"17",X"23",X"23",X"41",X"43",X"80",X"80",
		X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"07",X"1F",X"0F",X"3F",X"7F",X"7F",
		X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"01",X"01",X"01",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"40",X"40",X"20",X"10",X"10",X"08",X"04",X"02",X"04",X"04",X"02",X"02",X"02",X"01",
		X"80",X"80",X"40",X"20",X"18",X"04",X"08",X"08",X"04",X"04",X"02",X"04",X"02",X"02",X"01",X"01",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"01",X"02",X"04",X"04",X"02",X"04",X"08",X"08",X"10",X"20",X"40",X"40",X"80",X"80",
		X"01",X"01",X"02",X"02",X"04",X"04",X"06",X"08",X"10",X"20",X"10",X"20",X"20",X"40",X"80",X"80",
		X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"81",X"43",X"43",X"27",X"27",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"27",X"27",X"43",X"43",X"81",X"81",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"06",X"0C",X"0E",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"07",X"0D",X"0F",X"05",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"05",X"07",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"04",X"03",X"0F",X"05",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0E",X"04",X"03",X"02",X"06",X"0C",X"03",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"05",X"0F",X"05",X"02",X"03",X"07",X"0D",X"02",X"03",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"0F",X"05",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"0C",X"06",X"04",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"09",X"0D",X"07",X"05",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"02",X"0E",X"04",X"03",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"0F",X"05",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"06",X"04",X"0E",X"04",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"0F",X"05",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"03",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"03",X"02",X"06",X"0C",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"07",X"0D",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"06",X"04",X"03",X"02",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"04",X"03",X"02",X"03",X"07",X"05",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"09",X"05",X"02",X"03",X"02",X"03",X"02",X"03",X"0F",X"05",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"06",X"04",X"03",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"05",X"02",X"03",X"0F",X"05",X"02",X"03",X"0A",X"00",
		X"08",X"09",X"0D",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"06",X"00",
		X"02",X"03",X"02",X"06",X"0C",X"03",X"02",X"06",X"04",X"03",X"02",X"0E",X"04",X"03",X"07",X"0B",
		X"03",X"02",X"03",X"07",X"0D",X"02",X"03",X"07",X"05",X"02",X"03",X"0F",X"05",X"02",X"06",X"04",
		X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"07",X"05",
		X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"02",
		X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0A",X"00",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"09",X"0D",X"02",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"08",X"09",X"0D",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"08",X"02",X"06",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"06",X"0C",X"03",X"07",X"05",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"07",X"0D",X"02",X"0E",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"00",X"08",X"0A",X"08",X"09",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"08",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"06",X"04",X"03",X"02",X"03",X"0F",X"05",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"09",X"0D",X"07",X"05",X"02",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"06",X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"0B",X"09",X"0B",X"02",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"06",X"0C",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"08",X"09",X"0D",X"07",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"06",X"0C",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"08",X"02",X"03",X"07",X"0D",X"07",X"0B",X"0A",X"08",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"0E",X"04",X"0E",X"04",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"0F",X"05",X"0F",X"05",X"02",X"0E",X"0C",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"08",X"09",X"0D",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0B",X"0A",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"06",X"04",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"03",X"07",X"05",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"0C",X"06",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0D",X"07",X"0B",X"0A",X"00",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"0E",X"04",X"03",X"02",X"03",X"0A",X"08",X"0A",X"00",X"00",X"00",
		X"08",X"09",X"0D",X"02",X"03",X"0F",X"05",X"02",X"0E",X"04",X"03",X"02",X"03",X"0A",X"08",X"0A",
		X"02",X"03",X"02",X"03",X"02",X"06",X"04",X"03",X"0F",X"05",X"02",X"06",X"04",X"03",X"02",X"03",
		X"03",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"02",
		X"04",X"03",X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"03",X"0F",X"0B",X"09",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"04",X"0E",X"04",X"06",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"09",X"0B",X"09",X"05",X"07",X"05",X"0F",X"05",X"07",X"0D",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"04",X"06",X"0C",X"06",X"04",X"0E",X"04",X"06",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"05",X"07",X"0D",X"07",X"05",X"0F",X"05",X"07",X"0B",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"04",X"0E",X"04",X"06",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"05",X"0F",X"05",X"07",X"05",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"06",X"0C",X"06",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"0B",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"04",X"06",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"08",X"09",X"0B",X"09",X"05",X"0F",X"05",X"07",X"0D",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"04",X"06",X"04",X"06",X"04",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"05",X"07",X"05",X"07",X"05",X"07",X"0B",X"09",X"0B",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"04",X"0E",X"04",X"06",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"05",X"0F",X"05",X"07",X"05",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"0E",X"04",X"06",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"0F",X"05",X"07",X"0B",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"0C",X"06",X"04",X"03",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"08",X"09",X"0B",X"09",X"05",X"07",X"0D",X"07",X"05",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"04",X"06",X"04",X"0E",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"05",X"07",X"05",X"0F",X"05",X"0F",X"0B",X"09",X"0B",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"0C",X"06",X"04",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"0D",X"07",X"05",X"0F",X"05",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"06",X"04",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"0F",X"0B",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"04",X"06",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"08",X"09",X"0B",X"09",X"05",X"0F",X"05",X"07",X"0D",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"04",X"0E",X"04",X"0E",X"04",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"05",X"0F",X"05",X"0F",X"05",X"07",X"0B",X"09",X"0B",X"0A",X"00",
		X"00",X"00",X"00",X"04",X"0E",X"04",X"06",X"04",X"06",X"0C",X"06",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"09",X"05",X"0F",X"05",X"07",X"05",X"07",X"0D",X"07",X"05",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"03",X"02",X"06",X"04",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"02",X"03",X"07",X"0D",X"02",X"03",X"07",X"05",X"02",X"03",X"0F",X"0B",X"0A",X"00",
		X"08",X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"0A",
		X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0A",X"00",X"00",X"00",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"02",X"0E",X"00",X"08",X"09",X"0D",X"02",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"0A",X"00",X"0C",X"03",X"02",X"0E",X"00",X"08",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"02",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",X"0C",X"03",X"0F",X"0B",X"0A",X"00",
		X"00",X"0C",X"03",X"0F",X"0B",X"0A",X"08",X"02",X"0E",X"00",X"00",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"0E",X"0C",X"03",X"0F",X"0B",X"0A",X"08",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"0A",X"00",X"0C",X"0E",X"0C",X"0E",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"09",X"0D",X"02",X"0E",X"00",X"00",X"00",X"08",X"09",X"0D",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0A",X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"0E",X"00",X"00",X"00",X"08",X"02",X"0E",X"0C",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"0F",X"0B",X"0A",X"00",X"0C",X"03",X"0F",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"08",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"0A",X"08",X"02",X"03",X"02",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"0E",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"0C",X"0E",X"0C",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"0A",X"00",X"00",X"08",X"02",X"0E",X"00",X"08",X"09",X"0D",X"02",X"0E",X"00",
		X"00",X"08",X"02",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"0F",X"0B",X"0A",X"00",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"08",X"02",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0A",X"00",X"00",X"08",X"02",X"03",X"0A",X"00",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"0A",X"00",X"0C",X"03",X"02",X"0E",X"00",X"08",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"02",X"0E",X"00",X"08",X"02",X"03",X"0A",X"00",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"0E",X"00",X"08",X"02",X"0E",X"0C",X"03",X"09",X"0D",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"0F",X"0B",X"02",X"03",X"0F",X"0D",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"0E",X"0C",X"03",X"02",X"0E",X"0C",X"03",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"0A",X"00",X"0C",X"0E",X"00",X"08",X"02",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"09",X"0D",X"02",X"03",X"0A",X"00",X"00",X"08",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",X"0C",X"03",X"0F",X"0B",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",X"08",X"02",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"0E",X"00",X"00",X"0C",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"0E",X"00",X"08",X"09",X"0D",X"02",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"0F",X"0B",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"08",X"09",X"0D",X"02",X"06",X"04",X"03",X"02",X"03",X"0F",X"05",X"02",X"03",X"0F",X"0B",X"0A",
		X"02",X"06",X"04",X"03",X"07",X"05",X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",
		X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",
		X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"03",X"A0",X"00",X"A0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
