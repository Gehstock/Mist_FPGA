/*
  MIT License

  Copyright (c) 2019 Richard Eng

  Permission is hereby granted, free of charge, to any person obtaining a copy
  of this software and associated documentation files (the "Software"), to deal
  in the Software without restriction, including without limitation the rights
  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
  copies of the Software, and to permit persons to whom the Software is
  furnished to do so, subject to the following conditions:

  The above copyright notice and this permission notice shall be included in all
  copies or substantial portions of the Software.

  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
  SOFTWARE.
*/

/*
    inputs      outputs
    _s  _r      q   _q
    0   0       x   x
    0   1       1   0
    1   0       0   1
    1   1       q0  _q0
*/

module srlatch
(
    input wire mclk, _s, _r,
    output wire q,
    output wire _q
);

reg val;
initial val = 1'b0;

always @(posedge mclk) begin
    case({_s, _r})
        {1'b0, 1'b0}: val <= 1'bx;
        {1'b0, 1'b1}: val <= 1'b1;
        {1'b1, 1'b0}: val <= 1'b0;
        {1'b1, 1'b1}: val <= val;
    endcase
end

assign q = val;
assign _q = ~q;

endmodule
