library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"29",X"58",X"20",X"E1",X"74",X"20",X"2F",X"67",X"20",X"0C",X"7B",X"A9",X"14",X"85",X"91",X"46",
		X"9F",X"90",X"FC",X"A9",X"00",X"85",X"9F",X"20",X"3E",X"50",X"20",X"A6",X"50",X"A5",X"F2",X"29",
		X"40",X"D0",X"EC",X"4C",X"4B",X"7B",X"20",X"FB",X"55",X"20",X"5A",X"52",X"20",X"46",X"61",X"20",
		X"D0",X"53",X"20",X"21",X"53",X"20",X"58",X"54",X"20",X"32",X"51",X"4C",X"EE",X"59",X"A6",X"91",
		X"BD",X"4A",X"50",X"48",X"BD",X"49",X"50",X"48",X"60",X"D0",X"5A",X"0F",X"5B",X"25",X"50",X"6C",
		X"5D",X"E9",X"5B",X"1F",X"5C",X"81",X"5C",X"A9",X"5C",X"0B",X"5D",X"A1",X"5D",X"81",X"5A",X"B8",
		X"5A",X"3E",X"75",X"44",X"76",X"FF",X"76",X"85",X"77",X"9E",X"77",X"6C",X"50",X"A5",X"CA",X"29",
		X"03",X"D0",X"30",X"A4",X"AF",X"F0",X"02",X"C6",X"AF",X"D0",X"28",X"A5",X"92",X"85",X"91",X"C9",
		X"04",X"D0",X"20",X"A5",X"93",X"F0",X"1C",X"A9",X"00",X"20",X"49",X"6A",X"A9",X"06",X"20",X"49",
		X"6A",X"A9",X"1E",X"20",X"49",X"6A",X"A9",X"15",X"20",X"49",X"6A",X"A9",X"00",X"85",X"FA",X"85",
		X"95",X"85",X"94",X"4C",X"32",X"51",X"A5",X"93",X"D0",X"55",X"20",X"5D",X"5F",X"A5",X"66",X"F0",
		X"32",X"A0",X"00",X"C9",X"02",X"A5",X"F1",X"49",X"FF",X"29",X"18",X"F0",X"23",X"B0",X"05",X"29",
		X"10",X"B8",X"50",X"05",X"C8",X"C6",X"66",X"29",X"08",X"F0",X"03",X"C6",X"66",X"C8",X"98",X"85",
		X"AE",X"F0",X"0D",X"A0",X"FF",X"84",X"93",X"C8",X"84",X"68",X"A9",X"00",X"85",X"91",X"C6",X"AE",
		X"B8",X"50",X"12",X"A5",X"67",X"F0",X"0E",X"A5",X"91",X"C9",X"20",X"F0",X"08",X"C9",X"12",X"F0",
		X"04",X"A9",X"1E",X"85",X"91",X"A5",X"F3",X"29",X"03",X"D0",X"04",X"A9",X"02",X"85",X"66",X"E6",
		X"CA",X"A5",X"9F",X"D0",X"1C",X"A5",X"D4",X"F0",X"05",X"A4",X"B9",X"20",X"FC",X"5F",X"A5",X"D8",
		X"D0",X"0F",X"20",X"52",X"5A",X"A5",X"D7",X"49",X"01",X"85",X"D7",X"AA",X"BD",X"30",X"51",X"85",
		X"D8",X"A5",X"5F",X"F0",X"04",X"A9",X"F0",X"85",X"E0",X"A5",X"E0",X"F0",X"02",X"C6",X"E0",X"60",
		X"0A",X"32",X"A5",X"A6",X"F0",X"1E",X"A5",X"93",X"D0",X"06",X"20",X"55",X"51",X"B8",X"50",X"0E",
		X"A0",X"00",X"A5",X"95",X"84",X"95",X"85",X"B1",X"A5",X"94",X"84",X"94",X"85",X"B0",X"20",X"39",
		X"52",X"20",X"D3",X"64",X"60",X"A9",X"00",X"85",X"B1",X"85",X"B0",X"A6",X"D0",X"BD",X"65",X"01",
		X"D0",X"03",X"20",X"E7",X"51",X"A6",X"D0",X"BD",X"65",X"01",X"C5",X"A6",X"B0",X"05",X"A9",X"FE",
		X"B8",X"50",X"12",X"38",X"E5",X"A6",X"C9",X"0E",X"D0",X"05",X"A9",X"00",X"B8",X"50",X"06",X"A9",
		X"02",X"B0",X"02",X"A9",X"FE",X"85",X"B1",X"BD",X"18",X"06",X"85",X"98",X"BD",X"08",X"06",X"46",
		X"98",X"6A",X"46",X"98",X"6A",X"46",X"98",X"6A",X"46",X"98",X"6A",X"18",X"7D",X"30",X"01",X"C5",
		X"A5",X"B0",X"05",X"A9",X"FE",X"B8",X"50",X"09",X"D0",X"05",X"A9",X"00",X"B8",X"50",X"02",X"A9",
		X"02",X"85",X"B0",X"05",X"B1",X"D0",X"2F",X"A5",X"BC",X"C9",X"02",X"B0",X"29",X"A2",X"02",X"A5",
		X"A5",X"C9",X"60",X"B0",X"05",X"A2",X"00",X"B8",X"50",X"06",X"C9",X"A0",X"B0",X"02",X"A2",X"01",
		X"A5",X"BC",X"18",X"65",X"8E",X"C5",X"8C",X"B0",X"0D",X"20",X"BD",X"52",X"A0",X"00",X"84",X"B0",
		X"88",X"84",X"B1",X"20",X"E7",X"51",X"60",X"A6",X"D0",X"CA",X"10",X"02",X"A2",X"07",X"E4",X"D0",
		X"D0",X"01",X"60",X"BD",X"65",X"01",X"F0",X"F1",X"86",X"D0",X"60",X"A0",X"00",X"B5",X"B0",X"10",
		X"01",X"88",X"94",X"9D",X"A0",X"06",X"A5",X"FC",X"0A",X"A5",X"F4",X"29",X"08",X"6A",X"25",X"93",
		X"F0",X"01",X"C8",X"16",X"B0",X"36",X"9D",X"88",X"10",X"F9",X"B5",X"A3",X"18",X"75",X"B0",X"95",
		X"A3",X"B5",X"A5",X"75",X"9D",X"D5",X"A5",X"F0",X"0F",X"B4",X"9D",X"10",X"07",X"90",X"02",X"A9",
		X"00",X"B8",X"50",X"04",X"B0",X"02",X"A9",X"FF",X"60",X"A2",X"00",X"20",X"40",X"52",X"A2",X"01",
		X"20",X"FB",X"51",X"DD",X"56",X"52",X"B0",X"03",X"BD",X"56",X"52",X"DD",X"58",X"52",X"90",X"03",
		X"BD",X"58",X"52",X"95",X"A5",X"60",X"08",X"2D",X"F7",X"CE",X"A5",X"93",X"F0",X"57",X"A5",X"8D",
		X"05",X"8C",X"05",X"DB",X"05",X"DA",X"0D",X"6D",X"01",X"F0",X"47",X"A5",X"8F",X"18",X"65",X"BC",
		X"C9",X"10",X"B0",X"10",X"65",X"8C",X"18",X"65",X"DA",X"18",X"AE",X"6D",X"01",X"F0",X"01",X"38",
		X"65",X"90",X"C9",X"14",X"B0",X"1E",X"A2",X"02",X"A5",X"FA",X"3D",X"BA",X"52",X"F0",X"0F",X"B5",
		X"A0",X"F0",X"06",X"20",X"BD",X"52",X"B8",X"50",X"05",X"A9",X"80",X"20",X"EC",X"79",X"CA",X"10",
		X"E7",X"B8",X"50",X"0B",X"A5",X"FA",X"29",X"07",X"F0",X"05",X"A9",X"80",X"20",X"EC",X"79",X"B8",
		X"50",X"03",X"20",X"72",X"65",X"A9",X"00",X"85",X"FA",X"60",X"04",X"02",X"01",X"A0",X"07",X"B9",
		X"5D",X"01",X"D0",X"59",X"84",X"97",X"A9",X"00",X"99",X"4D",X"01",X"99",X"18",X"01",X"BD",X"E8",
		X"60",X"99",X"82",X"01",X"99",X"28",X"01",X"BD",X"F4",X"60",X"99",X"92",X"01",X"99",X"5D",X"01",
		X"A5",X"A5",X"99",X"A2",X"01",X"A5",X"A6",X"99",X"B2",X"01",X"20",X"7C",X"65",X"20",X"F6",X"58",
		X"A5",X"93",X"F0",X"14",X"B5",X"A0",X"C9",X"04",X"D0",X"09",X"8A",X"20",X"24",X"68",X"A9",X"01",
		X"B8",X"50",X"02",X"A9",X"04",X"20",X"EC",X"79",X"D6",X"A0",X"D0",X"08",X"A5",X"93",X"F0",X"04",
		X"8A",X"20",X"36",X"68",X"8A",X"A8",X"20",X"D1",X"67",X"98",X"AA",X"A0",X"00",X"88",X"10",X"9F",
		X"60",X"A5",X"B3",X"F0",X"05",X"C6",X"B3",X"B8",X"50",X"4E",X"A5",X"B2",X"18",X"65",X"B7",X"85",
		X"B2",X"A5",X"B3",X"65",X"B8",X"85",X"B3",X"A2",X"07",X"86",X"DC",X"A9",X"FF",X"85",X"BD",X"85",
		X"C2",X"A9",X"00",X"85",X"8C",X"85",X"DA",X"85",X"BE",X"A6",X"DC",X"BD",X"65",X"01",X"F0",X"1A",
		X"8A",X"18",X"69",X"08",X"85",X"97",X"BD",X"65",X"01",X"C5",X"BD",X"B0",X"02",X"85",X"BD",X"C5",
		X"BE",X"90",X"02",X"85",X"BE",X"25",X"93",X"20",X"79",X"53",X"C6",X"DC",X"10",X"DB",X"A4",X"8E",
		X"C0",X"0C",X"90",X"04",X"A9",X"FF",X"85",X"C2",X"60",X"A8",X"A5",X"D9",X"3D",X"F7",X"60",X"D0",
		X"13",X"C0",X"80",X"90",X"06",X"C0",X"A0",X"B0",X"02",X"86",X"C2",X"20",X"F7",X"66",X"20",X"11",
		X"54",X"B8",X"50",X"06",X"20",X"AC",X"77",X"20",X"0D",X"63",X"A6",X"DC",X"90",X"1D",X"A5",X"D9",
		X"3D",X"F7",X"60",X"F0",X"06",X"20",X"E9",X"7A",X"B8",X"50",X"07",X"A6",X"97",X"20",X"86",X"66",
		X"A6",X"DC",X"20",X"6B",X"58",X"20",X"9F",X"55",X"B8",X"50",X"14",X"A5",X"D9",X"3D",X"F7",X"60",
		X"D0",X"08",X"20",X"F0",X"66",X"E6",X"8C",X"B8",X"50",X"05",X"20",X"A8",X"77",X"E6",X"DA",X"60",
		X"A9",X"00",X"85",X"BC",X"A2",X"07",X"BD",X"5D",X"01",X"F0",X"32",X"86",X"97",X"A0",X"02",X"BD",
		X"82",X"01",X"C9",X"7B",X"D0",X"02",X"A0",X"06",X"84",X"D5",X"20",X"F7",X"66",X"20",X"11",X"54",
		X"90",X"0D",X"20",X"92",X"65",X"20",X"86",X"66",X"20",X"6B",X"58",X"A9",X"00",X"85",X"D5",X"C6",
		X"D5",X"10",X"E7",X"BD",X"5D",X"01",X"F0",X"05",X"20",X"F0",X"66",X"E6",X"BC",X"CA",X"10",X"C6",
		X"60",X"A4",X"97",X"B9",X"18",X"01",X"18",X"79",X"00",X"06",X"99",X"18",X"01",X"B9",X"28",X"01",
		X"79",X"10",X"06",X"99",X"28",X"01",X"B9",X"4D",X"01",X"18",X"79",X"20",X"06",X"99",X"4D",X"01",
		X"B9",X"5D",X"01",X"79",X"30",X"06",X"99",X"5D",X"01",X"D9",X"B2",X"01",X"F0",X"08",X"6A",X"59",
		X"30",X"06",X"10",X"02",X"38",X"60",X"B9",X"28",X"01",X"D9",X"A2",X"01",X"F0",X"08",X"6A",X"59",
		X"10",X"06",X"10",X"02",X"38",X"60",X"18",X"60",X"A4",X"B4",X"88",X"10",X"02",X"A0",X"04",X"84",
		X"B4",X"A5",X"8E",X"F0",X"4B",X"BE",X"B2",X"54",X"BD",X"6E",X"01",X"F0",X"3A",X"85",X"9C",X"FE",
		X"C2",X"01",X"BD",X"C2",X"01",X"29",X"7F",X"A8",X"C9",X"1B",X"90",X"16",X"BD",X"C2",X"01",X"30",
		X"05",X"C6",X"8F",X"B8",X"50",X"02",X"C6",X"90",X"C6",X"8E",X"A9",X"00",X"9D",X"6E",X"01",X"B8",
		X"50",X"15",X"BD",X"39",X"01",X"85",X"9B",X"B9",X"B7",X"54",X"85",X"B5",X"B9",X"B8",X"54",X"85",
		X"9A",X"20",X"71",X"5E",X"20",X"D4",X"54",X"CA",X"A4",X"B4",X"8A",X"D9",X"B1",X"54",X"D0",X"B8",
		X"60",X"FF",X"03",X"07",X"0B",X"0F",X"13",X"00",X"00",X"02",X"03",X"04",X"05",X"06",X"07",X"08",
		X"09",X"0A",X"0B",X"0C",X"0D",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"04",X"03",
		X"02",X"01",X"00",X"00",X"8A",X"48",X"A5",X"9A",X"85",X"D5",X"A0",X"08",X"A5",X"9C",X"C9",X"21",
		X"90",X"5E",X"B9",X"65",X"01",X"F0",X"56",X"85",X"9E",X"B9",X"30",X"01",X"85",X"9D",X"C0",X"08",
		X"D0",X"05",X"A9",X"06",X"B8",X"50",X"0E",X"A5",X"D9",X"39",X"F7",X"60",X"D0",X"05",X"A9",X"01",
		X"B8",X"50",X"02",X"A9",X"03",X"18",X"65",X"D5",X"85",X"9A",X"20",X"AB",X"58",X"B0",X"2E",X"98",
		X"48",X"18",X"69",X"08",X"85",X"97",X"C4",X"C2",X"D0",X"04",X"A9",X"FF",X"85",X"C2",X"C0",X"08",
		X"90",X"06",X"20",X"43",X"55",X"B8",X"50",X"10",X"A5",X"D9",X"39",X"F7",X"60",X"D0",X"06",X"20",
		X"50",X"55",X"B8",X"50",X"03",X"20",X"66",X"55",X"20",X"6B",X"58",X"68",X"A8",X"88",X"10",X"A2",
		X"68",X"AA",X"60",X"20",X"F8",X"7A",X"A9",X"00",X"85",X"C9",X"85",X"E3",X"A2",X"03",X"D0",X"20",
		X"C6",X"8C",X"20",X"7B",X"55",X"A6",X"97",X"20",X"86",X"66",X"A2",X"00",X"A4",X"97",X"B9",X"5D",
		X"01",X"C9",X"21",X"B0",X"0B",X"60",X"C6",X"DA",X"20",X"7B",X"55",X"20",X"E9",X"7A",X"A2",X"04",
		X"20",X"9F",X"5F",X"A4",X"B9",X"20",X"13",X"60",X"4C",X"EA",X"79",X"A4",X"97",X"B9",X"A2",X"01",
		X"48",X"A9",X"00",X"99",X"A2",X"01",X"68",X"A0",X"07",X"D9",X"AA",X"01",X"D0",X"01",X"60",X"88",
		X"10",X"F7",X"A0",X"09",X"88",X"D9",X"E2",X"60",X"D0",X"FA",X"A9",X"00",X"4C",X"47",X"58",X"A4",
		X"97",X"B9",X"A2",X"01",X"A0",X"09",X"88",X"D9",X"E2",X"60",X"D0",X"FA",X"A9",X"00",X"20",X"47",
		X"58",X"C0",X"06",X"90",X"21",X"A9",X"00",X"99",X"9A",X"00",X"B9",X"F1",X"60",X"49",X"E0",X"25",
		X"CD",X"C5",X"CD",X"F0",X"0E",X"85",X"CD",X"A9",X"02",X"20",X"EC",X"79",X"98",X"38",X"E9",X"06",
		X"20",X"36",X"68",X"B8",X"50",X"24",X"B9",X"F7",X"60",X"49",X"FC",X"A4",X"B9",X"39",X"C5",X"00",
		X"D9",X"C5",X"00",X"F0",X"15",X"99",X"C5",X"00",X"B9",X"C0",X"00",X"F0",X"06",X"38",X"E9",X"01",
		X"99",X"C0",X"00",X"E6",X"CF",X"A9",X"02",X"20",X"EC",X"79",X"60",X"A5",X"8D",X"05",X"DB",X"F0",
		X"76",X"A5",X"A7",X"0A",X"49",X"FF",X"38",X"69",X"CA",X"C9",X"B4",X"B0",X"02",X"A9",X"B4",X"C5",
		X"BE",X"90",X"64",X"A9",X"07",X"38",X"AE",X"6D",X"01",X"F0",X"01",X"18",X"E5",X"90",X"38",X"E5",
		X"8C",X"38",X"E5",X"DA",X"30",X"0B",X"85",X"DE",X"18",X"69",X"0C",X"38",X"E5",X"8F",X"38",X"E5",
		X"BC",X"30",X"44",X"C5",X"DE",X"B0",X"02",X"85",X"DE",X"20",X"FF",X"60",X"A5",X"DE",X"30",X"37",
		X"A5",X"DB",X"D0",X"06",X"20",X"78",X"56",X"B8",X"50",X"2D",X"A5",X"DA",X"C9",X"03",X"B0",X"24",
		X"18",X"65",X"8C",X"C9",X"05",X"B0",X"1A",X"A5",X"8D",X"D0",X"06",X"20",X"17",X"57",X"B8",X"50",
		X"10",X"AD",X"0A",X"40",X"29",X"03",X"D0",X"06",X"20",X"17",X"57",X"B8",X"50",X"03",X"20",X"78",
		X"56",X"B8",X"50",X"03",X"20",X"78",X"56",X"60",X"A2",X"FF",X"A5",X"8D",X"F0",X"2A",X"38",X"AD",
		X"6D",X"01",X"F0",X"01",X"18",X"A9",X"07",X"E5",X"DA",X"38",X"E5",X"DA",X"38",X"E5",X"8C",X"30",
		X"17",X"AA",X"E8",X"E0",X"04",X"90",X"02",X"A2",X"04",X"E4",X"8D",X"90",X"02",X"A6",X"8D",X"E6",
		X"DE",X"E4",X"DE",X"90",X"02",X"A6",X"DE",X"CA",X"86",X"DE",X"A6",X"DE",X"30",X"33",X"A5",X"A7",
		X"C9",X"02",X"90",X"1D",X"AD",X"6D",X"01",X"F0",X"18",X"A5",X"C9",X"C5",X"E1",X"90",X"12",X"AD",
		X"38",X"01",X"C9",X"30",X"90",X"0B",X"C9",X"D0",X"B0",X"07",X"A9",X"00",X"85",X"C9",X"4C",X"39",
		X"57",X"A5",X"A7",X"C9",X"01",X"90",X"07",X"A4",X"C2",X"30",X"03",X"4C",X"3B",X"57",X"4C",X"31",
		X"57",X"60",X"86",X"AC",X"20",X"82",X"57",X"A6",X"97",X"30",X"29",X"A9",X"DE",X"9D",X"65",X"01",
		X"9D",X"9A",X"01",X"AD",X"0A",X"40",X"A2",X"07",X"DD",X"8A",X"01",X"D0",X"05",X"AD",X"0A",X"40",
		X"A2",X"08",X"CA",X"10",X"F3",X"A6",X"97",X"9D",X"8A",X"01",X"9D",X"30",X"01",X"20",X"91",X"57",
		X"A9",X"FF",X"85",X"BE",X"A6",X"AC",X"60",X"20",X"E2",X"56",X"A6",X"97",X"30",X"12",X"20",X"D1",
		X"7A",X"E6",X"DA",X"C6",X"DB",X"E6",X"8D",X"C6",X"8C",X"A5",X"D9",X"1D",X"EF",X"60",X"85",X"D9",
		X"60",X"20",X"E2",X"56",X"C6",X"DE",X"10",X"F9",X"60",X"A0",X"08",X"A5",X"DE",X"C9",X"02",X"90",
		X"02",X"A9",X"02",X"85",X"DE",X"84",X"AC",X"20",X"82",X"57",X"A6",X"97",X"30",X"31",X"A4",X"AC",
		X"A9",X"00",X"C0",X"09",X"D0",X"0B",X"A5",X"C8",X"10",X"05",X"A9",X"FC",X"B8",X"50",X"02",X"A9",
		X"04",X"24",X"FC",X"50",X"02",X"49",X"FF",X"18",X"79",X"30",X"01",X"9D",X"30",X"01",X"9D",X"8A",
		X"01",X"B9",X"65",X"01",X"9D",X"65",X"01",X"9D",X"9A",X"01",X"20",X"91",X"57",X"C6",X"DE",X"10",
		X"C6",X"60",X"A2",X"07",X"BD",X"65",X"01",X"D0",X"04",X"86",X"97",X"A2",X"00",X"CA",X"10",X"F4",
		X"60",X"A6",X"B9",X"B5",X"C5",X"45",X"CB",X"35",X"C5",X"85",X"98",X"A5",X"CD",X"45",X"CC",X"25",
		X"CD",X"85",X"99",X"A4",X"CF",X"A5",X"CB",X"35",X"C5",X"10",X"01",X"C8",X"0A",X"D0",X"FA",X"C0",
		X"03",X"B0",X"1E",X"A0",X"00",X"A5",X"98",X"F0",X"06",X"20",X"1D",X"58",X"B8",X"50",X"0F",X"A0",
		X"06",X"A5",X"99",X"F0",X"06",X"20",X"1D",X"58",X"B8",X"50",X"03",X"20",X"0C",X"58",X"B8",X"50",
		X"0F",X"A0",X"06",X"A5",X"99",X"F0",X"06",X"20",X"1D",X"58",X"B8",X"50",X"03",X"20",X"17",X"58",
		X"A9",X"FF",X"20",X"47",X"58",X"A6",X"97",X"B9",X"E2",X"60",X"9D",X"AA",X"01",X"B9",X"EB",X"60",
		X"9D",X"BA",X"01",X"A9",X"00",X"9D",X"20",X"01",X"9D",X"55",X"01",X"BD",X"F7",X"60",X"49",X"FF",
		X"25",X"D9",X"85",X"D9",X"20",X"FA",X"58",X"C6",X"8D",X"E6",X"8C",X"60",X"AD",X"0A",X"40",X"4A",
		X"29",X"07",X"A8",X"90",X"01",X"C8",X"60",X"A0",X"00",X"A5",X"98",X"49",X"FF",X"48",X"A2",X"00",
		X"29",X"FF",X"10",X"01",X"E8",X"0A",X"D0",X"F8",X"86",X"98",X"AD",X"0A",X"40",X"3D",X"3E",X"58",
		X"C5",X"98",X"B0",X"F6",X"AA",X"68",X"88",X"0A",X"C8",X"90",X"FC",X"CA",X"10",X"F9",X"60",X"00",
		X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"85",X"98",X"84",X"99",X"A2",X"00",X"98",X"C9",X"06",
		X"90",X"06",X"38",X"E9",X"06",X"A8",X"A2",X"01",X"B9",X"F7",X"60",X"49",X"FF",X"35",X"CB",X"24",
		X"98",X"10",X"03",X"19",X"F7",X"60",X"95",X"CB",X"A4",X"99",X"60",X"86",X"AB",X"A6",X"97",X"BD",
		X"5D",X"01",X"C9",X"D2",X"B0",X"2A",X"A4",X"96",X"C6",X"96",X"10",X"04",X"A9",X"13",X"85",X"96",
		X"E6",X"8E",X"BD",X"28",X"01",X"99",X"39",X"01",X"BD",X"5D",X"01",X"99",X"6E",X"01",X"E0",X"08",
		X"90",X"07",X"E6",X"90",X"A9",X"80",X"B8",X"50",X"04",X"E6",X"8F",X"A9",X"00",X"99",X"C2",X"01",
		X"A9",X"00",X"9D",X"5D",X"01",X"9D",X"28",X"01",X"A6",X"AB",X"60",X"A5",X"9E",X"C5",X"9C",X"90",
		X"05",X"E5",X"9C",X"B8",X"50",X"05",X"A5",X"9C",X"38",X"E5",X"9E",X"C5",X"9A",X"B0",X"36",X"85",
		X"B1",X"A5",X"9D",X"C5",X"9B",X"90",X"05",X"E5",X"9B",X"B8",X"50",X"05",X"A5",X"9B",X"38",X"E5",
		X"9D",X"C5",X"9A",X"B0",X"20",X"C5",X"B1",X"B0",X"09",X"85",X"98",X"A5",X"B1",X"85",X"99",X"B8",
		X"50",X"06",X"85",X"99",X"A5",X"B1",X"85",X"98",X"A5",X"98",X"4A",X"18",X"65",X"98",X"4A",X"4A",
		X"18",X"65",X"99",X"C5",X"9A",X"60",X"84",X"97",X"10",X"06",X"8A",X"18",X"69",X"08",X"85",X"97",
		X"8A",X"48",X"98",X"48",X"A6",X"97",X"BD",X"B2",X"01",X"DD",X"5D",X"01",X"90",X"06",X"FD",X"5D",
		X"01",X"B8",X"50",X"07",X"BD",X"5D",X"01",X"38",X"FD",X"B2",X"01",X"85",X"B1",X"BD",X"A2",X"01",
		X"DD",X"28",X"01",X"90",X"06",X"FD",X"28",X"01",X"B8",X"50",X"07",X"BD",X"28",X"01",X"38",X"FD",
		X"A2",X"01",X"85",X"B0",X"A5",X"B0",X"C5",X"B1",X"B0",X"09",X"85",X"98",X"A5",X"B1",X"85",X"99",
		X"B8",X"50",X"06",X"85",X"99",X"A5",X"B1",X"85",X"98",X"A5",X"98",X"4A",X"18",X"65",X"98",X"4A",
		X"4A",X"18",X"65",X"99",X"90",X"02",X"A9",X"FF",X"85",X"98",X"A4",X"98",X"A5",X"B1",X"20",X"BB",
		X"59",X"A5",X"A9",X"9D",X"30",X"06",X"A5",X"AA",X"9D",X"20",X"06",X"A4",X"98",X"A5",X"B0",X"20",
		X"BB",X"59",X"A5",X"A9",X"9D",X"10",X"06",X"A5",X"AA",X"9D",X"00",X"06",X"BD",X"B2",X"01",X"DD",
		X"5D",X"01",X"B0",X"15",X"BD",X"20",X"06",X"49",X"FF",X"18",X"69",X"01",X"9D",X"20",X"06",X"BD",
		X"30",X"06",X"49",X"FF",X"69",X"00",X"9D",X"30",X"06",X"BD",X"A2",X"01",X"DD",X"28",X"01",X"B0",
		X"15",X"BD",X"00",X"06",X"49",X"FF",X"18",X"69",X"01",X"9D",X"00",X"06",X"BD",X"10",X"06",X"49",
		X"FF",X"69",X"00",X"9D",X"10",X"06",X"68",X"A8",X"68",X"AA",X"60",X"84",X"AD",X"86",X"AB",X"20",
		X"D0",X"59",X"86",X"A9",X"A2",X"00",X"86",X"A8",X"20",X"D4",X"59",X"86",X"AA",X"A6",X"AB",X"60",
		X"85",X"A8",X"A9",X"00",X"A0",X"07",X"26",X"A8",X"2A",X"90",X"05",X"E5",X"AD",X"38",X"B0",X"06",
		X"C5",X"AD",X"90",X"02",X"E5",X"AD",X"88",X"10",X"ED",X"26",X"A8",X"A6",X"A8",X"60",X"A4",X"B9",
		X"A5",X"A0",X"05",X"A1",X"05",X"A2",X"85",X"99",X"D0",X"24",X"B9",X"C5",X"00",X"F0",X"08",X"A5",
		X"CF",X"C9",X"03",X"90",X"02",X"A9",X"00",X"D0",X"15",X"A9",X"00",X"85",X"C9",X"85",X"8D",X"85",
		X"DB",X"AD",X"6D",X"01",X"05",X"BC",X"05",X"8E",X"D0",X"04",X"A9",X"08",X"85",X"91",X"A5",X"BC",
		X"05",X"8E",X"05",X"99",X"D0",X"04",X"A9",X"FF",X"85",X"BF",X"A5",X"BF",X"F0",X"0D",X"A9",X"00",
		X"85",X"C7",X"85",X"B3",X"85",X"B8",X"85",X"B7",X"20",X"72",X"65",X"A5",X"8D",X"05",X"BC",X"05",
		X"DB",X"05",X"8C",X"05",X"DA",X"0D",X"6D",X"01",X"05",X"8E",X"D0",X"04",X"A9",X"08",X"85",X"91",
		X"60",X"4D",X"A5",X"93",X"F0",X"03",X"4C",X"F0",X"65",X"A5",X"91",X"C9",X"04",X"D0",X"22",X"A0",
		X"00",X"A5",X"D7",X"D0",X"02",X"A0",X"40",X"84",X"B6",X"A2",X"05",X"86",X"AB",X"A5",X"B6",X"85",
		X"0B",X"A0",X"24",X"BD",X"E2",X"60",X"AA",X"A9",X"1C",X"20",X"00",X"66",X"A6",X"AB",X"CA",X"10",
		X"EA",X"60",X"A9",X"10",X"85",X"B3",X"A9",X"40",X"85",X"B2",X"A9",X"00",X"85",X"93",X"85",X"EC",
		X"A2",X"07",X"A9",X"0E",X"95",X"E4",X"CA",X"10",X"FB",X"20",X"86",X"69",X"A9",X"1C",X"20",X"51",
		X"6A",X"A9",X"1D",X"20",X"51",X"6A",X"A9",X"06",X"85",X"EA",X"A9",X"00",X"A2",X"13",X"9D",X"6E",
		X"01",X"CA",X"10",X"FA",X"A9",X"16",X"85",X"91",X"60",X"A5",X"B2",X"F0",X"05",X"C6",X"B2",X"B8",
		X"50",X"0E",X"C6",X"B3",X"D0",X"07",X"A9",X"00",X"85",X"91",X"B8",X"50",X"03",X"20",X"B3",X"62",
		X"60",X"20",X"2F",X"67",X"A9",X"40",X"85",X"CE",X"A5",X"93",X"F0",X"03",X"20",X"D6",X"5F",X"A9",
		X"00",X"85",X"DF",X"85",X"C1",X"85",X"C6",X"85",X"C3",X"85",X"C4",X"A9",X"01",X"85",X"A7",X"A6",
		X"AE",X"A5",X"F4",X"29",X"03",X"A8",X"B9",X"08",X"5B",X"95",X"C0",X"B9",X"0C",X"5B",X"95",X"C5",
		X"CA",X"10",X"F3",X"A9",X"02",X"85",X"91",X"60",X"06",X"04",X"05",X"07",X"FC",X"E8",X"F8",X"FC",
		X"A5",X"DF",X"85",X"B9",X"20",X"0C",X"7B",X"A9",X"10",X"20",X"EC",X"79",X"A5",X"93",X"D0",X"09",
		X"A0",X"01",X"84",X"A7",X"A9",X"12",X"B8",X"50",X"0B",X"A4",X"A7",X"C0",X"13",X"90",X"02",X"A0",
		X"13",X"B9",X"8F",X"60",X"85",X"8D",X"BE",X"C0",X"60",X"86",X"DB",X"A9",X"30",X"85",X"EC",X"20",
		X"1A",X"67",X"20",X"9E",X"5B",X"A9",X"FF",X"85",X"C2",X"A9",X"00",X"85",X"BF",X"85",X"96",X"85",
		X"8E",X"85",X"90",X"85",X"8F",X"85",X"DA",X"85",X"C9",X"85",X"D9",X"85",X"8C",X"85",X"D0",X"85",
		X"FA",X"85",X"B4",X"85",X"CC",X"85",X"CB",X"85",X"B3",X"85",X"CF",X"A2",X"AA",X"9D",X"17",X"01",
		X"CA",X"D0",X"FA",X"A9",X"E0",X"85",X"CD",X"A5",X"93",X"F0",X"03",X"20",X"CE",X"65",X"20",X"16",
		X"5F",X"A0",X"02",X"A9",X"0A",X"99",X"A0",X"00",X"20",X"6A",X"68",X"88",X"10",X"F5",X"20",X"5C",
		X"65",X"A9",X"04",X"85",X"92",X"A9",X"22",X"85",X"91",X"A9",X"1E",X"85",X"AF",X"60",X"A9",X"00",
		X"85",X"BA",X"85",X"BB",X"A5",X"A7",X"18",X"69",X"01",X"4A",X"C9",X"06",X"90",X"02",X"A9",X"06",
		X"85",X"DD",X"AA",X"F8",X"A5",X"BA",X"18",X"69",X"25",X"85",X"BA",X"A5",X"BB",X"69",X"00",X"85",
		X"BB",X"D8",X"CA",X"D0",X"EE",X"A4",X"A7",X"C0",X"0F",X"90",X"02",X"A0",X"0F",X"B9",X"A2",X"60",
		X"85",X"B7",X"B9",X"B1",X"60",X"85",X"B8",X"C0",X"08",X"90",X"02",X"A0",X"08",X"B9",X"D2",X"60",
		X"85",X"E1",X"B9",X"D9",X"60",X"85",X"E2",X"85",X"E3",X"60",X"20",X"37",X"5E",X"20",X"72",X"65",
		X"20",X"96",X"5F",X"A9",X"00",X"85",X"97",X"A2",X"10",X"A5",X"93",X"F0",X"20",X"A5",X"A0",X"05",
		X"A1",X"05",X"A2",X"F0",X"0A",X"A9",X"07",X"20",X"55",X"6A",X"A2",X"0A",X"B8",X"50",X"0E",X"A4",
		X"B9",X"B9",X"C5",X"00",X"F0",X"07",X"A9",X"07",X"20",X"55",X"6A",X"A2",X"0C",X"86",X"91",X"60",
		X"C6",X"B4",X"10",X"5D",X"A0",X"02",X"B9",X"A0",X"00",X"F0",X"3B",X"38",X"E9",X"01",X"99",X"A0",
		X"00",X"20",X"D1",X"67",X"20",X"BB",X"5F",X"A2",X"40",X"A0",X"80",X"A9",X"40",X"20",X"F6",X"6A",
		X"A9",X"82",X"49",X"FF",X"85",X"07",X"A5",X"97",X"0A",X"0A",X"18",X"69",X"7A",X"24",X"FC",X"50",
		X"02",X"49",X"FF",X"85",X"06",X"A9",X"E0",X"20",X"ED",X"67",X"E6",X"97",X"A9",X"05",X"85",X"B4",
		X"A9",X"08",X"20",X"EC",X"79",X"60",X"88",X"10",X"BD",X"A9",X"0C",X"85",X"92",X"A2",X"0F",X"A4",
		X"B9",X"B9",X"C5",X"00",X"F0",X"02",X"A2",X"00",X"86",X"AF",X"20",X"13",X"60",X"A9",X"22",X"85",
		X"91",X"60",X"A9",X"10",X"85",X"91",X"A4",X"B9",X"B9",X"C5",X"00",X"25",X"93",X"F0",X"0B",X"A2",
		X"00",X"0A",X"90",X"01",X"E8",X"C9",X"00",X"D0",X"F8",X"8A",X"F0",X"0D",X"86",X"97",X"A9",X"00",
		X"85",X"8D",X"A9",X"0E",X"85",X"91",X"20",X"96",X"5F",X"60",X"C6",X"B4",X"10",X"5D",X"A4",X"B9",
		X"B9",X"C5",X"00",X"85",X"98",X"A6",X"97",X"A0",X"06",X"88",X"A5",X"98",X"39",X"F7",X"60",X"F0",
		X"01",X"CA",X"E0",X"00",X"D0",X"F3",X"20",X"53",X"67",X"A2",X"03",X"20",X"A2",X"5F",X"A2",X"40",
		X"A0",X"60",X"A9",X"40",X"20",X"F6",X"6A",X"A5",X"8D",X"E6",X"8D",X"0A",X"0A",X"0A",X"0A",X"18",
		X"65",X"8D",X"18",X"69",X"80",X"AA",X"A0",X"60",X"A9",X"E4",X"20",X"95",X"67",X"A9",X"08",X"20",
		X"EC",X"79",X"A9",X"0A",X"85",X"B4",X"C6",X"97",X"D0",X"11",X"A9",X"10",X"85",X"92",X"A9",X"22",
		X"85",X"91",X"A9",X"0F",X"85",X"AF",X"A4",X"B9",X"20",X"13",X"60",X"60",X"A9",X"02",X"85",X"92",
		X"A9",X"00",X"85",X"AF",X"A9",X"22",X"85",X"91",X"20",X"ED",X"5D",X"A5",X"C0",X"05",X"C1",X"25",
		X"93",X"D0",X"07",X"A9",X"18",X"85",X"91",X"B8",X"50",X"42",X"A4",X"AE",X"F0",X"1D",X"A4",X"B9",
		X"B9",X"C0",X"00",X"D0",X"16",X"A9",X"07",X"20",X"49",X"6A",X"A9",X"09",X"20",X"49",X"6A",X"A9",
		X"0E",X"20",X"55",X"6A",X"20",X"48",X"5F",X"A9",X"0F",X"85",X"AF",X"A5",X"B9",X"85",X"DF",X"A4",
		X"AE",X"F0",X"10",X"C4",X"DF",X"D0",X"07",X"C6",X"DF",X"E6",X"A7",X"B8",X"50",X"02",X"E6",X"DF",
		X"B8",X"50",X"02",X"E6",X"A7",X"A4",X"DF",X"B9",X"C0",X"00",X"F0",X"E3",X"60",X"A2",X"1C",X"A5",
		X"93",X"F0",X"1E",X"A9",X"06",X"85",X"E4",X"85",X"E5",X"85",X"E6",X"85",X"E7",X"85",X"E9",X"85",
		X"EA",X"85",X"EB",X"A9",X"80",X"85",X"CE",X"20",X"E1",X"5F",X"A9",X"20",X"20",X"EC",X"79",X"A2",
		X"12",X"86",X"91",X"A0",X"00",X"8C",X"C3",X"01",X"84",X"AE",X"84",X"93",X"A0",X"01",X"8C",X"C2",
		X"01",X"60",X"AD",X"C2",X"01",X"85",X"B5",X"F0",X"3C",X"C9",X"6D",X"90",X"05",X"A9",X"6C",X"B8",
		X"50",X"1B",X"CD",X"C3",X"01",X"B0",X"06",X"38",X"E9",X"01",X"B8",X"50",X"10",X"18",X"69",X"01",
		X"48",X"C9",X"62",X"D0",X"05",X"A9",X"08",X"20",X"55",X"6A",X"C6",X"B5",X"68",X"8D",X"C2",X"01",
		X"85",X"9A",X"A4",X"B5",X"8C",X"C3",X"01",X"A9",X"80",X"85",X"9B",X"A9",X"73",X"85",X"9C",X"20",
		X"71",X"5E",X"B8",X"50",X"07",X"A9",X"1C",X"85",X"91",X"20",X"0C",X"7B",X"60",X"A5",X"93",X"F0",
		X"45",X"20",X"40",X"60",X"A4",X"B9",X"B6",X"C0",X"E0",X"06",X"90",X"02",X"A2",X"06",X"B9",X"C5",
		X"00",X"85",X"98",X"0A",X"90",X"01",X"CA",X"A8",X"D0",X"F9",X"8A",X"F0",X"29",X"86",X"DC",X"A4",
		X"B9",X"B9",X"C5",X"00",X"49",X"FC",X"A0",X"00",X"20",X"1D",X"58",X"A6",X"B9",X"B5",X"C5",X"19",
		X"F7",X"60",X"95",X"C5",X"C6",X"DC",X"D0",X"E7",X"A9",X"40",X"20",X"EC",X"79",X"A9",X"05",X"20",
		X"55",X"6A",X"A9",X"2D",X"85",X"AF",X"60",X"A5",X"8C",X"05",X"DA",X"F0",X"2C",X"A2",X"07",X"86",
		X"DC",X"A6",X"DC",X"BD",X"65",X"01",X"F0",X"1D",X"8A",X"18",X"69",X"08",X"85",X"97",X"A5",X"D9",
		X"3D",X"F7",X"60",X"D0",X"06",X"20",X"86",X"66",X"B8",X"50",X"0A",X"20",X"AC",X"77",X"A9",X"00",
		X"85",X"DA",X"20",X"E9",X"7A",X"C6",X"DC",X"10",X"D8",X"20",X"0C",X"7B",X"A9",X"0F",X"4C",X"49",
		X"6A",X"86",X"AC",X"A5",X"9A",X"C5",X"B5",X"F0",X"23",X"B0",X"12",X"A9",X"00",X"85",X"B6",X"20",
		X"9F",X"5E",X"A5",X"B5",X"C6",X"B5",X"C5",X"9A",X"D0",X"F5",X"B8",X"50",X"0F",X"A9",X"80",X"85",
		X"B6",X"20",X"9F",X"5E",X"A5",X"B5",X"C5",X"9A",X"E6",X"B5",X"90",X"F5",X"A6",X"AC",X"60",X"A6",
		X"B5",X"86",X"9D",X"A2",X"00",X"86",X"9E",X"20",X"CD",X"5E",X"A6",X"9D",X"A5",X"9E",X"86",X"9E",
		X"85",X"9D",X"20",X"CD",X"5E",X"E6",X"9D",X"A5",X"9D",X"85",X"9E",X"4A",X"18",X"65",X"9E",X"4A",
		X"4A",X"49",X"FF",X"38",X"65",X"B5",X"85",X"9D",X"C5",X"9E",X"B0",X"DB",X"60",X"A2",X"00",X"A5",
		X"9B",X"18",X"65",X"9D",X"85",X"B0",X"85",X"98",X"A5",X"9C",X"18",X"65",X"9E",X"49",X"FF",X"85",
		X"B1",X"A1",X"B0",X"29",X"20",X"05",X"B6",X"81",X"B0",X"A5",X"9B",X"38",X"E5",X"9D",X"85",X"B0",
		X"A1",X"B0",X"29",X"20",X"05",X"B6",X"81",X"B0",X"A5",X"9C",X"38",X"E5",X"9E",X"49",X"FF",X"85",
		X"B1",X"A1",X"B0",X"29",X"20",X"05",X"B6",X"81",X"B0",X"A5",X"98",X"85",X"B0",X"A1",X"B0",X"29",
		X"20",X"05",X"B6",X"81",X"B0",X"60",X"A5",X"93",X"F0",X"1D",X"20",X"48",X"5F",X"A9",X"06",X"20",
		X"55",X"6A",X"A5",X"DD",X"A2",X"40",X"86",X"0B",X"A2",X"58",X"A0",X"70",X"20",X"9D",X"6A",X"A9",
		X"1E",X"20",X"55",X"6A",X"B8",X"50",X"03",X"20",X"33",X"6C",X"A5",X"A7",X"C9",X"04",X"B0",X"05",
		X"A9",X"15",X"20",X"51",X"6A",X"4C",X"23",X"75",X"A9",X"00",X"20",X"55",X"6A",X"A5",X"B9",X"18",
		X"69",X"01",X"A2",X"40",X"86",X"0B",X"A2",X"9C",X"A0",X"90",X"4C",X"9D",X"6A",X"A5",X"CA",X"4A",
		X"B0",X"03",X"20",X"66",X"5F",X"60",X"20",X"8C",X"6B",X"A2",X"00",X"8A",X"29",X"3F",X"C9",X"3E",
		X"D0",X"08",X"38",X"7E",X"01",X"04",X"38",X"B8",X"50",X"0B",X"BD",X"03",X"04",X"4A",X"7E",X"01",
		X"04",X"BD",X"03",X"05",X"4A",X"7E",X"01",X"05",X"8A",X"18",X"69",X"40",X"AA",X"90",X"DC",X"E8",
		X"E8",X"E0",X"40",X"90",X"D6",X"60",X"A9",X"00",X"85",X"D1",X"85",X"D2",X"85",X"D3",X"60",X"20",
		X"96",X"5F",X"F8",X"A5",X"BA",X"18",X"65",X"D1",X"85",X"D1",X"A5",X"D2",X"65",X"BB",X"85",X"D2",
		X"A5",X"D3",X"69",X"00",X"85",X"D3",X"CA",X"10",X"EA",X"D8",X"60",X"A6",X"DD",X"F8",X"A9",X"05",
		X"18",X"65",X"D1",X"85",X"D1",X"A9",X"00",X"65",X"D2",X"85",X"D2",X"A5",X"D3",X"69",X"00",X"85",
		X"D3",X"CA",X"D0",X"EA",X"D8",X"60",X"A9",X"00",X"A2",X"05",X"9D",X"D6",X"01",X"CA",X"10",X"FA",
		X"60",X"A5",X"93",X"D0",X"0C",X"AD",X"D7",X"01",X"0D",X"D9",X"01",X"0D",X"DB",X"01",X"B8",X"50",
		X"02",X"A5",X"AE",X"F0",X"05",X"A0",X"01",X"20",X"FC",X"5F",X"A0",X"00",X"20",X"96",X"5F",X"20");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
