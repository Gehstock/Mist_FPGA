library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_spr_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_spr_bit2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"3C",X"3F",X"3F",X"3F",X"1F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"1F",X"3F",X"3F",X"3F",X"3C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"41",X"41",X"41",X"40",X"40",X"60",X"20",X"21",X"17",X"FE",X"FF",X"FF",X"E8",X"E0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"03",X"07",X"FF",X"FF",X"0F",X"07",X"00",
		X"00",X"E0",X"E8",X"FF",X"FF",X"FE",X"17",X"21",X"20",X"60",X"40",X"40",X"41",X"41",X"41",X"41",
		X"00",X"07",X"0F",X"FF",X"FF",X"07",X"03",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"83",X"83",X"83",X"83",X"C7",X"F7",X"FF",X"1F",X"3F",X"FE",X"FE",X"FE",X"EC",X"E0",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"13",X"19",X"78",X"D0",X"08",X"1B",X"77",X"C5",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"3F",X"3F",X"7E",X"FC",X"FC",X"D8",X"80",X"00",X"00",X"3F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"82",X"80",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"38",X"BC",X"7E",X"3E",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"13",X"19",X"78",X"D0",X"08",X"1B",X"77",X"C5",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"77",X"3F",X"7E",X"FC",X"F8",X"F0",X"80",X"00",X"00",X"3F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"82",X"80",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"70",X"F8",X"7C",X"3E",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"37",X"FF",X"38",X"31",X"33",X"63",X"C7",X"0D",X"0E",X"08",X"01",X"01",X"02",X"00",X"00",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"01",X"01",X"21",X"C1",X"F0",X"3C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"3F",X"47",X"43",X"7B",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"37",X"FF",X"38",X"31",X"33",X"63",X"C7",X"0D",X"0E",X"08",X"01",X"01",X"00",X"01",X"00",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"01",X"01",X"21",X"C1",X"F0",X"3C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"3F",X"47",X"43",X"7B",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"12",X"00",X"33",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"33",X"00",X"12",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"2D",X"00",X"4C",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"4C",X"00",X"2D",X"00",
		X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"80",X"40",X"30",X"08",X"18",X"F8",X"B8",X"18",X"18",X"18",X"18",X"30",X"70",X"B0",X"20",X"00",
		X"00",X"00",X"01",X"00",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"30",X"40",X"80",X"08",X"18",X"F8",X"B8",X"18",X"18",X"18",X"18",X"30",X"70",X"B0",X"20",X"00",
		X"1F",X"FF",X"FF",X"7F",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"FC",X"7C",X"3E",X"8E",X"CE",X"E7",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"01",X"19",X"98",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"98",X"19",X"01",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"0E",X"0E",X"0E",X"01",X"19",X"98",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"98",X"19",X"01",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"0F",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"CF",X"DF",X"FE",X"FC",X"FA",X"7F",X"3F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0B",X"1F",X"1F",X"0F",X"03",X"13",
		X"00",X"00",X"00",X"00",X"70",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"EF",
		X"81",X"01",X"03",X"03",X"01",X"0C",X"0E",X"87",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"3E",X"DE",X"FD",X"FB",X"FB",X"F6",X"C0",X"80",X"80",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"80",X"C0",
		X"81",X"01",X"03",X"03",X"01",X"0C",X"0E",X"87",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"E7",X"FB",X"FD",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"E1",X"9B",X"3C",X"24",X"24",X"24",X"24",X"3C",X"9B",X"E1",X"C0",X"C0",X"00",
		X"00",X"40",X"80",X"80",X"C0",X"70",X"00",X"00",X"00",X"00",X"70",X"C0",X"80",X"80",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"76",X"6F",X"FE",X"FD",X"FD",X"FD",X"FD",X"FE",X"6F",X"76",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"F0",X"D8",X"40",X"40",X"D8",X"F0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0E",X"0F",X"1F",X"3F",X"3F",X"1F",X"0F",X"0E",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"B0",X"A0",X"40",X"40",X"A0",X"B0",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"B0",X"EC",X"F4",X"E0",X"F4",X"EC",X"B0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"1E",X"3C",X"1E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"07",X"07",X"0F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"0F",X"07",X"07",X"07",X"01",
		X"80",X"D0",X"B0",X"78",X"F6",X"EE",X"E8",X"E8",X"E9",X"EF",X"F6",X"F8",X"70",X"B0",X"C0",X"80",
		X"00",X"00",X"20",X"60",X"F0",X"10",X"00",X"00",X"00",X"30",X"F0",X"60",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"00",X"00",X"00",
		X"1F",X"17",X"07",X"03",X"00",X"00",X"00",X"00",X"81",X"86",X"20",X"E0",X"01",X"17",X"1F",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"BF",X"3F",X"3E",X"3E",X"7E",X"78",X"38",X"70",X"E0",X"C0",X"80",X"00",X"00",
		X"60",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"38",X"B8",X"F8",X"FC",X"FE",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"60",X"40",X"00",X"40",X"40",X"80",X"00",X"10",X"30",
		X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"82",X"02",X"83",X"01",X"00",X"00",X"00",X"A0",X"F9",X"7F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"05",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FE",X"FC",X"FB",X"60",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"06",X"0C",X"0C",X"06",X"20",X"40",X"00",X"40",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FD",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"A0",X"E4",X"64",X"62",X"70",X"38",X"1F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"30",X"10",X"10",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"70",X"00",X"66",X"30",X"18",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"D0",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"18",X"3C",X"0E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"C0",X"E0",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"2F",X"20",X"30",X"34",X"22",X"20",X"01",X"01",X"03",X"02",X"00",
		X"FC",X"FC",X"F0",X"E0",X"F0",X"F8",X"38",X"10",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"18",X"30",X"38",X"30",X"30",X"72",X"62",X"64",X"70",X"70",X"78",X"78",X"7C",X"7C",
		X"40",X"C0",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"0E",X"76",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"60",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"03",X"07",X"03",X"31",X"78",X"78",X"78",X"7E",X"7F",X"7F",X"3F",X"03",X"01",
		X"FF",X"7F",X"7F",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"09",X"00",X"00",
		X"F8",X"D8",X"D8",X"98",X"38",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"CF",X"CF",X"86",X"81",X"9C",X"B8",X"F8",X"F8",X"F8",X"FC",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"20",X"60",X"40",X"C0",X"80",X"00",X"00",X"50",X"78",X"7C",X"FC",X"FC",X"FC",X"E8",X"E0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"41",X"E2",X"C6",X"C6",X"E4",X"C6",
		X"00",X"00",X"00",X"00",X"60",X"40",X"C0",X"80",X"82",X"06",X"04",X"0C",X"08",X"18",X"10",X"30",
		X"01",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"FF",X"C7",X"C3",X"C3",X"E3",X"E3",X"E3",X"C3",X"C7",X"FF",X"1F",X"0F",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"01",X"03",X"07",X"07",X"C7",X"E7",X"A7",X"87",X"C7",X"87",X"C3",X"80",X"E3",X"F7",X"F7",
		X"40",X"10",X"7E",X"7E",X"3F",X"1F",X"0E",X"06",X"1E",X"0E",X"16",X"DC",X"DC",X"EC",X"FC",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"F0",X"F0",X"60",X"81",X"C7",X"DC",X"F0",X"C0",X"C0",X"C0",X"40",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"17",X"07",X"07",X"03",X"03",X"03",X"01",X"01",
		X"CF",X"C5",X"C6",X"DA",X"C3",X"E1",X"61",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"60",X"20",X"00",X"00",X"00",X"00",
		X"FB",X"FB",X"FB",X"F9",X"FD",X"FD",X"FC",X"FC",X"FE",X"FE",X"FE",X"9E",X"9D",X"8E",X"CE",X"C7",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"60",X"60",X"60",X"60",X"40",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"08",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"30",X"70",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"ED",X"C7",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"1F",X"3F",
		X"00",X"00",X"00",X"01",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"64",X"4C",X"48",X"78",X"B0",X"08",X"0F",X"86",X"04",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"BF",X"6F",X"F6",X"D4",X"E0",X"F0",X"E0",X"E0",X"80",X"19",X"3F",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"3C",X"3F",X"3F",X"3F",X"1B",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"1B",X"3F",X"3F",X"3F",X"3C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"41",X"41",X"41",X"40",X"40",X"60",X"20",X"21",X"17",X"FE",X"FF",X"FF",X"F8",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"03",X"07",X"FF",X"FF",X"0B",X"03",X"00",
		X"00",X"F0",X"F8",X"FF",X"FF",X"FE",X"17",X"21",X"20",X"60",X"40",X"40",X"41",X"41",X"41",X"41",
		X"00",X"03",X"0B",X"FF",X"FF",X"07",X"03",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"83",X"83",X"83",X"83",X"C7",X"F7",X"FF",X"1F",X"3F",X"FE",X"FE",X"FE",X"FC",X"F0",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"FC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"82",X"E2",X"FA",X"FF",X"FF",X"FF",X"3F",X"0D",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"F7",X"E1",X"C0",X"F8",X"3E",X"0F",X"03",X"01",X"01",
		X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"02",X"02",
		X"F8",X"FC",X"7F",X"1F",X"37",X"62",X"43",X"C1",X"81",X"81",X"01",X"01",X"05",X"05",X"05",X"0D",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"FC",X"7C",X"66",X"C3",X"FF",X"FF",X"FF",X"FF",X"7F",X"1B",X"00",
		X"1C",X"1C",X"1C",X"38",X"38",X"38",X"78",X"F0",X"E0",X"F0",X"20",X"20",X"C0",X"80",X"C0",X"C0",
		X"C3",X"FB",X"3F",X"0F",X"07",X"C7",X"F6",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"00",X"C0",X"F0",X"F0",X"F8",X"FC",X"7C",X"3C",X"BE",X"FE",X"FE",X"0E",X"0E",X"0C",X"0E",X"0C",
		X"0E",X"0E",X"0E",X"0E",X"0D",X"0D",X"0D",X"03",X"07",X"07",X"03",X"02",X"00",X"00",X"00",X"00",
		X"9F",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0E",X"06",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"07",X"0F",X"0F",
		X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"C7",X"80",X"80",X"00",X"00",X"80",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"2F",X"FF",X"FF",X"F0",X"C0",X"E0",X"E0",X"A0",X"30",X"3F",X"3F",X"FF",
		X"F8",X"F8",X"F8",X"FC",X"7F",X"79",X"60",X"30",X"18",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"0C",X"08",X"DF",X"FF",X"3F",X"1B",X"F3",X"F1",X"FB",X"7F",X"7F",X"3F",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1C",X"38",X"78",X"78",X"F8",X"F8",X"F8",
		X"00",X"00",X"03",X"03",X"07",X"3F",X"FF",X"FF",X"08",X"0C",X"04",X"04",X"04",X"04",X"04",X"04",
		X"01",X"01",X"07",X"3F",X"F7",X"EF",X"EF",X"EF",X"E6",X"F1",X"FF",X"FF",X"FF",X"FF",X"BF",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"F8",X"F8",X"F8",X"F0",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"37",X"EF",X"EF",X"EF",X"E6",X"F1",X"FF",X"07",X"00",X"00",X"00",X"01",X"03",X"03",X"03",
		X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"10",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"CE",X"47",X"61",X"3F",X"1F",X"0F",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"0E",X"38",X"70",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"C3",X"8E",X"FD",X"FD",X"3C",X"7E",X"3F",X"FF",X"F7",
		X"FF",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"B0",X"70",X"E0",X"F8",X"F0",
		X"FC",X"8E",X"C3",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"B8",X"78",X"C8",X"00",X"18",X"38",X"78",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"7D",X"3D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"04",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"D7",X"7F",X"3F",X"E7",X"E7",X"7F",X"3D",X"00",
		X"7B",X"7B",X"7B",X"78",X"78",X"78",X"38",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"F8",X"00",
		X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"D7",X"09",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"E0",X"18",X"38",X"78",X"78",X"7B",X"7B",X"7B",
		X"31",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"79",X"7C",X"27",X"31",X"1F",X"07",X"03",X"00",
		X"1C",X"1F",X"1F",X"1F",X"1F",X"1F",X"1C",X"0C",X"3C",X"FC",X"FC",X"FC",X"F8",X"F0",X"BC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0C",X"19",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"3C",X"00",
		X"00",X"00",X"01",X"03",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"03",X"01",X"00",X"00",
		X"1C",X"7E",X"FE",X"0E",X"02",X"06",X"07",X"07",X"07",X"07",X"06",X"02",X"0E",X"FE",X"7E",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"7E",X"CE",X"82",X"86",X"87",X"87",X"86",X"82",X"CE",X"7E",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1E",X"36",X"36",X"36",X"36",X"36",X"36",X"1E",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0A",X"0A",X"0A",X"0A",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"A0",X"A0",X"B0",X"D0",X"40",X"4C",X"5F",X"7D",X"7C",X"3D",X"2F",X"07",X"03",
		X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"C0",X"F8",X"FF",X"FF",X"FF",X"FE",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"18",X"7C",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"F8",X"C0",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"7C",X"18",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"E0",X"E0",X"E0",X"FF",X"7F",X"7F",X"60",X"60",X"60",X"7F",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"80",
		X"7F",X"FE",X"FE",X"70",X"7F",X"7F",X"7F",X"60",X"60",X"E0",X"FF",X"FF",X"FF",X"E0",X"E0",X"E0",
		X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"03",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FE",
		X"03",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FE",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"22",X"22",X"22",X"1C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"3E",X"3E",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1A",X"3A",X"2E",X"26",X"36",X"12",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"14",X"3E",X"2A",X"22",X"36",X"14",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"3E",X"3E",X"34",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"2E",X"2A",X"3A",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"2E",X"2A",X"2A",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"2E",X"26",X"20",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"14",X"2E",X"2A",X"2A",X"3A",X"14",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"3E",X"2A",X"2A",X"3A",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"80",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"01",X"07",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"C0",X"00",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"06",X"03",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"60",X"00",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"06",X"07",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"06",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"60",X"E0",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"06",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"00",X"20",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"06",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"20",X"C0",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"06",X"07",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"C0",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"1C",X"00",X"02",X"02",X"02",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"2A",X"2A",X"12",X"00",X"1C",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"1C",X"00",X"2A",X"2A",X"3E",X"00",X"30",X"0C",X"02",X"0C",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"2A",X"2A",X"12",X"00",X"1E",X"24",X"24",X"1E",X"00",X"2E",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"00",X"3C",X"02",X"02",X"3C",X"00",X"1C",X"22",X"22",X"1C",X"00",X"3E",X"08",X"08",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"08",X"10",X"3E",X"00",X"1C",X"22",X"22",X"1C",X"00",X"20",X"3E",X"20",X"04",X"2A",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"1C",X"00",X"3E",X"00",X"3E",X"08",X"08",X"3E",X"00",X"22",X"22",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"22",X"22",X"1C",X"00",X"2E",X"2A",X"22",X"1C",X"00",X"1E",X"24",X"24",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"3E",X"08",X"10",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"30",X"08",X"0E",X"08",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"14",X"5C",X"0F",X"1B",X"77",X"94",X"20",X"84",X"10",X"42",X"90",X"05",X"20",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"80",X"12",X"40",X"08",X"21",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"20",X"05",X"90",X"42",X"10",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"21",X"08",X"40",X"12",X"80",X"00",
		X"20",X"68",X"F0",X"90",X"18",X"98",X"F0",X"50",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"7F",X"E0",X"C0",X"C0",X"C0",X"E0",X"7F",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"38",X"18",X"18",X"18",X"38",X"F0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"E7",X"C3",X"C3",X"C1",X"E1",X"F0",X"70",X"30",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",X"98",X"98",X"D8",X"F8",X"F8",X"78",X"18",
		X"00",X"00",X"00",X"00",X"00",X"38",X"7D",X"FF",X"EF",X"C6",X"C6",X"C6",X"E0",X"F0",X"70",X"30",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"38",X"18",X"18",X"18",X"38",X"78",X"70",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"3F",X"3F",X"3F",X"1F",X"07",X"07",X"03",X"01",
		X"6C",X"7E",X"FE",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"FC",X"F8",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"01",X"01",X"01",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"3F",X"29",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"29",X"3F",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"01",X"01",X"21",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"3F",X"29",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"29",X"3F",X"1E",
		X"00",X"C0",X"F0",X"FC",X"FF",X"7F",X"FF",X"87",X"87",X"FF",X"7F",X"FF",X"FC",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"81",X"81",X"81",X"80",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"7C",X"3F",X"03",X"01",X"00",X"00",X"00",X"00",
		X"7C",X"8C",X"86",X"F7",X"7F",X"3F",X"FF",X"7F",X"FF",X"FE",X"FC",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"1E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"03",X"06",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0A",X"40",X"40",X"80",X"80",X"00",X"C0",X"D0",X"70",
		X"3F",X"7F",X"FF",X"FF",X"7E",X"F8",X"E0",X"5F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"00",X"00",X"00",X"01",X"01",X"E3",X"FD",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"38",X"1C",X"3C",X"46",X"42",X"7B",X"3F",X"9F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"03",X"06",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0A",X"40",X"40",X"80",X"80",X"00",X"C0",X"D0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"01",X"01",X"21",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"28",X"01",X"01",X"41",X"03",X"02",X"02",X"03",X"41",X"01",X"01",X"28",X"3F",X"1F",
		X"80",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"1F",X"1F",X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"81",X"81",X"81",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"01",X"01",X"41",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"28",X"01",X"01",X"41",X"03",X"02",X"02",X"03",X"41",X"01",X"01",X"28",X"3F",X"1F",
		X"80",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"1F",X"1F",X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"81",X"81",X"81",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"07",X"0C",X"00",
		X"00",X"1F",X"3F",X"2A",X"02",X"03",X"01",X"04",X"03",X"00",X"40",X"C0",X"80",X"29",X"3F",X"1F",
		X"00",X"C0",X"F0",X"3C",X"1E",X"DF",X"FF",X"FF",X"FF",X"7F",X"77",X"7F",X"FF",X"FE",X"F0",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"81",X"81",X"81",X"01",X"00",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"06",X"0C",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"41",
		X"00",X"00",X"00",X"00",X"00",X"1F",X"3E",X"2E",X"03",X"01",X"04",X"03",X"00",X"40",X"E8",X"BE",
		X"EF",X"FF",X"FE",X"F8",X"C1",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"03",X"01",X"40",X"FC",X"FC",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"38",X"1C",X"DE",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"81",
		X"03",X"26",X"0C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"20",X"01",
		X"00",X"00",X"00",X"00",X"00",X"1F",X"3E",X"2A",X"03",X"01",X"04",X"03",X"00",X"40",X"E8",X"BE",
		X"EF",X"FF",X"FE",X"F8",X"C1",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"03",X"01",X"40",X"FC",X"FC",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"3C",X"1E",X"DF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"81",
		X"00",X"00",X"00",X"07",X"01",X"01",X"11",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"01",X"01",X"5D",X"3F",X"21",X"21",X"3F",X"5D",X"01",X"01",X"21",X"36",X"17",X"03",X"00",
		X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"E0",X"60",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"E0",
		X"00",X"00",X"00",X"0F",X"01",X"01",X"41",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2B",X"03",X"03",X"5F",X"3F",X"21",X"21",X"3F",X"5F",X"03",X"03",X"2B",X"3D",X"1E",X"03",X"00",
		X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"E0",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"07",X"0C",X"00",X"00",X"00",X"00",
		X"3F",X"23",X"21",X"3D",X"1F",X"0F",X"1B",X"43",X"C3",X"81",X"29",X"3E",X"1F",X"00",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"DE",X"BC",X"F8",X"E0",X"C3",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"7C",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"01",X"01",X"01",X"00",X"00",X"10",X"01",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",
		X"21",X"3D",X"1F",X"0F",X"5B",X"63",X"E3",X"85",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"9E",X"FE",X"FC",X"F8",X"E3",X"EF",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"01",X"40",X"7C",X"FC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"FC",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"41",X"03",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"21",X"3D",X"1F",X"0D",X"59",X"69",X"F9",X"9E",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"DE",X"FE",X"FC",X"F8",X"E3",X"EF",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"40",X"7C",X"FC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3D",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"15",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"50",X"7F",X"3F",X"00",
		X"C0",X"E0",X"FC",X"FF",X"FF",X"7F",X"FF",X"87",X"87",X"FF",X"7F",X"FC",X"F8",X"F0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"81",X"81",X"81",X"81",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"1F",X"17",X"40",X"40",X"80",X"80",X"00",X"00",X"28",X"38",
		X"3F",X"3F",X"7F",X"FF",X"FE",X"F8",X"E0",X"5F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"01",X"01",X"E3",X"FD",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"78",X"1C",X"3C",X"46",X"42",X"7B",X"3F",X"9F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"E7",X"E3",X"E3",X"E2",
		X"80",X"80",X"90",X"90",X"92",X"92",X"D0",X"B0",X"98",X"8C",X"8C",X"C8",X"A0",X"80",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"B8",X"9C",X"8F",X"87",X"C3",X"E3",X"91",X"88",X"80",X"80",X"E0",X"BC",X"9F",X"87",X"83",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"87",X"83",X"81",X"C0",X"E0",X"B8",X"9C",X"87",X"83",X"82",X"82",X"92",X"92",X"82",X"82",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"90",X"90",X"90",X"90",X"82",X"82",X"C2",X"A2",X"9A",X"8E",X"8F",X"CF",X"A7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F8",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"67",X"61",X"60",X"60",X"70",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"70",X"78",X"FE",X"FF",X"EF",X"E7",X"E1",X"60",X"60",X"70",X"78",X"FE",X"FF",X"FF",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"DC",X"FC",X"FC",X"FC",X"3F",X"1F",X"07",X"02",X"00",X"C0",
		X"FF",X"FF",X"FF",X"6F",X"67",X"63",X"63",X"63",X"E3",X"E3",X"63",X"63",X"63",X"63",X"63",X"61",
		X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"3E",X"1F",X"07",X"03",X"00",X"00",X"00",X"18",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"60",X"60",X"60",X"70",X"78",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7C",X"58",X"70",X"40",X"80",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"70",X"78",X"7C",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C6",X"C7",X"C7",X"C7",X"E7",X"F7",X"FE",X"FC",X"F8",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"18",X"08",X"08",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F3",X"F1",X"F1",X"D1",X"CD",X"CF",X"C7",X"C3",X"C3",X"C1",X"C0",X"C0",X"C0",X"C4",X"C4",
		X"04",X"80",X"C0",X"70",X"38",X"0E",X"07",X"81",X"C0",X"F0",X"F8",X"FE",X"F9",X"78",X"38",X"38",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"30",X"38",X"0C",X"04",X"80",X"C0",X"70",X"38",X"0E",X"07",X"01",X"00",X"30",X"38",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"1F",X"0F",X"87",X"C7",X"E3",X"11",X"00",X"00",X"00",X"F0",X"7F",X"3F",X"0F",X"07",X"01",
		X"00",X"80",X"C0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"FC",X"FE",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"39",X"19",X"09",X"09",X"C9",X"E1",X"F1",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"00",X"80",X"C0",X"F0",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"39",X"19",X"09",X"09",X"C9",X"E9",X"F9",X"F9",X"F9",
		X"FC",X"FC",X"FC",X"7C",X"3C",X"0E",X"07",X"01",X"00",X"00",X"10",X"18",X"18",X"18",X"08",X"00",
		X"F0",X"F8",X"F8",X"F9",X"F9",X"F9",X"F9",X"F9",X"79",X"39",X"19",X"09",X"87",X"C3",X"E3",X"F1",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FD",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"83",X"83",X"93",X"93",X"83",X"83",X"C3",X"E7",X"FF",X"9F",X"03",X"03",X"03",X"00",X"60",
		X"80",X"C0",X"E0",X"F8",X"FC",X"FE",X"FF",X"FE",X"FC",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"38",X"1C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
