library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_graphx_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_graphx_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"80",X"80",X"81",X"81",X"80",X"80",X"00",X"00",X"08",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"FB",X"FD",X"FB",X"F7",X"F7",X"FF",X"0F",X"1F",X"FF",X"BF",X"BF",X"BF",X"3F",X"7F",X"FF",
		X"FF",X"FE",X"FC",X"FE",X"FD",X"FD",X"FF",X"F8",X"F0",X"FF",X"EF",X"EF",X"EF",X"9F",X"7E",X"00",
		X"FF",X"3F",X"BF",X"7F",X"BF",X"BF",X"FF",X"1F",X"0F",X"FF",X"F7",X"F7",X"F7",X"FB",X"7B",X"00",
		X"00",X"7F",X"9F",X"EF",X"EF",X"EF",X"FF",X"F0",X"F8",X"FF",X"FD",X"FD",X"FE",X"FC",X"FF",X"FF",
		X"00",X"FD",X"FD",X"FB",X"F7",X"EF",X"EF",X"F7",X"F7",X"CF",X"BF",X"BF",X"7F",X"7F",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FD",X"FD",X"FD",X"FB",X"E7",X"F7",X"CF",X"BF",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"3F",X"DF",X"DF",X"EF",X"EF",X"F7",X"FB",X"FD",X"00",
		X"00",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"80",X"BF",X"BF",X"DF",X"DF",X"EF",X"DF",X"EF",X"F7",X"F7",X"FB",X"FB",X"F9",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",
		X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F0",X"F0",X"F8",X"F8",X"FC",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FE",X"FC",X"F8",X"F8",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"05",X"07",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"04",X"03",X"0F",X"05",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0E",X"04",X"03",X"02",X"06",X"0C",X"03",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"05",X"0F",X"05",X"02",X"03",X"07",X"0D",X"02",X"03",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"0F",X"05",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"0C",X"06",X"04",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"09",X"0D",X"07",X"05",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"02",X"0E",X"04",X"03",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"0F",X"05",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"06",X"04",X"0E",X"04",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"0F",X"05",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"03",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"03",X"02",X"06",X"0C",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"07",X"0D",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"06",X"04",X"03",X"02",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"04",X"03",X"02",X"03",X"07",X"05",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"09",X"05",X"02",X"03",X"02",X"03",X"02",X"03",X"0F",X"05",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"06",X"04",X"03",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"05",X"02",X"03",X"0F",X"05",X"02",X"03",X"0A",X"00",
		X"08",X"09",X"0D",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"06",X"00",
		X"02",X"03",X"02",X"06",X"0C",X"03",X"02",X"06",X"04",X"03",X"02",X"0E",X"04",X"03",X"07",X"0B",
		X"03",X"02",X"03",X"07",X"0D",X"02",X"03",X"07",X"05",X"02",X"03",X"0F",X"05",X"02",X"06",X"04",
		X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"07",X"05",
		X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"02",
		X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0A",X"00",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"09",X"0D",X"02",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"08",X"09",X"0D",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"08",X"02",X"06",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"06",X"0C",X"03",X"07",X"05",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"07",X"0D",X"02",X"0E",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"00",X"08",X"0A",X"08",X"09",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"08",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"06",X"04",X"03",X"02",X"03",X"0F",X"05",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"09",X"0D",X"07",X"05",X"02",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"06",X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"0B",X"09",X"0B",X"02",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"06",X"0C",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"08",X"09",X"0D",X"07",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"06",X"0C",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"08",X"02",X"03",X"07",X"0D",X"07",X"0B",X"0A",X"08",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"0E",X"04",X"0E",X"04",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"0F",X"05",X"0F",X"05",X"02",X"0E",X"0C",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"08",X"09",X"0D",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0B",X"0A",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"06",X"04",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"03",X"07",X"05",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"0C",X"06",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0D",X"07",X"0B",X"0A",X"00",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"0E",X"04",X"03",X"02",X"03",X"0A",X"08",X"0A",X"00",X"00",X"00",
		X"08",X"09",X"0D",X"02",X"03",X"0F",X"05",X"02",X"0E",X"04",X"03",X"02",X"03",X"0A",X"08",X"0A",
		X"02",X"03",X"02",X"03",X"02",X"06",X"04",X"03",X"0F",X"05",X"02",X"06",X"04",X"03",X"02",X"03",
		X"03",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"02",
		X"04",X"03",X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
