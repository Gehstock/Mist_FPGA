library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GALAXIAN_1K is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"82",X"82",X"82",X"82",X"7C",X"00",X"00",X"02",X"02",X"FE",X"42",X"02",X"00",X"00",
		X"00",X"62",X"92",X"8A",X"86",X"86",X"42",X"00",X"00",X"8C",X"D2",X"B2",X"92",X"82",X"84",X"00",
		X"00",X"08",X"FE",X"48",X"28",X"18",X"08",X"00",X"00",X"1C",X"A2",X"A2",X"A2",X"A6",X"E4",X"00",
		X"00",X"8C",X"92",X"92",X"92",X"52",X"3C",X"00",X"00",X"C0",X"A0",X"90",X"8E",X"80",X"80",X"00",
		X"00",X"6C",X"92",X"92",X"92",X"92",X"6C",X"00",X"00",X"7C",X"92",X"92",X"92",X"92",X"60",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0C",X"08",X"0C",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"18",X"42",X"24",X"81",X"81",X"24",X"42",X"18",
		X"40",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"18",X"00",X"00",X"81",X"81",X"00",X"00",X"18",X"00",X"40",X"20",X"10",X"08",X"04",X"02",X"00",
		X"3C",X"42",X"A5",X"A5",X"A5",X"99",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"1C",X"0E",X"07",X"02",
		X"00",X"0C",X"0C",X"0C",X"06",X"06",X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"00",
		X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"02",X"07",X"0E",X"1C",X"38",X"30",X"00",X"00",
		X"00",X"06",X"06",X"06",X"0C",X"0C",X"0C",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"00",
		X"00",X"00",X"06",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"E3",X"A1",X"CD",X"C2",X"F1",X"E7",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"1F",X"1F",X"0F",X"07",X"03",X"20",X"1D",X"01",X"01",X"01",X"01",X"01",X"01",
		X"3E",X"3F",X"FE",X"FE",X"FE",X"FE",X"3F",X"3E",X"01",X"01",X"01",X"01",X"01",X"01",X"1D",X"20",
		X"00",X"00",X"00",X"00",X"00",X"01",X"22",X"0C",X"08",X"10",X"20",X"40",X"80",X"00",X"00",X"00",
		X"08",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"08",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",
		X"0C",X"22",X"01",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1E",X"1E",X"1E",X"3E",X"3F",X"3E",X"FE",X"FE",X"FE",X"3E",X"3F",X"3E",X"3E",
		X"3F",X"3E",X"1E",X"1E",X"1E",X"1C",X"1C",X"1C",X"3E",X"3E",X"3F",X"3E",X"FE",X"FE",X"FE",X"3E",
		X"00",X"03",X"00",X"10",X"08",X"04",X"40",X"40",X"00",X"C0",X"00",X"08",X"10",X"20",X"02",X"02",
		X"40",X"40",X"04",X"08",X"10",X"00",X"03",X"00",X"02",X"02",X"20",X"10",X"08",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"CC",
		X"03",X"03",X"01",X"01",X"03",X"06",X"0C",X"00",X"98",X"B0",X"F0",X"F0",X"F0",X"F0",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"40",X"40",X"40",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"03",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"FC",X"FC",X"F8",X"F8",X"EC",X"C4",X"80",X"00",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"00",X"40",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"01",X"01",
		X"48",X"68",X"7E",X"70",X"60",X"40",X"40",X"40",X"09",X"0B",X"3F",X"07",X"03",X"01",X"01",X"01",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"11",X"F0",X"E0",X"C0",X"80",X"80",X"80",X"80",X"C4",
		X"11",X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"C4",X"C4",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"1F",X"80",X"80",X"80",X"80",X"C0",X"E0",X"E0",X"E0",
		X"1F",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"01",X"11",X"17",X"3F",X"00",X"00",X"00",X"00",X"80",X"80",X"A0",X"F0",
		X"3F",X"17",X"11",X"00",X"00",X"00",X"00",X"00",X"F0",X"A0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"03",X"07",X"0F",X"0F",X"0F",X"03",X"01",X"0F",X"0F",X"1F",X"1F",X"0F",X"07",X"03",X"01",
		X"7F",X"3F",X"3F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",X"07",X"0F",X"1F",X"1F",X"0F",
		X"7F",X"3F",X"1F",X"0F",X"1F",X"1F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"0F",X"0F",X"1F",X"3F",X"FF",X"1F",X"1F",X"3F",X"7F",X"3F",X"7F",X"FF",X"FF",
		X"FF",X"7F",X"7F",X"3F",X"7F",X"3F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"7F",X"60",X"C0",X"00",X"00",X"00",X"00",X"F8",X"FE",X"06",X"03",
		X"C0",X"C0",X"E0",X"FF",X"FF",X"7F",X"7F",X"1F",X"03",X"03",X"07",X"FF",X"FF",X"FE",X"FE",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"7E",X"63",X"C1",X"00",X"00",X"00",X"00",X"7F",X"7F",X"C0",X"80",
		X"C1",X"C1",X"E1",X"FF",X"FF",X"7F",X"7F",X"1F",X"80",X"80",X"80",X"FC",X"FE",X"FF",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"78",X"7E",X"C6",X"83",X"00",X"00",X"00",X"FC",X"FE",X"FF",X"FE",X"FC",
		X"83",X"83",X"87",X"FF",X"FF",X"FE",X"FE",X"F8",X"00",X"00",X"00",X"21",X"73",X"FB",X"73",X"21",
		X"00",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"E0",X"C0",X"C0",X"C0",X"FE",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"01",X"03",X"07",X"00",X"00",X"00",X"F8",X"FE",X"FF",X"FF",X"FF",
		X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"7F",X"1F",X"FE",X"FC",X"F0",X"E0",X"C0",X"80",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"06",X"09",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"10",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"08",X"10",X"10",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"20",
		X"10",X"10",X"08",X"07",X"00",X"00",X"00",X"00",X"20",X"20",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"08",X"10",X"10",X"10",X"00",X"00",X"F0",X"08",X"04",X"02",X"02",X"02",
		X"10",X"10",X"10",X"08",X"04",X"03",X"00",X"00",X"02",X"02",X"02",X"04",X"08",X"F0",X"00",X"00",
		X"0F",X"10",X"20",X"40",X"C0",X"80",X"82",X"82",X"E0",X"10",X"08",X"46",X"03",X"01",X"01",X"81",
		X"80",X"81",X"82",X"C0",X"48",X"20",X"10",X"0F",X"09",X"81",X"01",X"03",X"02",X"04",X"08",X"F0",
		X"00",X"00",X"20",X"19",X"08",X"00",X"20",X"03",X"00",X"00",X"00",X"60",X"00",X"10",X"00",X"20",
		X"07",X"23",X"15",X"55",X"02",X"00",X"00",X"00",X"80",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0B",X"07",X"03",X"27",X"00",X"00",X"00",X"20",X"40",X"00",X"80",X"C0",
		X"17",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"D0",X"90",X"90",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"10",X"08",X"04",X"25",X"17",X"15",X"00",X"10",X"20",X"40",X"60",X"E0",X"C8",X"C2",
		X"07",X"03",X"01",X"00",X"08",X"11",X"21",X"00",X"DC",X"C0",X"C8",X"E0",X"C8",X"44",X"00",X"00",
		X"08",X"08",X"08",X"04",X"14",X"03",X"01",X"03",X"00",X"80",X"84",X"98",X"A0",X"A0",X"80",X"C4",
		X"07",X"07",X"07",X"01",X"04",X"10",X"20",X"00",X"E2",X"CC",X"F0",X"88",X"40",X"44",X"40",X"40");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
