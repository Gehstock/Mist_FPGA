library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tn01 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tn01 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"C3",X"18",X"00",X"00",X"00",X"FB",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E5",X"D5",X"C5",X"F5",X"C3",X"D8",X"04",X"FF",X"31",X"00",X"24",X"CD",X"76",X"01",X"06",X"00",
		X"CD",X"BC",X"04",X"CD",X"C5",X"04",X"CD",X"D0",X"04",X"CD",X"4C",X"00",X"FB",X"AF",X"D3",X"03",
		X"D3",X"05",X"CD",X"BC",X"00",X"CD",X"BB",X"01",X"CD",X"C1",X"00",X"CD",X"24",X"01",X"CD",X"01",
		X"01",X"CD",X"BB",X"01",X"CD",X"55",X"00",X"D3",X"06",X"C3",X"2D",X"00",X"21",X"3C",X"09",X"CD",
		X"7B",X"1A",X"C3",X"35",X"1B",X"CD",X"BA",X"04",X"CD",X"C5",X"04",X"21",X"2F",X"20",X"34",X"21",
		X"E0",X"20",X"34",X"CD",X"52",X"1A",X"2E",X"06",X"06",X"12",X"70",X"2E",X"0A",X"70",X"2E",X"0E",
		X"70",X"2E",X"12",X"70",X"2E",X"16",X"70",X"2E",X"1A",X"70",X"21",X"35",X"20",X"AF",X"BE",X"C2",
		X"A5",X"00",X"CD",X"94",X"00",X"21",X"54",X"20",X"34",X"CD",X"DB",X"16",X"CD",X"18",X"12",X"D3",
		X"06",X"C3",X"7A",X"00",X"21",X"14",X"20",X"AF",X"BE",X"C0",X"3A",X"01",X"20",X"E6",X"7F",X"C0",
		X"23",X"23",X"36",X"01",X"C9",X"CD",X"9A",X"18",X"21",X"E0",X"20",X"36",X"00",X"CD",X"BA",X"04",
		X"CD",X"C5",X"04",X"C3",X"C1",X"00",X"3E",X"FF",X"32",X"DF",X"20",X"C9",X"AF",X"32",X"DF",X"20",
		X"C9",X"3E",X"50",X"C3",X"D5",X"14",X"21",X"05",X"26",X"11",X"D7",X"00",X"01",X"08",X"01",X"CD",
		X"D5",X"01",X"06",X"17",X"C3",X"60",X"02",X"3C",X"42",X"99",X"A5",X"A5",X"81",X"42",X"3C",X"1B",
		X"21",X"29",X"28",X"20",X"1B",X"13",X"00",X"08",X"13",X"0E",X"1B",X"02",X"0E",X"11",X"0F",X"0E",
		X"11",X"00",X"13",X"08",X"0E",X"0D",X"01",X"0E",X"0C",X"01",X"04",X"11",X"3E",X"20",X"C3",X"D5",
		X"14",X"CD",X"BB",X"01",X"CD",X"C6",X"00",X"CD",X"FC",X"00",X"21",X"11",X"2C",X"06",X"0C",X"11",
		X"18",X"01",X"CD",X"60",X"02",X"C3",X"C1",X"00",X"08",X"0D",X"12",X"04",X"11",X"13",X"1B",X"1B",
		X"02",X"0E",X"08",X"0D",X"11",X"A0",X"20",X"21",X"A0",X"46",X"06",X"15",X"CD",X"8B",X"03",X"CD",
		X"82",X"17",X"21",X"AA",X"20",X"34",X"3A",X"AA",X"20",X"A7",X"D3",X"06",X"C2",X"36",X"01",X"CD",
		X"FC",X"00",X"21",X"0C",X"2E",X"11",X"F6",X"00",X"06",X"06",X"CD",X"60",X"02",X"CD",X"C1",X"00",
		X"CD",X"C6",X"00",X"11",X"A0",X"20",X"21",X"81",X"18",X"06",X"15",X"CD",X"8B",X"03",X"CD",X"82",
		X"17",X"21",X"AA",X"20",X"34",X"3A",X"AA",X"20",X"A7",X"D3",X"06",X"C2",X"65",X"01",X"3E",X"80",
		X"CD",X"D5",X"14",X"C3",X"76",X"01",X"21",X"00",X"24",X"AF",X"77",X"23",X"7C",X"FE",X"40",X"DA",
		X"79",X"01",X"C9",X"21",X"1E",X"25",X"11",X"E0",X"43",X"06",X"1A",X"CD",X"60",X"02",X"21",X"1D",
		X"26",X"11",X"C3",X"20",X"CD",X"B1",X"01",X"21",X"1D",X"30",X"11",X"DC",X"20",X"CD",X"B1",X"01",
		X"3A",X"DA",X"20",X"A7",X"CA",X"B0",X"01",X"21",X"1D",X"39",X"11",X"C6",X"20",X"CD",X"B1",X"01",
		X"C9",X"22",X"D6",X"20",X"EB",X"22",X"D4",X"20",X"C3",X"A3",X"02",X"CD",X"76",X"01",X"CD",X"83",
		X"01",X"CD",X"23",X"03",X"CD",X"15",X"03",X"21",X"02",X"24",X"01",X"E0",X"01",X"3E",X"7F",X"C3",
		X"8D",X"08",X"01",X"20",X"03",X"C5",X"E5",X"1A",X"77",X"23",X"13",X"05",X"C2",X"D7",X"01",X"E1",
		X"01",X"20",X"00",X"09",X"C1",X"0D",X"C2",X"D5",X"01",X"C9",X"21",X"B0",X"04",X"11",X"D8",X"20",
		X"06",X"02",X"C3",X"8B",X"03",X"21",X"B2",X"04",X"C3",X"ED",X"01",X"21",X"E6",X"20",X"46",X"B0",
		X"D3",X"03",X"77",X"C9",X"21",X"E6",X"20",X"46",X"2F",X"A0",X"D3",X"03",X"77",X"C9",X"21",X"E5",
		X"20",X"46",X"B0",X"D3",X"05",X"77",X"C9",X"21",X"E5",X"20",X"46",X"2F",X"A0",X"D3",X"05",X"77",
		X"C9",X"21",X"C3",X"20",X"3A",X"D8",X"20",X"6F",X"2B",X"2B",X"22",X"C9",X"20",X"06",X"03",X"11",
		X"DC",X"20",X"AF",X"1A",X"BE",X"DA",X"41",X"02",X"96",X"C0",X"23",X"13",X"05",X"C2",X"33",X"02",
		X"C9",X"06",X"03",X"2A",X"C9",X"20",X"11",X"DC",X"20",X"7E",X"12",X"23",X"13",X"05",X"C2",X"49",
		X"02",X"21",X"1D",X"30",X"22",X"D6",X"20",X"2A",X"C9",X"20",X"22",X"D4",X"20",X"C3",X"A3",X"02",
		X"D5",X"1A",X"CD",X"2E",X"03",X"CD",X"45",X"03",X"D1",X"13",X"05",X"C2",X"60",X"02",X"C9",X"21",
		X"C2",X"20",X"11",X"C5",X"20",X"3A",X"D8",X"20",X"5F",X"CD",X"E1",X"02",X"13",X"23",X"06",X"03",
		X"CD",X"8B",X"03",X"21",X"C0",X"20",X"11",X"03",X"00",X"C3",X"64",X"03",X"3A",X"E4",X"20",X"A7",
		X"C8",X"CD",X"6F",X"02",X"21",X"D8",X"20",X"7E",X"3D",X"3D",X"2E",X"D4",X"77",X"2E",X"D9",X"7E",
		X"2E",X"D7",X"77",X"2A",X"D4",X"20",X"7E",X"23",X"22",X"D4",X"20",X"E6",X"0F",X"CD",X"D1",X"02",
		X"06",X"02",X"C5",X"2A",X"D4",X"20",X"7E",X"F5",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"CD",X"D1",
		X"02",X"F1",X"E6",X"0F",X"CD",X"D1",X"02",X"21",X"D4",X"20",X"34",X"C1",X"05",X"C2",X"B2",X"02",
		X"C9",X"C6",X"20",X"CD",X"2E",X"03",X"2A",X"D6",X"20",X"CD",X"45",X"03",X"21",X"D7",X"20",X"34",
		X"C9",X"06",X"03",X"AF",X"1A",X"8E",X"27",X"77",X"2B",X"1B",X"05",X"C2",X"E4",X"02",X"C9",X"1A",
		X"77",X"13",X"23",X"1A",X"77",X"13",X"23",X"23",X"23",X"7E",X"FE",X"FF",X"C2",X"EF",X"02",X"C9",
		X"06",X"06",X"C5",X"7D",X"12",X"13",X"7C",X"12",X"01",X"00",X"06",X"09",X"13",X"13",X"13",X"C1",
		X"05",X"C2",X"02",X"03",X"C9",X"3A",X"E7",X"20",X"C6",X"20",X"CD",X"2E",X"03",X"21",X"01",X"3E",
		X"C3",X"45",X"03",X"21",X"01",X"37",X"11",X"B4",X"04",X"06",X"06",X"C3",X"60",X"02",X"11",X"94",
		X"03",X"A7",X"C8",X"E5",X"21",X"00",X"00",X"C5",X"01",X"05",X"00",X"09",X"3D",X"C2",X"38",X"03",
		X"19",X"EB",X"C1",X"E1",X"C9",X"C5",X"06",X"05",X"D3",X"06",X"C5",X"1A",X"07",X"77",X"13",X"01",
		X"20",X"00",X"09",X"C1",X"05",X"C2",X"48",X"03",X"AF",X"77",X"01",X"20",X"00",X"09",X"77",X"09",
		X"77",X"09",X"C1",X"C9",X"AF",X"77",X"23",X"1B",X"BA",X"C2",X"65",X"03",X"BB",X"C2",X"65",X"03",
		X"C9",X"7D",X"E6",X"07",X"D3",X"02",X"C5",X"06",X"03",X"7C",X"1F",X"67",X"7D",X"1F",X"6F",X"05",
		X"C2",X"79",X"03",X"7C",X"E6",X"3F",X"F6",X"20",X"67",X"C1",X"C9",X"7E",X"12",X"23",X"13",X"05",
		X"C2",X"8B",X"03",X"C9",X"1F",X"24",X"44",X"24",X"1F",X"7F",X"49",X"49",X"49",X"36",X"3E",X"41",
		X"41",X"41",X"22",X"7F",X"41",X"41",X"41",X"3E",X"7F",X"49",X"49",X"49",X"41",X"7F",X"48",X"48",
		X"48",X"40",X"3E",X"41",X"41",X"45",X"47",X"7F",X"08",X"08",X"08",X"7F",X"00",X"41",X"7F",X"41",
		X"00",X"02",X"01",X"01",X"01",X"7E",X"7F",X"08",X"14",X"22",X"41",X"7F",X"01",X"01",X"01",X"01",
		X"7F",X"20",X"18",X"20",X"7F",X"7F",X"10",X"08",X"04",X"7F",X"3E",X"41",X"41",X"41",X"3E",X"7F",
		X"48",X"48",X"48",X"30",X"3E",X"41",X"45",X"42",X"3D",X"7F",X"48",X"4C",X"4A",X"31",X"32",X"49",
		X"49",X"49",X"26",X"40",X"40",X"7F",X"40",X"40",X"7E",X"01",X"01",X"01",X"7E",X"7C",X"02",X"01",
		X"02",X"7C",X"7F",X"02",X"0C",X"02",X"7F",X"63",X"14",X"08",X"14",X"63",X"60",X"10",X"0F",X"10",
		X"60",X"43",X"45",X"49",X"51",X"61",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"22",X"14",X"7F",X"14",X"22",X"08",X"14",X"22",X"41",X"00",X"00",
		X"41",X"22",X"14",X"08",X"3E",X"45",X"49",X"51",X"3E",X"00",X"21",X"7F",X"01",X"00",X"23",X"45",
		X"49",X"49",X"31",X"42",X"41",X"49",X"59",X"66",X"0C",X"14",X"24",X"7F",X"04",X"72",X"51",X"51",
		X"51",X"4E",X"1E",X"29",X"49",X"49",X"46",X"40",X"47",X"48",X"50",X"60",X"36",X"49",X"49",X"49",
		X"36",X"31",X"49",X"49",X"4A",X"3C",X"14",X"14",X"14",X"14",X"14",X"01",X"02",X"04",X"08",X"10",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"18",X"18",X"00",X"0F",
		X"14",X"12",X"07",X"1B",X"0E",X"0D",X"0B",X"18",X"1B",X"21",X"1B",X"0F",X"0B",X"00",X"18",X"04",
		X"11",X"12",X"1B",X"01",X"14",X"13",X"13",X"0E",X"0D",X"1B",X"21",X"1B",X"0E",X"11",X"1B",X"22",
		X"1B",X"0F",X"0B",X"00",X"18",X"04",X"11",X"12",X"1B",X"01",X"14",X"13",X"13",X"0E",X"0D",X"00",
		X"C5",X"26",X"C8",X"39",X"02",X"11",X"04",X"03",X"08",X"13",X"06",X"C0",X"21",X"00",X"46",X"11",
		X"00",X"20",X"C3",X"8B",X"03",X"06",X"50",X"11",X"00",X"21",X"21",X"00",X"47",X"C3",X"8B",X"03",
		X"06",X"50",X"11",X"00",X"22",X"C3",X"CA",X"04",X"21",X"00",X"20",X"35",X"23",X"34",X"CD",X"EC",
		X"13",X"DB",X"01",X"0F",X"DA",X"28",X"05",X"21",X"E8",X"20",X"7E",X"A7",X"CA",X"03",X"05",X"2B",
		X"7E",X"FE",X"09",X"D2",X"FF",X"04",X"C6",X"01",X"27",X"32",X"E7",X"20",X"CD",X"15",X"03",X"AF",
		X"32",X"E8",X"20",X"3A",X"DF",X"20",X"A7",X"C2",X"22",X"05",X"3A",X"E4",X"20",X"A7",X"C2",X"D3",
		X"08",X"3A",X"E7",X"20",X"A7",X"C2",X"2D",X"05",X"3A",X"E0",X"20",X"A7",X"C2",X"D3",X"08",X"CD",
		X"3D",X"17",X"F1",X"C1",X"D1",X"E1",X"FB",X"C9",X"3E",X"01",X"C3",X"00",X"05",X"3A",X"02",X"20",
		X"A7",X"C2",X"22",X"05",X"3E",X"01",X"32",X"02",X"20",X"31",X"00",X"24",X"FB",X"CD",X"B6",X"00",
		X"21",X"E0",X"20",X"36",X"00",X"2E",X"AA",X"36",X"00",X"CD",X"BB",X"01",X"21",X"13",X"30",X"11",
		X"7F",X"04",X"06",X"04",X"CD",X"60",X"02",X"3A",X"E7",X"20",X"3D",X"D3",X"06",X"21",X"11",X"27",
		X"06",X"16",X"C2",X"A7",X"07",X"11",X"83",X"04",X"CD",X"60",X"02",X"D3",X"06",X"DB",X"01",X"E6",
		X"04",X"CA",X"57",X"05",X"06",X"99",X"AF",X"32",X"DA",X"20",X"3A",X"E7",X"20",X"80",X"27",X"32",
		X"E7",X"20",X"CD",X"15",X"03",X"21",X"C3",X"20",X"11",X"06",X"00",X"CD",X"64",X"03",X"CD",X"BA",
		X"04",X"CD",X"C5",X"04",X"CD",X"D0",X"04",X"CD",X"BB",X"01",X"21",X"2F",X"20",X"34",X"2E",X"E4",
		X"34",X"CD",X"BC",X"00",X"21",X"01",X"01",X"22",X"E9",X"20",X"CD",X"18",X"1A",X"CD",X"0D",X"19",
		X"3E",X"20",X"CD",X"FB",X"01",X"CD",X"B6",X"00",X"CD",X"2A",X"1A",X"CD",X"0E",X"06",X"CD",X"BC",
		X"00",X"CD",X"78",X"1A",X"CD",X"18",X"12",X"D3",X"06",X"CD",X"6B",X"07",X"CD",X"A1",X"1A",X"21",
		X"35",X"20",X"AF",X"BE",X"C2",X"48",X"06",X"CD",X"E6",X"18",X"CD",X"FB",X"18",X"CD",X"F2",X"18",
		X"CD",X"04",X"19",X"CD",X"E9",X"05",X"C3",X"C4",X"05",X"2E",X"24",X"CD",X"52",X"1A",X"7E",X"FE",
		X"03",X"21",X"9B",X"20",X"D2",X"FA",X"05",X"36",X"00",X"C9",X"36",X"01",X"CD",X"07",X"13",X"7E",
		X"0F",X"0F",X"01",X"40",X"00",X"DA",X"FE",X"12",X"01",X"C0",X"FF",X"C3",X"FE",X"12",X"06",X"07",
		X"C5",X"CD",X"52",X"1A",X"21",X"1E",X"25",X"D2",X"1C",X"06",X"26",X"38",X"01",X"38",X"01",X"CD",
		X"24",X"14",X"3E",X"08",X"CD",X"D5",X"14",X"CD",X"52",X"1A",X"11",X"F3",X"43",X"21",X"1E",X"38",
		X"DA",X"38",X"06",X"11",X"E0",X"43",X"26",X"25",X"06",X"07",X"CD",X"60",X"02",X"3E",X"08",X"CD",
		X"D5",X"14",X"C1",X"05",X"C2",X"10",X"06",X"C9",X"CD",X"B6",X"00",X"E5",X"CD",X"4C",X"00",X"CD",
		X"0D",X"19",X"E1",X"CD",X"9A",X"18",X"3A",X"DA",X"20",X"A7",X"C2",X"91",X"06",X"CD",X"44",X"1A",
		X"35",X"CA",X"7A",X"07",X"CD",X"7A",X"06",X"CD",X"BA",X"04",X"CD",X"BB",X"01",X"21",X"2F",X"20",
		X"34",X"CD",X"FC",X"00",X"CD",X"BC",X"00",X"C3",X"B5",X"05",X"7E",X"3D",X"21",X"01",X"25",X"CA",
		X"88",X"06",X"24",X"24",X"3D",X"C2",X"82",X"06",X"01",X"10",X"01",X"CD",X"8C",X"08",X"C3",X"C1",
		X"00",X"CD",X"B6",X"00",X"3A",X"DB",X"20",X"0F",X"DA",X"C8",X"06",X"CD",X"44",X"1A",X"35",X"C2",
		X"F5",X"06",X"CD",X"5D",X"07",X"21",X"07",X"30",X"3E",X"21",X"CD",X"2E",X"03",X"CD",X"45",X"03",
		X"CD",X"21",X"02",X"CD",X"C1",X"00",X"21",X"DB",X"20",X"36",X"01",X"CD",X"44",X"1A",X"A7",X"C2",
		X"04",X"07",X"CD",X"1E",X"14",X"C3",X"7D",X"07",X"CD",X"44",X"1A",X"35",X"C2",X"46",X"07",X"CD",
		X"5D",X"07",X"21",X"07",X"30",X"3E",X"22",X"CD",X"2E",X"03",X"CD",X"45",X"03",X"CD",X"21",X"02",
		X"CD",X"C1",X"00",X"21",X"DB",X"20",X"36",X"00",X"CD",X"44",X"1A",X"A7",X"C2",X"38",X"07",X"CD",
		X"1E",X"14",X"C3",X"7D",X"07",X"CD",X"7A",X"06",X"21",X"DB",X"20",X"36",X"01",X"CD",X"44",X"1A",
		X"A7",X"CA",X"3E",X"07",X"CD",X"F5",X"01",X"CD",X"1E",X"14",X"CD",X"16",X"07",X"CD",X"EF",X"12",
		X"CD",X"B6",X"00",X"C3",X"67",X"06",X"3A",X"DB",X"20",X"0F",X"DA",X"33",X"07",X"AF",X"21",X"E5",
		X"20",X"77",X"F3",X"D3",X"05",X"06",X"0A",X"0E",X"00",X"0D",X"C2",X"29",X"07",X"05",X"C2",X"27",
		X"07",X"FB",X"C9",X"3E",X"20",X"C3",X"1E",X"07",X"CD",X"EA",X"01",X"C3",X"07",X"07",X"21",X"DB",
		X"20",X"36",X"00",X"C3",X"38",X"07",X"CD",X"7A",X"06",X"21",X"DB",X"20",X"36",X"00",X"CD",X"44",
		X"1A",X"A7",X"C2",X"38",X"07",X"21",X"DB",X"20",X"36",X"01",X"C3",X"04",X"07",X"21",X"07",X"28",
		X"11",X"D4",X"44",X"06",X"14",X"CD",X"60",X"02",X"C3",X"FC",X"00",X"CD",X"52",X"1A",X"2E",X"25",
		X"7E",X"FE",X"02",X"D8",X"21",X"54",X"20",X"36",X"01",X"C9",X"CD",X"21",X"02",X"21",X"00",X"00",
		X"22",X"DA",X"20",X"22",X"E4",X"20",X"22",X"E5",X"20",X"22",X"E9",X"20",X"21",X"DA",X"20",X"36",
		X"01",X"21",X"14",X"2D",X"11",X"DF",X"44",X"06",X"09",X"CD",X"60",X"02",X"3E",X"80",X"CD",X"D5",
		X"14",X"CD",X"EA",X"01",X"C3",X"2D",X"00",X"11",X"99",X"04",X"CD",X"60",X"02",X"DB",X"01",X"0F",
		X"0F",X"DA",X"BB",X"07",X"0F",X"DA",X"74",X"05",X"C3",X"57",X"05",X"3E",X"01",X"06",X"98",X"C3",
		X"77",X"05",X"21",X"05",X"20",X"AF",X"BE",X"C8",X"CD",X"77",X"08",X"22",X"07",X"20",X"2A",X"09",
		X"20",X"01",X"60",X"00",X"09",X"22",X"09",X"20",X"44",X"21",X"0B",X"20",X"AF",X"BE",X"C2",X"E7",
		X"07",X"78",X"FE",X"2B",X"D2",X"32",X"08",X"23",X"AF",X"BE",X"C2",X"F3",X"07",X"78",X"FE",X"31",
		X"D2",X"4D",X"08",X"23",X"AF",X"BE",X"C2",X"FF",X"07",X"78",X"FE",X"37",X"D2",X"5B",X"08",X"23");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
