library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"02",X"23",X"00",X"30",X"FF",X"02",X"21",X"12",X"33",X"00",X"FF",X"32",X"99",X"29",X"93",
		X"30",X"FF",X"38",X"AA",X"8A",X"A8",X"30",X"FF",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"D8",X"AD",
		X"8D",X"A8",X"D0",X"FF",X"77",X"24",X"44",X"27",X"70",X"FF",X"7E",X"44",X"45",X"47",X"E0",X"FF",
		X"02",X"35",X"56",X"32",X"00",X"FF",X"00",X"00",X"30",X"00",X"00",X"FF",X"00",X"03",X"13",X"00",
		X"00",X"FF",X"00",X"31",X"91",X"30",X"00",X"FF",X"03",X"19",X"A9",X"13",X"00",X"FF",X"33",X"19",
		X"A9",X"13",X"30",X"FF",X"03",X"21",X"91",X"23",X"00",X"FF",X"00",X"32",X"33",X"30",X"00",X"FF",
		X"00",X"06",X"06",X"00",X"00",X"FF",X"04",X"56",X"86",X"55",X"00",X"FF",X"00",X"02",X"23",X"00",
		X"30",X"FF",X"02",X"21",X"11",X"23",X"00",X"FF",X"32",X"99",X"29",X"92",X"30",X"FF",X"38",X"AA",
		X"8A",X"A8",X"30",X"FF",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",
		X"77",X"24",X"44",X"27",X"70",X"FF",X"7E",X"44",X"45",X"57",X"E0",X"FF",X"02",X"35",X"56",X"32",
		X"00",X"FF",X"00",X"02",X"92",X"00",X"00",X"FF",X"00",X"39",X"A9",X"30",X"00",X"FF",X"02",X"89",
		X"99",X"82",X"00",X"FF",X"02",X"89",X"99",X"82",X"00",X"FF",X"02",X"81",X"91",X"82",X"00",X"FF",
		X"30",X"28",X"08",X"30",X"30",X"FF",X"05",X"66",X"06",X"66",X"00",X"FF",X"00",X"02",X"23",X"00",
		X"30",X"FF",X"02",X"22",X"12",X"33",X"00",X"FF",X"32",X"99",X"29",X"93",X"30",X"FF",X"38",X"AA",
		X"8A",X"A8",X"30",X"FF",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",
		X"77",X"24",X"44",X"27",X"70",X"FF",X"7E",X"44",X"45",X"47",X"E0",X"FF",X"02",X"35",X"56",X"32",
		X"00",X"FF",X"00",X"02",X"12",X"00",X"00",X"FF",X"00",X"31",X"91",X"30",X"00",X"FF",X"83",X"1A",
		X"A9",X"13",X"80",X"FF",X"33",X"19",X"99",X"13",X"30",X"FF",X"03",X"51",X"11",X"53",X"00",X"FF",
		X"00",X"62",X"33",X"60",X"00",X"FF",X"00",X"80",X"00",X"80",X"00",X"FF",X"00",X"02",X"23",X"03",
		X"00",X"FF",X"02",X"22",X"12",X"23",X"00",X"FF",X"32",X"99",X"29",X"92",X"30",X"FF",X"38",X"AA",
		X"8A",X"A8",X"30",X"FF",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",
		X"77",X"24",X"44",X"27",X"70",X"FF",X"7E",X"44",X"85",X"47",X"E0",X"FF",X"02",X"35",X"56",X"32",
		X"00",X"FF",X"00",X"02",X"12",X"00",X"00",X"FF",X"00",X"3A",X"A9",X"30",X"00",X"FF",X"02",X"89",
		X"99",X"82",X"00",X"FF",X"03",X"89",X"99",X"83",X"00",X"FF",X"08",X"35",X"25",X"28",X"00",X"FF",
		X"00",X"84",X"34",X"80",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"30",X"32",X"23",X"30",
		X"00",X"FF",X"03",X"29",X"22",X"33",X"00",X"FF",X"33",X"22",X"23",X"1A",X"30",X"FF",X"33",X"32",
		X"88",X"AA",X"80",X"FF",X"33",X"38",X"88",X"AD",X"80",X"FF",X"33",X"33",X"88",X"AD",X"80",X"FF",
		X"33",X"37",X"73",X"34",X"00",X"FF",X"03",X"3E",X"73",X"36",X"40",X"FF",X"00",X"33",X"33",X"66",
		X"00",X"FF",X"00",X"00",X"30",X"00",X"00",X"FF",X"00",X"03",X"11",X"00",X"00",X"FF",X"00",X"83",
		X"1A",X"90",X"00",X"FF",X"88",X"23",X"19",X"90",X"00",X"FF",X"21",X"13",X"19",X"10",X"00",X"FF",
		X"03",X"31",X"11",X"00",X"00",X"FF",X"00",X"31",X"26",X"60",X"00",X"FF",X"00",X"06",X"00",X"00",
		X"00",X"FF",X"00",X"66",X"66",X"00",X"00",X"FF",X"30",X"21",X"22",X"30",X"00",X"FF",X"02",X"1A",
		X"12",X"33",X"00",X"FF",X"32",X"11",X"12",X"1A",X"30",X"FF",X"33",X"22",X"23",X"AA",X"80",X"FF",
		X"33",X"33",X"88",X"AD",X"80",X"FF",X"33",X"38",X"88",X"AD",X"80",X"FF",X"33",X"33",X"88",X"AD",
		X"80",X"FF",X"03",X"37",X"73",X"34",X"00",X"FF",X"00",X"3E",X"73",X"66",X"40",X"FF",X"00",X"00",
		X"30",X"00",X"00",X"FF",X"00",X"03",X"12",X"00",X"00",X"FF",X"08",X"33",X"19",X"10",X"00",X"FF",
		X"08",X"23",X"9A",X"90",X"00",X"FF",X"02",X"92",X"19",X"10",X"00",X"FF",X"00",X"31",X"11",X"00",
		X"00",X"FF",X"05",X"55",X"26",X"00",X"00",X"FF",X"00",X"00",X"05",X"00",X"00",X"FF",X"00",X"00",
		X"66",X"65",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"30",X"32",X"22",X"30",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"22",X"92",X"33",
		X"00",X"FF",X"00",X"00",X"02",X"08",X"33",X"22",X"23",X"1A",X"30",X"FF",X"00",X"00",X"32",X"88",
		X"33",X"32",X"88",X"AA",X"80",X"FF",X"00",X"00",X"21",X"28",X"33",X"38",X"88",X"AD",X"80",X"FF",
		X"00",X"03",X"21",X"28",X"33",X"33",X"88",X"AD",X"80",X"FF",X"30",X"88",X"32",X"12",X"33",X"37",
		X"73",X"34",X"00",X"FF",X"08",X"81",X"13",X"23",X"03",X"3E",X"73",X"36",X"40",X"FF",X"00",X"01",
		X"91",X"33",X"33",X"33",X"33",X"66",X"00",X"FF",X"00",X"04",X"81",X"11",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"44",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"04",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"30",X"22",X"23",X"30",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"19",
		X"23",X"33",X"00",X"FF",X"00",X"00",X"00",X"00",X"32",X"22",X"23",X"1A",X"30",X"FF",X"00",X"00",
		X"00",X"00",X"33",X"22",X"88",X"AA",X"80",X"FF",X"03",X"00",X"00",X"00",X"33",X"38",X"88",X"AD",
		X"80",X"FF",X"33",X"30",X"33",X"00",X"33",X"33",X"88",X"AD",X"80",X"FF",X"03",X"33",X"21",X"30",
		X"33",X"37",X"73",X"34",X"00",X"FF",X"00",X"01",X"33",X"33",X"03",X"3E",X"73",X"36",X"40",X"FF",
		X"00",X"01",X"13",X"33",X"11",X"33",X"33",X"66",X"00",X"FF",X"00",X"05",X"11",X"33",X"30",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"44",X"60",X"22",X"30",X"00",X"00",X"00",X"00",X"FF",X"00",X"46",
		X"00",X"88",X"23",X"00",X"00",X"00",X"00",X"FF",X"00",X"46",X"00",X"08",X"02",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",
		X"00",X"22",X"30",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"32",X"22",X"23",X"80",X"00",X"FF",
		X"00",X"00",X"00",X"03",X"22",X"2A",X"A3",X"AA",X"00",X"FF",X"00",X"00",X"00",X"03",X"28",X"8A",
		X"C8",X"CA",X"00",X"FF",X"02",X"00",X"00",X"03",X"88",X"8C",X"D8",X"DC",X"00",X"FF",X"33",X"20",
		X"00",X"03",X"38",X"8C",X"D8",X"DC",X"00",X"FF",X"03",X"33",X"32",X"22",X"17",X"74",X"4B",X"47",
		X"00",X"FF",X"00",X"00",X"23",X"29",X"2E",X"E4",X"44",X"87",X"00",X"FF",X"00",X"00",X"13",X"32",
		X"21",X"22",X"55",X"60",X"00",X"FF",X"00",X"05",X"1A",X"33",X"20",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"04",X"B1",X"33",X"30",X"00",X"00",X"00",X"00",X"FF",X"00",X"04",X"60",X"DD",X"32",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"05",X"80",X"0D",X"03",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"23",X"00",X"30",
		X"00",X"FF",X"00",X"00",X"00",X"03",X"22",X"12",X"23",X"00",X"00",X"FF",X"00",X"00",X"00",X"32",
		X"AA",X"2A",X"A2",X"30",X"00",X"FF",X"00",X"00",X"00",X"38",X"AC",X"8C",X"A8",X"30",X"00",X"FF",
		X"00",X"00",X"00",X"88",X"CD",X"8D",X"C8",X"80",X"00",X"FF",X"00",X"00",X"00",X"D8",X"CD",X"8D",
		X"C8",X"D0",X"00",X"FF",X"00",X"00",X"00",X"77",X"24",X"44",X"27",X"70",X"00",X"FF",X"00",X"00",
		X"00",X"7E",X"44",X"85",X"47",X"E0",X"00",X"FF",X"08",X"00",X"00",X"03",X"D5",X"56",X"32",X"00",
		X"00",X"FF",X"00",X"80",X"02",X"23",X"30",X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"33",X"12",
		X"13",X"00",X"00",X"00",X"00",X"FF",X"08",X"88",X"33",X"33",X"29",X"30",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"83",X"38",X"29",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"81",X"10",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"08",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"44",X"44",X"86",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"33",X"30",X"30",X"00",X"00",X"FF",X"00",X"00",X"00",X"32",
		X"21",X"22",X"30",X"00",X"00",X"FF",X"00",X"00",X"03",X"2A",X"A2",X"AA",X"23",X"00",X"00",X"FF",
		X"00",X"00",X"03",X"8A",X"C8",X"CA",X"83",X"00",X"00",X"FF",X"00",X"00",X"08",X"8C",X"D8",X"DC",
		X"88",X"00",X"00",X"FF",X"00",X"00",X"0D",X"8C",X"D8",X"DC",X"8D",X"00",X"00",X"FF",X"00",X"00",
		X"07",X"72",X"44",X"42",X"77",X"00",X"00",X"FF",X"00",X"00",X"07",X"E4",X"48",X"54",X"7E",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"33",X"55",X"63",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",
		X"D2",X"00",X"00",X"00",X"00",X"FF",X"00",X"03",X"32",X"11",X"21",X"30",X"00",X"00",X"00",X"FF",
		X"00",X"08",X"33",X"22",X"1A",X"90",X"00",X"00",X"00",X"FF",X"00",X"00",X"83",X"33",X"19",X"90",
		X"00",X"00",X"00",X"FF",X"00",X"20",X"08",X"32",X"19",X"10",X"60",X"00",X"00",X"FF",X"00",X"08",
		X"88",X"C1",X"41",X"16",X"00",X"00",X"00",X"FF",X"00",X"33",X"38",X"22",X"42",X"60",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"30",X"03",X"00",X"00",X"FF",X"00",X"00",X"00",X"32",X"12",X"22",
		X"30",X"00",X"00",X"FF",X"00",X"00",X"03",X"AA",X"3A",X"A2",X"23",X"00",X"00",X"FF",X"00",X"00",
		X"08",X"AA",X"8A",X"AA",X"83",X"00",X"00",X"FF",X"00",X"00",X"08",X"AD",X"8D",X"AA",X"88",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"AD",X"8D",X"AA",X"8D",X"00",X"00",X"FF",X"00",X"00",X"07",X"74",
		X"44",X"42",X"77",X"08",X"00",X"FF",X"00",X"00",X"0E",X"44",X"44",X"54",X"7E",X"38",X"00",X"FF",
		X"00",X"00",X"00",X"24",X"85",X"83",X"23",X"88",X"66",X"FF",X"00",X"00",X"00",X"00",X"6C",X"19",
		X"AA",X"28",X"06",X"FF",X"00",X"00",X"00",X"80",X"22",X"31",X"9A",X"92",X"66",X"FF",X"00",X"00",
		X"08",X"32",X"23",X"31",X"99",X"91",X"D4",X"FF",X"00",X"00",X"00",X"22",X"33",X"33",X"21",X"11",
		X"D4",X"FF",X"00",X"00",X"08",X"33",X"30",X"D8",X"33",X"33",X"44",X"FF",X"00",X"00",X"00",X"03",
		X"00",X"8D",X"D3",X"80",X"04",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"23",X"00",X"30",X"FF",X"02",X"21",X"12",X"33",
		X"00",X"FF",X"32",X"22",X"22",X"23",X"30",X"FF",X"32",X"11",X"21",X"12",X"30",X"FF",X"88",X"AA",
		X"8A",X"A8",X"80",X"FF",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",X"77",X"A4",X"44",X"A7",X"70",X"FF",
		X"7E",X"44",X"85",X"47",X"E0",X"FF",X"80",X"05",X"56",X"00",X"80",X"FF",X"83",X"31",X"91",X"33",
		X"80",X"FF",X"33",X"1A",X"A9",X"13",X"30",X"FF",X"33",X"19",X"99",X"13",X"30",X"FF",X"03",X"51",
		X"11",X"53",X"00",X"FF",X"00",X"62",X"33",X"60",X"00",X"FF",X"00",X"80",X"00",X"80",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"23",X"00",
		X"30",X"FF",X"02",X"22",X"23",X"33",X"00",X"FF",X"32",X"21",X"12",X"33",X"30",X"FF",X"32",X"22",
		X"22",X"23",X"30",X"FF",X"32",X"11",X"21",X"12",X"30",X"FF",X"88",X"99",X"89",X"98",X"80",X"FF",
		X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",X"77",X"25",X"45",X"28",X"70",X"FF",X"E3",X"38",X"45",X"33",
		X"E0",X"FF",X"03",X"35",X"86",X"33",X"00",X"FF",X"33",X"8A",X"A9",X"83",X"30",X"FF",X"38",X"49",
		X"99",X"48",X"30",X"FF",X"08",X"51",X"11",X"58",X"00",X"FF",X"00",X"62",X"33",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"09",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"02",X"23",X"00",X"30",X"FF",X"02",X"22",X"23",X"33",X"00",X"FF",X"32",X"21",
		X"12",X"33",X"3A",X"FF",X"32",X"22",X"22",X"23",X"30",X"FF",X"32",X"22",X"22",X"22",X"30",X"FF",
		X"82",X"23",X"83",X"22",X"80",X"FF",X"D8",X"31",X"81",X"38",X"D0",X"FF",X"71",X"11",X"41",X"11",
		X"70",X"FF",X"12",X"28",X"42",X"22",X"10",X"FF",X"23",X"35",X"86",X"23",X"20",X"FF",X"24",X"3A",
		X"AA",X"44",X"30",X"FF",X"04",X"59",X"99",X"55",X"00",X"FF",X"00",X"62",X"11",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0A",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"23",X"00",X"30",X"FF",X"02",X"21",
		X"12",X"33",X"00",X"FF",X"32",X"22",X"22",X"23",X"30",X"FF",X"32",X"22",X"22",X"22",X"30",X"FF",
		X"82",X"23",X"83",X"22",X"80",X"FF",X"D1",X"11",X"11",X"38",X"D0",X"FF",X"11",X"22",X"12",X"11",
		X"70",X"FF",X"12",X"28",X"43",X"22",X"10",X"FF",X"05",X"55",X"86",X"23",X"20",X"FF",X"05",X"5A",
		X"AA",X"33",X"30",X"FF",X"06",X"69",X"99",X"54",X"00",X"FF",X"00",X"32",X"11",X"60",X"00",X"FF",
		X"33",X"33",X"88",X"83",X"38",X"FF",X"04",X"01",X"9A",X"91",X"13",X"43",X"9A",X"A9",X"38",X"FF",
		X"05",X"00",X"11",X"10",X"00",X"45",X"9E",X"E9",X"80",X"FF",X"00",X"00",X"00",X"00",X"05",X"46",
		X"58",X"88",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"FF",X"00",X"00",X"80",X"00",
		X"00",X"03",X"22",X"23",X"00",X"FF",X"00",X"88",X"80",X"00",X"00",X"32",X"22",X"22",X"30",X"FF",
		X"08",X"83",X"30",X"00",X"03",X"32",X"1A",X"22",X"33",X"FF",X"00",X"00",X"22",X"28",X"03",X"32",
		X"22",X"22",X"33",X"FF",X"40",X"03",X"21",X"92",X"03",X"33",X"26",X"23",X"33",X"FF",X"44",X"51",
		X"32",X"12",X"33",X"33",X"88",X"83",X"33",X"FF",X"46",X"61",X"33",X"33",X"33",X"33",X"88",X"83",
		X"38",X"FF",X"40",X"01",X"93",X"33",X"13",X"43",X"9A",X"A9",X"38",X"FF",X"60",X"00",X"9A",X"10",
		X"00",X"45",X"97",X"79",X"80",X"FF",X"00",X"00",X"00",X"00",X"05",X"46",X"58",X"88",X"00",X"FF",
		X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"1D",
		X"00",X"FF",X"D1",X"13",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",X"33",X"13",X"13",X"13",
		X"13",X"11",X"D0",X"FF",X"D1",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"13",
		X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"0D",
		X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",
		X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",
		X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",
		X"11",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"13",X"13",X"13",
		X"11",X"D0",X"FF",X"D1",X"13",X"11",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",
		X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",
		X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",
		X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",X"11",X"13",X"13",X"13",X"13",X"13",
		X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"11",X"13",
		X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",
		X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"D0",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",
		X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",X"31",X"13",X"33",X"13",X"33",
		X"11",X"D0",X"FF",X"D1",X"31",X"31",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"31",X"31",
		X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"33",X"33",X"13",X"13",X"13",X"13",X"11",X"D0",
		X"FF",X"D1",X"11",X"31",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"0D",X"11",X"11",X"11",X"11",
		X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",
		X"1D",X"00",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",X"13",X"11",
		X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"13",X"13",X"13",X"11",X"D0",
		X"FF",X"D1",X"11",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"33",
		X"13",X"33",X"11",X"D0",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"D0",X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",X"33",
		X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",
		X"FF",X"D1",X"13",X"33",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"13",X"13",X"13",
		X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"0D",
		X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"D0",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",X"13",X"33",X"13",X"33",X"13",
		X"33",X"11",X"D0",X"FF",X"D1",X"33",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",
		X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",
		X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",
		X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",X"11",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"13",X"13",X"13",X"13",X"13",X"11",
		X"D0",X"FF",X"D1",X"13",X"11",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",
		X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"11",X"D0",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",
		X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",
		X"33",X"13",X"33",X"11",X"D0",X"FF",X"D1",X"11",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"11",
		X"D0",X"FF",X"D1",X"13",X"33",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"11",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",
		X"33",X"13",X"33",X"11",X"D0",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",
		X"00",X"FF",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"00",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"1D",X"00",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"11",
		X"D0",X"FF",X"D1",X"13",X"11",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",
		X"33",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"11",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"11",X"D0",X"FF",X"D1",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"11",
		X"D0",X"FF",X"0D",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1D",X"00",X"FF",X"00",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"FF",X"55",X"25",X"25",X"25",X"50",X"00",X"00",X"00",X"FF",X"55",X"55",X"55",X"55",
		X"50",X"00",X"00",X"00",X"FF",X"55",X"25",X"25",X"25",X"50",X"00",X"00",X"00",X"FF",X"55",X"55",
		X"55",X"55",X"50",X"00",X"00",X"00",X"FF",X"55",X"25",X"25",X"25",X"50",X"00",X"00",X"00",X"FF",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"FF",X"05",X"25",X"25",X"25",X"00",X"00",X"00",
		X"00",X"FF",X"05",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"FF",X"05",X"25",X"25",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"52",
		X"52",X"52",X"54",X"00",X"00",X"00",X"00",X"FF",X"55",X"55",X"55",X"54",X"50",X"00",X"00",X"00",
		X"FF",X"05",X"25",X"25",X"25",X"45",X"00",X"00",X"00",X"FF",X"00",X"55",X"55",X"55",X"54",X"50",
		X"00",X"00",X"FF",X"00",X"05",X"25",X"25",X"25",X"45",X"00",X"00",X"FF",X"00",X"00",X"55",X"55",
		X"55",X"45",X"00",X"00",X"FF",X"00",X"00",X"05",X"52",X"52",X"55",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"05",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"01",X"37",X"85",X"00",X"FF",X"13",X"33",X"9A",X"50",X"FF",X"02",X"44",X"46",X"00",X"FF",X"00",
		X"24",X"60",X"00",X"FF",X"00",X"04",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"FF",
		X"44",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",
		X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"46",X"64",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"20",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"01",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"10",X"01",
		X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",
		X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"05",X"46",X"67",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"25",X"45",
		X"66",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"03",
		X"22",X"45",X"46",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"32",X"25",X"45",X"66",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"22",X"45",X"46",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"25",X"46",X"67",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"33",X"45",X"66",X"70",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"45",X"46",X"67",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"46",X"64",X"20",X"32",X"25",
		X"45",X"66",X"70",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"20",X"40",X"00",
		X"03",X"22",X"45",X"46",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"01",X"11",
		X"00",X"00",X"00",X"32",X"25",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"10",X"01",
		X"C1",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",
		X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"45",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"45",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"45",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"45",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"22",X"45",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"22",X"45",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"45",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"45",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"32",X"45",X"66",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"22",X"45",X"66",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"46",X"64",X"20",X"22",X"45",
		X"66",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"20",X"40",X"00",
		X"22",X"45",X"66",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"01",X"11",
		X"00",X"00",X"22",X"45",X"66",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"10",X"01",
		X"C1",X"00",X"00",X"00",X"22",X"45",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",
		X"01",X"11",X"00",X"00",X"00",X"00",X"22",X"00",X"FF",X"22",X"22",X"22",X"FF",X"27",X"77",X"77",
		X"FF",X"00",X"55",X"00",X"FF",X"00",X"55",X"00",X"FF",X"00",X"55",X"00",X"FF",X"00",X"55",X"00",
		X"FF",X"00",X"55",X"00",X"FF",X"00",X"55",X"00",X"FF",X"00",X"02",X"00",X"00",X"FF",X"00",X"27",
		X"20",X"00",X"FF",X"02",X"77",X"00",X"00",X"FF",X"27",X"75",X"50",X"00",X"FF",X"07",X"00",X"55",
		X"00",X"FF",X"00",X"00",X"05",X"50",X"FF",X"00",X"00",X"00",X"55",X"FF",X"00",X"00",X"00",X"05",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"22",X"00",X"00",X"00",X"FF",X"27",X"00",X"00",X"00",X"FF",
		X"27",X"55",X"55",X"55",X"FF",X"27",X"55",X"55",X"55",X"FF",X"27",X"00",X"00",X"00",X"FF",X"27",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"B1",X"B0",X"FF",X"00",X"BB",X"B0",
		X"FF",X"00",X"0A",X"00",X"FF",X"0A",X"0A",X"0A",X"FF",X"00",X"AA",X"A0",X"FF",X"02",X"22",X"22",
		X"FF",X"00",X"22",X"20",X"FF",X"00",X"22",X"20",X"FF",X"00",X"0B",X"00",X"00",X"FF",X"00",X"1B",
		X"00",X"00",X"FF",X"0B",X"BA",X"0A",X"00",X"FF",X"00",X"00",X"AA",X"20",X"FF",X"00",X"0A",X"A2",
		X"22",X"FF",X"00",X"00",X"22",X"22",X"FF",X"00",X"00",X"02",X"20",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"0A",X"02",X"00",X"FF",X"BB",X"00",X"A2",X"22",X"FF",
		X"1B",X"AA",X"A2",X"22",X"FF",X"BB",X"00",X"A2",X"22",X"FF",X"00",X"0A",X"02",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"08",X"CC",X"EE",X"00",X"FF",X"08",X"CD",
		X"EE",X"88",X"FF",X"08",X"CD",X"EE",X"0C",X"FF",X"08",X"CD",X"EE",X"0C",X"FF",X"08",X"CD",X"EE",
		X"0C",X"FF",X"08",X"CD",X"EE",X"C0",X"FF",X"08",X"CD",X"EE",X"00",X"FF",X"08",X"CD",X"EE",X"00",
		X"FF",X"00",X"08",X"CC",X"C0",X"00",X"FF",X"00",X"CC",X"80",X"0C",X"00",X"FF",X"0C",X"ED",X"C8",
		X"00",X"E0",X"FF",X"CE",X"EE",X"DD",X"80",X"E0",X"FF",X"0E",X"EE",X"ED",X"C8",X"00",X"FF",X"00",
		X"EE",X"ED",X"DC",X"80",X"FF",X"00",X"0E",X"EE",X"ED",X"00",X"FF",X"00",X"00",X"EE",X"E0",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"08",X"88",X"80",X"00",X"FF",X"0E",X"00",X"0C",X"00",X"FF",
		X"CC",X"CC",X"CC",X"C0",X"FF",X"DD",X"DD",X"DD",X"D0",X"FF",X"EE",X"EE",X"EE",X"E0",X"FF",X"EE",
		X"EE",X"EE",X"E0",X"FF",X"EE",X"EE",X"EE",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"7E",X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",X"82",X"88",X"00",X"0D",X"70",X"00",X"FF",X"00",
		X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"E0",X"00",X"FF",X"00",X"00",X"EE",X"ED",X"65",X"50",
		X"00",X"EE",X"EE",X"00",X"FF",X"00",X"88",X"88",X"EE",X"DD",X"50",X"0E",X"89",X"88",X"E0",X"FF",
		X"02",X"88",X"88",X"8E",X"EE",X"EE",X"E8",X"21",X"28",X"8E",X"FF",X"01",X"26",X"99",X"9C",X"CC",
		X"70",X"08",X"86",X"68",X"8E",X"FF",X"02",X"84",X"68",X"8C",X"97",X"77",X"08",X"86",X"48",X"80",
		X"FF",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"FF",X"70",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"0C",X"C0",X"FF",X"00",X"08",X"80",
		X"FF",X"02",X"CC",X"D0",X"FF",X"0C",X"0C",X"D0",X"FF",X"0C",X"0C",X"D0",X"FF",X"02",X"CC",X"D0",
		X"FF",X"00",X"0C",X"D0",X"FF",X"00",X"C1",X"C0",X"FF",X"0C",X"C2",X"CC",X"FF",X"CC",X"00",X"00",
		X"00",X"FF",X"D8",X"00",X"00",X"00",X"FF",X"0D",X"C0",X"00",X"00",X"FF",X"0C",X"DC",X"00",X"00",
		X"FF",X"02",X"0D",X"C0",X"00",X"FF",X"00",X"CC",X"DC",X"CC",X"FF",X"00",X"00",X"C1",X"C0",X"FF",
		X"00",X"00",X"CC",X"00",X"FF",X"00",X"00",X"C0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"FF",X"00",X"00",X"00",X"0C",X"C0",X"FF",X"C8",X"CC",X"CC",X"C1",
		X"C0",X"FF",X"C8",X"DD",X"DD",X"DC",X"C0",X"FF",X"00",X"C0",X"0C",X"00",X"C0",X"FF",X"00",X"2C",
		X"C2",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"C1",X"00",X"FF",X"0C",
		X"DD",X"DD",X"20",X"FF",X"CC",X"C0",X"0C",X"CC",X"FF",X"00",X"0C",X"C0",X"00",X"FF",X"00",X"C1",
		X"1C",X"00",X"FF",X"0C",X"13",X"31",X"C0",X"FF",X"C2",X"C1",X"1C",X"CC",X"FF",X"DD",X"DD",X"DD",
		X"DD",X"FF",X"00",X"01",X"2C",X"C0",X"00",X"FF",X"00",X"CD",X"CC",X"00",X"00",X"FF",X"0C",X"D0",
		X"C0",X"00",X"00",X"FF",X"CD",X"0C",X"CC",X"CC",X"00",X"FF",X"CC",X"CC",X"31",X"CC",X"D0",X"FF",
		X"CC",X"0C",X"31",X"CD",X"00",X"FF",X"C0",X"0C",X"CC",X"D0",X"00",X"FF",X"00",X"0C",X"2D",X"00",
		X"00",X"FF",X"00",X"00",X"D0",X"00",X"00",X"FF",X"00",X"C0",X"00",X"CD",X"FF",X"02",X"C0",X"0C",
		X"CD",X"FF",X"1D",X"C0",X"C1",X"CD",X"FF",X"CD",X"0C",X"13",X"1D",X"FF",X"CD",X"0C",X"13",X"1D",
		X"FF",X"CD",X"C0",X"C1",X"CD",X"FF",X"0C",X"C0",X"0C",X"2D",X"FF",X"00",X"C0",X"00",X"CD",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"10",X"FF",X"22",X"CC",X"22",X"01",X"FF",X"11",
		X"11",X"11",X"01",X"FF",X"01",X"11",X"10",X"10",X"FF",X"00",X"77",X"00",X"00",X"FF",X"11",X"11",
		X"11",X"10",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"00",X"FF",X"00",X"00",X"20",
		X"10",X"FF",X"00",X"0C",X"10",X"10",X"FF",X"00",X"C1",X"11",X"00",X"FF",X"02",X"11",X"10",X"01",
		X"FF",X"21",X"11",X"10",X"10",X"FF",X"01",X"11",X"71",X"00",X"FF",X"00",X"00",X"10",X"00",X"FF",
		X"00",X"01",X"00",X"00",X"FF",X"00",X"10",X"00",X"00",X"FF",X"11",X"10",X"00",X"FF",X"10",X"01",
		X"01",X"FF",X"02",X"10",X"01",X"FF",X"02",X"11",X"01",X"FF",X"0C",X"11",X"71",X"FF",X"0C",X"11",
		X"71",X"FF",X"02",X"11",X"01",X"FF",X"02",X"10",X"01",X"FF",X"ED",X"00",X"FF",X"00",X"00",X"EE",
		X"E0",X"00",X"FF",X"00",X"04",X"44",X"50",X"00",X"FF",X"00",X"43",X"23",X"45",X"00",X"FF",X"00",
		X"42",X"31",X"75",X"00",X"FF",X"00",X"53",X"33",X"45",X"00",X"FF",X"00",X"05",X"33",X"59",X"A0",
		X"FF",X"53",X"44",X"56",X"00",X"00",X"FF",X"42",X"23",X"43",X"50",X"00",X"FF",X"53",X"34",X"33",
		X"50",X"00",X"FF",X"06",X"54",X"45",X"00",X"00",X"FF",X"77",X"66",X"60",X"00",X"00",X"FF",X"00",
		X"0A",X"00",X"00",X"00",X"FF",X"00",X"99",X"A0",X"00",X"00",X"FF",X"00",X"04",X"44",X"50",X"00",
		X"FF",X"00",X"43",X"23",X"45",X"00",X"FF",X"00",X"42",X"31",X"75",X"00",X"FF",X"00",X"53",X"33",
		X"45",X"00",X"FF",X"00",X"05",X"33",X"59",X"A0",X"FF",X"65",X"44",X"56",X"00",X"00",X"FF",X"53",
		X"22",X"43",X"50",X"00",X"FF",X"53",X"34",X"33",X"50",X"00",X"FF",X"06",X"54",X"45",X"00",X"00",
		X"FF",X"00",X"66",X"60",X"00",X"00",X"FF",X"08",X"A7",X"00",X"00",X"00",X"FF",X"00",X"99",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",X"23",X"17",X"50",X"FF",X"00",
		X"04",X"22",X"34",X"50",X"FF",X"00",X"05",X"33",X"33",X"5A",X"FF",X"05",X"44",X"54",X"45",X"00",
		X"FF",X"53",X"22",X"34",X"50",X"00",X"FF",X"53",X"34",X"33",X"50",X"00",X"FF",X"06",X"54",X"45",
		X"50",X"00",X"FF",X"00",X"66",X"66",X"00",X"00",X"FF",X"09",X"9A",X"70",X"00",X"00",X"FF",X"00",
		X"07",X"77",X"00",X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",X"22",X"11",X"50",
		X"FF",X"00",X"04",X"22",X"17",X"50",X"FF",X"00",X"65",X"33",X"24",X"59",X"FF",X"32",X"26",X"54",
		X"44",X"A0",X"FF",X"53",X"22",X"56",X"60",X"00",X"FF",X"53",X"33",X"53",X"34",X"00",X"FF",X"05",
		X"55",X"43",X"35",X"00",X"FF",X"00",X"05",X"55",X"50",X"00",X"FF",X"00",X"0A",X"A0",X"00",X"00",
		X"FF",X"00",X"00",X"98",X"00",X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",X"22",
		X"11",X"50",X"FF",X"00",X"04",X"22",X"17",X"50",X"FF",X"00",X"05",X"33",X"24",X"59",X"FF",X"00",
		X"66",X"54",X"44",X"90",X"FF",X"00",X"32",X"56",X"60",X"00",X"FF",X"03",X"23",X"53",X"30",X"00",
		X"FF",X"02",X"55",X"43",X"30",X"00",X"FF",X"00",X"A5",X"55",X"50",X"00",X"FF",X"00",X"0A",X"00",
		X"00",X"00",X"FF",X"04",X"40",X"74",X"44",X"50",X"FF",X"03",X"37",X"42",X"11",X"45",X"FF",X"54",
		X"46",X"42",X"17",X"35",X"FF",X"45",X"55",X"43",X"33",X"37",X"FF",X"44",X"34",X"54",X"43",X"50",
		X"FF",X"A4",X"32",X"46",X"0A",X"00",X"FF",X"05",X"45",X"60",X"00",X"00",X"FF",X"00",X"A0",X"00",
		X"00",X"00",X"FF",X"0A",X"00",X"44",X"00",X"00",X"FF",X"00",X"45",X"33",X"00",X"00",X"FF",X"04",
		X"32",X"55",X"00",X"00",X"FF",X"A3",X"32",X"46",X"55",X"50",X"FF",X"64",X"43",X"64",X"33",X"46",
		X"FF",X"65",X"34",X"A9",X"37",X"15",X"FF",X"56",X"55",X"53",X"33",X"35",X"FF",X"35",X"60",X"64",
		X"73",X"46",X"FF",X"00",X"00",X"06",X"55",X"60",X"FF",X"00",X"0A",X"00",X"A0",X"FF",X"05",X"55",
		X"45",X"00",X"FF",X"55",X"53",X"53",X"50",X"FF",X"43",X"54",X"53",X"30",X"FF",X"32",X"43",X"32",
		X"30",X"FF",X"25",X"43",X"35",X"20",X"FF",X"06",X"65",X"55",X"60",X"FF",X"00",X"64",X"33",X"46",
		X"FF",X"00",X"51",X"31",X"15",X"FF",X"00",X"57",X"37",X"15",X"FF",X"00",X"64",X"33",X"46",X"FF",
		X"00",X"06",X"55",X"60",X"FF",X"00",X"04",X"43",X"50",X"00",X"FF",X"00",X"41",X"21",X"15",X"00",
		X"FF",X"00",X"47",X"37",X"14",X"00",X"FF",X"00",X"43",X"83",X"35",X"00",X"FF",X"04",X"62",X"A2",
		X"46",X"40",X"FF",X"33",X"45",X"55",X"56",X"32",X"FF",X"54",X"55",X"23",X"55",X"45",X"FF",X"05",
		X"63",X"22",X"36",X"50",X"FF",X"00",X"05",X"44",X"50",X"00",X"FF",X"00",X"00",X"80",X"90",X"00",
		X"FF",X"00",X"00",X"A0",X"A0",X"00",X"FF",X"00",X"44",X"35",X"00",X"FF",X"04",X"12",X"11",X"50",
		X"FF",X"04",X"73",X"71",X"40",X"FF",X"04",X"38",X"33",X"50",X"FF",X"06",X"2A",X"24",X"60",X"FF",
		X"54",X"55",X"55",X"65",X"FF",X"42",X"52",X"35",X"34",X"FF",X"52",X"42",X"24",X"25",X"FF",X"00",
		X"54",X"45",X"00",X"FF",X"00",X"0A",X"0A",X"00",X"FF",X"00",X"03",X"34",X"40",X"FF",X"00",X"33",
		X"23",X"44",X"FF",X"00",X"33",X"71",X"37",X"FF",X"00",X"33",X"33",X"94",X"FF",X"00",X"42",X"39",
		X"9A",X"FF",X"00",X"65",X"34",X"A0",X"FF",X"06",X"23",X"54",X"56",X"FF",X"03",X"33",X"52",X"45",
		X"FF",X"05",X"45",X"44",X"63",X"FF",X"00",X"65",X"66",X"00",X"FF",X"00",X"99",X"0A",X"00",X"FF",
		X"00",X"00",X"88",X"A0",X"FF",X"00",X"33",X"34",X"00",X"FF",X"03",X"32",X"23",X"40",X"FF",X"03",
		X"73",X"37",X"40",X"FF",X"03",X"13",X"31",X"40",X"FF",X"04",X"39",X"93",X"40",X"FF",X"00",X"4A",
		X"A4",X"00",X"FF",X"06",X"55",X"55",X"60",X"FF",X"05",X"33",X"34",X"50",X"FF",X"35",X"43",X"35",
		X"53",X"FF",X"00",X"55",X"55",X"00",X"FF",X"00",X"AA",X"0A",X"00",X"FF",X"0A",X"9A",X"AA",X"A0",
		X"FF",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"02",X"EE",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"23",X"EE",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"3E",
		X"EE",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"07",X"CC",X"CC",
		X"CB",X"00",X"00",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",X"73",X"3E",X"EE",X"E3",
		X"00",X"7C",X"54",X"DD",X"DD",X"45",X"00",X"00",X"02",X"00",X"FF",X"CC",X"CC",X"CC",X"CA",X"67",
		X"55",X"CC",X"44",X"44",X"5C",X"77",X"00",X"03",X"00",X"FF",X"CC",X"CC",X"CC",X"C6",X"45",X"63",
		X"3C",X"CC",X"BB",X"C5",X"66",X"70",X"06",X"00",X"FF",X"73",X"EE",X"E7",X"65",X"63",X"32",X"22",
		X"2E",X"EE",X"EE",X"E3",X"67",X"04",X"00",X"FF",X"73",X"EE",X"E7",X"66",X"33",X"22",X"22",X"22",
		X"22",X"22",X"2E",X"36",X"05",X"00",X"FF",X"07",X"EE",X"33",X"63",X"22",X"11",X"12",X"22",X"22",
		X"11",X"22",X"E3",X"60",X"00",X"FF",X"07",X"3E",X"33",X"EE",X"22",X"55",X"66",X"66",X"33",X"E1",
		X"12",X"23",X"49",X"E0",X"FF",X"00",X"76",X"33",X"EE",X"E5",X"6E",X"33",X"33",X"3E",X"A1",X"12",
		X"23",X"48",X"80",X"FF",X"00",X"66",X"73",X"33",X"56",X"E3",X"33",X"33",X"EA",X"71",X"12",X"E3",
		X"50",X"00",X"FF",X"00",X"05",X"67",X"64",X"43",X"63",X"33",X"3E",X"A7",X"22",X"22",X"E6",X"5D",
		X"00",X"FF",X"00",X"00",X"56",X"5D",X"43",X"66",X"3E",X"AA",X"73",X"22",X"EE",X"65",X"04",X"00",
		X"FF",X"00",X"00",X"05",X"44",X"D4",X"77",X"77",X"77",X"63",X"3E",X"E6",X"50",X"08",X"00",X"FF",
		X"00",X"00",X"00",X"D4",X"44",X"45",X"57",X"75",X"66",X"66",X"75",X"00",X"08",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"D4",X"44",X"45",X"55",X"54",X"44",X"00",X"00",X"09",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"FF",X"0D",X"00",X"0D",
		X"00",X"FF",X"DC",X"00",X"0C",X"D0",X"FF",X"0D",X"C4",X"CD",X"00",X"FF",X"00",X"08",X"00",X"00",
		X"FF",X"00",X"C4",X"C0",X"00",X"FF",X"0C",X"40",X"4C",X"00",X"FF",X"D4",X"00",X"04",X"D0",X"FF",
		X"D4",X"00",X"04",X"D0",X"FF",X"0C",X"00",X"0C",X"00",X"FF",X"00",X"DD",X"C0",X"00",X"00",X"FF",
		X"00",X"0C",X"D0",X"00",X"00",X"FF",X"D0",X"00",X"D0",X"00",X"00",X"FF",X"DC",X"08",X"CC",X"CD",
		X"00",X"FF",X"CD",X"DC",X"04",X"44",X"D0",X"FF",X"00",X"0C",X"40",X"04",X"C0",X"FF",X"00",X"0C",
		X"40",X"00",X"C0",X"FF",X"00",X"0D",X"44",X"00",X"00",X"FF",X"00",X"00",X"DC",X"C0",X"00",X"FF",
		X"0D",X"00",X"00",X"DD",X"00",X"FF",X"DC",X"D0",X"0C",X"44",X"C0",X"FF",X"00",X"C0",X"C4",X"00",
		X"00",X"FF",X"00",X"48",X"40",X"00",X"00",X"FF",X"00",X"C0",X"C4",X"00",X"00",X"FF",X"DC",X"D0",
		X"0C",X"44",X"C0",X"FF",X"0D",X"00",X"00",X"DD",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"09",X"00",X"00",X"FF",X"08",X"89",X"98",X"80",X"FF",X"81",X"38",X"88",X"88",X"FF",X"82",
		X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"88",X"FF",X"08",X"88",X"88",X"80",X"FF",X"08",X"88",
		X"8A",X"80",X"FF",X"00",X"8A",X"AA",X"00",X"FF",X"00",X"88",X"80",X"00",X"FF",X"08",X"88",X"88",
		X"80",X"FF",X"08",X"88",X"88",X"AA",X"FF",X"09",X"88",X"88",X"8A",X"FF",X"99",X"88",X"88",X"8A",
		X"FF",X"08",X"38",X"88",X"88",X"FF",X"08",X"12",X"88",X"80",X"FF",X"00",X"88",X"80",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"90",X"08",X"88",X"00",X"FF",X"09",X"98",X"88",X"80",X"FF",X"83",
		X"88",X"88",X"80",X"FF",X"81",X"38",X"88",X"88",X"FF",X"88",X"88",X"88",X"AA",X"FF",X"08",X"88",
		X"8A",X"AA",X"FF",X"00",X"08",X"AA",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",X"01",
		X"11",X"00",X"00",X"FF",X"10",X"08",X"88",X"0E",X"E0",X"FF",X"01",X"01",X"11",X"E0",X"E0",X"FF",
		X"01",X"01",X"11",X"00",X"E0",X"FF",X"01",X"11",X"11",X"E0",X"E0",X"FF",X"00",X"01",X"11",X"0E",
		X"00",X"FF",X"00",X"01",X"11",X"00",X"00",X"FF",X"00",X"00",X"0E",X"E0",X"FF",X"01",X"11",X"0E",
		X"0E",X"FF",X"01",X"18",X"1E",X"0E",X"FF",X"01",X"81",X"11",X"0E",X"FF",X"00",X"11",X"11",X"10",
		X"FF",X"10",X"01",X"11",X"11",X"FF",X"01",X"11",X"11",X"10",X"FF",X"00",X"10",X"01",X"00",X"FF",
		X"00",X"EE",X"EE",X"00",X"FF",X"00",X"E0",X"00",X"E0",X"FF",X"00",X"0E",X"0E",X"00",X"FF",X"01",
		X"81",X"11",X"11",X"FF",X"11",X"81",X"11",X"11",X"FF",X"01",X"81",X"11",X"11",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"00",X"01",X"11",X"00",X"FF",X"00",X"0B",X"00",X"FF",X"00",X"05",X"00",X"FF",
		X"00",X"05",X"00",X"FF",X"00",X"55",X"50",X"FF",X"00",X"11",X"50",X"FF",X"00",X"11",X"50",X"FF",
		X"00",X"11",X"50",X"FF",X"00",X"55",X"50",X"FF",X"00",X"55",X"50",X"FF",X"00",X"00",X"00",X"FF",
		X"B0",X"00",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"FF",X"00",X"55",X"00",X"00",X"F0",X"00",
		X"55",X"50",X"00",X"FF",X"00",X"51",X"55",X"00",X"FF",X"00",X"01",X"15",X"50",X"FF",X"00",X"00",
		X"15",X"50",X"FF",X"00",X"00",X"05",X"50",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"05",X"55",X"55",X"50",X"FF",
		X"B5",X"55",X"11",X"15",X"50",X"FF",X"00",X"05",X"11",X"15",X"50",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"09",X"90",X"90",
		X"00",X"FF",X"00",X"99",X"99",X"00",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",X"EE",X"E9",X"EE",X"E0",
		X"FF",X"99",X"99",X"99",X"90",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",
		X"00",X"90",X"E0",X"00",X"FF",X"90",X"9E",X"EE",X"00",X"FF",X"99",X"9E",X"E9",X"E0",X"FF",X"0E",
		X"E9",X"9E",X"EE",X"FF",X"EE",X"E9",X"9E",X"E0",X"FF",X"0E",X"9E",X"E9",X"00",X"FF",X"00",X"EE",
		X"E0",X"00",X"FF",X"00",X"0E",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"9E",
		X"E0",X"FF",X"09",X"EE",X"9E",X"E0",X"FF",X"99",X"EE",X"9E",X"E0",X"FF",X"09",X"99",X"99",X"90",
		X"FF",X"99",X"EE",X"9E",X"E0",X"FF",X"90",X"EE",X"9E",X"E0",X"FF",X"00",X"EE",X"9E",X"E0",X"FF",
		X"0B",X"DE",X"DD",X"DB",X"FF",X"00",X"BE",X"DD",X"B0",X"FF",X"00",X"0B",X"DB",X"00",X"FF",X"00",
		X"00",X"B0",X"00",X"FF",X"00",X"00",X"B0",X"00",X"FF",X"00",X"00",X"B0",X"00",X"FF",X"00",X"00",
		X"B0",X"00",X"FF",X"00",X"00",X"B0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",
		X"EE",X"01",X"10",X"FF",X"AA",X"AA",X"AA",X"10",X"01",X"FF",X"AA",X"AA",X"AA",X"00",X"01",X"FF",
		X"AA",X"AA",X"AA",X"00",X"01",X"FF",X"AA",X"AA",X"AA",X"11",X"10",X"FF",X"AA",X"AA",X"AA",X"00",
		X"00",X"FF",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"FF",X"00",X"00",
		X"E0",X"10",X"01",X"FF",X"00",X"0E",X"AA",X"10",X"01",X"FF",X"00",X"EA",X"AA",X"A0",X"10",X"FF",
		X"0E",X"AA",X"AA",X"AA",X"10",X"FF",X"EA",X"AA",X"AA",X"AA",X"A0",X"FF",X"0A",X"AA",X"AA",X"AA",
		X"00",X"FF",X"00",X"AA",X"AA",X"A0",X"00",X"FF",X"00",X"0A",X"AA",X"00",X"00",X"FF",X"00",X"00",
		X"A0",X"00",X"00",X"FF",X"00",X"11",X"10",X"00",X"FF",X"01",X"00",X"01",X"00",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"00",X"10",X"01",X"00",X"FF",X"0E",X"AA",X"AA",X"AA",X"FF",X"0E",X"AA",X"AA",
		X"AA",X"FF",X"0E",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"FF",X"00",X"08",
		X"00",X"FF",X"00",X"88",X"80",X"FF",X"08",X"88",X"88",X"FF",X"0E",X"EE",X"EB",X"FF",X"0E",X"EE",
		X"EB",X"FF",X"0E",X"EE",X"EB",X"FF",X"0E",X"EE",X"EB",X"FF",X"0E",X"EE",X"EB",X"FF",X"0E",X"EE",
		X"EB",X"FF",X"0C",X"BB",X"BC",X"FF",X"80",X"00",X"00",X"00",X"00",X"FF",X"08",X"88",X"80",X"00",
		X"00",X"FF",X"08",X"8E",X"EB",X"00",X"00",X"FF",X"08",X"EE",X"EB",X"B0",X"00",X"FF",X"08",X"EE",
		X"EE",X"BB",X"00",X"FF",X"00",X"EE",X"EE",X"EB",X"C0",X"FF",X"00",X"0E",X"EE",X"EB",X"00",X"FF",
		X"00",X"00",X"EE",X"B0",X"00",X"FF",X"00",X"00",X"0C",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"8B",X"BB",X"BB",X"BC",X"FF",
		X"00",X"08",X"8E",X"EE",X"EE",X"EB",X"FF",X"08",X"88",X"8E",X"EE",X"EE",X"EB",X"FF",X"00",X"08",
		X"8E",X"EE",X"EE",X"EB",X"FF",X"00",X"00",X"8E",X"EE",X"EE",X"EC",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",X"0D",X"DD",X"00",
		X"10",X"FF",X"BB",X"BB",X"BB",X"B1",X"01",X"FF",X"0B",X"BB",X"BB",X"B0",X"01",X"FF",X"00",X"BB",
		X"BB",X"B1",X"11",X"FF",X"00",X"BB",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"00",X"10",X"FF",X"00",
		X"00",X"01",X"01",X"FF",X"00",X"00",X"B1",X"01",X"FF",X"00",X"1D",X"BB",X"01",X"FF",X"00",X"DB",
		X"BB",X"B0",X"FF",X"00",X"BB",X"BB",X"BB",X"FF",X"0B",X"BB",X"BB",X"B0",X"FF",X"BB",X"BB",X"BB",
		X"00",X"FF",X"00",X"00",X"B0",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"11",X"10",X"FF",
		X"01",X"00",X"10",X"FF",X"00",X"10",X"10",X"FF",X"00",X"BB",X"BB",X"FF",X"0D",X"BB",X"BB",X"FF",
		X"1D",X"BB",X"BB",X"FF",X"0D",X"BB",X"BB",X"FF",X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"00",X"FF",
		X"00",X"B0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"00",X"00",X"FF",
		X"00",X"99",X"99",X"99",X"00",X"FF",X"18",X"88",X"88",X"88",X"81",X"FF",X"19",X"99",X"99",X"99",
		X"11",X"FF",X"09",X"99",X"99",X"99",X"90",X"FF",X"09",X"99",X"99",X"99",X"90",X"FF",X"00",X"99",
		X"99",X"99",X"00",X"FF",X"00",X"00",X"98",X"10",X"FF",X"00",X"19",X"81",X"10",X"FF",X"01",X"98",
		X"99",X"90",X"FF",X"09",X"89",X"99",X"90",X"FF",X"98",X"99",X"99",X"90",X"FF",X"89",X"99",X"99",
		X"00",X"FF",X"19",X"99",X"90",X"00",X"FF",X"00",X"99",X"00",X"00",X"FF",X"00",X"11",X"00",X"00",
		X"FF",X"00",X"81",X"99",X"00",X"FF",X"09",X"89",X"99",X"90",X"FF",X"09",X"89",X"99",X"90",X"FF",
		X"19",X"89",X"99",X"90",X"FF",X"19",X"89",X"99",X"90",X"FF",X"09",X"89",X"99",X"90",X"FF",X"09",
		X"89",X"99",X"90",X"FF",X"00",X"89",X"99",X"00",X"FF",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"98",X"89",X"90",X"09",X"88",X"88",X"90",X"00",
		X"00",X"0B",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"09",X"88",X"88",
		X"8B",X"98",X"88",X"88",X"9B",X"00",X"00",X"B8",X"88",X"B0",X"BB",X"BB",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"98",X"88",X"89",X"9B",X"B8",X"88",X"88",X"9B",X"BB",X"B0",X"B8",X"88",X"8B",
		X"88",X"88",X"BB",X"00",X"00",X"FF",X"00",X"00",X"99",X"88",X"88",X"98",X"88",X"8B",X"98",X"89",
		X"88",X"B8",X"8B",X"88",X"88",X"88",X"88",X"88",X"88",X"B0",X"00",X"FF",X"00",X"09",X"88",X"88",
		X"89",X"88",X"88",X"88",X"B9",X"88",X"88",X"B8",X"88",X"88",X"88",X"88",X"88",X"99",X"98",X"8B",
		X"00",X"FF",X"00",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"B9",X"98",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"89",X"9B",X"B0",X"FF",X"0B",X"88",X"8B",X"88",X"88",X"88",X"88",X"88",
		X"B8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"9B",X"FF",X"0B",X"88",
		X"8B",X"88",X"88",X"88",X"88",X"88",X"B8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"9B",X"FF",X"0B",X"88",X"8B",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"9B",X"FF",X"00",X"B8",X"89",X"BB",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"9B",X"FF",
		X"00",X"B9",X"9B",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"89",X"88",X"88",X"89",X"B0",X"FF",X"00",X"B9",X"9B",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"98",X"88",X"98",X"88",X"89",X"98",X"89",X"9B",X"00",X"FF",X"00",X"0B",X"B9",X"98",
		X"9B",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"89",X"88",X"88",X"99",X"99",X"BB",X"B0",
		X"00",X"FF",X"00",X"00",X"B9",X"99",X"9B",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",
		X"98",X"89",X"9B",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"BB",X"9B",X"88",X"88",X"89",
		X"88",X"88",X"88",X"88",X"89",X"99",X"99",X"BB",X"B0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"B9",X"B8",X"88",X"88",X"98",X"88",X"88",X"89",X"9B",X"BB",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",X"98",X"98",X"89",X"98",X"88",X"88",X"99",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"99",X"99",X"9B",X"88",X"8B",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"B0",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"B0",X"00",X"00",
		X"00",X"B9",X"9B",X"00",X"00",X"00",X"FF",X"00",X"00",X"09",X"99",X"B0",X"99",X"89",X"9B",X"00",
		X"0B",X"BB",X"B8",X"88",X"BB",X"00",X"00",X"FF",X"00",X"00",X"98",X"88",X"9B",X"88",X"88",X"9B",
		X"B0",X"B8",X"88",X"88",X"99",X"99",X"B0",X"00",X"FF",X"00",X"09",X"88",X"88",X"89",X"B8",X"9B",
		X"B8",X"9B",X"88",X"88",X"88",X"88",X"88",X"9B",X"00",X"FF",X"00",X"98",X"88",X"88",X"88",X"B9",
		X"88",X"88",X"8B",X"88",X"88",X"98",X"88",X"88",X"8B",X"00",X"FF",X"00",X"98",X"88",X"88",X"88",
		X"99",X"98",X"88",X"9B",X"88",X"88",X"88",X"89",X"88",X"99",X"B0",X"FF",X"00",X"98",X"8B",X"98",
		X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"88",X"90",X"FF",X"00",X"98",X"89",
		X"98",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"99",X"FF",X"09",X"89",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"9B",X"FF",X"98",
		X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"89",X"9B",X"FF",
		X"0B",X"B9",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"B0",
		X"FF",X"00",X"00",X"B9",X"98",X"98",X"89",X"88",X"88",X"88",X"88",X"88",X"98",X"89",X"99",X"9B",
		X"00",X"FF",X"00",X"00",X"B9",X"99",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"BB",
		X"00",X"00",X"FF",X"00",X"00",X"0B",X"98",X"89",X"8B",X"88",X"88",X"88",X"88",X"89",X"B9",X"9B",
		X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"99",X"9B",X"98",X"88",X"88",X"88",X"99",X"BB",
		X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0B",X"99",X"99",X"B9",X"88",X"88",X"99",X"BB",
		X"BB",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"BB",X"B9",X"9B",X"99",X"99",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"7E",
		X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",X"82",X"88",X"00",X"0D",X"70",X"00",X"FF",X"00",X"00",
		X"00",X"08",X"88",X"88",X"80",X"00",X"E0",X"00",X"FF",X"00",X"00",X"EE",X"7D",X"69",X"50",X"00",
		X"EE",X"EE",X"00",X"FF",X"00",X"21",X"28",X"EE",X"DD",X"50",X"0E",X"88",X"21",X"E0",X"FF",X"08",
		X"82",X"88",X"8E",X"EE",X"EE",X"E8",X"88",X"81",X"2E",X"FF",X"08",X"86",X"6B",X"B7",X"77",X"C0",
		X"08",X"86",X"68",X"8E",X"FF",X"08",X"84",X"68",X"8C",X"DD",X"D0",X"08",X"86",X"48",X"80",X"FF",
		X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",
		X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",
		X"22",X"34",X"50",X"FF",X"00",X"04",X"27",X"77",X"70",X"FF",X"00",X"05",X"33",X"37",X"70",X"FF",
		X"53",X"44",X"53",X"35",X"9A",X"FF",X"42",X"23",X"43",X"50",X"00",X"FF",X"53",X"34",X"33",X"60",
		X"00",X"FF",X"06",X"54",X"45",X"00",X"00",X"FF",X"77",X"66",X"60",X"00",X"00",X"FF",X"00",X"0A",
		X"00",X"00",X"00",X"FF",X"00",X"99",X"A0",X"00",X"00",X"FF",X"00",X"04",X"44",X"50",X"00",X"FF",
		X"00",X"43",X"23",X"45",X"00",X"FF",X"00",X"42",X"77",X"77",X"00",X"FF",X"00",X"53",X"33",X"77",
		X"00",X"FF",X"00",X"05",X"33",X"59",X"A0",X"FF",X"65",X"44",X"56",X"00",X"00",X"FF",X"53",X"22",
		X"43",X"50",X"00",X"FF",X"53",X"34",X"33",X"50",X"00",X"FF",X"06",X"54",X"45",X"00",X"00",X"FF",
		X"00",X"66",X"60",X"00",X"00",X"FF",X"08",X"A7",X"00",X"00",X"00",X"FF",X"00",X"99",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",X"27",X"77",X"70",X"FF",X"00",X"04",
		X"22",X"37",X"70",X"FF",X"00",X"05",X"33",X"33",X"5A",X"FF",X"05",X"44",X"54",X"45",X"00",X"FF",
		X"53",X"22",X"34",X"50",X"00",X"FF",X"53",X"34",X"33",X"50",X"00",X"FF",X"06",X"54",X"45",X"50",
		X"00",X"FF",X"00",X"66",X"66",X"00",X"00",X"FF",X"09",X"9A",X"70",X"00",X"00",X"FF",X"00",X"07",
		X"77",X"00",X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",X"27",X"77",X"70",X"FF",
		X"00",X"04",X"22",X"17",X"70",X"FF",X"00",X"65",X"33",X"24",X"59",X"FF",X"32",X"26",X"54",X"44",
		X"A0",X"FF",X"53",X"22",X"56",X"60",X"00",X"FF",X"53",X"33",X"53",X"34",X"00",X"FF",X"05",X"55",
		X"43",X"35",X"00",X"FF",X"00",X"05",X"55",X"50",X"00",X"FF",X"00",X"0A",X"A0",X"00",X"00",X"FF",
		X"00",X"00",X"98",X"00",X"00",X"FF",X"00",X"00",X"44",X"45",X"00",X"FF",X"00",X"04",X"27",X"77",
		X"70",X"FF",X"00",X"04",X"22",X"47",X"70",X"FF",X"00",X"05",X"33",X"24",X"59",X"FF",X"00",X"66",
		X"54",X"44",X"90",X"FF",X"00",X"32",X"56",X"60",X"00",X"FF",X"03",X"23",X"53",X"30",X"00",X"FF",
		X"02",X"55",X"43",X"30",X"00",X"FF",X"00",X"A5",X"55",X"50",X"00",X"FF",X"00",X"0A",X"00",X"00",
		X"00",X"FF",X"00",X"04",X"33",X"50",X"00",X"FF",X"00",X"41",X"71",X"75",X"00",X"FF",X"00",X"71",
		X"11",X"15",X"00",X"FF",X"00",X"77",X"77",X"77",X"00",X"FF",X"04",X"67",X"7A",X"77",X"40",X"FF",
		X"33",X"45",X"55",X"56",X"32",X"FF",X"54",X"55",X"23",X"55",X"45",X"FF",X"05",X"63",X"22",X"36",
		X"50",X"FF",X"00",X"05",X"44",X"50",X"00",X"FF",X"00",X"00",X"80",X"90",X"00",X"FF",X"00",X"00",
		X"A0",X"A0",X"00",X"FF",X"00",X"44",X"35",X"00",X"FF",X"04",X"17",X"17",X"50",X"FF",X"07",X"11",
		X"11",X"70",X"FF",X"07",X"77",X"77",X"70",X"FF",X"06",X"77",X"A7",X"70",X"FF",X"54",X"55",X"55",
		X"65",X"FF",X"42",X"52",X"35",X"34",X"FF",X"52",X"42",X"24",X"25",X"FF",X"00",X"54",X"45",X"00",
		X"FF",X"00",X"0A",X"0A",X"00",X"FF",X"00",X"03",X"34",X"40",X"FF",X"00",X"43",X"23",X"44",X"FF",
		X"00",X"77",X"77",X"77",X"FF",X"00",X"33",X"77",X"97",X"FF",X"00",X"42",X"39",X"9A",X"FF",X"00",
		X"65",X"34",X"A0",X"FF",X"06",X"23",X"54",X"56",X"FF",X"03",X"33",X"52",X"45",X"FF",X"05",X"45",
		X"44",X"63",X"FF",X"00",X"65",X"66",X"00",X"FF",X"00",X"99",X"0A",X"00",X"FF",X"00",X"00",X"88",
		X"A0",X"FF",X"00",X"33",X"34",X"00",X"FF",X"03",X"32",X"23",X"40",X"FF",X"07",X"77",X"77",X"70",
		X"FF",X"07",X"77",X"37",X"70",X"FF",X"04",X"39",X"93",X"40",X"FF",X"00",X"4A",X"A4",X"00",X"FF",
		X"06",X"55",X"55",X"60",X"FF",X"05",X"33",X"34",X"50",X"FF",X"35",X"43",X"35",X"53",X"FF",X"00",
		X"55",X"55",X"00",X"FF",X"00",X"AA",X"0A",X"00",X"FF",X"0A",X"9A",X"AA",X"A0",X"FF",X"00",X"AA",
		X"0A",X"00",X"FF",X"0A",X"9A",X"AA",X"A0",X"FF",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"08",X"58",
		X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"86",X"46",X"60",X"00",X"FF",X"00",X"00",X"00",X"08",
		X"65",X"45",X"57",X"00",X"FF",X"00",X"00",X"00",X"09",X"A5",X"51",X"15",X"70",X"FF",X"00",X"00",
		X"00",X"87",X"65",X"11",X"19",X"70",X"FF",X"00",X"00",X"00",X"9A",X"65",X"51",X"1A",X"3A",X"FF",
		X"00",X"00",X"00",X"87",X"75",X"45",X"62",X"2C",X"FF",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",
		X"2C",X"FF",X"00",X"00",X"00",X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",X"A6",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"86",X"64",X"40",X"00",X"FF",X"00",X"00",X"00",X"00",X"9A",X"3E",X"20",X"00",X"FF",X"08",
		X"70",X"00",X"09",X"68",X"D5",X"40",X"00",X"FF",X"00",X"09",X"00",X"58",X"A3",X"DE",X"50",X"00",
		X"FF",X"00",X"00",X"69",X"00",X"86",X"76",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"07",X"60",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"77",X"66",X"55",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"08",X"58",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"86",
		X"46",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"08",X"65",X"45",X"57",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"09",X"A5",X"51",X"15",X"70",X"FF",X"00",X"00",X"00",X"00",X"87",X"65",X"11",X"19",
		X"70",X"FF",X"00",X"00",X"00",X"00",X"9A",X"65",X"51",X"1A",X"3A",X"FF",X"00",X"00",X"00",X"00",
		X"87",X"75",X"45",X"62",X"2C",X"FF",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",X"2C",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"60",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"9A",X"54",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"9A",X"3D",X"22",X"00",
		X"00",X"FF",X"08",X"79",X"00",X"09",X"7A",X"EC",X"D4",X"90",X"00",X"FF",X"00",X"00",X"69",X"58",
		X"A6",X"55",X"CD",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"86",X"55",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"77",X"66",
		X"55",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"58",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"86",X"46",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"08",X"65",X"45",X"57",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"09",X"A5",X"51",X"15",X"70",X"FF",X"00",X"00",X"00",X"00",X"87",X"65",
		X"11",X"19",X"70",X"FF",X"00",X"00",X"00",X"00",X"9A",X"65",X"51",X"1A",X"3A",X"FF",X"00",X"00",
		X"00",X"00",X"87",X"75",X"45",X"62",X"2C",X"FF",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",
		X"2C",X"FF",X"00",X"00",X"00",X"00",X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"96",X"70",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"09",X"97",X"63",X"D9",X"00",X"00",X"FF",X"87",X"96",X"95",X"97",X"6E",X"54",
		X"33",X"99",X"00",X"FF",X"00",X"00",X"00",X"8A",X"54",X"2C",X"03",X"30",X"00",X"FF",X"00",X"00",
		X"00",X"08",X"54",X"50",X"00",X"E3",X"00",X"FF",X"00",X"00",X"00",X"00",X"76",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"07",X"76",X"65",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"58",
		X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"46",X"60",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"08",X"65",X"45",X"57",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"A5",
		X"51",X"15",X"70",X"FF",X"00",X"00",X"00",X"00",X"00",X"87",X"65",X"11",X"19",X"70",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"9A",X"65",X"51",X"1A",X"3A",X"FF",X"00",X"00",X"00",X"00",X"00",X"87",
		X"75",X"45",X"62",X"2C",X"FF",X"00",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",X"2C",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",X"79",
		X"79",X"00",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"5A",X"5A",X"79",X"77",X"00",X"00",
		X"FF",X"08",X"79",X"69",X"69",X"5E",X"4E",X"44",X"54",X"00",X"00",X"FF",X"00",X"00",X"00",X"64",
		X"26",X"24",X"3C",X"40",X"00",X"00",X"FF",X"00",X"00",X"09",X"44",X"87",X"60",X"53",X"90",X"00",
		X"00",X"FF",X"00",X"00",X"05",X"59",X"00",X"00",X"03",X"90",X"00",X"00",X"FF",X"00",X"00",X"90",
		X"00",X"00",X"00",X"0C",X"C0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"58",X"50",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"86",X"46",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",
		X"65",X"45",X"57",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"A5",X"51",X"15",X"70",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"87",X"65",X"11",X"19",X"70",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"9A",X"65",X"51",X"1A",X"3A",X"FF",X"00",X"00",X"00",X"00",X"00",X"87",X"75",X"45",X"62",X"2C",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",X"2C",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"07",X"97",X"90",X"08",X"60",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"86",X"A4",X"A7",X"97",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"95",X"22",X"54",X"44",X"00",X"00",X"00",X"FF",X"08",X"70",X"09",X"86",X"42",X"73",X"C2",X"00",
		X"00",X"00",X"FF",X"00",X"09",X"50",X"08",X"59",X"03",X"90",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"07",X"44",X"43",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"90",X"39",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"75",
		X"00",X"70",X"00",X"FF",X"00",X"00",X"00",X"68",X"57",X"80",X"00",X"FF",X"00",X"00",X"07",X"65",
		X"54",X"70",X"00",X"FF",X"00",X"00",X"76",X"11",X"55",X"67",X"00",X"FF",X"00",X"0A",X"71",X"19",
		X"14",X"51",X"00",X"FF",X"00",X"07",X"76",X"1A",X"14",X"61",X"00",X"FF",X"00",X"09",X"A6",X"55",
		X"CC",X"AC",X"00",X"FF",X"00",X"08",X"77",X"C2",X"22",X"22",X"C0",X"FF",X"00",X"00",X"AE",X"C2",
		X"22",X"22",X"C0",X"FF",X"00",X"00",X"09",X"7C",X"C9",X"9C",X"00",X"FF",X"00",X"00",X"79",X"79",
		X"80",X"00",X"00",X"FF",X"00",X"0A",X"6A",X"66",X"79",X"00",X"00",X"FF",X"00",X"09",X"52",X"26",
		X"64",X"60",X"00",X"FF",X"80",X"98",X"64",X"23",X"64",X"56",X"00",X"FF",X"79",X"50",X"85",X"93",
		X"30",X"56",X"00",X"FF",X"00",X"00",X"74",X"24",X"00",X"07",X"70",X"FF",X"00",X"00",X"00",X"09",
		X"00",X"00",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"07",X"00",X"00",X"07",X"00",X"FF",X"00",X"07",X"60",X"00",X"67",X"00",X"FF",
		X"00",X"07",X"54",X"45",X"57",X"00",X"FF",X"00",X"06",X"15",X"45",X"16",X"00",X"FF",X"00",X"61",
		X"91",X"59",X"11",X"60",X"FF",X"00",X"66",X"A1",X"6A",X"15",X"60",X"FF",X"0E",X"65",X"22",X"92",
		X"24",X"5E",X"FF",X"06",X"52",X"22",X"22",X"22",X"66",X"FF",X"00",X"E5",X"22",X"B2",X"26",X"E0",
		X"FF",X"00",X"00",X"00",X"80",X"00",X"00",X"FF",X"00",X"00",X"06",X"55",X"60",X"00",X"FF",X"00",
		X"00",X"65",X"44",X"55",X"00",X"FF",X"00",X"00",X"DA",X"22",X"4A",X"60",X"FF",X"00",X"00",X"36",
		X"42",X"46",X"77",X"FF",X"00",X"02",X"2A",X"44",X"4A",X"08",X"FF",X"08",X"00",X"96",X"65",X"60",
		X"00",X"FF",X"00",X"96",X"06",X"08",X"00",X"00",X"FF",X"00",X"00",X"65",X"45",X"86",X"00",X"FF",
		X"00",X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"07",X"50",X"07",X"00",X"FF",X"00",X"00",
		X"06",X"85",X"78",X"00",X"FF",X"00",X"00",X"76",X"55",X"47",X"00",X"FF",X"00",X"07",X"61",X"15",
		X"56",X"70",X"FF",X"00",X"77",X"11",X"19",X"45",X"10",X"FF",X"00",X"77",X"51",X"1A",X"46",X"10",
		X"FF",X"00",X"9A",X"65",X"5C",X"CA",X"C0",X"FF",X"00",X"87",X"7C",X"C2",X"22",X"2C",X"FF",X"00",
		X"0A",X"EC",X"22",X"22",X"2C",X"FF",X"00",X"00",X"77",X"CC",X"99",X"C0",X"FF",X"00",X"00",X"00",
		X"80",X"00",X"00",X"FF",X"00",X"00",X"09",X"A6",X"00",X"00",X"FF",X"00",X"00",X"86",X"64",X"40",
		X"00",X"FF",X"00",X"00",X"9A",X"3E",X"20",X"00",X"FF",X"00",X"09",X"68",X"D5",X"40",X"00",X"FF",
		X"00",X"08",X"A3",X"DE",X"50",X"00",X"FF",X"00",X"50",X"86",X"76",X"00",X"00",X"FF",X"09",X"78",
		X"07",X"60",X"00",X"00",X"FF",X"00",X"00",X"77",X"66",X"55",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"70",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"87",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"57",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"A5",X"DD",X"45",X"60",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"05",X"5D",X"DB",X"54",X"56",X"77",X"FF",X"00",X"00",X"00",X"00",X"0A",X"25",X"B9",
		X"65",X"45",X"70",X"FF",X"00",X"00",X"00",X"00",X"06",X"22",X"25",X"9B",X"D6",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"22",X"92",X"BD",X"D6",X"00",X"FF",X"00",X"00",X"04",X"00",X"00",X"0B",
		X"22",X"5D",X"5A",X"00",X"FF",X"00",X"00",X"04",X"43",X"75",X"68",X"22",X"25",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"9A",X"54",X"25",X"06",X"26",X"A0",X"00",X"FF",X"87",X"00",X"95",X"95",X"44",
		X"25",X"00",X"00",X"00",X"00",X"FF",X"00",X"96",X"00",X"A6",X"54",X"56",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"06",X"57",X"65",X"A3",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"87",X"08",
		X"79",X"94",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"07",X"50",X"04",X"40",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"80",X"00",X"00",X"00",X"6A",
		X"70",X"00",X"00",X"FF",X"09",X"00",X"40",X"00",X"0E",X"55",X"66",X"00",X"00",X"FF",X"06",X"00",
		X"44",X"00",X"05",X"25",X"6D",X"67",X"77",X"FF",X"07",X"90",X"04",X"60",X"02",X"22",X"BD",X"B5",
		X"60",X"FF",X"06",X"67",X"6A",X"56",X"02",X"22",X"99",X"54",X"00",X"FF",X"08",X"04",X"42",X"45",
		X"8B",X"29",X"65",X"44",X"00",X"FF",X"05",X"54",X"22",X"45",X"02",X"22",X"99",X"55",X"00",X"FF",
		X"07",X"04",X"44",X"56",X"02",X"22",X"BD",X"B5",X"60",X"FF",X"07",X"07",X"6A",X"50",X"06",X"24",
		X"5D",X"67",X"77",X"FF",X"00",X"00",X"76",X"00",X"0E",X"65",X"66",X"00",X"00",X"FF",X"00",X"08",
		X"70",X"00",X"00",X"69",X"70",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"05",X"60",X"00",X"FF",X"05",X"44",X"45",X"60",X"FF",X"54",X"21",X"24",X"56",X"FF",X"54",
		X"21",X"24",X"56",X"FF",X"65",X"52",X"45",X"66",X"FF",X"06",X"62",X"46",X"60",X"FF",X"00",X"04",
		X"60",X"00",X"FF",X"00",X"05",X"60",X"00",X"FF",X"04",X"44",X"50",X"FF",X"42",X"12",X"45",X"FF",
		X"42",X"12",X"45",X"FF",X"65",X"24",X"56",X"FF",X"00",X"24",X"00",X"FF",X"00",X"11",X"10",X"FF",
		X"01",X"11",X"11",X"FF",X"00",X"01",X"00",X"FF",X"00",X"07",X"00",X"00",X"07",X"00",X"FF",X"00",
		X"07",X"60",X"00",X"67",X"00",X"FF",X"00",X"07",X"54",X"45",X"57",X"00",X"FF",X"00",X"06",X"15",
		X"45",X"16",X"00",X"FF",X"00",X"61",X"91",X"59",X"11",X"60",X"FF",X"00",X"66",X"A1",X"6A",X"15",
		X"60",X"FF",X"0E",X"65",X"22",X"92",X"24",X"5E",X"FF",X"06",X"52",X"22",X"22",X"22",X"66",X"FF",
		X"00",X"E5",X"22",X"B2",X"26",X"E0",X"FF",X"00",X"22",X"50",X"00",X"00",X"00",X"FF",X"00",X"44",
		X"50",X"00",X"00",X"00",X"FF",X"00",X"07",X"87",X"77",X"87",X"00",X"FF",X"00",X"07",X"69",X"A9",
		X"67",X"00",X"FF",X"00",X"87",X"54",X"45",X"57",X"80",X"FF",X"00",X"86",X"15",X"45",X"16",X"80",
		X"FF",X"00",X"61",X"19",X"51",X"91",X"60",X"FF",X"00",X"66",X"1A",X"61",X"A5",X"60",X"FF",X"0E",
		X"65",X"22",X"92",X"24",X"5E",X"FF",X"06",X"52",X"22",X"22",X"22",X"66",X"FF",X"00",X"E5",X"22",
		X"B2",X"26",X"E0",X"FF",X"00",X"22",X"50",X"00",X"06",X"60",X"FF",X"00",X"44",X"50",X"00",X"05",
		X"60",X"FF",X"00",X"00",X"00",X"00",X"05",X"50",X"FF",X"00",X"00",X"00",X"00",X"02",X"50",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"08",X"58",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"86",X"46",X"60",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"08",X"65",X"45",X"57",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",X"A5",X"51",
		X"19",X"70",X"FF",X"00",X"00",X"00",X"00",X"87",X"65",X"11",X"1E",X"70",X"FF",X"00",X"00",X"00",
		X"00",X"9A",X"65",X"51",X"11",X"3A",X"FF",X"00",X"00",X"00",X"00",X"87",X"75",X"45",X"62",X"2C",
		X"FF",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",X"2C",X"FF",X"00",X"00",X"00",X"00",X"08",
		X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"08",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"9A",X"52",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"9A",X"54",X"63",X"90",X"00",X"FF",X"00",X"00",X"00",
		X"09",X"7A",X"E3",X"37",X"29",X"00",X"FF",X"00",X"00",X"69",X"58",X"A3",X"36",X"50",X"64",X"00",
		X"FF",X"08",X"79",X"00",X"00",X"84",X"56",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"07",X"43",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"95",X"33",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"08",X"58",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"86",X"46",X"60",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"08",X"65",X"45",X"57",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",
		X"A5",X"51",X"19",X"70",X"FF",X"00",X"00",X"00",X"00",X"87",X"65",X"11",X"1A",X"70",X"FF",X"00",
		X"00",X"00",X"00",X"9A",X"65",X"51",X"11",X"3A",X"FF",X"00",X"00",X"00",X"00",X"87",X"75",X"45",
		X"62",X"2C",X"FF",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",X"2C",X"FF",X"00",X"00",X"00",
		X"00",X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"69",X"6A",X"79",X"77",X"00",X"00",X"FF",X"00",X"00",X"69",X"69",X"4E",
		X"44",X"54",X"00",X"00",X"FF",X"00",X"09",X"00",X"8A",X"23",X"35",X"49",X"00",X"00",X"FF",X"09",
		X"80",X"09",X"33",X"46",X"50",X"C4",X"90",X"00",X"FF",X"00",X"00",X"03",X"39",X"80",X"00",X"0C",
		X"40",X"00",X"FF",X"00",X"00",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"58",X"50",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"86",X"46",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"65",
		X"45",X"57",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"A5",X"51",X"11",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"87",X"65",X"11",X"1A",X"70",X"FF",X"00",X"00",X"00",X"00",X"00",X"9A",
		X"65",X"51",X"19",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"87",X"75",X"45",X"52",X"2A",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"9A",X"E5",X"45",X"22",X"2C",X"FF",X"08",X"70",X"00",X"00",X"79",
		X"08",X"77",X"66",X"39",X"90",X"FF",X"00",X"09",X"00",X"08",X"59",X"79",X"00",X"80",X"00",X"00",
		X"FF",X"00",X"00",X"69",X"6A",X"A7",X"5A",X"79",X"77",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",
		X"24",X"A7",X"44",X"54",X"00",X"00",X"FF",X"00",X"00",X"88",X"44",X"55",X"24",X"3C",X"40",X"00",
		X"00",X"FF",X"00",X"00",X"84",X"86",X"88",X"65",X"53",X"90",X"00",X"00",X"FF",X"00",X"96",X"68",
		X"00",X"00",X"00",X"73",X"90",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"C9",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"06",X"06",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"85",X"85",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"08",X"64",X"66",X"00",X"00",X"FF",X"00",X"00",X"00",X"86",X"54",X"55",X"70",X"00",X"FF",
		X"00",X"00",X"00",X"9A",X"55",X"11",X"57",X"00",X"FF",X"00",X"00",X"08",X"76",X"51",X"11",X"97",
		X"00",X"FF",X"00",X"00",X"09",X"A6",X"55",X"11",X"A3",X"A0",X"FF",X"00",X"00",X"08",X"77",X"54",
		X"56",X"22",X"C0",X"FF",X"00",X"00",X"09",X"AE",X"54",X"52",X"22",X"C0",X"FF",X"00",X"00",X"00",
		X"87",X"76",X"63",X"99",X"00",X"FF",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"FF",X"00",
		X"00",X"00",X"00",X"9A",X"68",X"88",X"82",X"FF",X"00",X"00",X"00",X"08",X"66",X"42",X"22",X"20",
		X"FF",X"00",X"00",X"00",X"09",X"AE",X"54",X"00",X"00",X"FF",X"87",X"00",X"00",X"96",X"64",X"54",
		X"00",X"00",X"FF",X"00",X"90",X"05",X"8A",X"E5",X"55",X"00",X"00",X"FF",X"00",X"06",X"90",X"08",
		X"67",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"07",X"76",X"65",X"50",X"00",X"FF",X"00",X"07",X"00",X"00",X"07",X"00",X"FF",X"00",X"07",
		X"60",X"00",X"67",X"00",X"FF",X"00",X"07",X"54",X"45",X"57",X"00",X"FF",X"00",X"06",X"15",X"45",
		X"16",X"00",X"FF",X"00",X"61",X"91",X"59",X"11",X"60",X"FF",X"00",X"66",X"A1",X"6A",X"15",X"60",
		X"FF",X"0E",X"65",X"22",X"92",X"24",X"5E",X"FF",X"06",X"52",X"22",X"22",X"22",X"66",X"FF",X"00",
		X"E5",X"22",X"B2",X"26",X"E0",X"FF",X"00",X"77",X"00",X"00",X"07",X"70",X"FF",X"00",X"55",X"00",
		X"00",X"05",X"50",X"FF",X"00",X"22",X"00",X"00",X"02",X"20",X"FF",X"00",X"02",X"00",X"00",X"02",
		X"00",X"FF",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"02",X"EE",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"23",X"EE",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",
		X"3E",X"EE",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"07",X"CC",
		X"CC",X"CB",X"00",X"00",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",X"73",X"3E",X"EE",
		X"E3",X"00",X"7C",X"54",X"DD",X"DD",X"45",X"00",X"00",X"00",X"00",X"FF",X"CC",X"CC",X"CC",X"CA",
		X"67",X"55",X"CC",X"44",X"44",X"5C",X"77",X"00",X"00",X"00",X"FF",X"CC",X"CC",X"CC",X"C6",X"45",
		X"63",X"3C",X"CC",X"BB",X"C5",X"66",X"70",X"00",X"00",X"FF",X"73",X"EE",X"E7",X"65",X"63",X"32",
		X"22",X"2E",X"EE",X"EE",X"E3",X"67",X"00",X"00",X"FF",X"73",X"EE",X"E7",X"66",X"33",X"22",X"22",
		X"22",X"22",X"22",X"2E",X"36",X"00",X"00",X"FF",X"07",X"EE",X"33",X"63",X"22",X"11",X"12",X"22",
		X"22",X"11",X"22",X"E3",X"60",X"00",X"FF",X"07",X"3E",X"33",X"EE",X"22",X"55",X"66",X"66",X"33",
		X"E1",X"12",X"23",X"48",X"80",X"FF",X"00",X"76",X"33",X"EE",X"E5",X"6E",X"33",X"33",X"3E",X"A1",
		X"12",X"23",X"49",X"E0",X"FF",X"00",X"66",X"73",X"33",X"56",X"E3",X"33",X"33",X"EA",X"71",X"12",
		X"E3",X"50",X"00",X"FF",X"00",X"05",X"67",X"64",X"43",X"63",X"33",X"3E",X"A7",X"22",X"22",X"E6",
		X"50",X"00",X"FF",X"00",X"00",X"56",X"5D",X"43",X"66",X"3E",X"AA",X"73",X"22",X"EE",X"65",X"00",
		X"00",X"FF",X"00",X"00",X"05",X"44",X"D4",X"77",X"77",X"77",X"63",X"3E",X"E6",X"50",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"D4",X"44",X"45",X"57",X"75",X"66",X"66",X"75",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"D4",X"44",X"45",X"55",X"54",X"44",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"7E",X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",X"83",X"88",X"00",
		X"0D",X"70",X"00",X"FF",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"E0",X"00",X"FF",X"00",
		X"00",X"EE",X"ED",X"69",X"50",X"00",X"EE",X"EE",X"00",X"FF",X"00",X"88",X"88",X"EE",X"D6",X"50",
		X"0E",X"88",X"88",X"E0",X"FF",X"08",X"88",X"88",X"2E",X"77",X"7E",X"E8",X"88",X"88",X"8E",X"FF",
		X"08",X"86",X"4C",X"CE",X"66",X"80",X"08",X"84",X"68",X"8E",X"FF",X"08",X"86",X"68",X"8D",X"DD",
		X"D0",X"08",X"86",X"68",X"80",X"FF",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"31",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"7E",X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"83",X"88",X"00",X"0D",X"70",X"00",X"FF",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"E0",
		X"00",X"FF",X"00",X"00",X"EE",X"ED",X"69",X"50",X"00",X"EE",X"EE",X"00",X"FF",X"00",X"88",X"88",
		X"EE",X"D6",X"50",X"0E",X"88",X"88",X"E0",X"FF",X"08",X"88",X"88",X"DE",X"77",X"7E",X"E8",X"88",
		X"88",X"8E",X"FF",X"08",X"86",X"4C",X"CE",X"66",X"80",X"08",X"84",X"68",X"8E",X"FF",X"08",X"86",
		X"68",X"8D",X"DD",X"D0",X"08",X"D6",X"68",X"80",X"FF",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"D8",X"88",X"00",X"FF",X"03",X"00",X"22",X"30",X"00",X"FF",X"00",X"31",X"22",X"23",X"80",X"FF",
		X"03",X"19",X"22",X"AA",X"3A",X"FF",X"03",X"22",X"88",X"AB",X"3B",X"FF",X"03",X"38",X"88",X"BD",
		X"3D",X"FF",X"03",X"33",X"88",X"BD",X"3D",X"FF",X"08",X"33",X"77",X"24",X"45",X"FF",X"00",X"83",
		X"E7",X"44",X"44",X"FF",X"00",X"08",X"82",X"66",X"60",X"FF",X"00",X"00",X"08",X"00",X"00",X"FF",
		X"00",X"03",X"12",X"30",X"00",X"FF",X"02",X"32",X"19",X"13",X"33",X"FF",X"21",X"22",X"11",X"11",
		X"20",X"FF",X"21",X"32",X"22",X"33",X"00",X"FF",X"83",X"33",X"38",X"00",X"00",X"FF",X"08",X"88",
		X"80",X"00",X"00",X"FF",X"00",X"60",X"00",X"00",X"00",X"FF",X"06",X"66",X"60",X"00",X"00",X"FF",
		X"00",X"80",X"22",X"30",X"00",X"FF",X"00",X"81",X"22",X"23",X"80",X"FF",X"02",X"92",X"2A",X"A3",
		X"AA",X"FF",X"03",X"28",X"8A",X"B8",X"AB",X"FF",X"03",X"88",X"8B",X"D8",X"BD",X"FF",X"03",X"38",
		X"8B",X"D8",X"BD",X"FF",X"08",X"17",X"74",X"44",X"57",X"FF",X"00",X"3E",X"E4",X"44",X"4E",X"FF",
		X"00",X"08",X"82",X"66",X"60",X"FF",X"00",X"00",X"08",X"00",X"00",X"FF",X"00",X"82",X"11",X"30",
		X"00",X"FF",X"03",X"32",X"11",X"91",X"33",X"FF",X"31",X"22",X"21",X"22",X"20",X"FF",X"22",X"32",
		X"22",X"33",X"00",X"FF",X"03",X"53",X"38",X"00",X"00",X"FF",X"00",X"58",X"80",X"00",X"00",X"FF",
		X"05",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"30",X"00",X"FF",X"00",X"22",X"11",X"12",
		X"30",X"FF",X"03",X"29",X"92",X"99",X"23",X"FF",X"03",X"8A",X"A8",X"AA",X"83",X"FF",X"08",X"8A",
		X"D8",X"DA",X"88",X"FF",X"0D",X"8A",X"D8",X"DA",X"8D",X"FF",X"07",X"72",X"44",X"42",X"77",X"FF",
		X"07",X"E4",X"44",X"55",X"7E",X"FF",X"00",X"23",X"55",X"63",X"20",X"FF",X"00",X"00",X"08",X"80",
		X"00",X"FF",X"00",X"03",X"33",X"30",X"00",X"FF",X"01",X"12",X"11",X"92",X"33",X"FF",X"31",X"22",
		X"21",X"11",X"20",X"FF",X"83",X"32",X"22",X"33",X"00",X"FF",X"08",X"86",X"38",X"00",X"00",X"FF",
		X"00",X"55",X"56",X"00",X"00",X"FF",X"00",X"00",X"22",X"30",X"08",X"FF",X"00",X"22",X"11",X"12",
		X"30",X"FF",X"03",X"29",X"92",X"99",X"23",X"FF",X"03",X"8A",X"A8",X"AA",X"83",X"FF",X"08",X"8A",
		X"D8",X"DA",X"88",X"FF",X"0D",X"8A",X"D8",X"DA",X"8D",X"FF",X"07",X"72",X"44",X"42",X"77",X"FF",
		X"07",X"E4",X"48",X"55",X"7E",X"FF",X"00",X"23",X"55",X"63",X"80",X"FF",X"00",X"00",X"08",X"80",
		X"00",X"FF",X"00",X"00",X"33",X"30",X"00",X"FF",X"02",X"12",X"21",X"93",X"33",X"FF",X"21",X"22",
		X"11",X"11",X"20",X"FF",X"32",X"22",X"22",X"33",X"00",X"FF",X"08",X"23",X"23",X"00",X"00",X"FF",
		X"00",X"88",X"60",X"00",X"00",X"FF",X"00",X"06",X"66",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",
		X"00",X"88",X"44",X"55",X"24",X"3C",X"40",X"00",X"00",X"FF",X"00",X"00",X"84",X"86",X"88",X"65",
		X"53",X"90",X"00",X"00",X"FF",X"00",X"96",X"68",X"00",X"00",X"00",X"73",X"90",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"C9",X"00",X"00",X"FF",X"00",X"00",X"00",X"09",X"09",
		X"00",X"90",X"FF",X"00",X"00",X"09",X"03",X"34",X"44",X"00",X"FF",X"00",X"09",X"03",X"34",X"67",
		X"55",X"C0",X"FF",X"00",X"00",X"34",X"46",X"66",X"5C",X"E0",X"FF",X"00",X"00",X"45",X"32",X"34",
		X"44",X"E4",X"FF",X"08",X"03",X"57",X"61",X"22",X"24",X"43",X"FF",X"00",X"35",X"24",X"65",X"12",
		X"62",X"30",X"FF",X"00",X"01",X"18",X"9A",X"11",X"9E",X"00",X"FF",X"00",X"00",X"08",X"9A",X"E0",
		X"88",X"E0",X"FF",X"00",X"00",X"00",X"09",X"09",X"00",X"90",X"FF",X"00",X"00",X"09",X"03",X"34",
		X"44",X"00",X"FF",X"00",X"09",X"03",X"34",X"67",X"55",X"C0",X"FF",X"00",X"00",X"34",X"23",X"66",
		X"5C",X"E0",X"FF",X"00",X"00",X"47",X"55",X"34",X"44",X"E4",X"FF",X"00",X"02",X"56",X"65",X"22",
		X"24",X"43",X"FF",X"08",X"04",X"38",X"9A",X"12",X"62",X"30",X"FF",X"00",X"22",X"18",X"9A",X"19",
		X"AE",X"00",X"FF",X"00",X"00",X"EE",X"E0",X"08",X"90",X"00",X"FF",X"00",X"00",X"00",X"09",X"09",
		X"00",X"90",X"FF",X"00",X"00",X"09",X"03",X"34",X"44",X"00",X"FF",X"00",X"09",X"03",X"45",X"67",
		X"55",X"E0",X"FF",X"00",X"00",X"34",X"55",X"66",X"5C",X"E0",X"FF",X"00",X"00",X"46",X"63",X"34",
		X"44",X"C4",X"FF",X"00",X"03",X"36",X"75",X"22",X"24",X"43",X"FF",X"09",X"05",X"24",X"44",X"19",
		X"A2",X"30",X"FF",X"00",X"33",X"18",X"9A",X"19",X"A1",X"10",X"FF",X"00",X"00",X"E8",X"9A",X"00",
		X"01",X"10",X"FF",X"00",X"00",X"00",X"08",X"09",X"09",X"00",X"FF",X"00",X"00",X"08",X"03",X"44",
		X"44",X"00",X"FF",X"00",X"00",X"83",X"67",X"54",X"EC",X"4E",X"FF",X"00",X"00",X"35",X"76",X"54",
		X"EC",X"4E",X"FF",X"00",X"00",X"45",X"63",X"33",X"CC",X"4C",X"FF",X"00",X"02",X"55",X"37",X"52",
		X"44",X"43",X"FF",X"08",X"03",X"14",X"3A",X"A1",X"23",X"30",X"FF",X"00",X"12",X"18",X"8A",X"A1",
		X"11",X"10",X"FF",X"00",X"00",X"E8",X"8E",X"E0",X"01",X"10",X"FF",X"00",X"00",X"08",X"09",X"09",
		X"00",X"FF",X"00",X"00",X"03",X"44",X"56",X"43",X"FF",X"00",X"08",X"45",X"5E",X"C5",X"EC",X"FF",
		X"00",X"84",X"54",X"6E",X"C4",X"EC",X"FF",X"00",X"34",X"54",X"5C",X"C4",X"CC",X"FF",X"00",X"46",
		X"43",X"55",X"66",X"54",X"FF",X"81",X"33",X"64",X"23",X"44",X"30",X"FF",X"01",X"88",X"A9",X"11",
		X"11",X"10",X"FF",X"00",X"01",X"A9",X"11",X"08",X"80",X"FF",X"00",X"00",X"80",X"90",X"00",X"FF",
		X"00",X"03",X"44",X"44",X"30",X"FF",X"00",X"35",X"CC",X"5C",X"C3",X"FF",X"05",X"46",X"EC",X"5E",
		X"C4",X"FF",X"06",X"46",X"EC",X"5E",X"C4",X"FF",X"04",X"35",X"56",X"65",X"53",X"FF",X"83",X"33",
		X"45",X"54",X"3E",X"FF",X"11",X"A9",X"22",X"22",X"89",X"FF",X"01",X"A9",X"11",X"E8",X"9A",X"FF",
		X"00",X"00",X"00",X"00",X"31",X"80",X"FF",X"00",X"00",X"00",X"03",X"30",X"00",X"FF",X"00",X"00",
		X"0A",X"A3",X"53",X"90",X"FF",X"00",X"00",X"E9",X"45",X"54",X"00",X"FF",X"00",X"00",X"88",X"65",
		X"54",X"39",X"FF",X"0A",X"98",X"11",X"12",X"66",X"30",X"FF",X"00",X"12",X"66",X"65",X"66",X"30",
		X"FF",X"03",X"22",X"32",X"55",X"67",X"49",X"FF",X"04",X"EC",X"46",X"24",X"55",X"40",X"FF",X"00",
		X"EC",X"44",X"44",X"44",X"00",X"FF",X"00",X"CC",X"44",X"44",X"30",X"90",X"FF",X"00",X"02",X"23",
		X"20",X"00",X"00",X"FF",X"00",X"00",X"90",X"09",X"00",X"00",X"FF",X"00",X"00",X"09",X"00",X"90",
		X"00",X"00",X"FF",X"08",X"09",X"03",X"33",X"44",X"09",X"00",X"FF",X"01",X"03",X"44",X"66",X"75",
		X"40",X"00",X"FF",X"03",X"35",X"55",X"66",X"65",X"43",X"00",X"FF",X"00",X"33",X"55",X"25",X"54",
		X"44",X"09",X"FF",X"00",X"0A",X"46",X"16",X"52",X"44",X"20",X"FF",X"00",X"0A",X"98",X"16",X"26",
		X"44",X"30",X"FF",X"00",X"00",X"E8",X"16",X"34",X"44",X"29",X"FF",X"00",X"00",X"00",X"82",X"2C",
		X"CC",X"20",X"FF",X"00",X"00",X"00",X"91",X"2E",X"EC",X"00",X"FF",X"00",X"00",X"00",X"A0",X"34",
		X"00",X"00",X"FF",X"80",X"00",X"00",X"00",X"FF",X"02",X"40",X"00",X"00",X"FF",X"01",X"53",X"00",
		X"00",X"FF",X"E1",X"25",X"39",X"00",X"FF",X"E1",X"25",X"50",X"00",X"FF",X"88",X"47",X"54",X"90",
		X"FF",X"99",X"66",X"44",X"00",X"FF",X"AA",X"54",X"46",X"39",X"FF",X"0E",X"12",X"56",X"30",X"FF",
		X"EE",X"22",X"67",X"49",X"FF",X"89",X"65",X"55",X"30",X"FF",X"89",X"25",X"54",X"30",X"FF",X"00",
		X"34",X"CC",X"39",X"FF",X"00",X"14",X"EE",X"C0",X"FF",X"00",X"01",X"50",X"00",X"FF",X"00",X"80",
		X"00",X"00",X"FF",X"02",X"00",X"00",X"00",X"FF",X"02",X"53",X"00",X"00",X"FF",X"13",X"35",X"39",
		X"00",X"FF",X"E1",X"25",X"50",X"00",X"FF",X"18",X"87",X"64",X"90",X"FF",X"09",X"96",X"74",X"00",
		X"FF",X"0A",X"A4",X"46",X"39",X"FF",X"0E",X"12",X"56",X"30",X"FF",X"89",X"22",X"67",X"49",X"FF",
		X"8A",X"65",X"55",X"30",X"FF",X"08",X"25",X"54",X"30",X"FF",X"08",X"34",X"CC",X"39",X"FF",X"00",
		X"24",X"EE",X"C0",X"FF",X"00",X"02",X"50",X"00",X"FF",X"00",X"80",X"00",X"00",X"FF",X"02",X"00",
		X"00",X"00",X"FF",X"02",X"43",X"00",X"00",X"FF",X"03",X"65",X"30",X"00",X"FF",X"02",X"25",X"59",
		X"00",X"FF",X"02",X"26",X"64",X"00",X"FF",X"88",X"47",X"64",X"90",X"FF",X"99",X"57",X"46",X"30",
		X"FF",X"AA",X"42",X"56",X"39",X"FF",X"02",X"96",X"64",X"40",X"FF",X"02",X"A6",X"63",X"39",X"FF",
		X"18",X"33",X"34",X"30",X"FF",X"11",X"34",X"CC",X"39",X"FF",X"00",X"24",X"EE",X"40",X"FF",X"00",
		X"02",X"50",X"00",X"FF",X"00",X"00",X"00",X"90",X"90",X"80",X"FF",X"00",X"00",X"90",X"33",X"43",
		X"30",X"FF",X"00",X"90",X"33",X"46",X"75",X"53",X"FF",X"00",X"03",X"44",X"33",X"66",X"43",X"FF",
		X"00",X"35",X"56",X"63",X"55",X"43",X"FF",X"80",X"56",X"76",X"62",X"22",X"30",X"FF",X"03",X"32",
		X"66",X"51",X"26",X"20",X"FF",X"00",X"11",X"89",X"A1",X"19",X"E0",X"FF",X"0E",X"E0",X"89",X"AE",
		X"08",X"8E",X"FF",X"00",X"00",X"09",X"23",X"09",X"FF",X"00",X"02",X"22",X"25",X"20",X"FF",X"00",
		X"24",X"94",X"45",X"52",X"FF",X"02",X"46",X"66",X"54",X"63",X"FF",X"02",X"46",X"77",X"64",X"63",
		X"FF",X"02",X"56",X"97",X"64",X"23",X"FF",X"02",X"35",X"66",X"54",X"11",X"FF",X"00",X"11",X"28",
		X"9A",X"19",X"FF",X"00",X"89",X"08",X"9A",X"00",X"FF",X"00",X"22",X"22",X"00",X"FF",X"02",X"49",
		X"54",X"20",X"FF",X"02",X"46",X"75",X"20",X"FF",X"24",X"59",X"55",X"42",X"FF",X"25",X"22",X"22",
		X"42",X"FF",X"22",X"49",X"44",X"22",X"FF",X"24",X"66",X"65",X"42",X"FF",X"34",X"69",X"76",X"52",
		X"FF",X"35",X"67",X"76",X"52",X"FF",X"24",X"56",X"65",X"42",X"FF",X"E3",X"49",X"43",X"2E",X"FF",
		X"89",X"A0",X"08",X"9A",X"FF",X"00",X"00",X"22",X"00",X"00",X"FF",X"00",X"0C",X"55",X"C0",X"88",
		X"FF",X"08",X"2E",X"94",X"E2",X"A9",X"FF",X"09",X"24",X"67",X"52",X"62",X"FF",X"03",X"45",X"95",
		X"54",X"30",X"FF",X"03",X"52",X"44",X"44",X"30",X"FF",X"00",X"33",X"94",X"42",X"30",X"FF",X"08",
		X"36",X"66",X"53",X"00",X"FF",X"09",X"36",X"97",X"63",X"00",X"FF",X"00",X"36",X"77",X"63",X"00",
		X"FF",X"00",X"03",X"96",X"40",X"00",X"FF",X"00",X"03",X"56",X"30",X"00",X"FF",X"00",X"00",X"35",
		X"00",X"00",X"FF",X"00",X"00",X"02",X"00",X"00",X"FF",X"00",X"00",X"00",X"80",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"43",X"00",X"FF",X"00",X"00",X"00",X"90",X"CE",X"E3",X"00",X"FF",X"00",
		X"00",X"00",X"02",X"CC",X"C5",X"21",X"FF",X"00",X"00",X"00",X"23",X"44",X"44",X"41",X"FF",X"00",
		X"09",X"09",X"33",X"57",X"7A",X"3E",X"FF",X"00",X"00",X"35",X"66",X"55",X"69",X"20",X"FF",X"00",
		X"03",X"55",X"67",X"72",X"33",X"20",X"FF",X"08",X"04",X"62",X"24",X"54",X"33",X"00",X"FF",X"00",
		X"22",X"32",X"28",X"9A",X"20",X"00",X"FF",X"00",X"00",X"00",X"08",X"9A",X"00",X"00",X"FF",X"00",
		X"80",X"00",X"00",X"00",X"FF",X"02",X"00",X"00",X"00",X"00",X"FF",X"02",X"43",X"09",X"00",X"00",
		X"FF",X"03",X"65",X"30",X"00",X"00",X"FF",X"02",X"25",X"59",X"00",X"00",X"FF",X"02",X"26",X"63",
		X"20",X"90",X"FF",X"88",X"47",X"63",X"32",X"00",X"FF",X"99",X"57",X"55",X"4C",X"C0",X"FF",X"AA",
		X"42",X"57",X"4C",X"E0",X"FF",X"02",X"33",X"67",X"4C",X"E4",X"FF",X"00",X"33",X"9A",X"45",X"33",
		X"FF",X"00",X"02",X"23",X"42",X"00",X"FF",X"00",X"00",X"0E",X"11",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"34",X"43",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"62",X"24",X"32",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"34",X"23",X"52",X"42",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"13",X"42",X"36",X"43",X"23",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"03",X"42",X"35",X"73",X"23",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"42",X"52",X"54",X"43",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"22",X"22",X"43",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"32",X"44",X"21",X"30",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"23",X"03",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"04",X"44",X"44",X"44",X"40",X"00",X"FF",X"00",X"00",X"44",X"88",X"88",X"88",X"44",X"00",
		X"FF",X"00",X"04",X"48",X"88",X"88",X"88",X"84",X"40",X"FF",X"00",X"04",X"88",X"88",X"85",X"55",
		X"84",X"45",X"FF",X"00",X"04",X"88",X"85",X"55",X"45",X"58",X"44",X"FF",X"08",X"04",X"48",X"85",
		X"54",X"76",X"58",X"44",X"FF",X"40",X"04",X"48",X"85",X"45",X"63",X"58",X"44",X"FF",X"00",X"00",
		X"44",X"88",X"74",X"47",X"55",X"45",X"FF",X"00",X"40",X"04",X"48",X"85",X"64",X"55",X"85",X"FF",
		X"00",X"00",X"00",X"44",X"45",X"03",X"58",X"85",X"FF",X"05",X"40",X"00",X"00",X"00",X"35",X"48",
		X"50",X"FF",X"00",X"54",X"00",X"00",X"47",X"44",X"48",X"00",X"FF",X"00",X"55",X"74",X"43",X"44",
		X"48",X"80",X"04",X"FF",X"00",X"05",X"55",X"44",X"48",X"80",X"00",X"00",X"FF",X"00",X"00",X"05",
		X"50",X"50",X"00",X"70",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"54",X"44",X"55",X"50",X"00",X"00",X"FF",X"00",X"04",X"44",X"44",X"48",X"85",
		X"00",X"00",X"FF",X"00",X"44",X"48",X"88",X"55",X"88",X"80",X"00",X"FF",X"04",X"48",X"85",X"55",
		X"55",X"54",X"48",X"00",X"FF",X"04",X"88",X"55",X"63",X"74",X"35",X"48",X"00",X"FF",X"04",X"88",
		X"54",X"76",X"46",X"03",X"44",X"80",X"FF",X"44",X"88",X"55",X"45",X"45",X"50",X"7A",X"80",X"FF",
		X"44",X"88",X"85",X"54",X"78",X"40",X"44",X"45",X"FF",X"44",X"88",X"85",X"55",X"88",X"40",X"03",
		X"40",X"FF",X"04",X"88",X"88",X"88",X"84",X"40",X"04",X"45",X"FF",X"04",X"48",X"88",X"88",X"44",
		X"00",X"04",X"55",X"FF",X"00",X"44",X"88",X"44",X"40",X"00",X"07",X"50",X"FF",X"00",X"04",X"44",
		X"44",X"00",X"00",X"45",X"50",X"FF",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"00",X"FF",X"00",
		X"00",X"00",X"04",X"00",X"05",X"00",X"00",X"FF",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"40",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",X"44",X"44",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"44",X"44",X"44",X"44",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"44",X"44",X"88",X"88",X"84",X"44",X"00",X"00",X"FF",X"00",X"00",X"04",
		X"44",X"88",X"88",X"88",X"84",X"45",X"48",X"00",X"FF",X"00",X"00",X"04",X"48",X"88",X"88",X"88",
		X"88",X"44",X"50",X"80",X"FF",X"00",X"00",X"44",X"48",X"88",X"98",X"88",X"88",X"84",X"40",X"00",
		X"FF",X"00",X"00",X"44",X"48",X"88",X"87",X"63",X"78",X"84",X"44",X"00",X"FF",X"00",X"00",X"54",
		X"88",X"88",X"74",X"44",X"37",X"88",X"44",X"00",X"FF",X"00",X"00",X"54",X"88",X"87",X"54",X"34",
		X"43",X"88",X"44",X"00",X"FF",X"00",X"00",X"04",X"88",X"87",X"55",X"33",X"47",X"88",X"84",X"00",
		X"FF",X"00",X"08",X"04",X"88",X"89",X"33",X"39",X"43",X"88",X"84",X"00",X"FF",X"00",X"00",X"00",
		X"48",X"88",X"73",X"38",X"57",X"48",X"45",X"00",X"FF",X"00",X"00",X"00",X"55",X"88",X"88",X"88",
		X"78",X"88",X"85",X"00",X"FF",X"00",X"08",X"07",X"05",X"58",X"88",X"00",X"07",X"88",X"55",X"80",
		X"FF",X"00",X"00",X"04",X"70",X"00",X"00",X"00",X"48",X"85",X"45",X"00",X"FF",X"00",X"00",X"00",
		X"44",X"07",X"77",X"07",X"78",X"44",X"50",X"00",X"FF",X"00",X"00",X"40",X"00",X"44",X"44",X"66",
		X"84",X"4A",X"40",X"00",X"FF",X"00",X"00",X"04",X"70",X"07",X"88",X"44",X"44",X"54",X"00",X"00",
		X"FF",X"00",X"00",X"04",X"44",X"44",X"44",X"44",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"54",X"44",X"45",X"55",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"08",X"00",X"44",X"44",X"45",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"04",
		X"54",X"44",X"48",X"84",X"85",X"45",X"40",X"00",X"FF",X"00",X"00",X"45",X"44",X"48",X"88",X"88",
		X"88",X"54",X"A4",X"00",X"FF",X"00",X"00",X"44",X"48",X"88",X"88",X"84",X"88",X"84",X"45",X"00",
		X"FF",X"00",X"04",X"44",X"88",X"87",X"37",X"37",X"87",X"88",X"44",X"50",X"FF",X"00",X"04",X"88",
		X"88",X"73",X"44",X"45",X"70",X"47",X"84",X"50",X"FF",X"00",X"44",X"88",X"88",X"34",X"43",X"98",
		X"80",X"07",X"64",X"45",X"FF",X"00",X"44",X"88",X"88",X"64",X"33",X"33",X"80",X"00",X"64",X"45",
		X"FF",X"00",X"44",X"88",X"88",X"74",X"45",X"33",X"88",X"07",X"48",X"45",X"FF",X"00",X"44",X"88",
		X"89",X"87",X"55",X"37",X"88",X"07",X"48",X"44",X"FF",X"00",X"44",X"48",X"88",X"88",X"77",X"98",
		X"88",X"07",X"47",X"44",X"FF",X"00",X"04",X"48",X"88",X"88",X"88",X"88",X"85",X"00",X"40",X"44",
		X"FF",X"00",X"04",X"44",X"88",X"88",X"88",X"88",X"55",X"04",X"00",X"44",X"FF",X"00",X"00",X"44",
		X"44",X"48",X"88",X"84",X"50",X"74",X"07",X"45",X"FF",X"00",X"00",X"04",X"44",X"44",X"44",X"40",
		X"07",X"40",X"04",X"40",X"FF",X"00",X"00",X"00",X"04",X"45",X"50",X"00",X"00",X"00",X"40",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"02",X"23",X"00",X"30",X"FF",X"02",X"21",X"12",X"33",X"00",X"FF",X"32",X"99",X"29",
		X"93",X"30",X"FF",X"38",X"AA",X"8A",X"A8",X"30",X"FF",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"D8",
		X"AD",X"8D",X"A8",X"D0",X"FF",X"77",X"24",X"44",X"27",X"70",X"FF",X"7E",X"44",X"85",X"47",X"E0",
		X"FF",X"02",X"35",X"56",X"32",X"00",X"FF",X"00",X"00",X"30",X"00",X"00",X"FF",X"00",X"03",X"13",
		X"00",X"00",X"FF",X"00",X"31",X"91",X"30",X"00",X"FF",X"02",X"23",X"A2",X"23",X"00",X"FF",X"02",
		X"28",X"A8",X"23",X"00",X"FF",X"03",X"81",X"91",X"83",X"00",X"FF",X"00",X"32",X"33",X"30",X"00",
		X"FF",X"04",X"56",X"06",X"00",X"00",X"FF",X"00",X"56",X"86",X"55",X"00",X"FF",X"06",X"00",X"00",
		X"FF",X"00",X"05",X"56",X"65",X"56",X"00",X"FF",X"00",X"80",X"22",X"30",X"00",X"00",X"FF",X"00",
		X"81",X"22",X"23",X"80",X"00",X"FF",X"02",X"92",X"2A",X"B3",X"AB",X"00",X"FF",X"03",X"28",X"8B",
		X"D8",X"BD",X"00",X"FF",X"03",X"88",X"8B",X"D8",X"BD",X"00",X"FF",X"03",X"38",X"8A",X"A8",X"AA",
		X"00",X"FF",X"08",X"17",X"74",X"44",X"57",X"00",X"FF",X"00",X"3E",X"E4",X"44",X"4E",X"00",X"FF",
		X"00",X"08",X"82",X"66",X"60",X"00",X"0F",X"00",X"00",X"00",X"80",X"01",X"20",X"FF",X"00",X"00",
		X"32",X"92",X"23",X"28",X"FF",X"08",X"08",X"32",X"23",X"31",X"80",X"0F",X"00",X"88",X"22",X"33",
		X"98",X"80",X"0F",X"00",X"08",X"33",X"29",X"98",X"00",X"FF",X"00",X"00",X"88",X"99",X"30",X"00",
		X"0F",X"00",X"00",X"06",X"0D",X"00",X"00",X"FF",X"00",X"05",X"56",X"D5",X"56",X"00",X"FF",X"08",
		X"02",X"23",X"00",X"00",X"00",X"FF",X"08",X"12",X"22",X"38",X"00",X"00",X"FF",X"29",X"22",X"AB",
		X"3A",X"B0",X"00",X"FF",X"32",X"88",X"BD",X"8B",X"D0",X"00",X"FF",X"38",X"88",X"BD",X"8B",X"D0",
		X"00",X"FF",X"33",X"88",X"AA",X"8A",X"A0",X"00",X"FF",X"81",X"77",X"44",X"45",X"70",X"00",X"FF",
		X"03",X"EE",X"44",X"44",X"E0",X"88",X"FF",X"00",X"88",X"26",X"66",X"D8",X"80",X"FF",X"00",X"00",
		X"80",X"02",X"18",X"80",X"FF",X"00",X"32",X"11",X"21",X"28",X"00",X"FF",X"08",X"31",X"13",X"32",
		X"80",X"00",X"FF",X"88",X"22",X"33",X"98",X"80",X"00",X"FF",X"08",X"33",X"29",X"98",X"00",X"00",
		X"FF",X"00",X"88",X"99",X"36",X"60",X"00",X"FF",X"00",X"06",X"00",X"00",X"00",X"00",X"FF",X"05",
		X"56",X"D0",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"23",X"00",X"30",X"FF",X"00",X"02",X"21",
		X"12",X"33",X"00",X"FF",X"00",X"32",X"99",X"29",X"93",X"30",X"FF",X"00",X"38",X"AA",X"8A",X"A8",
		X"30",X"FF",X"00",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"00",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",
		X"00",X"77",X"24",X"44",X"27",X"70",X"FF",X"00",X"7E",X"44",X"45",X"47",X"E0",X"FF",X"00",X"02",
		X"35",X"56",X"32",X"00",X"FF",X"00",X"00",X"00",X"30",X"00",X"00",X"FF",X"03",X"33",X"33",X"13",
		X"33",X"33",X"FF",X"00",X"33",X"31",X"91",X"33",X"30",X"FF",X"00",X"03",X"19",X"A9",X"13",X"00",
		X"FF",X"00",X"00",X"19",X"A9",X"10",X"00",X"FF",X"00",X"00",X"21",X"91",X"20",X"00",X"FF",X"00",
		X"00",X"02",X"33",X"30",X"00",X"FF",X"00",X"00",X"06",X"00",X"60",X"00",X"FF",X"00",X"05",X"56",
		X"00",X"56",X"D0",X"FF",X"00",X"00",X"02",X"23",X"00",X"30",X"FF",X"00",X"02",X"21",X"12",X"33",
		X"00",X"FF",X"00",X"32",X"99",X"29",X"93",X"30",X"FF",X"00",X"38",X"AA",X"8A",X"A8",X"30",X"FF",
		X"00",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"00",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",X"00",X"77",
		X"24",X"44",X"27",X"70",X"FF",X"00",X"7E",X"44",X"45",X"47",X"E0",X"FF",X"00",X"00",X"85",X"55",
		X"22",X"38",X"FF",X"83",X"33",X"31",X"23",X"33",X"80",X"FF",X"08",X"33",X"19",X"92",X"38",X"00",
		X"FF",X"00",X"81",X"9A",X"99",X"30",X"00",X"FF",X"00",X"01",X"9A",X"91",X"20",X"00",X"FF",X"00",
		X"03",X"19",X"12",X"30",X"00",X"FF",X"00",X"00",X"33",X"33",X"00",X"00",X"FF",X"00",X"00",X"60",
		X"06",X"00",X"00",X"FF",X"00",X"55",X"60",X"05",X"6D",X"00",X"FF",X"00",X"00",X"02",X"23",X"00",
		X"30",X"FF",X"00",X"02",X"21",X"12",X"33",X"00",X"FF",X"00",X"32",X"99",X"29",X"93",X"30",X"FF",
		X"00",X"38",X"AA",X"8A",X"A8",X"30",X"FF",X"00",X"88",X"AD",X"8D",X"A8",X"80",X"FF",X"00",X"D8",
		X"AD",X"8D",X"A8",X"D0",X"FF",X"00",X"77",X"24",X"44",X"27",X"70",X"FF",X"00",X"7E",X"44",X"45",
		X"47",X"E0",X"FF",X"00",X"02",X"35",X"56",X"32",X"00",X"FF",X"00",X"00",X"00",X"30",X"00",X"00",
		X"FF",X"03",X"33",X"33",X"13",X"33",X"33",X"FF",X"00",X"33",X"31",X"91",X"33",X"30",X"FF",X"00",
		X"03",X"19",X"A9",X"13",X"00",X"FF",X"00",X"00",X"19",X"A9",X"10",X"D0",X"FF",X"00",X"00",X"21",
		X"91",X"20",X"60",X"FF",X"00",X"00",X"02",X"33",X"D6",X"50",X"FF",X"00",X"00",X"06",X"00",X"00",
		X"60",X"FF",X"00",X"05",X"56",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"02",X"23",X"00",X"30",X"FF",X"00",X"02",X"21",X"12",X"33",X"00",X"FF",X"00",X"32",
		X"22",X"22",X"23",X"30",X"FF",X"00",X"38",X"AA",X"8A",X"A8",X"30",X"FF",X"00",X"88",X"AB",X"8B",
		X"A8",X"80",X"FF",X"00",X"D8",X"AD",X"8D",X"A8",X"D0",X"FF",X"00",X"77",X"24",X"44",X"27",X"70",
		X"FF",X"00",X"7E",X"43",X"43",X"47",X"E0",X"FF",X"00",X"02",X"33",X"53",X"32",X"00",X"FF",X"00",
		X"00",X"33",X"33",X"33",X"00",X"FF",X"00",X"03",X"33",X"13",X"33",X"30",X"FF",X"00",X"03",X"33",
		X"91",X"33",X"30",X"FF",X"00",X"02",X"39",X"A9",X"12",X"00",X"FF",X"00",X"00",X"29",X"A9",X"10",
		X"00",X"FF",X"00",X"00",X"22",X"22",X"20",X"00",X"FF",X"00",X"06",X"00",X"00",X"60",X"00",X"FF",
		X"66",X"60",X"00",X"06",X"66",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"02",X"23",X"08",X"00",X"FF",X"02",X"21",X"12",X"38",X"00",X"FF",X"32",
		X"22",X"22",X"23",X"30",X"FF",X"32",X"22",X"22",X"22",X"30",X"FF",X"32",X"22",X"32",X"23",X"30",
		X"FF",X"D8",X"AA",X"8A",X"A8",X"D0",X"FF",X"78",X"CD",X"8D",X"C8",X"70",X"FF",X"77",X"24",X"44",
		X"27",X"70",X"FF",X"08",X"64",X"44",X"68",X"00",X"FF",X"03",X"86",X"56",X"83",X"00",X"FF",X"33",
		X"1A",X"A9",X"13",X"30",X"FF",X"33",X"19",X"A9",X"13",X"30",X"FF",X"03",X"21",X"91",X"23",X"00",
		X"FF",X"00",X"32",X"33",X"30",X"00",X"FF",X"00",X"06",X"06",X"00",X"00",X"FF",X"04",X"56",X"86",
		X"55",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"03",X"33",X"00",X"00",X"FF",X"00",X"03",X"21",
		X"12",X"33",X"00",X"FF",X"80",X"32",X"19",X"91",X"23",X"30",X"8F",X"08",X"32",X"19",X"11",X"23",
		X"38",X"8F",X"08",X"32",X"21",X"12",X"23",X"38",X"FF",X"08",X"33",X"22",X"22",X"23",X"38",X"FF",
		X"08",X"83",X"32",X"22",X"33",X"80",X"FF",X"00",X"88",X"33",X"33",X"38",X"80",X"FF",X"00",X"08",
		X"65",X"45",X"68",X"00",X"FF",X"00",X"03",X"26",X"56",X"23",X"00",X"FF",X"00",X"00",X"19",X"99",
		X"10",X"00",X"FF",X"00",X"00",X"06",X"06",X"00",X"00",X"FF",X"00",X"04",X"56",X"86",X"55",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"FF",X"00",X"55",X"D5",X"34",X"D5",X"30",X"00",X"FF",
		X"00",X"4D",X"DD",X"2D",X"DD",X"20",X"00",X"FF",X"04",X"48",X"81",X"21",X"88",X"22",X"00",X"FF",
		X"05",X"55",X"55",X"45",X"55",X"32",X"00",X"FF",X"5E",X"E4",X"54",X"34",X"53",X"33",X"20",X"FF",
		X"54",X"43",X"33",X"33",X"33",X"33",X"20",X"FF",X"44",X"2E",X"E2",X"22",X"EE",X"2A",X"32",X"FF",
		X"42",X"E1",X"EE",X"7E",X"E1",X"E2",X"AA",X"FF",X"BB",X"77",X"17",X"77",X"17",X"7C",X"CB",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"CC",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"7C",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",X"FF",X"11",X"22",X"99",X"99",X"22",X"11",X"1C",X"FF",
		X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"FF",X"00",X"55",X"D5",X"34",X"D5",X"30",X"00",X"FF",
		X"00",X"4D",X"DD",X"2D",X"DD",X"20",X"00",X"FF",X"04",X"48",X"81",X"21",X"88",X"22",X"00",X"FF",
		X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"FF",X"00",X"55",X"D5",X"34",X"D5",X"30",X"00",X"FF",
		X"00",X"4D",X"DD",X"2D",X"DD",X"20",X"00",X"FF",X"04",X"48",X"81",X"21",X"88",X"22",X"00",X"FF",
		X"05",X"55",X"55",X"45",X"55",X"32",X"00",X"FF",X"5E",X"E4",X"54",X"34",X"53",X"33",X"20",X"FF",
		X"54",X"43",X"33",X"33",X"33",X"33",X"20",X"FF",X"44",X"2E",X"E2",X"22",X"EE",X"2A",X"32",X"FF",
		X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"FF",X"00",X"55",X"D5",X"34",X"D5",X"30",X"00",X"FF",
		X"00",X"4D",X"DD",X"2D",X"DD",X"20",X"00",X"FF",X"04",X"48",X"81",X"21",X"88",X"22",X"00",X"FF",
		X"05",X"55",X"55",X"45",X"55",X"32",X"00",X"FF",X"5E",X"E4",X"54",X"34",X"53",X"33",X"20",X"FF",
		X"54",X"43",X"33",X"33",X"33",X"33",X"20",X"FF",X"44",X"2E",X"E2",X"22",X"EE",X"2A",X"32",X"FF",
		X"42",X"E1",X"EE",X"7E",X"E1",X"E2",X"AA",X"FF",X"BB",X"77",X"17",X"77",X"17",X"7C",X"CB",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"CC",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"7C",X"FF",
		X"00",X"55",X"D5",X"34",X"D5",X"30",X"00",X"FF",X"00",X"4D",X"DD",X"2D",X"DD",X"20",X"00",X"FF",
		X"04",X"48",X"81",X"21",X"88",X"22",X"00",X"FF",X"05",X"55",X"55",X"45",X"55",X"32",X"00",X"FF",
		X"5E",X"E4",X"54",X"34",X"53",X"33",X"20",X"FF",X"54",X"43",X"33",X"33",X"33",X"33",X"20",X"FF",
		X"44",X"2E",X"E2",X"22",X"EE",X"2A",X"32",X"FF",X"42",X"E1",X"EE",X"7E",X"E1",X"E2",X"AA",X"FF",
		X"BB",X"77",X"17",X"77",X"17",X"7C",X"CB",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"CC",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"7C",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",X"FF",
		X"11",X"22",X"99",X"99",X"22",X"11",X"1C",X"FF",X"C7",X"77",X"EE",X"8E",X"77",X"77",X"7B",X"FF",
		X"00",X"00",X"00",X"55",X"50",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"5D",X"53",X"4D",
		X"53",X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"D2",X"DD",X"D2",X"00",X"00",X"FF",X"00",X"00",
		X"44",X"88",X"12",X"18",X"82",X"20",X"00",X"FF",X"00",X"00",X"55",X"55",X"54",X"55",X"53",X"20",
		X"00",X"FF",X"00",X"05",X"EE",X"45",X"43",X"45",X"33",X"32",X"00",X"FF",X"00",X"05",X"44",X"33",
		X"33",X"33",X"33",X"32",X"00",X"FF",X"00",X"54",X"42",X"EE",X"22",X"2E",X"E2",X"A3",X"20",X"FF",
		X"00",X"44",X"2E",X"1E",X"E7",X"EE",X"1E",X"2A",X"A0",X"FF",X"0A",X"3B",X"B7",X"71",X"77",X"71",
		X"77",X"CC",X"BA",X"FF",X"03",X"B7",X"77",X"77",X"77",X"77",X"77",X"7C",X"CB",X"FF",X"0B",X"C7",
		X"77",X"77",X"77",X"77",X"77",X"77",X"CB",X"FF",X"0B",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"CB",X"FF",X"0B",X"C1",X"12",X"29",X"99",X"92",X"21",X"11",X"CB",X"FF",X"0B",X"BC",X"77",X"7E",
		X"E8",X"E7",X"77",X"77",X"BA",X"FF",X"02",X"BB",X"E7",X"77",X"AA",X"A7",X"77",X"EB",X"A0",X"FF",
		X"0D",X"44",X"BB",X"BC",X"77",X"7C",X"CB",X"AA",X"20",X"FF",X"02",X"22",X"AA",X"BB",X"EE",X"7B",
		X"BA",X"A2",X"30",X"FF",X"00",X"03",X"43",X"3A",X"AA",X"AE",X"26",X"26",X"20",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"20",
		X"00",X"FF",X"00",X"00",X"00",X"55",X"50",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"5D",
		X"53",X"4D",X"53",X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"D2",X"DD",X"D2",X"00",X"00",X"FF",
		X"00",X"00",X"44",X"DD",X"D2",X"DD",X"D2",X"20",X"00",X"FF",X"00",X"00",X"55",X"67",X"64",X"57",
		X"63",X"20",X"00",X"FF",X"00",X"05",X"6E",X"76",X"43",X"45",X"54",X"32",X"00",X"FF",X"00",X"05",
		X"64",X"33",X"33",X"33",X"34",X"42",X"00",X"FF",X"00",X"54",X"42",X"EE",X"32",X"3E",X"E2",X"A3",
		X"20",X"FF",X"00",X"44",X"2E",X"11",X"E7",X"E1",X"1E",X"2A",X"A0",X"FF",X"0A",X"3B",X"B7",X"7C",
		X"77",X"7C",X"77",X"CC",X"BA",X"FF",X"03",X"B7",X"77",X"77",X"77",X"77",X"77",X"7C",X"CB",X"FF",
		X"0B",X"C7",X"7E",X"EE",X"EE",X"EE",X"EE",X"77",X"CB",X"FF",X"0B",X"C1",X"DD",X"8D",X"88",X"D8",
		X"8D",X"D1",X"CB",X"FF",X"0B",X"C1",X"12",X"99",X"99",X"99",X"21",X"11",X"CB",X"FF",X"0B",X"CC",
		X"7E",X"EE",X"E8",X"E7",X"77",X"77",X"CA",X"FF",X"00",X"BC",X"CE",X"E7",X"AA",X"A7",X"77",X"CB",
		X"A0",X"FF",X"02",X"2A",X"BC",X"C7",X"77",X"77",X"CC",X"AA",X"20",X"FF",X"0D",X"45",X"AA",X"BC",
		X"EE",X"7C",X"BA",X"A2",X"30",X"FF",X"02",X"22",X"42",X"AA",X"AA",X"AA",X"22",X"44",X"40",X"FF",
		X"0D",X"45",X"65",X"55",X"43",X"45",X"55",X"66",X"70",X"FF",X"00",X"22",X"E7",X"76",X"55",X"56",
		X"67",X"7E",X"E0",X"FF",X"00",X"0E",X"EE",X"77",X"65",X"64",X"24",X"24",X"20",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"20",
		X"00",X"FF",X"00",X"00",X"00",X"55",X"50",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"5D",
		X"53",X"4D",X"53",X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"D2",X"DD",X"D2",X"00",X"00",X"FF",
		X"00",X"00",X"44",X"DD",X"D2",X"DD",X"D2",X"20",X"00",X"FF",X"00",X"00",X"55",X"67",X"64",X"57",
		X"63",X"20",X"00",X"FF",X"00",X"05",X"6E",X"44",X"43",X"45",X"54",X"32",X"00",X"FF",X"00",X"05",
		X"63",X"EE",X"23",X"2E",X"E3",X"42",X"00",X"FF",X"00",X"54",X"4E",X"11",X"E2",X"E1",X"1E",X"A3",
		X"20",X"FF",X"00",X"4B",X"7E",X"E7",X"77",X"77",X"77",X"CB",X"A0",X"FF",X"0A",X"B7",X"E7",X"7C",
		X"CC",X"77",X"77",X"7C",X"BA",X"FF",X"03",X"CE",X"7D",X"88",X"88",X"CC",X"CC",X"7C",X"CB",X"FF",
		X"0B",X"C7",X"D8",X"88",X"D8",X"D8",X"8D",X"C7",X"CB",X"FF",X"0B",X"7D",X"D1",X"12",X"22",X"22",
		X"11",X"DD",X"CB",X"FF",X"0B",X"C1",X"12",X"99",X"99",X"99",X"21",X"11",X"CB",X"FF",X"0B",X"CC",
		X"ED",X"DD",X"DD",X"DD",X"DD",X"E7",X"CA",X"FF",X"07",X"B7",X"EE",X"EE",X"EE",X"EE",X"EE",X"CB",
		X"A0",X"FF",X"02",X"2A",X"BE",X"77",X"AA",X"A7",X"CC",X"AA",X"20",X"FF",X"05",X"53",X"AA",X"C7",
		X"77",X"77",X"CA",X"A2",X"40",X"FF",X"02",X"22",X"55",X"AA",X"EE",X"EA",X"34",X"45",X"50",X"FF",
		X"04",X"76",X"66",X"55",X"43",X"45",X"55",X"66",X"70",X"FF",X"00",X"22",X"E7",X"76",X"55",X"56",
		X"67",X"7E",X"E0",X"FF",X"00",X"0E",X"EE",X"77",X"65",X"66",X"7E",X"EE",X"E0",X"FF",X"00",X"01",
		X"EE",X"77",X"65",X"67",X"EE",X"E1",X"E0",X"FF",X"00",X"0E",X"EE",X"76",X"55",X"54",X"24",X"24",
		X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"20",X"00",X"FF",X"00",X"00",X"00",X"55",X"50",X"55",X"50",X"00",X"00",X"FF",
		X"00",X"00",X"04",X"4D",X"43",X"4D",X"43",X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"D2",X"DD",
		X"D2",X"00",X"00",X"FF",X"00",X"00",X"44",X"88",X"12",X"88",X"12",X"20",X"00",X"FF",X"00",X"00",
		X"45",X"55",X"54",X"55",X"53",X"20",X"00",X"FF",X"00",X"04",X"55",X"EE",X"43",X"4E",X"E5",X"32",
		X"00",X"FF",X"00",X"05",X"5E",X"11",X"E3",X"E1",X"1E",X"42",X"00",X"FF",X"00",X"55",X"B7",X"77",
		X"77",X"77",X"77",X"B3",X"20",X"FF",X"00",X"AC",X"77",X"7C",X"CC",X"C7",X"77",X"CB",X"A0",X"FF",
		X"0B",X"C7",X"7C",X"C8",X"88",X"8C",X"C7",X"7C",X"BA",X"FF",X"0C",X"77",X"CD",X"88",X"88",X"88",
		X"8D",X"C7",X"CB",X"FF",X"0B",X"EC",X"DE",X"11",X"11",X"11",X"1D",X"8C",X"CB",X"FF",X"0E",X"7D",
		X"11",X"12",X"22",X"22",X"21",X"1D",X"CB",X"FF",X"07",X"71",X"12",X"99",X"99",X"99",X"22",X"11",
		X"CB",X"FF",X"0C",X"77",X"ED",X"D8",X"88",X"D8",X"DD",X"E7",X"CA",X"FF",X"00",X"B7",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"CB",X"A0",X"FF",X"00",X"66",X"BE",X"77",X"AA",X"A7",X"CC",X"AA",X"20",X"FF",
		X"00",X"22",X"AA",X"C7",X"77",X"77",X"CA",X"A2",X"40",X"FF",X"04",X"5E",X"55",X"AA",X"EE",X"EA",
		X"34",X"45",X"50",X"FF",X"02",X"22",X"66",X"55",X"43",X"45",X"55",X"66",X"70",X"FF",X"05",X"55",
		X"E7",X"76",X"55",X"56",X"67",X"7E",X"E0",X"FF",X"00",X"22",X"EE",X"77",X"65",X"66",X"7E",X"EE",
		X"E0",X"FF",X"00",X"01",X"EE",X"77",X"65",X"67",X"EE",X"E1",X"E0",X"FF",X"00",X"0E",X"EE",X"76",
		X"55",X"54",X"24",X"24",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"20",X"00",X"FF",X"00",X"00",X"00",X"55",X"50",X"55",
		X"50",X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"43",X"DD",X"43",X"00",X"00",X"FF",X"00",X"00",
		X"04",X"DD",X"D2",X"88",X"14",X"00",X"00",X"FF",X"00",X"00",X"34",X"88",X"12",X"88",X"14",X"30",
		X"00",X"FF",X"00",X"00",X"35",X"55",X"54",X"55",X"55",X"53",X"00",X"FF",X"00",X"03",X"5E",X"E3",
		X"43",X"EE",X"46",X"65",X"00",X"FF",X"00",X"03",X"E1",X"1E",X"4E",X"11",X"E4",X"55",X"30",X"FF",
		X"00",X"35",X"B7",X"77",X"77",X"77",X"7E",X"B4",X"40",X"FF",X"00",X"AC",X"7D",X"D8",X"88",X"87",
		X"7E",X"77",X"43",X"FF",X"0B",X"C7",X"D8",X"8D",X"8D",X"88",X"8C",X"C7",X"7A",X"FF",X"0C",X"7D",
		X"D8",X"11",X"11",X"1D",X"88",X"8C",X"7B",X"FF",X"0C",X"ED",X"D1",X"11",X"11",X"11",X"1D",X"88",
		X"7B",X"FF",X"0C",X"7D",X"11",X"22",X"12",X"22",X"11",X"1D",X"7B",X"FF",X"0C",X"71",X"12",X"99",
		X"22",X"99",X"21",X"11",X"CB",X"FF",X"0C",X"C7",X"29",X"99",X"99",X"99",X"9D",X"E7",X"7A",X"FF",
		X"00",X"77",X"7E",X"D8",X"88",X"8D",X"DE",X"77",X"A0",X"FF",X"00",X"07",X"77",X"EE",X"EE",X"EE",
		X"77",X"7A",X"20",X"FF",X"00",X"34",X"77",X"77",X"BA",X"B7",X"77",X"A2",X"40",X"FF",X"00",X"22",
		X"24",X"7E",X"EE",X"77",X"74",X"45",X"50",X"FF",X"04",X"57",X"76",X"5E",X"EE",X"E5",X"55",X"66",
		X"70",X"FF",X"02",X"22",X"27",X"76",X"55",X"56",X"67",X"7E",X"E0",X"FF",X"00",X"45",X"5E",X"77",
		X"65",X"66",X"7E",X"EE",X"E0",X"FF",X"00",X"22",X"2E",X"77",X"65",X"67",X"EE",X"E1",X"E0",X"FF",
		X"00",X"0E",X"EE",X"76",X"55",X"54",X"24",X"24",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"20",X"00",X"FF",X"00",X"00",
		X"00",X"55",X"40",X"45",X"50",X"00",X"00",X"FF",X"00",X"00",X"04",X"4D",X"43",X"4D",X"43",X"00",
		X"00",X"FF",X"00",X"00",X"34",X"DD",X"D2",X"DD",X"D2",X"00",X"00",X"FF",X"00",X"03",X"44",X"88",
		X"12",X"88",X"12",X"00",X"00",X"FF",X"00",X"04",X"55",X"55",X"54",X"35",X"53",X"20",X"00",X"FF",
		X"00",X"35",X"7E",X"77",X"55",X"35",X"54",X"32",X"00",X"FF",X"00",X"47",X"E6",X"55",X"5E",X"E2",
		X"54",X"EE",X"00",X"FF",X"03",X"37",X"65",X"BB",X"71",X"17",X"BE",X"11",X"E0",X"FF",X"03",X"56",
		X"5B",X"BE",X"E7",X"77",X"77",X"CB",X"A0",X"FF",X"03",X"55",X"BB",X"7E",X"E7",X"77",X"77",X"7C",
		X"BA",X"FF",X"05",X"5B",X"B7",X"E7",X"77",X"D8",X"88",X"DD",X"D3",X"FF",X"04",X"5B",X"7E",X"77",
		X"DD",X"21",X"11",X"11",X"D3",X"FF",X"05",X"BC",X"E7",X"CD",X"99",X"22",X"21",X"11",X"1D",X"FF",
		X"03",X"BC",X"EE",X"D9",X"99",X"99",X"92",X"21",X"D3",X"FF",X"03",X"3C",X"77",X"ED",X"DD",X"DD",
		X"DD",X"DD",X"DA",X"FF",X"00",X"3B",X"C7",X"7E",X"EE",X"EE",X"EE",X"77",X"A0",X"FF",X"00",X"2A",
		X"BC",X"C7",X"7C",X"CA",X"AA",X"AA",X"30",X"FF",X"04",X"77",X"AA",X"BC",X"C7",X"77",X"7B",X"23",
		X"00",X"FF",X"02",X"22",X"55",X"AB",X"BC",X"CE",X"EB",X"34",X"00",X"FF",X"47",X"77",X"66",X"55",
		X"43",X"43",X"35",X"55",X"00",X"FF",X"22",X"22",X"E7",X"76",X"55",X"56",X"66",X"67",X"00",X"FF",
		X"04",X"77",X"EE",X"77",X"65",X"66",X"67",X"7E",X"00",X"FF",X"02",X"22",X"EE",X"77",X"65",X"66",
		X"7E",X"E1",X"00",X"FF",X"00",X"EE",X"EE",X"76",X"55",X"E2",X"52",X"52",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"D2",X"42",X"D2",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"D2",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"04",X"57",X"40",X"45",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"45",X"77",X"76",X"47",X"73",X"00",X"00",X"FF",X"00",X"00",X"04",X"57",X"5D",X"D6",X"4D",X"D5",
		X"00",X"00",X"FF",X"00",X"00",X"35",X"54",X"88",X"16",X"48",X"81",X"00",X"00",X"FF",X"00",X"03",
		X"45",X"44",X"55",X"54",X"35",X"53",X"20",X"00",X"FF",X"00",X"05",X"55",X"7E",X"77",X"55",X"35",
		X"54",X"32",X"00",X"FF",X"00",X"35",X"57",X"EE",X"75",X"5E",X"EE",X"E4",X"EE",X"00",X"FF",X"00",
		X"56",X"67",X"77",X"53",X"35",X"11",X"E3",X"61",X"B0",X"FF",X"03",X"56",X"67",X"55",X"3C",X"C7",
		X"77",X"77",X"CB",X"A0",X"FF",X"04",X"55",X"66",X"63",X"CE",X"EE",X"77",X"77",X"7C",X"BA",X"FF",
		X"05",X"75",X"66",X"3C",X"EE",X"EE",X"77",X"77",X"EE",X"E3",X"FF",X"06",X"77",X"55",X"3E",X"EE",
		X"88",X"E7",X"7E",X"88",X"B2",X"FF",X"06",X"75",X"54",X"C7",X"EE",X"88",X"E7",X"E2",X"11",X"14",
		X"FF",X"05",X"54",X"54",X"CE",X"7E",X"EE",X"77",X"E9",X"91",X"D2",X"FF",X"05",X"54",X"43",X"3C",
		X"E7",X"77",X"7C",X"77",X"EE",X"EA",X"FF",X"04",X"53",X"33",X"33",X"CC",X"CC",X"CE",X"EE",X"77",
		X"A0",X"FF",X"65",X"E5",X"45",X"54",X"33",X"CC",X"EE",X"7C",X"00",X"00",X"FF",X"22",X"26",X"66",
		X"55",X"43",X"22",X"EE",X"C0",X"00",X"00",X"FF",X"66",X"77",X"77",X"65",X"43",X"43",X"33",X"40",
		X"00",X"00",X"FF",X"22",X"2E",X"E7",X"76",X"55",X"55",X"55",X"40",X"00",X"00",X"FF",X"44",X"EE",
		X"EE",X"76",X"55",X"66",X"66",X"60",X"00",X"00",X"FF",X"22",X"E1",X"EE",X"76",X"55",X"77",X"7E",
		X"E0",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"77",X"57",X"25",X"25",X"20",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"04",X"24",X"24",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"35",X"77",X"42",X"45",X"30",X"00",X"00",
		X"FF",X"00",X"00",X"02",X"34",X"77",X"77",X"74",X"47",X"70",X"00",X"00",X"FF",X"00",X"00",X"23",
		X"45",X"77",X"66",X"77",X"47",X"70",X"00",X"00",X"FF",X"00",X"02",X"43",X"55",X"76",X"44",X"11",
		X"76",X"10",X"00",X"00",X"FF",X"00",X"04",X"43",X"56",X"66",X"66",X"77",X"15",X"12",X"20",X"00",
		X"FF",X"00",X"34",X"54",X"56",X"65",X"54",X"46",X"77",X"54",X"32",X"00",X"FF",X"03",X"34",X"56",
		X"55",X"55",X"77",X"6E",X"54",X"EE",X"4E",X"E0",X"FF",X"03",X"47",X"67",X"76",X"57",X"45",X"55",
		X"4E",X"E1",X"E6",X"B0",X"FF",X"04",X"57",X"EE",X"75",X"54",X"5B",X"C7",X"77",X"77",X"5B",X"A0",
		X"FF",X"04",X"36",X"EE",X"65",X"4A",X"B7",X"EE",X"EE",X"77",X"77",X"BA",X"FF",X"05",X"35",X"66",
		X"55",X"AB",X"C7",X"E8",X"8E",X"E7",X"77",X"EE",X"FF",X"05",X"43",X"55",X"54",X"AC",X"77",X"E8",
		X"8E",X"EE",X"7E",X"12",X"FF",X"06",X"54",X"35",X"54",X"AA",X"C7",X"EE",X"EE",X"8E",X"E1",X"91",
		X"FF",X"45",X"E5",X"43",X"33",X"33",X"CC",X"77",X"7E",X"E7",X"7E",X"12",X"FF",X"22",X"22",X"44",
		X"33",X"43",X"3C",X"CC",X"CC",X"7B",X"77",X"EE",X"FF",X"45",X"E6",X"65",X"44",X"33",X"33",X"3B",
		X"BB",X"BB",X"BB",X"A0",X"FF",X"22",X"2E",X"E5",X"55",X"53",X"44",X"33",X"20",X"00",X"00",X"00",
		X"FF",X"45",X"EE",X"E7",X"76",X"35",X"53",X"55",X"40",X"00",X"00",X"00",X"FF",X"22",X"EE",X"EE",
		X"76",X"55",X"66",X"56",X"60",X"00",X"00",X"00",X"FF",X"0E",X"E1",X"EE",X"76",X"56",X"77",X"7E",
		X"E0",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"75",X"62",X"52",X"42",X"E0",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"02",X"42",X"42",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"D2",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"50",X"55",X"50",
		X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"43",X"DD",X"43",X"00",X"00",X"FF",X"00",X"00",X"04",
		X"81",X"82",X"81",X"84",X"00",X"00",X"FF",X"00",X"00",X"34",X"44",X"42",X"44",X"44",X"30",X"00",
		X"FF",X"00",X"00",X"35",X"EE",X"54",X"5E",X"E5",X"53",X"00",X"FF",X"00",X"03",X"5E",X"11",X"E3",
		X"E1",X"1E",X"65",X"00",X"FF",X"00",X"03",X"47",X"77",X"77",X"77",X"E4",X"55",X"30",X"FF",X"00",
		X"34",X"78",X"88",X"88",X"77",X"7E",X"B4",X"40",X"FF",X"00",X"47",X"D8",X"D8",X"8D",X"88",X"7E",
		X"77",X"43",X"FF",X"0B",X"C7",X"D8",X"11",X"11",X"18",X"8C",X"C7",X"7A",X"FF",X"0C",X"7D",X"D1",
		X"11",X"11",X"11",X"18",X"DC",X"7B",X"FF",X"0C",X"ED",X"11",X"11",X"11",X"11",X"11",X"DD",X"7B",
		X"FF",X"0C",X"7D",X"11",X"22",X"12",X"22",X"11",X"1D",X"7B",X"FF",X"0C",X"71",X"12",X"99",X"99",
		X"99",X"21",X"11",X"CB",X"FF",X"03",X"C7",X"EE",X"EE",X"EE",X"EE",X"EE",X"E7",X"7A",X"FF",X"00",
		X"37",X"77",X"7C",X"AA",X"BC",X"77",X"77",X"A0",X"FF",X"00",X"55",X"77",X"7E",X"EE",X"E7",X"77",
		X"A2",X"40",X"FF",X"00",X"22",X"44",X"7E",X"EE",X"77",X"74",X"45",X"50",X"FF",X"03",X"66",X"E6",
		X"54",X"44",X"45",X"55",X"66",X"70",X"FF",X"02",X"22",X"27",X"76",X"55",X"56",X"67",X"7E",X"E0",
		X"FF",X"00",X"35",X"5E",X"77",X"65",X"66",X"7E",X"EE",X"E0",X"FF",X"00",X"22",X"2E",X"77",X"65",
		X"67",X"EE",X"E1",X"E0",X"FF",X"00",X"0E",X"EE",X"76",X"55",X"54",X"24",X"24",X"20",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"20",X"00",X"FF",X"00",X"00",X"00",X"33",X"30",X"33",X"20",X"00",X"00",X"FF",X"00",X"00",X"0B",
		X"CC",X"33",X"3C",X"CB",X"00",X"00",X"FF",X"00",X"00",X"2C",X"17",X"74",X"77",X"1C",X"20",X"00",
		X"FF",X"00",X"00",X"27",X"7E",X"EE",X"EE",X"77",X"30",X"00",X"FF",X"00",X"02",X"77",X"EB",X"BB",
		X"BB",X"E7",X"73",X"00",X"FF",X"00",X"02",X"7E",X"B8",X"D8",X"D8",X"BE",X"73",X"00",X"FF",X"00",
		X"57",X"EB",X"D8",X"D8",X"D8",X"DB",X"E7",X"40",X"FF",X"00",X"77",X"EB",X"D1",X"11",X"11",X"DB",
		X"E7",X"50",X"FF",X"07",X"8E",X"BD",X"11",X"22",X"21",X"1D",X"EE",X"E5",X"FF",X"07",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"87",X"FF",X"05",X"EE",X"E7",X"77",X"BA",X"B7",X"77",X"77",X"E7",
		X"FF",X"0A",X"C7",X"77",X"77",X"77",X"77",X"77",X"77",X"7C",X"FF",X"0A",X"BC",X"77",X"CA",X"AA",
		X"AA",X"AC",X"77",X"CB",X"FF",X"00",X"AB",X"7C",X"AB",X"BB",X"BA",X"AA",X"C7",X"C0",X"FF",X"00",
		X"AA",X"BC",X"AB",X"BB",X"BB",X"AA",X"CC",X"C0",X"FF",X"00",X"0A",X"BA",X"AB",X"BB",X"BB",X"AA",
		X"AC",X"20",X"FF",X"00",X"03",X"AA",X"BB",X"BB",X"BB",X"B4",X"AA",X"20",X"FF",X"00",X"03",X"A4",
		X"4B",X"BB",X"B4",X"44",X"A2",X"40",X"FF",X"00",X"05",X"44",X"44",X"44",X"44",X"44",X"45",X"50",
		X"FF",X"00",X"22",X"26",X"54",X"44",X"45",X"55",X"66",X"70",X"FF",X"05",X"55",X"57",X"76",X"55",
		X"56",X"67",X"7E",X"E0",X"FF",X"02",X"22",X"2E",X"77",X"65",X"66",X"7E",X"EE",X"E0",X"FF",X"00",
		X"45",X"5E",X"77",X"65",X"67",X"EE",X"E1",X"E0",X"FF",X"00",X"22",X"2E",X"76",X"55",X"54",X"24",
		X"24",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"20",X"00",X"FF",X"00",X"00",X"03",X"3E",X"EE",X"32",X"00",X"00",X"FF",
		X"00",X"00",X"BC",X"E1",X"11",X"EC",X"B0",X"00",X"FF",X"00",X"0E",X"E7",X"1D",X"DD",X"17",X"CC",
		X"00",X"FF",X"00",X"E8",X"E7",X"77",X"77",X"77",X"EC",X"C0",X"FF",X"00",X"EE",X"77",X"EE",X"EE",
		X"77",X"EE",X"E0",X"FF",X"00",X"77",X"77",X"CB",X"BA",X"C7",X"77",X"E0",X"FF",X"05",X"77",X"7C",
		X"55",X"55",X"AC",X"77",X"7C",X"FF",X"07",X"77",X"7C",X"56",X"55",X"3C",X"C7",X"CC",X"FF",X"0C",
		X"77",X"7C",X"56",X"55",X"AB",X"BC",X"CC",X"FF",X"0C",X"77",X"CC",X"56",X"55",X"AA",X"BB",X"CC",
		X"FF",X"0C",X"CC",X"C5",X"66",X"55",X"AA",X"BB",X"BB",X"FF",X"0B",X"BB",X"B5",X"66",X"55",X"AA",
		X"BB",X"BB",X"FF",X"0B",X"BB",X"55",X"66",X"55",X"5A",X"AB",X"BB",X"FF",X"03",X"BB",X"56",X"66",
		X"55",X"5A",X"AB",X"BB",X"FF",X"02",X"A5",X"56",X"66",X"55",X"5A",X"3A",X"BB",X"FF",X"00",X"2A",
		X"5C",X"66",X"55",X"4A",X"AA",X"BB",X"FF",X"00",X"23",X"AA",X"C6",X"54",X"AA",X"AA",X"AB",X"FF",
		X"00",X"2A",X"AA",X"A6",X"4A",X"AA",X"AA",X"A3",X"FF",X"04",X"64",X"43",X"AA",X"AA",X"44",X"44",
		X"5A",X"FF",X"02",X"26",X"65",X"33",X"44",X"55",X"56",X"67",X"FF",X"35",X"5E",X"77",X"63",X"35",
		X"66",X"77",X"EE",X"FF",X"22",X"2E",X"E7",X"76",X"56",X"67",X"EE",X"EE",X"FF",X"04",X"5E",X"E7",
		X"76",X"56",X"7E",X"EE",X"1E",X"FF",X"02",X"2E",X"E7",X"65",X"55",X"42",X"42",X"42",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"D2",X"42",X"D2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"D2",X"00",
		X"FF",X"00",X"00",X"00",X"05",X"65",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"56",X"66",X"50",
		X"00",X"00",X"FF",X"00",X"00",X"66",X"66",X"66",X"66",X"60",X"00",X"FF",X"00",X"06",X"EE",X"66",
		X"76",X"6E",X"86",X"00",X"FF",X"00",X"6E",X"8E",X"7E",X"E7",X"7E",X"8E",X"60",X"FF",X"00",X"6E",
		X"EE",X"CE",X"EE",X"7E",X"EE",X"60",X"FF",X"00",X"77",X"77",X"CC",X"CC",X"7C",X"77",X"60",X"FF",
		X"00",X"76",X"7C",X"CB",X"54",X"CC",X"76",X"70",X"FF",X"0C",X"77",X"CC",X"C6",X"45",X"4C",X"C7",
		X"7C",X"FF",X"0C",X"CC",X"CC",X"C6",X"45",X"4C",X"CC",X"CC",X"FF",X"0C",X"CC",X"CC",X"66",X"45",
		X"4B",X"BC",X"CC",X"FF",X"0C",X"CC",X"CC",X"66",X"45",X"A4",X"BB",X"CC",X"FF",X"0C",X"CC",X"CC",
		X"66",X"45",X"A4",X"BB",X"BB",X"FF",X"0B",X"BB",X"BC",X"66",X"45",X"A4",X"BB",X"B3",X"FF",X"03",
		X"BB",X"C6",X"66",X"44",X"5A",X"43",X"32",X"FF",X"02",X"3B",X"66",X"66",X"44",X"5A",X"43",X"22",
		X"FF",X"02",X"3C",X"66",X"66",X"45",X"55",X"34",X"21",X"FF",X"00",X"24",X"CC",X"66",X"44",X"55",
		X"44",X"43",X"FF",X"00",X"14",X"44",X"C6",X"45",X"44",X"45",X"55",X"FF",X"00",X"26",X"55",X"4C",
		X"44",X"44",X"56",X"66",X"FF",X"00",X"76",X"66",X"54",X"44",X"55",X"67",X"77",X"FF",X"04",X"EE",
		X"75",X"64",X"45",X"56",X"77",X"EE",X"FF",X"42",X"EE",X"E7",X"65",X"55",X"67",X"EE",X"EE",X"FF",
		X"24",X"1E",X"E7",X"76",X"56",X"7E",X"EE",X"1E",X"FF",X"32",X"5E",X"EE",X"76",X"57",X"EE",X"EE",
		X"EE",X"FF",X"25",X"52",X"EE",X"75",X"57",X"42",X"42",X"42",X"FF",X"04",X"20",X"00",X"00",X"00",
		X"D2",X"42",X"D2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"D2",X"00",X"FF",X"00",X"00",X"00",
		X"55",X"50",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"55",X"53",X"45",X"53",X"00",X"00",
		X"FF",X"00",X"00",X"04",X"DD",X"52",X"58",X"82",X"00",X"00",X"FF",X"00",X"00",X"44",X"DD",X"D2",
		X"88",X"82",X"20",X"00",X"FF",X"00",X"00",X"43",X"38",X"13",X"18",X"83",X"20",X"00",X"FF",X"00",
		X"03",X"44",X"55",X"53",X"45",X"55",X"32",X"00",X"FF",X"00",X"35",X"54",X"32",X"25",X"52",X"23",
		X"44",X"30",X"FF",X"03",X"65",X"56",X"EE",X"62",X"6E",X"E5",X"45",X"54",X"FF",X"06",X"76",X"EE",
		X"11",X"E7",X"E1",X"1E",X"35",X"76",X"FF",X"05",X"6B",X"B7",X"31",X"77",X"71",X"37",X"CC",X"B5",
		X"FF",X"04",X"BC",X"77",X"77",X"77",X"77",X"77",X"7C",X"CB",X"FF",X"0B",X"77",X"CE",X"EE",X"EE",
		X"EE",X"EE",X"C7",X"76",X"FF",X"06",X"8E",X"6D",X"88",X"D8",X"88",X"D8",X"E6",X"8E",X"FF",X"06",
		X"EE",X"61",X"11",X"22",X"21",X"11",X"D6",X"76",X"FF",X"0B",X"77",X"C8",X"D2",X"99",X"92",X"D8",
		X"EC",X"BA",X"FF",X"00",X"BB",X"7E",X"E8",X"8D",X"88",X"EE",X"CB",X"A0",X"FF",X"00",X"2A",X"BB",
		X"BE",X"EE",X"EE",X"CB",X"AA",X"20",X"FF",X"04",X"42",X"AA",X"BB",X"77",X"7B",X"BA",X"A2",X"30",
		X"FF",X"02",X"22",X"22",X"AA",X"AA",X"AA",X"22",X"44",X"40",X"FF",X"00",X"46",X"65",X"55",X"43",
		X"45",X"55",X"66",X"50",X"FF",X"00",X"22",X"26",X"66",X"55",X"56",X"67",X"76",X"60",X"FF",X"00",
		X"0E",X"E7",X"76",X"65",X"66",X"7E",X"EE",X"E0",X"FF",X"00",X"01",X"EE",X"77",X"65",X"67",X"EE",
		X"E1",X"E0",X"FF",X"00",X"0E",X"E7",X"76",X"55",X"54",X"24",X"24",X"20",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"20",X"00",
		X"FF",X"00",X"00",X"00",X"55",X"50",X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"55",X"53",
		X"45",X"53",X"00",X"00",X"FF",X"00",X"00",X"04",X"DD",X"52",X"5D",X"D2",X"00",X"00",X"FF",X"00",
		X"00",X"44",X"DD",X"D2",X"DD",X"82",X"20",X"00",X"FF",X"00",X"00",X"43",X"38",X"13",X"18",X"83",
		X"20",X"00",X"FF",X"00",X"03",X"44",X"55",X"53",X"45",X"55",X"32",X"00",X"FF",X"00",X"35",X"54",
		X"32",X"25",X"52",X"23",X"44",X"30",X"FF",X"03",X"65",X"56",X"77",X"62",X"67",X"75",X"45",X"54",
		X"FF",X"06",X"76",X"7E",X"11",X"E7",X"E1",X"17",X"35",X"76",X"FF",X"05",X"6B",X"B7",X"31",X"77",
		X"71",X"37",X"BB",X"B5",X"FF",X"04",X"BC",X"77",X"77",X"77",X"77",X"77",X"77",X"CB",X"FF",X"0A",
		X"C7",X"EE",X"77",X"77",X"77",X"7E",X"E7",X"7C",X"FF",X"0B",X"CE",X"88",X"75",X"D8",X"D5",X"78",
		X"8E",X"7B",X"FF",X"0B",X"CE",X"8E",X"71",X"12",X"11",X"78",X"EE",X"7A",X"FF",X"0A",X"C7",X"EE",
		X"71",X"29",X"21",X"7E",X"E7",X"CA",X"FF",X"00",X"BB",X"77",X"75",X"88",X"D5",X"77",X"CC",X"A0",
		X"FF",X"00",X"2A",X"BB",X"B7",X"55",X"57",X"CB",X"AA",X"20",X"FF",X"05",X"76",X"AA",X"BB",X"77",
		X"7B",X"BA",X"A2",X"30",X"FF",X"02",X"22",X"25",X"AA",X"AA",X"AA",X"22",X"44",X"40",X"FF",X"00",
		X"76",X"65",X"55",X"43",X"45",X"55",X"66",X"50",X"FF",X"00",X"22",X"26",X"66",X"55",X"56",X"67",
		X"76",X"60",X"FF",X"00",X"07",X"77",X"76",X"65",X"66",X"7E",X"EE",X"E0",X"FF",X"00",X"01",X"EE",
		X"77",X"65",X"67",X"EE",X"E1",X"E0",X"FF",X"00",X"0E",X"EE",X"76",X"55",X"54",X"24",X"24",X"20",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"20",X"00",X"FF",X"00",X"00",X"00",X"03",X"33",X"34",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"04",X"43",X"44",X"43",X"43",X"00",X"00",X"FF",X"00",X"00",X"45",X"55",X"34",X"36",X"54",
		X"30",X"00",X"FF",X"00",X"00",X"45",X"DD",X"53",X"5D",X"84",X"30",X"00",X"FF",X"00",X"04",X"55",
		X"DD",X"D3",X"D8",X"85",X"43",X"00",X"FF",X"00",X"04",X"57",X"58",X"13",X"18",X"57",X"74",X"00",
		X"FF",X"00",X"44",X"47",X"55",X"53",X"55",X"67",X"44",X"30",X"FF",X"00",X"45",X"64",X"22",X"33",
		X"32",X"24",X"44",X"30",X"FF",X"04",X"66",X"56",X"65",X"32",X"35",X"65",X"55",X"43",X"FF",X"04",
		X"44",X"44",X"44",X"32",X"34",X"45",X"55",X"43",X"FF",X"03",X"4B",X"BB",X"EE",X"32",X"3E",X"E5",
		X"55",X"33",X"FF",X"04",X"BC",X"CE",X"11",X"E2",X"E1",X"1E",X"AA",X"3A",X"FF",X"0B",X"C7",X"77",
		X"A1",X"EB",X"E1",X"AE",X"BC",X"BA",X"FF",X"0B",X"7E",X"E7",X"77",X"77",X"77",X"77",X"EE",X"CB",
		X"FF",X"03",X"E8",X"EE",X"E7",X"CC",X"77",X"7E",X"E8",X"EC",X"FF",X"0B",X"3E",X"8E",X"6C",X"77",
		X"7C",X"7E",X"8E",X"EC",X"FF",X"00",X"3C",X"C6",X"57",X"E1",X"E7",X"C5",X"CC",X"C0",X"FF",X"04",
		X"63",X"3C",X"CE",X"11",X"1E",X"CC",X"C3",X"30",X"FF",X"02",X"22",X"43",X"AC",X"E1",X"EC",X"33",
		X"33",X"30",X"FF",X"00",X"44",X"65",X"55",X"43",X"43",X"33",X"33",X"30",X"FF",X"00",X"22",X"76",
		X"66",X"55",X"56",X"67",X"76",X"60",X"FF",X"00",X"0E",X"E7",X"76",X"65",X"66",X"7E",X"EE",X"E0",
		X"FF",X"00",X"01",X"EE",X"77",X"65",X"67",X"EE",X"E1",X"E0",X"FF",X"00",X"0E",X"E7",X"76",X"55",
		X"54",X"24",X"24",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"24",X"2D",X"20",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"20",X"00",X"FF",X"00",X"00",X"00",X"35",X"32",X"34",X"30",
		X"00",X"00",X"FF",X"00",X"00",X"03",X"55",X"53",X"44",X"43",X"00",X"00",X"FF",X"00",X"00",X"33",
		X"44",X"33",X"34",X"43",X"30",X"00",X"FF",X"00",X"00",X"34",X"55",X"43",X"45",X"54",X"30",X"00",
		X"FF",X"00",X"04",X"45",X"55",X"44",X"57",X"75",X"43",X"00",X"FF",X"00",X"03",X"56",X"66",X"52",
		X"7E",X"77",X"43",X"00",X"FF",X"00",X"04",X"56",X"E7",X"63",X"55",X"46",X"44",X"00",X"FF",X"00",
		X"34",X"66",X"DD",X"D4",X"58",X"86",X"54",X"30",X"FF",X"00",X"34",X"62",X"28",X"14",X"18",X"22",
		X"74",X"40",X"FF",X"00",X"44",X"67",X"44",X"44",X"44",X"47",X"55",X"40",X"FF",X"00",X"46",X"66",
		X"64",X"44",X"44",X"66",X"66",X"43",X"FF",X"00",X"36",X"63",X"33",X"23",X"23",X"33",X"66",X"43",
		X"FF",X"00",X"44",X"44",X"44",X"32",X"34",X"46",X"66",X"44",X"FF",X"03",X"4A",X"AA",X"77",X"32",
		X"37",X"7A",X"AA",X"AA",X"FF",X"04",X"BC",X"C7",X"E7",X"72",X"77",X"E7",X"BB",X"B3",X"FF",X"0B",
		X"C7",X"77",X"11",X"7B",X"71",X"17",X"CC",X"B3",X"FF",X"0C",X"77",X"77",X"A2",X"77",X"72",X"A7",
		X"77",X"77",X"FF",X"0C",X"77",X"77",X"E7",X"77",X"77",X"77",X"77",X"77",X"FF",X"0C",X"77",X"7E",
		X"E7",X"CC",X"77",X"7E",X"77",X"77",X"FF",X"0B",X"C7",X"EE",X"EC",X"77",X"7C",X"CE",X"E7",X"70",
		X"FF",X"00",X"43",X"CC",X"BE",X"EE",X"EE",X"CC",X"B3",X"30",X"FF",X"00",X"04",X"43",X"A1",X"EE",
		X"E1",X"33",X"33",X"30",X"FF",X"00",X"0E",X"65",X"55",X"11",X"14",X"24",X"24",X"20",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"26",X"2D",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"33",X"30",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"34",X"44",X"43",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"02",X"34",X"46",X"66",X"54",X"33",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"23",X"46",X"66",
		X"66",X"65",X"44",X"32",X"00",X"00",X"FF",X"00",X"00",X"02",X"34",X"66",X"88",X"76",X"55",X"55",
		X"44",X"20",X"00",X"FF",X"00",X"00",X"23",X"45",X"68",X"87",X"65",X"55",X"55",X"54",X"42",X"00",
		X"FF",X"00",X"00",X"24",X"55",X"77",X"76",X"55",X"55",X"55",X"55",X"43",X"00",X"FF",X"00",X"02",
		X"34",X"56",X"66",X"55",X"55",X"55",X"54",X"44",X"43",X"20",X"FF",X"00",X"02",X"34",X"66",X"66",
		X"55",X"55",X"54",X"44",X"44",X"44",X"30",X"FF",X"00",X"03",X"46",X"68",X"86",X"65",X"55",X"44",
		X"44",X"44",X"44",X"30",X"FF",X"00",X"23",X"46",X"88",X"66",X"55",X"54",X"44",X"43",X"33",X"33",
		X"32",X"FF",X"00",X"23",X"56",X"88",X"66",X"55",X"44",X"44",X"33",X"33",X"23",X"32",X"FF",X"00",
		X"23",X"58",X"86",X"65",X"55",X"44",X"43",X"33",X"22",X"23",X"22",X"FF",X"00",X"23",X"58",X"87",
		X"65",X"54",X"44",X"43",X"32",X"22",X"22",X"22",X"FF",X"00",X"23",X"58",X"87",X"65",X"54",X"44",
		X"33",X"32",X"22",X"22",X"22",X"FF",X"00",X"23",X"58",X"87",X"65",X"54",X"44",X"33",X"32",X"22",
		X"22",X"22",X"FF",X"00",X"23",X"56",X"87",X"65",X"54",X"44",X"33",X"32",X"22",X"24",X"22",X"FF",
		X"00",X"03",X"55",X"87",X"65",X"54",X"44",X"43",X"33",X"22",X"24",X"20",X"FF",X"00",X"02",X"35",
		X"67",X"66",X"55",X"44",X"43",X"33",X"32",X"42",X"20",X"FF",X"00",X"02",X"35",X"67",X"76",X"55",
		X"44",X"44",X"43",X"33",X"43",X"10",X"FF",X"00",X"00",X"34",X"56",X"77",X"65",X"54",X"44",X"44",
		X"44",X"32",X"00",X"FF",X"00",X"00",X"13",X"45",X"67",X"76",X"55",X"44",X"44",X"44",X"31",X"00",
		X"FF",X"00",X"00",X"03",X"44",X"56",X"76",X"55",X"55",X"44",X"43",X"20",X"00",X"FF",X"00",X"00",
		X"01",X"34",X"45",X"55",X"55",X"55",X"55",X"53",X"10",X"00",X"FF",X"00",X"00",X"00",X"13",X"44",
		X"45",X"55",X"55",X"55",X"32",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"33",X"44",X"44",X"44",
		X"33",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"12",X"33",X"33",X"33",X"21",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"13",X"33",X"32",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"01",X"22",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"64",X"10",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"34",X"60",
		X"00",X"00",X"54",X"30",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"56",X"00",X"00",X"00",X"65",
		X"44",X"32",X"00",X"00",X"FF",X"00",X"02",X"45",X"68",X"80",X"00",X"00",X"15",X"55",X"44",X"20",
		X"00",X"FF",X"00",X"34",X"56",X"88",X"00",X"60",X"00",X"01",X"55",X"54",X"42",X"00",X"FF",X"02",
		X"45",X"57",X"70",X"08",X"87",X"10",X"00",X"55",X"55",X"43",X"00",X"FF",X"03",X"45",X"66",X"00",
		X"88",X"75",X"50",X"00",X"14",X"44",X"43",X"20",X"FF",X"23",X"46",X"66",X"01",X"07",X"55",X"50",
		X"00",X"04",X"44",X"44",X"30",X"FF",X"34",X"06",X"80",X"06",X"65",X"51",X"00",X"00",X"01",X"44",
		X"44",X"30",X"FF",X"34",X"68",X"06",X"66",X"65",X"11",X"00",X"00",X"00",X"13",X"03",X"32",X"FF",
		X"30",X"00",X"66",X"88",X"61",X"10",X"50",X"00",X"00",X"01",X"20",X"32",X"FF",X"30",X"00",X"08",
		X"86",X"65",X"55",X"00",X"00",X"00",X"00",X"10",X"22",X"FF",X"00",X"05",X"68",X"86",X"65",X"00",
		X"04",X"00",X"00",X"00",X"01",X"22",X"FF",X"00",X"05",X"88",X"06",X"55",X"10",X"40",X"30",X"00",
		X"00",X"00",X"12",X"FF",X"00",X"05",X"88",X"06",X"55",X"41",X"44",X"31",X"02",X"20",X"00",X"12",
		X"FF",X"00",X"05",X"88",X"70",X"55",X"44",X"43",X"10",X"02",X"22",X"00",X"12",X"FF",X"00",X"00",
		X"80",X"00",X"05",X"44",X"43",X"00",X"12",X"20",X"00",X"20",X"FF",X"00",X"00",X"68",X"06",X"00",
		X"40",X"03",X"11",X"22",X"20",X"00",X"00",X"FF",X"00",X"00",X"08",X"06",X"00",X"00",X"04",X"33",
		X"32",X"00",X"00",X"42",X"FF",X"00",X"00",X"06",X"70",X"65",X"54",X"44",X"33",X"30",X"00",X"00",
		X"43",X"FF",X"20",X"00",X"00",X"70",X"06",X"64",X"44",X"44",X"00",X"00",X"04",X"32",X"FF",X"21",
		X"60",X"00",X"67",X"06",X"65",X"00",X"00",X"00",X"00",X"44",X"31",X"FF",X"35",X"67",X"00",X"06",
		X"00",X"05",X"11",X"10",X"00",X"04",X"43",X"20",X"FF",X"22",X"56",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"53",X"10",X"FF",X"12",X"40",X"67",X"00",X"55",X"50",X"05",X"50",X"05",X"55",
		X"32",X"00",X"FF",X"03",X"44",X"56",X"00",X"04",X"50",X"00",X"00",X"44",X"33",X"20",X"00",X"FF",
		X"01",X"34",X"45",X"05",X"50",X"00",X"00",X"03",X"33",X"21",X"00",X"00",X"FF",X"00",X"13",X"44",
		X"40",X"50",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"FF",X"00",X"01",X"33",X"40",X"00",X"00",
		X"00",X"22",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"12",X"33",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"13",X"30",X"90",X"00",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"01",X"20",X"09",X"00",X"00",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",X"FF",X"00",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"FF",X"00",X"AA",X"A4",X"44",X"44",
		X"44",X"44",X"44",X"4A",X"AA",X"A0",X"FF",X"0A",X"AE",X"43",X"33",X"32",X"22",X"22",X"22",X"23",
		X"6A",X"A8",X"FF",X"0A",X"A4",X"33",X"22",X"11",X"11",X"11",X"11",X"12",X"36",X"AA",X"FF",X"8A",
		X"94",X"32",X"22",X"22",X"22",X"22",X"22",X"11",X"26",X"AA",X"FF",X"AA",X"54",X"32",X"22",X"22",
		X"22",X"22",X"22",X"22",X"26",X"AA",X"FF",X"AA",X"54",X"32",X"22",X"34",X"44",X"44",X"44",X"44",
		X"6A",X"A8",X"FF",X"AA",X"54",X"32",X"22",X"45",X"55",X"55",X"55",X"54",X"AA",X"A0",X"FF",X"AA",
		X"54",X"32",X"22",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",
		X"AA",X"AA",X"AA",X"A8",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",
		X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"AA",X"AA",X"80",X"00",X"00",X"00",X"FF",X"AA",
		X"54",X"32",X"12",X"66",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"34",
		X"44",X"44",X"6A",X"AA",X"00",X"00",X"FF",X"AA",X"54",X"32",X"21",X"22",X"22",X"22",X"36",X"AA",
		X"80",X"00",X"FF",X"AA",X"54",X"32",X"22",X"11",X"11",X"11",X"13",X"6A",X"A0",X"00",X"FF",X"AA",
		X"54",X"32",X"22",X"22",X"22",X"22",X"12",X"6A",X"A0",X"00",X"FF",X"AA",X"54",X"32",X"22",X"22",
		X"22",X"22",X"22",X"6A",X"A0",X"00",X"FF",X"AA",X"54",X"32",X"22",X"23",X"33",X"33",X"46",X"AA",
		X"80",X"00",X"FF",X"AA",X"54",X"32",X"22",X"35",X"55",X"55",X"4A",X"AA",X"00",X"00",X"FF",X"AA",
		X"54",X"32",X"12",X"44",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",
		X"AA",X"AA",X"80",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",
		X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"AA",X"94",X"31",X"22",X"6A",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",X"8A",
		X"E5",X"43",X"34",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"0A",X"AA",X"55",X"5A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"8A",X"AA",X"AA",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"08",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"08",X"AA",
		X"AA",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"FF",X"0A",X"AE",X"44",X"44",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"8A",X"94",X"32",X"23",X"6A",X"80",X"00",X"00",X"00",X"00",X"FF",X"AA",
		X"54",X"21",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"31",X"12",X"6A",X"A0",
		X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",
		X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",
		X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",
		X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",
		X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",
		X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",
		X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",
		X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",
		X"32",X"12",X"6A",X"A0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A8",X"00",
		X"00",X"00",X"00",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"AA",X"AA",X"A8",X"00",X"00",X"FF",X"AA",
		X"54",X"32",X"21",X"26",X"AA",X"AA",X"AA",X"A0",X"00",X"FF",X"AA",X"54",X"32",X"21",X"22",X"64",
		X"44",X"6A",X"AA",X"00",X"FF",X"AA",X"54",X"32",X"22",X"11",X"12",X"22",X"26",X"AA",X"80",X"FF",
		X"AA",X"54",X"33",X"22",X"22",X"21",X"11",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"33",X"32",X"22",
		X"22",X"22",X"21",X"6A",X"A0",X"FF",X"AA",X"E5",X"33",X"33",X"33",X"33",X"32",X"21",X"6A",X"A0",
		X"FF",X"8A",X"A9",X"54",X"44",X"44",X"44",X"33",X"16",X"AA",X"80",X"FF",X"0A",X"AA",X"E5",X"55",
		X"55",X"55",X"46",X"6A",X"AA",X"00",X"FF",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"00",X"FF",X"00",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",X"FF",X"00",X"08",X"AA",
		X"A8",X"00",X"00",X"FF",X"08",X"AA",X"AA",X"AA",X"A8",X"00",X"FF",X"0A",X"A9",X"E4",X"46",X"AA",
		X"00",X"FF",X"8A",X"5E",X"32",X"23",X"6A",X"80",X"FF",X"AA",X"54",X"31",X"12",X"6A",X"A0",X"FF",
		X"AA",X"54",X"31",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",
		X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",
		X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",
		X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",
		X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",
		X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"12",X"6A",
		X"A0",X"FF",X"AA",X"54",X"32",X"22",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"22",X"6A",X"A0",X"FF",
		X"AA",X"54",X"32",X"22",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"22",X"6A",X"A0",X"FF",X"AA",X"54",
		X"32",X"22",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"22",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"22",
		X"6A",X"A0",X"FF",X"8A",X"A5",X"43",X"34",X"AA",X"80",X"FF",X"0A",X"AA",X"55",X"44",X"AA",X"00",
		X"FF",X"08",X"AA",X"AA",X"AA",X"A8",X"00",X"FF",X"00",X"08",X"33",X"38",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"08",X"AA",X"AA",X"AA",X"A8",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",X"00",X"FF",X"00",X"00",X"AA",X"A6",X"44",X"44",X"44",
		X"4A",X"AA",X"A0",X"00",X"00",X"FF",X"00",X"0A",X"AE",X"59",X"93",X"33",X"33",X"66",X"6A",X"A8",
		X"00",X"00",X"FF",X"00",X"AA",X"E5",X"43",X"33",X"22",X"11",X"12",X"26",X"AA",X"00",X"00",X"FF",
		X"00",X"AA",X"54",X"33",X"22",X"22",X"22",X"21",X"22",X"6A",X"A0",X"00",X"FF",X"0A",X"AE",X"54",
		X"32",X"22",X"22",X"22",X"22",X"12",X"26",X"A8",X"00",X"FF",X"0A",X"A5",X"43",X"32",X"22",X"44",
		X"44",X"32",X"21",X"26",X"AA",X"00",X"FF",X"8A",X"85",X"43",X"22",X"24",X"AA",X"A5",X"43",X"21",
		X"22",X"6A",X"A0",X"FF",X"8A",X"95",X"33",X"22",X"4A",X"AA",X"AA",X"54",X"32",X"12",X"6A",X"A0",
		X"FF",X"AA",X"54",X"32",X"22",X"6A",X"80",X"8A",X"59",X"44",X"44",X"6A",X"A0",X"FF",X"AA",X"54",
		X"32",X"23",X"AA",X"00",X"0A",X"A5",X"55",X"55",X"AA",X"80",X"FF",X"A9",X"54",X"32",X"26",X"AA",
		X"00",X"08",X"AA",X"AA",X"AA",X"A8",X"00",X"FF",X"A5",X"54",X"22",X"26",X"A8",X"00",X"00",X"8A",
		X"AA",X"A8",X"00",X"00",X"FF",X"A5",X"54",X"22",X"26",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"A5",X"54",X"22",X"26",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"A5",
		X"54",X"22",X"26",X"A8",X"00",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"FF",X"A9",X"54",X"32",X"26",
		X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"A8",X"00",X"FF",X"AA",X"54",X"32",X"26",X"AA",X"00",X"0A",
		X"A9",X"44",X"44",X"AA",X"80",X"FF",X"AA",X"54",X"32",X"24",X"AA",X"80",X"8A",X"54",X"33",X"33",
		X"4A",X"A0",X"FF",X"8A",X"95",X"42",X"22",X"AA",X"AA",X"AA",X"54",X"32",X"12",X"6A",X"A0",X"FF",
		X"8A",X"85",X"43",X"22",X"4A",X"AA",X"A5",X"43",X"21",X"22",X"6A",X"80",X"FF",X"0A",X"A5",X"43",
		X"22",X"23",X"44",X"43",X"32",X"21",X"26",X"AA",X"00",X"FF",X"0A",X"AE",X"54",X"32",X"22",X"23",
		X"32",X"22",X"12",X"6A",X"A8",X"00",X"FF",X"00",X"AA",X"54",X"33",X"22",X"22",X"22",X"22",X"23",
		X"6A",X"A0",X"00",X"FF",X"00",X"AA",X"E5",X"44",X"33",X"22",X"22",X"22",X"36",X"AA",X"00",X"00",
		X"FF",X"00",X"0A",X"AE",X"55",X"44",X"44",X"44",X"36",X"6A",X"A8",X"00",X"00",X"FF",X"00",X"00",
		X"AA",X"AE",X"55",X"55",X"5A",X"6A",X"AA",X"A0",X"00",X"00",X"FF",X"00",X"00",X"08",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A8",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"AA",X"AA",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"AA",X"80",X"00",X"00",X"00",X"08",X"AA",X"AA",X"00",
		X"FF",X"08",X"AA",X"AA",X"AA",X"80",X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"FF",X"0A",X"A5",X"44",
		X"9A",X"A0",X"00",X"0A",X"A5",X"44",X"AA",X"A0",X"FF",X"AA",X"59",X"31",X"3A",X"A8",X"00",X"AA",
		X"54",X"33",X"66",X"AA",X"FF",X"AA",X"54",X"32",X"16",X"AA",X"0A",X"A5",X"43",X"31",X"26",X"AA",
		X"FF",X"AA",X"54",X"32",X"16",X"AA",X"AA",X"54",X"32",X"21",X"26",X"A8",X"FF",X"AA",X"54",X"32",
		X"16",X"AA",X"A5",X"43",X"22",X"21",X"6A",X"A0",X"FF",X"AA",X"54",X"32",X"16",X"AA",X"54",X"32",
		X"22",X"12",X"6A",X"80",X"FF",X"AA",X"54",X"32",X"16",X"A5",X"43",X"22",X"21",X"26",X"AA",X"00",
		X"FF",X"AA",X"54",X"32",X"16",X"54",X"32",X"22",X"12",X"6A",X"A0",X"00",X"FF",X"AA",X"54",X"32",
		X"13",X"43",X"22",X"21",X"26",X"AA",X"00",X"00",X"FF",X"AA",X"54",X"32",X"22",X"32",X"22",X"22",
		X"6A",X"A0",X"00",X"00",X"FF",X"AA",X"54",X"32",X"22",X"22",X"22",X"26",X"6A",X"00",X"00",X"00",
		X"FF",X"AA",X"54",X"32",X"22",X"22",X"22",X"22",X"6A",X"80",X"00",X"00",X"FF",X"AA",X"54",X"32",
		X"22",X"22",X"22",X"22",X"6A",X"A0",X"00",X"00",X"FF",X"AA",X"54",X"32",X"22",X"22",X"22",X"22",
		X"26",X"A0",X"00",X"00",X"FF",X"AA",X"54",X"32",X"22",X"26",X"42",X"21",X"26",X"A8",X"00",X"00",
		X"FF",X"AA",X"54",X"32",X"22",X"65",X"54",X"21",X"26",X"AA",X"00",X"00",X"FF",X"AA",X"54",X"32",
		X"26",X"AA",X"54",X"22",X"12",X"6A",X"00",X"00",X"FF",X"AA",X"54",X"32",X"26",X"AA",X"A5",X"42",
		X"12",X"6A",X"80",X"00",X"FF",X"AA",X"54",X"32",X"16",X"AA",X"A5",X"42",X"21",X"6A",X"A0",X"00",
		X"FF",X"AA",X"54",X"32",X"16",X"AA",X"AA",X"52",X"21",X"26",X"A0",X"00",X"FF",X"AA",X"54",X"32",
		X"16",X"AA",X"8A",X"54",X"21",X"26",X"AA",X"00",X"FF",X"AA",X"54",X"32",X"16",X"AA",X"0A",X"A5",
		X"22",X"16",X"AA",X"80",X"FF",X"AA",X"54",X"32",X"16",X"AA",X"0A",X"A5",X"42",X"12",X"6A",X"A0",
		X"FF",X"AA",X"59",X"31",X"26",X"AA",X"08",X"A5",X"42",X"22",X"6A",X"A0",X"FF",X"8A",X"E5",X"42",
		X"46",X"A8",X"00",X"AA",X"54",X"23",X"9A",X"80",X"FF",X"0A",X"AE",X"55",X"9A",X"A0",X"00",X"AA",
		X"E5",X"55",X"AA",X"00",X"FF",X"08",X"AA",X"AA",X"AA",X"80",X"00",X"0A",X"AA",X"AA",X"A8",X"00",
		X"FF",X"00",X"08",X"AA",X"80",X"00",X"00",X"00",X"8A",X"AA",X"80",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8A",X"AA",X"80",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A5",
		X"44",X"AA",X"A0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"59",X"33",X"6A",X"A0",
		X"FF",X"00",X"00",X"8A",X"AA",X"80",X"00",X"08",X"A5",X"43",X"12",X"36",X"A8",X"FF",X"00",X"0A",
		X"AA",X"AA",X"AA",X"00",X"0A",X"A5",X"42",X"11",X"36",X"AA",X"FF",X"00",X"AA",X"A5",X"44",X"AA",
		X"A0",X"0A",X"A5",X"42",X"21",X"36",X"AA",X"FF",X"00",X"AA",X"54",X"33",X"4A",X"A0",X"0A",X"A5",
		X"42",X"21",X"36",X"AA",X"FF",X"0A",X"A5",X"43",X"21",X"36",X"A8",X"0A",X"A5",X"42",X"21",X"36",
		X"AA",X"FF",X"0A",X"A5",X"43",X"11",X"36",X"AA",X"0A",X"A5",X"42",X"21",X"36",X"AA",X"FF",X"0A",
		X"A5",X"43",X"11",X"36",X"AA",X"0A",X"A5",X"42",X"21",X"36",X"AA",X"FF",X"0A",X"A5",X"43",X"21",
		X"36",X"AA",X"0A",X"A5",X"42",X"21",X"36",X"AA",X"FF",X"0A",X"A5",X"43",X"21",X"36",X"AA",X"0A",
		X"A5",X"42",X"21",X"36",X"AA",X"FF",X"0A",X"A5",X"43",X"22",X"23",X"6A",X"AA",X"A5",X"42",X"22",
		X"36",X"AA",X"FF",X"00",X"A5",X"43",X"22",X"23",X"6A",X"AA",X"A5",X"32",X"22",X"36",X"AA",X"FF",
		X"00",X"AA",X"54",X"32",X"22",X"36",X"AA",X"A5",X"32",X"22",X"36",X"AA",X"FF",X"00",X"AA",X"54",
		X"32",X"22",X"23",X"6A",X"A5",X"32",X"22",X"36",X"AA",X"FF",X"00",X"0A",X"A5",X"43",X"22",X"22",
		X"36",X"95",X"32",X"22",X"36",X"AA",X"FF",X"00",X"0A",X"A5",X"43",X"22",X"22",X"23",X"33",X"22",
		X"22",X"36",X"AA",X"FF",X"00",X"00",X"AA",X"54",X"32",X"22",X"22",X"22",X"22",X"22",X"36",X"AA",
		X"FF",X"00",X"00",X"AA",X"54",X"43",X"32",X"22",X"22",X"22",X"22",X"E6",X"A8",X"FF",X"00",X"00",
		X"0A",X"A5",X"54",X"44",X"32",X"22",X"22",X"23",X"6A",X"A0",X"FF",X"00",X"00",X"00",X"AA",X"A5",
		X"59",X"43",X"22",X"22",X"23",X"6A",X"A0",X"FF",X"00",X"00",X"00",X"0A",X"AA",X"A5",X"54",X"32",
		X"22",X"23",X"6A",X"80",X"FF",X"00",X"00",X"00",X"00",X"08",X"AA",X"54",X"32",X"22",X"23",X"6A",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"8E",X"AA",X"54",X"32",X"22",X"36",X"AA",X"00",X"FF",X"00",
		X"00",X"AA",X"AA",X"AA",X"A5",X"43",X"22",X"12",X"36",X"A0",X"00",X"FF",X"00",X"AA",X"AA",X"44",
		X"95",X"54",X"32",X"21",X"13",X"6A",X"A0",X"00",X"FF",X"0A",X"A4",X"44",X"44",X"44",X"43",X"22",
		X"11",X"23",X"6A",X"00",X"00",X"FF",X"AA",X"93",X"33",X"33",X"33",X"32",X"21",X"11",X"36",X"AA",
		X"00",X"00",X"FF",X"A5",X"32",X"22",X"22",X"22",X"22",X"11",X"14",X"6A",X"A0",X"00",X"00",X"FF",
		X"A5",X"32",X"22",X"22",X"22",X"22",X"22",X"46",X"AA",X"80",X"00",X"00",X"FF",X"AA",X"54",X"44",
		X"44",X"44",X"44",X"44",X"6A",X"A8",X"00",X"00",X"00",X"FF",X"0A",X"A5",X"55",X"55",X"55",X"9E",
		X"66",X"A8",X"00",X"00",X"00",X"00",X"FF",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"AA",X"A0",X"00",
		X"FF",X"00",X"00",X"00",X"0A",X"A3",X"AA",X"00",X"FF",X"00",X"00",X"00",X"AA",X"EE",X"3A",X"A0",
		X"FF",X"00",X"00",X"00",X"A3",X"A9",X"A5",X"A0",X"FF",X"00",X"00",X"00",X"A3",X"99",X"33",X"A0",
		X"FF",X"00",X"00",X"44",X"AA",X"3E",X"3A",X"A0",X"FF",X"00",X"00",X"9E",X"4A",X"A4",X"AA",X"A0",
		X"FF",X"00",X"00",X"35",X"DD",X"65",X"5D",X"A0",X"FF",X"0C",X"00",X"33",X"35",X"9E",X"45",X"50",
		X"FF",X"00",X"0B",X"00",X"01",X"19",X"EB",X"55",X"FF",X"01",X"00",X"94",X"41",X"1B",X"3E",X"45",
		X"FF",X"00",X"1C",X"33",X"44",X"BB",X"33",X"5C",X"FF",X"0B",X"12",X"B2",X"DD",X"DD",X"77",X"DD",
		X"FF",X"0D",X"77",X"88",X"89",X"88",X"77",X"8A",X"FF",X"0D",X"77",X"88",X"89",X"88",X"77",X"8A",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"AA",X"A0",X"00",
		X"FF",X"00",X"00",X"00",X"0A",X"A3",X"AA",X"00",X"FF",X"00",X"00",X"00",X"AA",X"EE",X"3A",X"A0",
		X"FF",X"00",X"00",X"00",X"A3",X"A9",X"A5",X"A0",X"FF",X"00",X"00",X"00",X"A3",X"99",X"33",X"A0",
		X"FF",X"00",X"04",X"40",X"AA",X"3E",X"3A",X"A0",X"FF",X"00",X"09",X"EE",X"AA",X"A4",X"AA",X"A0",
		X"FF",X"00",X"04",X"30",X"DD",X"65",X"5D",X"A0",X"FF",X"00",X"00",X"33",X"35",X"9E",X"45",X"50",
		X"FF",X"00",X"0B",X"00",X"01",X"19",X"EB",X"55",X"FF",X"00",X"00",X"94",X"41",X"1B",X"3E",X"45",
		X"FF",X"00",X"2E",X"33",X"44",X"BB",X"33",X"5C",X"FF",X"0B",X"19",X"11",X"DD",X"DD",X"28",X"DD",
		X"FF",X"0C",X"77",X"81",X"89",X"88",X"77",X"8A",X"FF",X"0D",X"77",X"88",X"89",X"88",X"77",X"8A",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"33",X"33",X"30",X"00",X"00",
		X"FF",X"00",X"03",X"66",X"36",X"63",X"00",X"00",X"FF",X"00",X"36",X"61",X"31",X"66",X"30",X"00",
		X"FF",X"00",X"36",X"61",X"31",X"66",X"30",X"00",X"FF",X"00",X"36",X"67",X"77",X"66",X"90",X"00",
		X"FF",X"00",X"33",X"77",X"77",X"73",X"99",X"00",X"FF",X"00",X"93",X"35",X"55",X"33",X"99",X"00",
		X"FF",X"00",X"93",X"A6",X"66",X"A3",X"99",X"00",X"FF",X"00",X"9A",X"66",X"66",X"6A",X"99",X"00",
		X"FF",X"00",X"9A",X"66",X"66",X"66",X"99",X"90",X"FF",X"00",X"92",X"2D",X"66",X"6D",X"22",X"00",
		X"FF",X"09",X"92",X"22",X"DD",X"D2",X"22",X"09",X"FF",X"00",X"00",X"22",X"22",X"22",X"99",X"99",
		X"FF",X"00",X"00",X"02",X"22",X"20",X"09",X"90",X"FF",X"00",X"00",X"00",X"09",X"00",X"09",X"00",
		X"FF",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"FF",X"00",X"00",X"33",X"33",X"30",X"00",X"00",
		X"FF",X"00",X"03",X"66",X"36",X"63",X"00",X"00",X"FF",X"00",X"36",X"66",X"36",X"66",X"30",X"00",
		X"FF",X"00",X"36",X"61",X"31",X"66",X"30",X"00",X"FF",X"00",X"36",X"67",X"77",X"66",X"90",X"00",
		X"FF",X"00",X"33",X"77",X"77",X"73",X"99",X"00",X"FF",X"00",X"93",X"35",X"55",X"33",X"99",X"00",
		X"FF",X"00",X"99",X"A6",X"66",X"A9",X"99",X"00",X"FF",X"00",X"99",X"66",X"66",X"69",X"99",X"00",
		X"FF",X"00",X"99",X"96",X"66",X"69",X"99",X"00",X"FF",X"00",X"09",X"96",X"66",X"99",X"20",X"00",
		X"FF",X"00",X"02",X"2A",X"DD",X"C2",X"20",X"00",X"FF",X"00",X"00",X"22",X"22",X"24",X"90",X"09",
		X"FF",X"00",X"00",X"02",X"22",X"20",X"99",X"94",X"FF",X"00",X"00",X"00",X"94",X"00",X"99",X"00",
		X"FF",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"03",X"33",X"33",X"00",X"00",X"FF",X"00",X"00",X"36",X"63",X"66",X"30",X"00",
		X"FF",X"00",X"03",X"66",X"63",X"66",X"63",X"00",X"FF",X"00",X"03",X"66",X"13",X"16",X"63",X"00",
		X"FF",X"00",X"03",X"66",X"77",X"76",X"63",X"00",X"FF",X"00",X"43",X"37",X"77",X"77",X"39",X"40",
		X"FF",X"00",X"89",X"33",X"55",X"53",X"39",X"40",X"FF",X"00",X"99",X"9A",X"66",X"6A",X"99",X"40",
		X"FF",X"00",X"99",X"99",X"66",X"69",X"99",X"40",X"FF",X"00",X"09",X"99",X"96",X"99",X"99",X"00",
		X"FF",X"00",X"02",X"99",X"99",X"99",X"93",X"00",X"FF",X"00",X"02",X"AD",X"DD",X"DC",X"33",X"00",
		X"FF",X"00",X"00",X"22",X"CC",X"C2",X"20",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"90",X"00",
		X"FF",X"00",X"89",X"99",X"90",X"00",X"90",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",X"99",X"90",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"03",X"33",X"33",X"00",X"00",X"FF",X"00",X"00",X"36",X"63",X"66",X"30",X"00",
		X"FF",X"00",X"03",X"66",X"13",X"16",X"63",X"00",X"FF",X"00",X"03",X"66",X"13",X"16",X"63",X"00",
		X"FF",X"00",X"03",X"66",X"77",X"76",X"63",X"00",X"FF",X"00",X"03",X"37",X"77",X"77",X"39",X"40",
		X"FF",X"00",X"09",X"33",X"55",X"53",X"39",X"40",X"FF",X"00",X"89",X"9A",X"66",X"6A",X"99",X"40",
		X"FF",X"00",X"89",X"96",X"66",X"66",X"99",X"40",X"FF",X"00",X"09",X"96",X"66",X"66",X"99",X"00",
		X"FF",X"00",X"08",X"9D",X"66",X"6D",X"99",X"00",X"FF",X"00",X"00",X"8A",X"D6",X"DC",X"42",X"00",
		X"FF",X"00",X"00",X"42",X"AA",X"A3",X"20",X"00",X"FF",X"00",X"99",X"99",X"22",X"22",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"89",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"99",X"99",X"90",
		X"FF",X"00",X"00",X"30",X"00",X"00",X"FF",X"00",X"06",X"56",X"00",X"00",X"FF",X"85",X"A5",X"85",
		X"30",X"00",X"FF",X"65",X"32",X"21",X"23",X"80",X"FF",X"08",X"3A",X"A2",X"AA",X"38",X"FF",X"03",
		X"8A",X"A8",X"AA",X"83",X"FF",X"08",X"8A",X"D8",X"DA",X"88",X"FF",X"0D",X"8A",X"D8",X"DA",X"8D",
		X"FF",X"07",X"78",X"44",X"48",X"77",X"FF",X"07",X"E4",X"4D",X"44",X"7E",X"FF",X"00",X"83",X"44",
		X"43",X"80",X"FF",X"00",X"00",X"03",X"00",X"00",X"FF",X"08",X"23",X"24",X"23",X"28",X"FF",X"00",
		X"82",X"9A",X"92",X"80",X"FF",X"00",X"01",X"AA",X"A1",X"00",X"FF",X"00",X"02",X"4A",X"12",X"40",
		X"FF",X"00",X"00",X"22",X"24",X"40",X"FF",X"00",X"00",X"40",X"00",X"40",X"FF",X"00",X"04",X"44",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"68",X"00",X"00",X"FF",X"00",
		X"02",X"56",X"00",X"00",X"FF",X"85",X"A5",X"85",X"30",X"00",X"FF",X"65",X"32",X"11",X"23",X"80",
		X"FF",X"08",X"32",X"22",X"22",X"38",X"FF",X"03",X"8A",X"A8",X"AA",X"83",X"FF",X"08",X"8A",X"A8",
		X"AA",X"88",X"FF",X"03",X"8A",X"D8",X"DA",X"83",X"FF",X"07",X"78",X"44",X"48",X"77",X"FF",X"07",
		X"E4",X"34",X"34",X"7E",X"FF",X"00",X"02",X"2C",X"33",X"00",X"FF",X"00",X"01",X"39",X"23",X"00",
		X"FF",X"00",X"03",X"8A",X"82",X"00",X"FF",X"00",X"08",X"8A",X"88",X"00",X"FF",X"00",X"03",X"3A",
		X"32",X"00",X"FF",X"00",X"00",X"28",X"30",X"00",X"FF",X"00",X"00",X"40",X"40",X"00",X"FF",X"00",
		X"04",X"44",X"44",X"00",X"FF",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"02",X"32",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"19",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"FF",X"00",X"01",X"51",
		X"51",X"00",X"00",X"00",X"FF",X"00",X"91",X"11",X"11",X"90",X"00",X"00",X"FF",X"00",X"09",X"13",
		X"19",X"00",X"00",X"90",X"FF",X"00",X"00",X"08",X"00",X"00",X"00",X"90",X"FF",X"00",X"00",X"11",
		X"10",X"00",X"00",X"90",X"FF",X"00",X"01",X"33",X"D1",X"00",X"00",X"90",X"FF",X"01",X"10",X"3D",
		X"11",X"00",X"00",X"90",X"FF",X"00",X"03",X"8D",X"D3",X"00",X"77",X"77",X"FF",X"00",X"D8",X"DD",
		X"8D",X"D0",X"AA",X"CC",X"FF",X"00",X"00",X"10",X"90",X"00",X"66",X"CC",X"FF",X"0B",X"BB",X"1B",
		X"99",X"BB",X"66",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"FF",X"00",X"02",X"32",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"FF",X"00",X"01",X"11",
		X"11",X"00",X"00",X"00",X"FF",X"00",X"91",X"51",X"51",X"90",X"00",X"00",X"FF",X"00",X"09",X"13",
		X"19",X"00",X"00",X"10",X"FF",X"00",X"00",X"08",X"00",X"00",X"00",X"90",X"FF",X"00",X"00",X"11",
		X"10",X"00",X"00",X"90",X"FF",X"00",X"01",X"D3",X"31",X"10",X"00",X"90",X"FF",X"00",X"01",X"1D",
		X"D0",X"00",X"00",X"90",X"FF",X"00",X"03",X"D8",X"D8",X"D0",X"77",X"77",X"FF",X"00",X"0D",X"8D",
		X"8D",X"00",X"AA",X"CC",X"FF",X"00",X"00",X"90",X"10",X"00",X"66",X"CC",X"FF",X"0B",X"B1",X"1B",
		X"1B",X"BB",X"66",X"CC",X"FF",X"00",X"00",X"02",X"12",X"20",X"00",X"00",X"FF",X"00",X"02",X"29",
		X"99",X"22",X"00",X"00",X"FF",X"00",X"00",X"61",X"11",X"12",X"00",X"00",X"FF",X"00",X"00",X"37",
		X"11",X"91",X"20",X"00",X"FF",X"00",X"03",X"44",X"42",X"19",X"22",X"20",X"FF",X"00",X"00",X"D1",
		X"52",X"22",X"22",X"20",X"FF",X"00",X"00",X"45",X"56",X"22",X"22",X"00",X"FF",X"00",X"03",X"99",
		X"44",X"45",X"50",X"00",X"FF",X"00",X"44",X"44",X"43",X"55",X"40",X"00",X"FF",X"09",X"46",X"53",
		X"35",X"45",X"54",X"CC",X"FF",X"0C",X"34",X"54",X"35",X"4C",X"64",X"4C",X"FF",X"0C",X"C3",X"95",
		X"35",X"46",X"64",X"CC",X"FF",X"0C",X"CC",X"95",X"45",X"66",X"4C",X"CC",X"FF",X"0B",X"BB",X"E5",
		X"55",X"6B",X"BB",X"BB",X"FF",X"0B",X"BE",X"88",X"88",X"88",X"BB",X"BB",X"FF",X"0A",X"AA",X"E8",
		X"88",X"8E",X"AA",X"AA",X"FF",X"0A",X"AA",X"44",X"58",X"44",X"AA",X"AA",X"FF",X"01",X"11",X"44",
		X"56",X"54",X"61",X"11",X"FF",X"00",X"00",X"02",X"12",X"20",X"00",X"00",X"FF",X"00",X"02",X"21",
		X"19",X"22",X"00",X"00",X"FF",X"00",X"00",X"51",X"19",X"92",X"20",X"00",X"FF",X"00",X"00",X"36",
		X"11",X"91",X"22",X"00",X"FF",X"00",X"03",X"44",X"22",X"99",X"22",X"20",X"FF",X"00",X"00",X"D1",
		X"52",X"22",X"22",X"00",X"FF",X"00",X"00",X"45",X"56",X"22",X"20",X"00",X"FF",X"00",X"00",X"33",
		X"44",X"45",X"30",X"00",X"FF",X"00",X"04",X"44",X"43",X"55",X"43",X"00",X"FF",X"00",X"44",X"33",
		X"35",X"45",X"53",X"9C",X"FF",X"0C",X"55",X"B6",X"35",X"46",X"54",X"3C",X"FF",X"0C",X"C4",X"96",
		X"35",X"45",X"53",X"CC",X"FF",X"0C",X"CC",X"45",X"45",X"56",X"4C",X"CC",X"FF",X"0B",X"BB",X"E5",
		X"55",X"56",X"BB",X"BB",X"FF",X"0B",X"BB",X"B8",X"88",X"88",X"8B",X"BB",X"FF",X"0A",X"AA",X"A8",
		X"88",X"88",X"5A",X"AA",X"FF",X"0A",X"AA",X"A5",X"54",X"84",X"4A",X"AA",X"FF",X"01",X"11",X"14",
		X"56",X"54",X"41",X"11",X"FF",X"22",X"22",X"22",X"00",X"FF",X"27",X"77",X"77",X"00",X"FF",X"00",
		X"55",X"00",X"00",X"FF",X"00",X"55",X"00",X"00",X"FF",X"00",X"55",X"00",X"00",X"FF",X"00",X"55",
		X"00",X"00",X"FF",X"00",X"55",X"00",X"00",X"FF",X"00",X"55",X"00",X"00",X"FF",X"00",X"02",X"00",
		X"00",X"FF",X"00",X"27",X"20",X"00",X"FF",X"02",X"77",X"00",X"00",X"FF",X"27",X"75",X"50",X"00",
		X"FF",X"07",X"00",X"55",X"00",X"FF",X"00",X"00",X"05",X"50",X"FF",X"00",X"00",X"00",X"55",X"FF",
		X"00",X"00",X"00",X"05",X"FF",X"00",X"00",X"00",X"00",X"FF",X"22",X"00",X"00",X"00",X"FF",X"27",
		X"00",X"00",X"00",X"FF",X"27",X"55",X"55",X"55",X"FF",X"27",X"55",X"55",X"55",X"FF",X"27",X"00",
		X"00",X"00",X"FF",X"27",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"B1",X"B0",
		X"00",X"FF",X"00",X"BB",X"B0",X"00",X"FF",X"00",X"0A",X"00",X"00",X"FF",X"0A",X"0A",X"0A",X"00",
		X"FF",X"00",X"AA",X"A0",X"00",X"FF",X"02",X"22",X"22",X"00",X"FF",X"00",X"22",X"20",X"00",X"FF",
		X"00",X"22",X"20",X"00",X"FF",X"00",X"0B",X"00",X"00",X"FF",X"00",X"1B",X"00",X"00",X"FF",X"0B",
		X"BA",X"0A",X"00",X"FF",X"00",X"00",X"AA",X"20",X"FF",X"00",X"0A",X"A2",X"22",X"FF",X"00",X"00",
		X"22",X"22",X"FF",X"00",X"00",X"02",X"20",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"0A",X"02",X"00",X"FF",X"BB",X"00",X"A2",X"22",X"FF",X"1B",X"AA",X"A2",X"22",
		X"FF",X"BB",X"00",X"A2",X"22",X"FF",X"00",X"0A",X"02",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"08",X"CC",X"EE",X"00",X"00",X"FF",X"08",X"CD",X"EE",X"88",X"00",
		X"FF",X"08",X"CD",X"EE",X"0C",X"00",X"FF",X"08",X"CD",X"EE",X"0C",X"00",X"FF",X"08",X"CD",X"EE",
		X"0C",X"00",X"FF",X"08",X"CD",X"EE",X"C0",X"00",X"FF",X"08",X"CD",X"EE",X"00",X"00",X"FF",X"08",
		X"CD",X"EE",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"08",X"CC",X"C0",X"00",X"FF",X"00",X"CC",X"80",X"0C",X"00",X"FF",X"0C",X"ED",X"C8",
		X"00",X"E0",X"FF",X"CE",X"EE",X"DD",X"80",X"E0",X"FF",X"0E",X"EE",X"ED",X"C8",X"00",X"FF",X"00",
		X"EE",X"ED",X"DC",X"80",X"FF",X"00",X"0E",X"EE",X"ED",X"00",X"FF",X"00",X"00",X"EE",X"E0",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"08",X"88",X"80",X"00",X"00",X"FF",X"0E",X"00",X"0C",
		X"00",X"00",X"FF",X"CC",X"CC",X"CC",X"C0",X"00",X"FF",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"EE",
		X"EE",X"EE",X"E0",X"00",X"FF",X"EE",X"EE",X"EE",X"E0",X"00",X"FF",X"EE",X"EE",X"EE",X"E0",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0C",X"C0",
		X"00",X"00",X"FF",X"00",X"08",X"80",X"00",X"00",X"FF",X"02",X"CC",X"D0",X"00",X"00",X"FF",X"0C",
		X"0C",X"D0",X"00",X"00",X"FF",X"0C",X"0C",X"D0",X"00",X"00",X"FF",X"02",X"CC",X"D0",X"00",X"00",
		X"FF",X"00",X"0C",X"D0",X"00",X"00",X"FF",X"00",X"C1",X"C0",X"00",X"00",X"FF",X"0C",X"C2",X"CC",
		X"00",X"00",X"FF",X"CC",X"00",X"00",X"00",X"00",X"FF",X"D8",X"00",X"00",X"00",X"00",X"FF",X"0D",
		X"C0",X"00",X"00",X"00",X"FF",X"0C",X"DC",X"00",X"00",X"00",X"FF",X"02",X"0D",X"C0",X"00",X"00",
		X"FF",X"00",X"CC",X"DC",X"CC",X"00",X"FF",X"00",X"00",X"C1",X"C0",X"00",X"FF",X"00",X"00",X"CC",
		X"00",X"00",X"FF",X"00",X"00",X"C0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"C0",X"FF",X"00",X"00",X"00",X"0C",X"C0",X"FF",X"C8",X"CC",X"CC",X"C1",X"C0",
		X"FF",X"C8",X"DD",X"DD",X"DC",X"C0",X"FF",X"00",X"C0",X"0C",X"00",X"C0",X"FF",X"00",X"2C",X"C2",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"C1",X"00",X"00",X"FF",X"0C",X"DD",X"DD",X"20",X"00",
		X"FF",X"CC",X"C0",X"0C",X"CC",X"00",X"FF",X"00",X"0C",X"C0",X"00",X"00",X"FF",X"00",X"C1",X"1C",
		X"00",X"00",X"FF",X"0C",X"13",X"31",X"C0",X"00",X"FF",X"C2",X"C1",X"1C",X"CC",X"00",X"FF",X"DD",
		X"DD",X"DD",X"DD",X"00",X"FF",X"00",X"01",X"2C",X"C0",X"00",X"FF",X"00",X"CD",X"CC",X"00",X"00",
		X"FF",X"0C",X"D0",X"C0",X"00",X"00",X"FF",X"CD",X"0C",X"CC",X"CC",X"00",X"FF",X"CC",X"CC",X"31",
		X"CC",X"D0",X"FF",X"CC",X"0C",X"31",X"CD",X"00",X"FF",X"C0",X"0C",X"CC",X"D0",X"00",X"FF",X"00",
		X"0C",X"2D",X"00",X"00",X"FF",X"00",X"00",X"D0",X"00",X"00",X"FF",X"00",X"C0",X"00",X"CD",X"00",
		X"FF",X"02",X"C0",X"0C",X"CD",X"00",X"FF",X"1D",X"C0",X"C1",X"CD",X"00",X"FF",X"CD",X"0C",X"13",
		X"1D",X"00",X"FF",X"CD",X"0C",X"13",X"1D",X"00",X"FF",X"CD",X"C0",X"C1",X"CD",X"00",X"FF",X"0C",
		X"C0",X"0C",X"2D",X"00",X"FF",X"00",X"C0",X"00",X"CD",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"10",X"FF",X"22",X"CC",X"22",X"01",X"FF",X"11",
		X"11",X"11",X"01",X"FF",X"01",X"11",X"10",X"10",X"FF",X"00",X"77",X"00",X"00",X"FF",X"11",X"11",
		X"11",X"10",X"FF",X"00",X"00",X"11",X"00",X"FF",X"00",X"00",X"20",X"10",X"FF",X"00",X"0C",X"10",
		X"10",X"FF",X"00",X"C1",X"11",X"00",X"FF",X"02",X"11",X"10",X"01",X"FF",X"21",X"11",X"10",X"10",
		X"FF",X"01",X"11",X"71",X"00",X"FF",X"00",X"00",X"10",X"00",X"FF",X"00",X"01",X"00",X"00",X"FF",
		X"00",X"10",X"00",X"00",X"FF",X"11",X"10",X"00",X"00",X"FF",X"10",X"01",X"01",X"00",X"FF",X"02",
		X"10",X"01",X"00",X"FF",X"02",X"11",X"01",X"00",X"FF",X"0C",X"11",X"71",X"00",X"FF",X"0C",X"11",
		X"71",X"00",X"FF",X"02",X"11",X"01",X"00",X"FF",X"02",X"10",X"01",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"09",X"00",X"09",X"00",X"00",X"FF",X"98",X"00",X"08",
		X"90",X"00",X"FF",X"09",X"85",X"89",X"00",X"00",X"FF",X"00",X"0C",X"00",X"00",X"00",X"FF",X"00",
		X"85",X"80",X"00",X"00",X"FF",X"08",X"55",X"58",X"00",X"00",X"FF",X"95",X"00",X"05",X"90",X"00",
		X"FF",X"95",X"00",X"05",X"90",X"00",X"FF",X"08",X"00",X"08",X"00",X"00",X"FF",X"00",X"99",X"80",
		X"00",X"00",X"FF",X"00",X"08",X"90",X"00",X"00",X"FF",X"90",X"00",X"90",X"00",X"00",X"FF",X"98",
		X"0C",X"88",X"89",X"00",X"FF",X"89",X"98",X"05",X"55",X"90",X"FF",X"00",X"08",X"50",X"05",X"80",
		X"FF",X"00",X"08",X"50",X"00",X"80",X"FF",X"00",X"09",X"55",X"00",X"00",X"FF",X"00",X"00",X"98",
		X"80",X"00",X"FF",X"09",X"00",X"00",X"99",X"00",X"FF",X"98",X"90",X"08",X"55",X"80",X"FF",X"00",
		X"80",X"85",X"00",X"00",X"FF",X"00",X"5C",X"50",X"00",X"00",X"FF",X"00",X"80",X"85",X"00",X"00",
		X"FF",X"98",X"90",X"08",X"55",X"80",X"FF",X"09",X"00",X"00",X"99",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"09",X"00",X"00",X"FF",X"08",X"89",
		X"98",X"80",X"FF",X"81",X"38",X"88",X"88",X"FF",X"82",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",
		X"88",X"FF",X"08",X"88",X"88",X"80",X"FF",X"08",X"88",X"8A",X"80",X"FF",X"00",X"8A",X"AA",X"00",
		X"FF",X"00",X"88",X"80",X"00",X"FF",X"08",X"88",X"88",X"80",X"FF",X"08",X"88",X"88",X"AA",X"FF",
		X"09",X"88",X"88",X"8A",X"FF",X"99",X"88",X"88",X"8A",X"FF",X"08",X"38",X"88",X"88",X"FF",X"08",
		X"12",X"88",X"80",X"FF",X"00",X"88",X"80",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"90",X"08",
		X"88",X"00",X"FF",X"09",X"98",X"88",X"80",X"FF",X"83",X"88",X"88",X"80",X"FF",X"81",X"38",X"88",
		X"88",X"FF",X"88",X"88",X"88",X"AA",X"FF",X"08",X"88",X"8A",X"AA",X"FF",X"00",X"08",X"AA",X"00",
		X"FF",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",X"01",X"11",X"00",X"00",X"FF",X"10",X"08",X"88",
		X"0E",X"E0",X"FF",X"01",X"01",X"11",X"E0",X"E0",X"FF",X"01",X"01",X"11",X"00",X"E0",X"FF",X"01",
		X"11",X"11",X"E0",X"E0",X"FF",X"00",X"01",X"11",X"0E",X"00",X"FF",X"00",X"01",X"11",X"00",X"00",
		X"FF",X"00",X"00",X"0E",X"E0",X"00",X"FF",X"01",X"11",X"0E",X"0E",X"00",X"FF",X"01",X"18",X"1E",
		X"0E",X"00",X"FF",X"01",X"81",X"11",X"0E",X"00",X"FF",X"00",X"11",X"11",X"10",X"00",X"FF",X"10",
		X"01",X"11",X"11",X"00",X"FF",X"01",X"11",X"11",X"10",X"00",X"FF",X"00",X"10",X"01",X"00",X"00",
		X"FF",X"00",X"EE",X"EE",X"00",X"00",X"FF",X"00",X"E0",X"00",X"E0",X"00",X"FF",X"00",X"0E",X"0E",
		X"00",X"00",X"FF",X"01",X"81",X"11",X"11",X"00",X"FF",X"11",X"81",X"11",X"11",X"00",X"FF",X"01",
		X"81",X"11",X"11",X"00",X"FF",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"01",X"11",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0B",X"00",X"00",X"00",X"FF",X"00",X"05",X"00",
		X"00",X"00",X"FF",X"00",X"05",X"00",X"00",X"00",X"FF",X"00",X"55",X"50",X"00",X"00",X"FF",X"00",
		X"11",X"50",X"00",X"00",X"FF",X"00",X"11",X"50",X"00",X"00",X"FF",X"00",X"11",X"50",X"00",X"00",
		X"FF",X"00",X"55",X"50",X"00",X"00",X"FF",X"00",X"55",X"50",X"00",X"00",X"FF",X"B0",X"00",X"00",
		X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"00",X"FF",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",
		X"55",X"50",X"00",X"00",X"FF",X"00",X"51",X"55",X"00",X"00",X"FF",X"00",X"01",X"15",X"50",X"00",
		X"FF",X"00",X"00",X"15",X"50",X"00",X"FF",X"00",X"00",X"05",X"50",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"05",X"55",X"55",X"50",
		X"FF",X"B5",X"55",X"11",X"15",X"50",X"FF",X"00",X"05",X"11",X"15",X"50",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"09",X"90",X"90",X"00",X"FF",X"00",
		X"99",X"99",X"00",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",X"99",X"99",
		X"99",X"90",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",X"EE",X"E9",X"EE",X"E0",X"FF",X"00",X"90",X"E0",
		X"00",X"FF",X"90",X"9E",X"EE",X"00",X"FF",X"99",X"9E",X"E9",X"E0",X"FF",X"0E",X"E9",X"9E",X"EE",
		X"FF",X"EE",X"E9",X"9E",X"E0",X"FF",X"0E",X"9E",X"E9",X"00",X"FF",X"00",X"EE",X"E0",X"00",X"FF",
		X"00",X"0E",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"9E",X"E0",X"FF",X"09",
		X"EE",X"9E",X"E0",X"FF",X"99",X"EE",X"9E",X"E0",X"FF",X"09",X"99",X"99",X"90",X"FF",X"99",X"EE",
		X"9E",X"E0",X"FF",X"90",X"EE",X"9E",X"E0",X"FF",X"00",X"EE",X"9E",X"E0",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"11",X"00",X"00",X"FF",X"00",X"99",X"99",X"99",X"00",X"FF",X"18",X"88",X"88",X"88",X"81",
		X"FF",X"19",X"99",X"99",X"99",X"11",X"FF",X"09",X"99",X"99",X"99",X"90",X"FF",X"09",X"99",X"99",
		X"99",X"90",X"FF",X"00",X"99",X"99",X"99",X"00",X"FF",X"00",X"00",X"98",X"10",X"00",X"FF",X"00",
		X"19",X"81",X"10",X"00",X"FF",X"01",X"98",X"99",X"90",X"00",X"FF",X"09",X"89",X"99",X"90",X"00",
		X"FF",X"98",X"99",X"99",X"90",X"00",X"FF",X"89",X"99",X"99",X"00",X"00",X"FF",X"19",X"99",X"90",
		X"00",X"00",X"FF",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"11",X"00",X"00",X"00",X"FF",X"00",X"81",X"99",X"00",X"00",
		X"FF",X"09",X"89",X"99",X"90",X"00",X"FF",X"09",X"89",X"99",X"90",X"00",X"FF",X"19",X"89",X"99",
		X"90",X"00",X"FF",X"19",X"89",X"99",X"90",X"00",X"FF",X"09",X"89",X"99",X"90",X"00",X"FF",X"09",
		X"89",X"99",X"90",X"00",X"FF",X"00",X"89",X"99",X"00",X"00",X"FF",X"00",X"11",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"01",X"10",X"FF",X"AA",X"AA",X"AA",X"10",X"01",X"FF",X"AA",
		X"AA",X"AA",X"00",X"01",X"FF",X"AA",X"AA",X"AA",X"00",X"01",X"FF",X"AA",X"AA",X"AA",X"11",X"10",
		X"FF",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"01",X"10",X"FF",X"00",X"00",X"E0",X"10",X"01",X"FF",X"00",X"0E",X"AA",X"10",X"01",X"FF",X"00",
		X"EA",X"AA",X"A0",X"10",X"FF",X"0E",X"AA",X"AA",X"AA",X"10",X"FF",X"EA",X"AA",X"AA",X"AA",X"A0",
		X"FF",X"0A",X"AA",X"AA",X"AA",X"00",X"FF",X"00",X"AA",X"AA",X"A0",X"00",X"FF",X"00",X"0A",X"AA",
		X"00",X"00",X"FF",X"00",X"00",X"A0",X"00",X"00",X"FF",X"00",X"11",X"10",X"00",X"00",X"FF",X"01",
		X"00",X"01",X"00",X"00",X"FF",X"01",X"00",X"01",X"00",X"00",X"FF",X"00",X"10",X"01",X"00",X"00",
		X"FF",X"0E",X"AA",X"AA",X"AA",X"00",X"FF",X"0E",X"AA",X"AA",X"AA",X"00",X"FF",X"0E",X"AA",X"AA",
		X"AA",X"00",X"FF",X"0E",X"AA",X"AA",X"AA",X"00",X"FF",X"0E",X"AA",X"AA",X"AA",X"00",X"FF",X"0E",
		X"AA",X"AA",X"AA",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"08",X"00",X"00",X"00",X"00",X"FF",X"00",X"88",X"80",X"00",X"00",X"00",
		X"FF",X"08",X"88",X"88",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EB",X"00",X"00",X"00",X"FF",X"0E",
		X"EE",X"EB",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EB",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EB",
		X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EB",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EB",X"00",X"00",
		X"00",X"FF",X"0C",X"BB",X"BC",X"00",X"00",X"00",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"08",X"88",X"80",X"00",X"00",X"00",X"FF",X"08",X"8E",X"EB",X"00",X"00",X"00",X"FF",X"08",X"EE",
		X"EB",X"B0",X"00",X"00",X"FF",X"08",X"EE",X"EE",X"BB",X"00",X"00",X"FF",X"00",X"EE",X"EE",X"EB",
		X"C0",X"00",X"FF",X"00",X"0E",X"EE",X"EB",X"00",X"00",X"FF",X"00",X"00",X"EE",X"B0",X"00",X"00",
		X"FF",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"8B",X"BB",X"BB",X"BC",X"FF",X"00",X"08",X"8E",X"EE",X"EE",
		X"EB",X"FF",X"08",X"88",X"8E",X"EE",X"EE",X"EB",X"FF",X"00",X"08",X"8E",X"EE",X"EE",X"EB",X"FF",
		X"00",X"00",X"8E",X"EE",X"EE",X"EC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",
		X"0D",X"DD",X"00",X"10",X"FF",X"BB",X"BB",X"BB",X"B1",X"01",X"FF",X"0B",X"BB",X"BB",X"B0",X"01",
		X"FF",X"00",X"BB",X"BB",X"B1",X"11",X"FF",X"00",X"BB",X"BB",X"B0",X"00",X"FF",X"00",X"00",X"00",
		X"10",X"00",X"FF",X"00",X"00",X"01",X"01",X"00",X"FF",X"00",X"00",X"B1",X"01",X"00",X"FF",X"00",
		X"1D",X"BB",X"01",X"00",X"FF",X"00",X"DB",X"BB",X"B0",X"00",X"FF",X"00",X"BB",X"BB",X"BB",X"00",
		X"FF",X"0B",X"BB",X"BB",X"B0",X"00",X"FF",X"BB",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"B0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"11",X"10",X"00",X"00",X"FF",X"01",
		X"00",X"10",X"00",X"00",X"FF",X"00",X"10",X"10",X"00",X"00",X"FF",X"00",X"BB",X"BB",X"00",X"00",
		X"FF",X"0D",X"BB",X"BB",X"00",X"00",X"FF",X"1D",X"BB",X"BB",X"00",X"00",X"FF",X"0D",X"BB",X"BB",
		X"00",X"00",X"FF",X"00",X"BB",X"BB",X"00",X"00",X"FF",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",
		X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"08",X"CC",X"EE",X"00",X"00",X"FF",X"08",X"CD",X"EE",X"88",X"00",X"FF",X"08",X"CD",X"EE",
		X"0C",X"00",X"FF",X"08",X"CD",X"EE",X"0C",X"00",X"FF",X"08",X"CD",X"EE",X"0C",X"00",X"FF",X"08",
		X"CD",X"EE",X"C0",X"00",X"FF",X"08",X"CD",X"EE",X"00",X"00",X"FF",X"08",X"CD",X"EE",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"CC",
		X"C0",X"00",X"FF",X"00",X"CC",X"80",X"0C",X"00",X"FF",X"0C",X"ED",X"C8",X"00",X"E0",X"FF",X"CE",
		X"EE",X"DD",X"80",X"E0",X"FF",X"0E",X"EE",X"ED",X"C8",X"00",X"FF",X"00",X"EE",X"ED",X"DC",X"80",
		X"FF",X"00",X"0E",X"EE",X"ED",X"00",X"FF",X"00",X"00",X"EE",X"E0",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"08",X"88",X"80",X"00",X"00",X"FF",X"0E",X"00",X"0C",X"00",X"00",X"FF",X"CC",
		X"CC",X"CC",X"C0",X"00",X"FF",X"DD",X"DD",X"DD",X"D0",X"00",X"FF",X"EE",X"EE",X"EE",X"E0",X"00",
		X"FF",X"EE",X"EE",X"EE",X"E0",X"00",X"FF",X"EE",X"EE",X"EE",X"E0",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
