library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_sp_bits_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"22",X"77",X"00",
		X"00",X"22",X"77",X"00",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"77",X"77",X"00",X"22",X"77",X"77",X"00",X"22",
		X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"77",X"66",X"66",X"00",X"77",X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"22",X"62",X"66",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"22",X"66",X"22",X"22",X"22",X"66",
		X"00",X"77",X"77",X"22",X"00",X"72",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",
		X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"77",X"77",X"00",X"22",X"77",X"77",X"00",X"22",
		X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"77",X"66",X"66",X"00",X"77",X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"22",X"62",X"66",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"22",X"66",X"22",X"22",X"22",X"66",
		X"00",X"77",X"77",X"22",X"00",X"72",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",
		X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"CC",X"77",X"00",X"00",X"0C",
		X"77",X"00",X"00",X"00",X"77",X"CC",X"00",X"00",X"C7",X"77",X"CC",X"00",X"CC",X"77",X"CC",X"00",
		X"00",X"22",X"77",X"C0",X"00",X"22",X"77",X"C0",X"CC",X"22",X"77",X"C0",X"CC",X"22",X"77",X"C0",
		X"77",X"22",X"22",X"00",X"77",X"22",X"22",X"00",X"22",X"22",X"22",X"C0",X"22",X"72",X"77",X"C0",
		X"77",X"77",X"72",X"77",X"77",X"77",X"22",X"77",X"77",X"22",X"22",X"CC",X"77",X"22",X"22",X"CC",
		X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"77",X"22",X"22",X"CC",X"77",X"72",X"22",X"CC",
		X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"55",X"00",X"CC",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"AA",X"A0",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"BB",X"C0",X"00",X"00",X"BB",X"C0",X"00",
		X"00",X"BB",X"C0",X"00",X"00",X"BB",X"C0",X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"2A",X"00",X"10",X"11",X"23",X"00",X"11",X"21",X"33",X"00",X"11",X"A1",X"33",X"00",X"13",
		X"21",X"13",X"00",X"13",X"21",X"23",X"00",X"13",X"21",X"13",X"00",X"13",X"A1",X"A3",X"11",X"13",
		X"21",X"13",X"DD",X"13",X"21",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"A1",X"A3",X"DD",X"13",
		X"21",X"13",X"DD",X"13",X"21",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"21",X"A3",X"22",X"13",
		X"A1",X"13",X"32",X"13",X"21",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"21",X"A3",X"33",X"13",
		X"21",X"13",X"33",X"13",X"A1",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"21",X"13",X"32",X"13",
		X"21",X"13",X"22",X"13",X"A1",X"D2",X"DD",X"13",X"21",X"11",X"11",X"13",X"21",X"00",X"00",X"13",
		X"A1",X"00",X"00",X"13",X"21",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"10",
		X"11",X"11",X"11",X"10",X"DD",X"DD",X"DD",X"11",X"33",X"33",X"33",X"31",X"11",X"11",X"11",X"11",
		X"22",X"22",X"2A",X"A2",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"11",X"13",X"33",X"22",X"10",
		X"11",X"11",X"32",X"00",X"00",X"DD",X"33",X"00",X"00",X"DD",X"3D",X"00",X"00",X"DD",X"3D",X"00",
		X"00",X"DD",X"33",X"00",X"00",X"DD",X"3D",X"00",X"A0",X"DD",X"3D",X"00",X"10",X"DD",X"33",X"00",
		X"12",X"12",X"32",X"00",X"33",X"33",X"22",X"00",X"33",X"33",X"33",X"00",X"12",X"12",X"12",X"00",
		X"10",X"DD",X"DD",X"00",X"A0",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"11",X"11",X"11",X"00",
		X"13",X"33",X"33",X"10",X"33",X"33",X"33",X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"2A",X"A2",
		X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"31",X"DD",X"DD",X"DD",X"11",X"11",X"11",X"11",X"10",
		X"55",X"00",X"00",X"55",X"CC",X"00",X"00",X"A5",X"CC",X"00",X"00",X"5C",X"CC",X"00",X"00",X"5C",
		X"6C",X"00",X"00",X"5C",X"CC",X"00",X"00",X"55",X"CC",X"00",X"00",X"A5",X"CC",X"22",X"00",X"5C",
		X"CC",X"22",X"22",X"5C",X"6C",X"2C",X"22",X"5C",X"CC",X"C7",X"22",X"55",X"CC",X"C7",X"22",X"A5",
		X"CC",X"77",X"C2",X"5C",X"CC",X"77",X"7C",X"5C",X"6C",X"75",X"77",X"5C",X"CC",X"55",X"77",X"55",
		X"CC",X"55",X"57",X"A5",X"CC",X"55",X"55",X"5C",X"CC",X"55",X"55",X"5C",X"6C",X"55",X"55",X"5C",
		X"CC",X"55",X"55",X"55",X"CC",X"55",X"57",X"A5",X"CC",X"55",X"77",X"5C",X"CC",X"75",X"7C",X"5C",
		X"6C",X"77",X"7C",X"5C",X"CC",X"CC",X"CC",X"55",X"CC",X"22",X"70",X"A5",X"CC",X"22",X"70",X"5C",
		X"CC",X"77",X"70",X"55",X"C5",X"C0",X"70",X"55",X"55",X"00",X"70",X"50",X"55",X"00",X"70",X"05",
		X"2C",X"55",X"C2",X"55",X"2C",X"55",X"C2",X"55",X"CC",X"5C",X"C5",X"25",X"55",X"A5",X"55",X"55",
		X"C6",X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"A6",X"66",X"6C",X"5C",X"CC",X"CC",X"C5",
		X"55",X"55",X"CC",X"50",X"00",X"55",X"77",X"00",X"00",X"55",X"55",X"00",X"00",X"5C",X"55",X"77",
		X"00",X"C7",X"55",X"27",X"00",X"77",X"55",X"27",X"00",X"C7",X"55",X"27",X"00",X"7C",X"55",X"27",
		X"00",X"7C",X"55",X"27",X"00",X"C7",X"55",X"27",X"00",X"77",X"55",X"27",X"00",X"C7",X"55",X"27",
		X"00",X"5C",X"55",X"77",X"00",X"55",X"55",X"00",X"00",X"55",X"77",X"00",X"05",X"55",X"CC",X"50",
		X"55",X"CC",X"CC",X"C5",X"CC",X"A6",X"66",X"6C",X"CC",X"CC",X"CC",X"CC",X"C6",X"CC",X"6C",X"CC",
		X"55",X"A5",X"55",X"55",X"CC",X"5C",X"C5",X"25",X"2C",X"55",X"C2",X"55",X"CC",X"55",X"CC",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"A0",X"33",X"00",
		X"00",X"AF",X"33",X"00",X"00",X"AA",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"35",X"39",X"00",
		X"00",X"3A",X"93",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"93",X"00",
		X"00",X"99",X"33",X"00",X"00",X"39",X"35",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"A9",X"00",
		X"00",X"3F",X"AA",X"00",X"00",X"30",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"0E",X"00",X"32",X"00",X"EE",X"EE",X"23",X"22",X"EE",X"E0",X"32",
		X"22",X"EE",X"00",X"20",X"22",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"02",X"00",X"00",
		X"23",X"22",X"00",X"00",X"03",X"22",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"20",X"00",X"00",X"02",X"22",X"00",X"00",X"02",X"02",X"00",X"00",X"02",X"02",X"00",
		X"00",X"02",X"02",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"20",X"00",X"00",X"A6",X"20",X"00",X"00",X"26",X"00",
		X"00",X"00",X"26",X"70",X"00",X"00",X"27",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"7A",X"70",
		X"00",X"00",X"7A",X"00",X"00",X"00",X"AA",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"22",X"00",X"00",X"70",X"00",X"00",X"02",X"03",X"00",X"00",X"02",X"22",X"00",
		X"00",X"02",X"22",X"00",X"00",X"20",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"EE",X"00",X"00",X"2D",X"EB",X"00",X"00",
		X"22",X"DD",X"00",X"00",X"22",X"ED",X"00",X"00",X"72",X"ED",X"00",X"00",X"D7",X"DD",X"00",X"00",
		X"DD",X"EB",X"00",X"00",X"0D",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"02",X"22",X"00",
		X"00",X"02",X"22",X"00",X"00",X"00",X"03",X"00",X"00",X"07",X"70",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FC",X"70",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",
		X"00",X"00",X"C7",X"FF",X"00",X"00",X"FC",X"70",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",
		X"00",X"00",X"C7",X"7F",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"7F",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"7F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"2C",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"70",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",
		X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"FF",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"70",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"70",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"F7",X"00",X"00",X"FF",X"77",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"70",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"F7",X"00",X"00",X"FF",X"77",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"77",X"0F",X"00",X"00",X"77",X"FF",X"00",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F7",X"00",X"00",X"FC",X"F7",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",
		X"CC",X"77",X"FF",X"00",X"77",X"77",X"FC",X"F0",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F7",
		X"00",X"00",X"C7",X"F7",X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"00",X"00",X"00",X"7F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"7F",X"00",
		X"00",X"00",X"FC",X"00",X"00",X"00",X"C7",X"00",X"77",X"07",X"7C",X"00",X"CC",X"7F",X"7C",X"70",
		X"CC",X"7F",X"7C",X"70",X"77",X"07",X"7C",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"FC",X"00",
		X"00",X"00",X"7F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"99",X"30",X"33",X"99",X"99",X"93",
		X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"EE",X"44",X"E9",X"99",X"99",X"44",X"9E",X"99",X"99",
		X"C4",X"9E",X"99",X"33",X"44",X"E9",X"9E",X"EE",X"33",X"99",X"9E",X"99",X"00",X"99",X"39",X"33",
		X"00",X"33",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"33",X"00",X"00",
		X"EE",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",
		X"33",X"33",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"33",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"99",X"99",X"EE",X"33",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"99",X"44",X"E9",X"99",X"93",X"44",X"9E",X"99",X"30",
		X"C4",X"9E",X"99",X"30",X"44",X"E9",X"9E",X"93",X"33",X"99",X"9E",X"99",X"00",X"99",X"39",X"99",
		X"00",X"33",X"03",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"03",X"EE",X"00",X"00",
		X"39",X"9E",X"00",X"00",X"3E",X"39",X"00",X"00",X"E9",X"03",X"00",X"00",X"99",X"00",X"00",X"00",
		X"93",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"33",X"00",X"00",
		X"99",X"E9",X"00",X"00",X"33",X"E9",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E9",X"EE",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"4E",X"99",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"4E",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"EE",X"EE",X"00",X"EE",X"CC",X"C9",X"00",
		X"EE",X"EE",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"9E",X"CC",X"11",X"F9",X"9E",X"CC",X"11",X"F9",
		X"9E",X"CC",X"11",X"F9",X"99",X"CC",X"11",X"F9",X"CC",X"CC",X"AC",X"00",X"EE",X"EE",X"CC",X"00",
		X"EE",X"CC",X"C9",X"00",X"99",X"EE",X"EE",X"00",X"99",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"E9",X"00",X"00",X"EE",X"E9",X"00",
		X"00",X"EC",X"E9",X"00",X"00",X"EC",X"E9",X"00",X"00",X"EC",X"E9",X"00",X"00",X"EC",X"E9",X"00",
		X"00",X"EC",X"C0",X"00",X"00",X"EC",X"C0",X"00",X"00",X"EC",X"C0",X"00",X"00",X"EC",X"CF",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"CA",X"CE",X"00",X"00",X"CC",X"9E",X"00",X"00",X"CC",X"90",X"00",X"00",X"C1",X"E0",X"00",
		X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F4",X"00",X"00",X"FF",X"77",X"77",X"00",X"77",X"CC",X"C4",X"00",
		X"77",X"77",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"F4",X"CC",X"44",X"44",X"F4",X"CC",X"44",X"44",
		X"F4",X"CC",X"44",X"44",X"FF",X"CC",X"44",X"44",X"CC",X"CC",X"CC",X"00",X"77",X"77",X"CC",X"00",
		X"77",X"CC",X"C4",X"00",X"FF",X"77",X"77",X"00",X"FF",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"7F",X"00",X"00",X"77",X"7F",X"00",
		X"00",X"7C",X"7F",X"00",X"00",X"7C",X"7F",X"00",X"00",X"7C",X"7F",X"00",X"00",X"7C",X"7F",X"00",
		X"00",X"7C",X"C0",X"00",X"00",X"7C",X"C0",X"00",X"00",X"7C",X"C0",X"00",X"00",X"7C",X"CF",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"CC",X"C7",X"00",X"00",X"CC",X"C4",X"00",
		X"00",X"CC",X"C7",X"00",X"00",X"CC",X"47",X"00",X"00",X"CC",X"40",X"00",X"00",X"C4",X"70",X"00",
		X"00",X"CC",X"70",X"00",X"00",X"CC",X"70",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"31",X"31",X"31",X"03",X"13",X"13",X"13",X"11",X"31",X"31",X"30",X"11",X"11",X"11",X"10",
		X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"35",X"35",X"35",X"30",
		X"53",X"53",X"53",X"50",X"35",X"35",X"35",X"30",X"53",X"53",X"53",X"50",X"35",X"35",X"35",X"30",
		X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"B0",X"DB",X"DB",X"DB",X"D0",X"BD",X"BD",X"BD",X"B0",
		X"DB",X"DB",X"DB",X"D0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",
		X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"DF",X"DF",X"DF",X"D0",X"0D",X"FD",X"FD",X"FD",X"0F",X"DF",X"DF",X"DF",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"40",
		X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"50",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F5",X"00",X"EA",X"00",X"00",X"00",X"09",X"00",X"FA",X"75",X"A0",
		X"00",X"05",X"07",X"09",X"A0",X"00",X"00",X"97",X"AF",X"00",X"0F",X"00",X"00",X"B0",X"F0",X"00",
		X"40",X"09",X"09",X"00",X"0A",X"A0",X"90",X"00",X"20",X"0B",X"00",X"A5",X"00",X"E0",X"00",X"00",
		X"00",X"02",X"9A",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"0A",X"00",X"90",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"92",X"00",X"00",
		X"09",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"B2",X"00",X"00",X"05",X"0B",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"E3",X"00",X"00",
		X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"04",X"44",X"44",X"00",X"00",
		X"44",X"04",X"00",X"00",X"44",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"07",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"93",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"07",X"77",X"55",X"00",X"05",X"55",
		X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",
		X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",
		X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"55",X"05",X"00",X"55",X"00",X"5C",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"CC",X"55",X"CC",X"C5",
		X"CC",X"00",X"5C",X"C5",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"50",
		X"00",X"00",X"50",X"C5",X"00",X"00",X"50",X"C5",X"00",X"00",X"50",X"CC",X"00",X"00",X"50",X"CC",
		X"00",X"00",X"50",X"CC",X"00",X"00",X"50",X"CC",X"00",X"00",X"50",X"C5",X"00",X"00",X"50",X"C5",
		X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
