`define BUILD_DATE "181123"
`define BUILD_TIME "011223"
