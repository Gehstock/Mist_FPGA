library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_bg_bits_2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"55",X"55",X"55",X"59",X"95",X"55",X"55",X"15",X"55",X"56",X"A5",X"5A",X"A9",X"55",X"55",
		X"55",X"55",X"66",X"56",X"55",X"AA",X"55",X"65",X"55",X"95",X"51",X"65",X"45",X"66",X"95",X"55",
		X"55",X"55",X"55",X"04",X"11",X"6A",X"56",X"55",X"56",X"54",X"41",X"15",X"45",X"69",X"69",X"55",
		X"55",X"11",X"54",X"14",X"54",X"59",X"66",X"95",X"55",X"44",X"50",X"05",X"55",X"64",X"5A",X"95",
		X"55",X"15",X"11",X"10",X"69",X"A5",X"56",X"95",X"55",X"51",X"55",X"54",X"6A",X"85",X"12",X"65",
		X"55",X"55",X"00",X"50",X"16",X"61",X"4A",X"95",X"55",X"51",X"51",X"66",X"55",X"50",X"19",X"95",
		X"55",X"55",X"45",X"9A",X"55",X"61",X"5A",X"55",X"55",X"55",X"56",X"55",X"55",X"54",X"55",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"12",X"65",X"55",X"55",X"55",X"5A",X"A5",
		X"56",X"55",X"6A",X"55",X"D9",X"95",X"59",X"69",X"55",X"46",X"5A",X"5A",X"A9",X"65",X"65",X"69",
		X"54",X"43",X"96",X"51",X"AA",X"55",X"51",X"A6",X"55",X"44",X"4A",X"65",X"56",X"A5",X"06",X"6A",
		X"57",X"14",X"56",X"81",X"51",X"A6",X"21",X"29",X"56",X"05",X"55",X"15",X"45",X"69",X"5A",X"69",
		X"59",X"11",X"16",X"05",X"55",X"6A",X"41",X"A5",X"56",X"21",X"4B",X"05",X"15",X"1A",X"56",X"55",
		X"54",X"51",X"99",X"90",X"50",X"5A",X"51",X"55",X"55",X"72",X"55",X"42",X"55",X"99",X"75",X"55",
		X"55",X"55",X"54",X"59",X"13",X"A5",X"55",X"55",X"55",X"55",X"55",X"54",X"45",X"A5",X"55",X"55",
		X"55",X"55",X"55",X"56",X"16",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"2A",X"59",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"65",X"55",
		X"55",X"57",X"55",X"55",X"59",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"56",X"55",X"57",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"56",X"55",X"55",X"75",X"55",
		X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"0D",X"D7",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"DD",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"03",X"75",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"0F",X"7D",X"DD",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"37",X"77",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"57",X"7C",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"57",X"DF",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"F7",X"C0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"77",X"DF",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"DF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"00",X"55",X"55",X"55",
		X"55",X"55",X"55",X"40",X"00",X"04",X"55",X"55",X"55",X"55",X"55",X"55",X"44",X"00",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",
		X"00",X"00",X"00",X"00",X"10",X"41",X"00",X"04",X"00",X"04",X"00",X"41",X"00",X"04",X"44",X"11",
		X"41",X"10",X"51",X"00",X"11",X"01",X"15",X"45",X"10",X"11",X"44",X"45",X"05",X"C5",X"51",X"55",
		X"44",X"41",X"11",X"44",X"55",X"54",X"55",X"55",X"45",X"14",X"45",X"15",X"51",X"5D",X"55",X"55",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D1",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"45",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"55",X"56",X"55",X"65",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"59",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"54",X"00",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"01",X"15",X"55",
		X"55",X"55",X"55",X"55",X"51",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"37",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"03",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"37",X"75",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"03",X"75",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"03",X"77",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"FC",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"57",X"F0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"5F",X"FC",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"FC",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",
		X"00",X"00",X"00",X"00",X"10",X"41",X"00",X"04",X"00",X"04",X"00",X"41",X"00",X"04",X"44",X"11",
		X"41",X"10",X"51",X"00",X"11",X"01",X"15",X"45",X"10",X"11",X"44",X"45",X"05",X"C5",X"51",X"55",
		X"44",X"41",X"11",X"44",X"55",X"54",X"55",X"55",X"45",X"14",X"45",X"15",X"51",X"5D",X"55",X"55",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D1",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"45",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"55",X"56",X"55",X"65",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"37",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"03",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"37",X"75",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"03",X"75",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"03",X"77",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"FC",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"57",X"F0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"5F",X"FC",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"FC",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"54",X"00",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"01",X"15",X"55",
		X"55",X"55",X"55",X"55",X"51",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",
		X"00",X"00",X"00",X"00",X"10",X"41",X"00",X"04",X"00",X"04",X"00",X"41",X"00",X"04",X"44",X"11",
		X"41",X"10",X"51",X"00",X"11",X"01",X"15",X"45",X"10",X"11",X"44",X"45",X"05",X"C5",X"51",X"55",
		X"44",X"41",X"11",X"44",X"55",X"54",X"55",X"55",X"45",X"14",X"45",X"15",X"51",X"5D",X"55",X"55",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D1",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"45",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"55",X"56",X"55",X"65",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"47",X"56",X"44",X"A9",X"55",X"55",X"50",X"00",X"07",X"D6",X"52",X"55",X"55",X"55",X"54",X"30",
		X"0D",X"5A",X"55",X"55",X"55",X"55",X"54",X"00",X"0F",X"66",X"55",X"55",X"75",X"55",X"54",X"00",
		X"0D",X"5A",X"A8",X"55",X"DF",X"55",X"54",X"30",X"05",X"5A",X"A9",X"45",X"75",X"55",X"54",X"10",
		X"04",X"7A",X"66",X"54",X"5D",X"D7",X"54",X"40",X"15",X"4A",X"A5",X"95",X"57",X"55",X"50",X"00",
		X"05",X"36",X"AA",X"A5",X"45",X"5D",X"50",X"0C",X"14",X"99",X"B5",X"59",X"55",X"D5",X"41",X"00",
		X"11",X"A6",X"AB",X"6A",X"55",X"75",X"50",X"C0",X"10",X"49",X"2D",X"96",X"95",X"77",X"40",X"00",
		X"00",X"69",X"AB",X"99",X"A7",X"55",X"07",X"00",X"01",X"99",X"5A",X"B5",X"EA",X"5C",X"00",X"00",
		X"06",X"16",X"6A",X"AB",X"69",X"50",X"40",X"00",X"05",X"49",X"56",X"9D",X"DD",X"44",X"0C",X"00",
		X"05",X"66",X"5A",X"BD",X"75",X"5C",X"00",X"00",X"09",X"55",X"56",X"BD",X"D7",X"40",X"30",X"00",
		X"05",X"55",X"67",X"DF",X"F5",X"10",X"00",X"00",X"0F",X"65",X"55",X"5F",X"C5",X"13",X"00",X"00",
		X"07",X"56",X"5D",X"D7",X"75",X"40",X"00",X"00",X"03",X"F5",X"57",X"33",X"C0",X"00",X"00",X"00",
		X"00",X"F9",X"55",X"10",X"04",X"43",X"00",X"00",X"00",X"F5",X"54",X"40",X"00",X"40",X"00",X"00",
		X"00",X"F7",X"75",X"01",X"04",X"40",X"00",X"00",X"00",X"3D",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3D",X"D4",X"03",X"00",X"0C",X"00",X"00",X"00",X"0F",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"40",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"0C",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"30",X"00",X"00",X"00",X"00",X"00",X"30",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"54",X"03",X"C0",X"4C",X"00",X"00",X"03",X"01",X"15",X"00",X"04",X"03",X"00",X"00",
		X"00",X"05",X"55",X"C3",X"C0",X"00",X"00",X"00",X"00",X"15",X"55",X"40",X"11",X"00",X"C0",X"00",
		X"30",X"15",X"55",X"43",X"04",X"50",X"00",X"C0",X"00",X"55",X"45",X"00",X"05",X"40",X"00",X"00",
		X"00",X"55",X"45",X"40",X"05",X"40",X"C0",X"00",X"01",X"55",X"55",X"50",X"15",X"44",X"00",X"30",
		X"01",X"44",X"45",X"54",X"15",X"40",X"30",X"00",X"0D",X"55",X"55",X"50",X"15",X"50",X"00",X"00",
		X"05",X"45",X"55",X"54",X"55",X"50",X"00",X"30",X"07",X"14",X"55",X"54",X"55",X"54",X"00",X"00",
		X"01",X"55",X"55",X"55",X"55",X"50",X"30",X"30",X"14",X"15",X"56",X"95",X"55",X"54",X"00",X"00",
		X"14",X"51",X"59",X"57",X"55",X"54",X"0C",X"00",X"10",X"55",X"65",X"55",X"55",X"54",X"00",X"00",
		X"54",X"51",X"66",X"55",X"55",X"54",X"40",X"03",X"49",X"55",X"55",X"55",X"45",X"54",X"03",X"00",
		X"55",X"95",X"66",X"A4",X"55",X"55",X"00",X"03",X"26",X"59",X"95",X"95",X"55",X"55",X"00",X"00",
		X"16",X"95",X"5A",X"54",X"55",X"55",X"50",X"00",X"3A",X"A6",X"66",X"51",X"55",X"55",X"00",X"C0",
		X"06",X"99",X"A9",X"15",X"55",X"55",X"10",X"00",X"0E",X"A6",X"A8",X"45",X"55",X"55",X"50",X"00",
		X"0D",X"6A",X"A5",X"14",X"55",X"55",X"50",X"0C",X"01",X"AA",X"A1",X"55",X"54",X"55",X"54",X"00",
		X"03",X"6A",X"D4",X"45",X"51",X"55",X"50",X"40",X"03",X"5A",X"51",X"11",X"15",X"55",X"54",X"00",
		X"55",X"55",X"55",X"55",X"6A",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A5",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5A",X"91",X"55",X"55",X"55",X"55",X"55",X"45",X"52",X"95",X"44",X"55",
		X"55",X"55",X"55",X"51",X"56",X"91",X"55",X"55",X"55",X"55",X"44",X"54",X"5A",X"54",X"45",X"45",
		X"55",X"54",X"51",X"15",X"56",X"55",X"54",X"55",X"55",X"55",X"15",X"15",X"55",X"51",X"55",X"55",
		X"55",X"55",X"01",X"54",X"65",X"51",X"52",X"55",X"55",X"55",X"41",X"46",X"95",X"54",X"0A",X"95",
		X"55",X"15",X"50",X"55",X"65",X"11",X"5A",X"95",X"55",X"55",X"51",X"55",X"95",X"55",X"12",X"55",
		X"51",X"11",X"55",X"45",X"59",X"45",X"55",X"95",X"54",X"55",X"55",X"54",X"55",X"55",X"41",X"59",
		X"54",X"55",X"51",X"45",X"5A",X"95",X"55",X"59",X"55",X"05",X"55",X"54",X"59",X"95",X"55",X"69",
		X"55",X"55",X"56",X"45",X"66",X"51",X"56",X"65",X"55",X"55",X"55",X"51",X"56",X"55",X"55",X"65",
		X"54",X"55",X"46",X"64",X"59",X"15",X"45",X"85",X"55",X"44",X"54",X"56",X"59",X"51",X"56",X"55",
		X"55",X"55",X"41",X"9A",X"A5",X"11",X"59",X"92",X"11",X"54",X"40",X"9A",X"95",X"55",X"45",X"69",
		X"54",X"54",X"52",X"5A",X"A4",X"11",X"45",X"65",X"15",X"56",X"15",X"5A",X"A9",X"54",X"55",X"95",
		X"45",X"46",X"85",X"6A",X"54",X"14",X"12",X"51",X"11",X"5A",X"A4",X"A5",X"56",X"15",X"55",X"15",
		X"44",X"5A",X"5A",X"95",X"55",X"84",X"49",X"85",X"A1",X"29",X"55",X"55",X"55",X"62",X"55",X"82",
		X"5A",X"95",X"55",X"55",X"55",X"59",X"86",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"C3",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"04",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"00",X"10",X"00",X"00",X"10",X"04",X"44",
		X"01",X"10",X"45",X"01",X"10",X"00",X"41",X"01",X"55",X"55",X"40",X"10",X"01",X"04",X"54",X"51",
		X"15",X"54",X"51",X"00",X"45",X"55",X"55",X"54",X"55",X"51",X"54",X"44",X"11",X"15",X"55",X"55",
		X"55",X"55",X"55",X"00",X"54",X"54",X"55",X"55",X"55",X"55",X"54",X"44",X"55",X"55",X"45",X"55",
		X"55",X"55",X"55",X"15",X"5D",X"51",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"15",X"55",
		X"55",X"54",X"00",X"00",X"00",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"54",X"55",X"65",X"51",X"95",X"51",X"51",X"55",X"55",X"55",X"59",X"95",X"59",X"55",
		X"15",X"51",X"55",X"55",X"55",X"55",X"5A",X"55",X"51",X"55",X"51",X"15",X"56",X"55",X"55",X"55",
		X"55",X"95",X"55",X"55",X"55",X"55",X"91",X"65",X"55",X"59",X"51",X"51",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"15",X"55",X"55",X"99",X"55",X"55",X"5A",X"91",X"45",X"55",X"55",X"65",X"55",
		X"59",X"A9",X"96",X"11",X"56",X"55",X"96",X"55",X"55",X"6A",X"55",X"45",X"59",X"54",X"55",X"55",
		X"55",X"59",X"55",X"9A",X"A9",X"15",X"59",X"95",X"45",X"56",X"55",X"56",X"A5",X"45",X"15",X"59",
		X"55",X"56",X"51",X"65",X"95",X"51",X"66",X"59",X"55",X"5A",X"55",X"56",X"66",X"44",X"55",X"55",
		X"45",X"59",X"45",X"55",X"65",X"55",X"69",X"55",X"55",X"59",X"54",X"59",X"95",X"A9",X"95",X"15",
		X"11",X"59",X"41",X"56",X"91",X"6A",X"51",X"55",X"45",X"5A",X"54",X"66",X"16",X"6A",X"A5",X"45",
		X"54",X"6A",X"91",X"56",X"59",X"AA",X"68",X"55",X"46",X"AA",X"A4",X"9A",X"46",X"A9",X"66",X"55",
		X"56",X"A9",X"61",X"6A",X"9A",X"65",X"55",X"85",X"56",X"95",X"58",X"A9",X"65",X"55",X"55",X"65",
		X"6A",X"55",X"56",X"95",X"55",X"55",X"55",X"65",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"59",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",X"55",
		X"59",X"59",X"55",X"55",X"55",X"69",X"55",X"55",X"65",X"56",X"55",X"51",X"15",X"59",X"51",X"55",
		X"55",X"55",X"59",X"55",X"55",X"99",X"55",X"55",X"54",X"55",X"59",X"54",X"55",X"99",X"14",X"55",
		X"55",X"55",X"59",X"15",X"55",X"65",X"51",X"45",X"55",X"69",X"69",X"55",X"55",X"A5",X"55",X"55",
		X"15",X"59",X"55",X"45",X"55",X"95",X"61",X"15",X"55",X"5A",X"A5",X"54",X"59",X"55",X"58",X"55",
		X"55",X"55",X"91",X"55",X"65",X"55",X"54",X"95",X"11",X"55",X"55",X"55",X"55",X"55",X"56",X"85",
		X"55",X"45",X"64",X"55",X"55",X"55",X"56",X"99",X"54",X"55",X"61",X"51",X"54",X"55",X"55",X"A5",
		X"55",X"55",X"94",X"45",X"55",X"55",X"55",X"69",X"5A",X"55",X"A5",X"95",X"55",X"15",X"55",X"65",
		X"69",X"56",X"AA",X"95",X"55",X"55",X"95",X"69",X"69",X"55",X"9A",X"65",X"51",X"5A",X"45",X"55",
		X"65",X"55",X"6A",X"A5",X"55",X"6A",X"51",X"65",X"55",X"55",X"69",X"A5",X"45",X"59",X"44",X"55",
		X"55",X"15",X"5A",X"55",X"15",X"55",X"51",X"55",X"51",X"55",X"59",X"55",X"55",X"55",X"50",X"55",
		X"55",X"55",X"59",X"15",X"15",X"15",X"55",X"55",X"45",X"15",X"65",X"55",X"45",X"55",X"15",X"55",
		X"51",X"55",X"65",X"55",X"41",X"55",X"55",X"55",X"55",X"19",X"94",X"55",X"A4",X"45",X"51",X"55",
		X"44",X"65",X"51",X"59",X"59",X"54",X"15",X"15",X"51",X"55",X"44",X"55",X"56",X"95",X"55",X"55",
		X"44",X"55",X"51",X"51",X"51",X"54",X"11",X"55",X"51",X"51",X"55",X"15",X"45",X"55",X"55",X"15",
		X"55",X"15",X"55",X"54",X"51",X"55",X"44",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"DC",
		X"55",X"55",X"55",X"5D",X"F7",X"DF",X"00",X"00",X"77",X"7D",X"F7",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"40",X"00",X"04",X"55",X"55",X"55",X"55",X"55",X"55",X"44",X"00",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"0D",X"D7",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"DD",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"03",X"75",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"0F",X"7D",X"DD",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"37",X"77",X"55",X"00",X"00",X"00",X"00",X"00",X"0D",X"DD",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"57",X"7C",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"57",X"DF",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"F7",X"C0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"77",X"DF",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"DF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"00",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"44",X"50",X"00",X"10",
		X"01",X"10",X"54",X"45",X"15",X"45",X"14",X"45",X"10",X"45",X"31",X"55",X"47",X"55",X"45",X"55",
		X"45",X"54",X"55",X"11",X"55",X"55",X"55",X"75",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"45",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"C0",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"01",X"04",X"04",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"00",X"C0",X"00",X"11",X"11",X"44",X"40",
		X"00",X"00",X"00",X"04",X"41",X"55",X"01",X"10",X"00",X"C0",X"00",X"00",X"15",X"55",X"15",X"00",
		X"00",X"00",X"00",X"11",X"15",X"55",X"54",X"44",X"00",X"0C",X"00",X"00",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"10",X"05",X"55",X"55",X"55",X"00",X"00",X"10",X"41",X"55",X"55",X"5D",X"55",
		X"00",X"00",X"00",X"04",X"55",X"55",X"55",X"55",X"30",X"00",X"00",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"0D",X"D7",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"DD",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"03",X"75",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"0F",X"7D",X"DD",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"37",X"77",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"D5",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"57",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"57",X"DF",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"F7",X"C0",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"77",X"DF",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"DF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"11",X"55",X"55",X"55",X"55",
		X"55",X"55",X"50",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"04",X"55",X"55",
		X"55",X"55",X"55",X"55",X"44",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"95",X"55",X"44",X"55",X"55",X"55",X"55",X"55",X"95",X"59",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"55",X"95",X"55",X"59",X"95",X"55",X"56",X"44",X"56",X"59",X"55",X"55",X"95",
		X"55",X"56",X"55",X"55",X"65",X"45",X"55",X"59",X"55",X"56",X"14",X"55",X"58",X"55",X"51",X"59",
		X"55",X"56",X"45",X"55",X"95",X"51",X"55",X"56",X"55",X"58",X"54",X"55",X"64",X"14",X"54",X"55",
		X"55",X"59",X"45",X"45",X"54",X"55",X"55",X"55",X"55",X"58",X"51",X"15",X"94",X"54",X"55",X"65",
		X"55",X"56",X"24",X"55",X"55",X"15",X"51",X"55",X"55",X"55",X"9A",X"55",X"55",X"85",X"96",X"55",
		X"55",X"55",X"56",X"45",X"55",X"64",X"6A",X"65",X"55",X"55",X"55",X"A8",X"56",X"65",X"5A",X"55",
		X"55",X"55",X"55",X"56",X"15",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"95",X"56",X"65",X"55",
		X"55",X"55",X"55",X"55",X"91",X"45",X"56",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"99",X"51",
		X"55",X"55",X"55",X"58",X"55",X"51",X"64",X"55",X"55",X"55",X"55",X"58",X"51",X"56",X"65",X"51",
		X"55",X"55",X"55",X"56",X"11",X"15",X"A6",X"55",X"55",X"55",X"55",X"55",X"84",X"59",X"95",X"11",
		X"55",X"55",X"55",X"55",X"91",X"46",X"A1",X"55",X"55",X"55",X"55",X"55",X"85",X"69",X"65",X"15",
		X"55",X"55",X"55",X"55",X"69",X"95",X"68",X"45",X"55",X"55",X"55",X"55",X"56",X"55",X"59",X"11",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"40",X"00",X"00",
		X"15",X"14",X"11",X"04",X"04",X"00",X"04",X"00",X"45",X"50",X"55",X"44",X"41",X"00",X"40",X"10",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"04",X"14",X"55",X"55",X"44",X"15",X"55",X"45",X"50",
		X"55",X"55",X"55",X"55",X"5D",X"50",X"54",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"4C",X"44",
		X"75",X"55",X"55",X"55",X"55",X"55",X"51",X"51",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"54",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",
		X"44",X"50",X"40",X"10",X"40",X"40",X"00",X"40",X"15",X"54",X"11",X"04",X"04",X"00",X"04",X"00",
		X"45",X"55",X"55",X"44",X"51",X"14",X"40",X"10",X"55",X"55",X"55",X"15",X"15",X"55",X"11",X"04",
		X"15",X"55",X"55",X"45",X"55",X"55",X"45",X"50",X"55",X"55",X"55",X"55",X"5D",X"55",X"54",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"45",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"C0",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"10",X"40",X"00",X"00",X"00",
		X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"44",X"44",X"00",X"03",X"00",X"00",
		X"04",X"40",X"55",X"41",X"10",X"00",X"00",X"00",X"00",X"54",X"55",X"54",X"00",X"00",X"00",X"00",
		X"11",X"15",X"55",X"54",X"44",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"30",X"00",
		X"55",X"55",X"55",X"50",X"04",X"00",X"00",X"00",X"55",X"75",X"55",X"55",X"41",X"04",X"00",X"00",
		X"55",X"55",X"55",X"55",X"10",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"44",X"50",X"40",X"10",X"40",X"40",X"00",X"40",
		X"15",X"54",X"11",X"04",X"04",X"00",X"04",X"00",X"45",X"55",X"55",X"44",X"51",X"14",X"40",X"10",
		X"55",X"55",X"55",X"15",X"15",X"55",X"11",X"04",X"15",X"55",X"55",X"45",X"55",X"55",X"45",X"50",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"54",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"45",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5A",X"56",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"A6",X"AA",X"95",
		X"55",X"55",X"55",X"55",X"65",X"AA",X"AA",X"65",X"55",X"55",X"45",X"55",X"55",X"6A",X"AA",X"95",
		X"54",X"55",X"51",X"45",X"59",X"6A",X"A9",X"55",X"55",X"55",X"45",X"55",X"55",X"96",X"AA",X"95",
		X"55",X"45",X"51",X"55",X"46",X"56",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"95",
		X"55",X"15",X"55",X"44",X"55",X"5A",X"A9",X"55",X"55",X"55",X"55",X"51",X"45",X"6A",X"A9",X"55",
		X"55",X"15",X"55",X"44",X"15",X"6A",X"A5",X"55",X"94",X"51",X"55",X"54",X"55",X"A9",X"55",X"55",
		X"65",X"95",X"55",X"68",X"11",X"A5",X"55",X"55",X"59",X"A5",X"51",X"AA",X"56",X"95",X"55",X"55",
		X"59",X"59",X"56",X"65",X"A9",X"55",X"55",X"55",X"55",X"6A",X"5A",X"A5",X"55",X"55",X"55",X"55",
		X"55",X"96",X"AA",X"95",X"55",X"55",X"55",X"55",X"56",X"56",X"AA",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"14",X"55",X"AA",X"95",X"55",X"55",X"55",X"55",
		X"54",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"A9",X"95",X"55",X"55",X"55",X"55",
		X"15",X"06",X"A6",X"55",X"55",X"55",X"55",X"55",X"56",X"A6",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"45",X"45",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5C",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"44",X"54",X"55",X"11",X"55",X"55",X"55",X"75",
		X"01",X"05",X"31",X"55",X"47",X"55",X"55",X"55",X"04",X"40",X"54",X"45",X"15",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",X"00",X"04",X"04",X"11",X"00",X"05",X"05",X"45",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"45",X"55",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5C",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"44",X"54",X"55",X"11",X"55",X"55",X"55",X"75",
		X"01",X"05",X"31",X"55",X"47",X"55",X"55",X"55",X"04",X"40",X"54",X"45",X"15",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",X"00",X"04",X"04",X"11",X"00",X"05",X"05",X"45",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"41",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"04",X"03",X"00",X"00",X"00",X"10",X"01",X"01",X"50",X"40",X"00",X"00",
		X"00",X"00",X"00",X"05",X"55",X"00",X"00",X"40",X"01",X"00",X"44",X"55",X"55",X"54",X"10",X"00",
		X"10",X"10",X"01",X"11",X"51",X"10",X"00",X"10",X"55",X"54",X"54",X"55",X"55",X"54",X"11",X"00",
		X"05",X"45",X"55",X"55",X"55",X"55",X"41",X"40",X"55",X"15",X"15",X"55",X"51",X"55",X"50",X"55",
		X"51",X"55",X"55",X"55",X"55",X"51",X"45",X"54",X"15",X"55",X"54",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"55",X"55",
		X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"54",X"54",X"55",X"11",X"55",X"55",X"55",X"75",
		X"01",X"05",X"31",X"55",X"47",X"55",X"55",X"55",X"44",X"40",X"54",X"45",X"15",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",X"01",X"04",X"04",X"11",X"00",X"05",X"05",X"45",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"45",X"55",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"54",X"54",X"55",X"11",X"55",X"55",X"55",X"75",X"01",X"05",X"31",X"55",X"47",X"55",X"55",X"55",
		X"44",X"40",X"54",X"45",X"15",X"45",X"55",X"55",X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",
		X"01",X"04",X"04",X"11",X"00",X"05",X"05",X"45",X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",
		X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"14",X"54",X"55",X"55",X"55",X"55",X"55",X"75",X"45",X"05",X"31",X"55",X"57",X"55",X"55",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"40",X"40",X"40",X"10",X"00",X"41",X"01",X"01",X"11",X"04",X"11",X"04",X"04",X"10",X"10",X"44",
		X"44",X"10",X"50",X"44",X"41",X"00",X"44",X"11",X"45",X"45",X"05",X"11",X"10",X"44",X"11",X"05",
		X"15",X"55",X"55",X"44",X"15",X"51",X"55",X"54",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"14",X"54",X"55",X"55",X"55",X"55",X"55",X"75",
		X"45",X"05",X"31",X"55",X"57",X"55",X"55",X"55",X"04",X"40",X"54",X"45",X"55",X"55",X"55",X"55",
		X"00",X"00",X"01",X"04",X"54",X"55",X"55",X"55",X"11",X"04",X"04",X"11",X"10",X"45",X"45",X"55",
		X"00",X"10",X"00",X"00",X"01",X"00",X"51",X"55",X"00",X"00",X"00",X"40",X"10",X"11",X"05",X"54",
		X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"45",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"44",X"44",
		X"00",X"00",X"00",X"11",X"10",X"00",X"01",X"01",X"00",X"00",X"00",X"10",X"01",X"04",X"54",X"11",
		X"00",X"00",X"51",X"00",X"45",X"54",X"45",X"54",X"00",X"01",X"44",X"44",X"11",X"15",X"54",X"45",
		X"00",X"10",X"41",X"10",X"54",X"44",X"15",X"55",X"00",X"45",X"51",X"44",X"45",X"55",X"45",X"55",
		X"00",X"14",X"44",X"55",X"5D",X"50",X"55",X"75",X"01",X"D5",X"5D",X"5D",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"15",X"55",X"55",X"55",X"5D",X"55",X"55",X"51",X"55",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"05",X"51",X"45",X"55",X"55",X"D5",X"75",X"55",X"04",X"44",X"55",X"15",X"55",X"55",X"55",X"75",
		X"00",X"05",X"31",X"55",X"57",X"55",X"55",X"55",X"00",X"40",X"54",X"45",X"55",X"55",X"55",X"55",
		X"00",X"00",X"01",X"04",X"54",X"55",X"55",X"55",X"00",X"00",X"04",X"11",X"10",X"45",X"45",X"55",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"55",X"00",X"00",X"00",X"40",X"10",X"11",X"05",X"54",
		X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"45",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"04",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"04",X"00",X"00",X"44",X"50",X"44",X"10",X"50",X"41",X"01",X"01",
		X"15",X"15",X"11",X"44",X"05",X"10",X"10",X"44",X"55",X"55",X"55",X"44",X"41",X"41",X"44",X"11",
		X"55",X"55",X"55",X"55",X"14",X"54",X"51",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"30",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"01",X"1D",X"5D",X"75",X"75",X"55",X"57",X"55",X"0D",X"5D",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"05",X"45",X"55",X"55",X"55",X"55",X"55",X"75",X"04",X"55",X"55",X"55",X"57",X"55",X"55",X"55",
		X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5D",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"14",X"54",X"55",X"55",X"55",X"55",X"55",X"75",X"45",X"05",X"31",X"55",X"57",X"55",X"55",X"55",
		X"04",X"40",X"54",X"45",X"55",X"55",X"55",X"55",X"00",X"00",X"01",X"04",X"54",X"55",X"55",X"55",
		X"11",X"04",X"04",X"11",X"10",X"45",X"45",X"55",X"00",X"10",X"00",X"00",X"01",X"00",X"51",X"55",
		X"00",X"00",X"00",X"40",X"10",X"11",X"05",X"54",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"45",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"FC",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"57",X"F0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"5F",X"FC",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"FC",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"75",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"57",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"56",X"45",X"55",X"55",X"55",X"55",X"54",
		X"55",X"56",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"59",X"15",X"55",X"55",X"15",X"54",X"55",
		X"55",X"58",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"58",X"55",X"55",X"55",X"55",X"55",X"54",
		X"55",X"56",X"45",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"91",X"55",X"45",X"45",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"15",X"15",X"55",X"55",X"55",X"95",X"55",X"51",X"51",X"55",X"15",
		X"55",X"56",X"15",X"15",X"55",X"51",X"55",X"55",X"55",X"58",X"55",X"55",X"55",X"15",X"45",X"15",
		X"55",X"58",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"56",X"04",X"55",X"55",X"55",X"15",X"54",
		X"55",X"55",X"95",X"55",X"55",X"55",X"51",X"65",X"55",X"55",X"64",X"51",X"55",X"51",X"55",X"55",
		X"55",X"55",X"61",X"15",X"55",X"55",X"55",X"56",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"15",X"55",X"54",X"55",X"54",X"56",X"55",X"56",X"11",X"45",X"51",X"15",X"55",X"55",
		X"55",X"56",X"04",X"55",X"54",X"55",X"45",X"15",X"55",X"55",X"85",X"55",X"51",X"15",X"54",X"55",
		X"55",X"55",X"91",X"55",X"54",X"55",X"55",X"55",X"55",X"56",X"54",X"51",X"55",X"55",X"44",X"45",
		X"55",X"56",X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"59",X"55",X"15",X"51",X"55",X"51",X"41",
		X"55",X"65",X"55",X"54",X"55",X"55",X"51",X"55",X"55",X"59",X"55",X"55",X"54",X"55",X"55",X"15",
		X"55",X"5A",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"04",X"50",X"00",X"00",X"00",X"01",X"00",X"44",X"44",X"00",X"04",X"00",X"00",
		X"10",X"10",X"01",X"11",X"51",X"10",X"00",X"00",X"55",X"54",X"54",X"55",X"15",X"54",X"00",X"00",
		X"05",X"45",X"45",X"14",X"55",X"00",X"40",X"00",X"55",X"15",X"15",X"51",X"51",X"45",X"10",X"00",
		X"51",X"55",X"55",X"55",X"55",X"00",X"01",X"00",X"15",X"55",X"54",X"55",X"45",X"11",X"40",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"44",X"55",X"55",X"55",X"55",X"55",X"51",X"40",X"00",
		X"55",X"55",X"55",X"55",X"5D",X"15",X"44",X"50",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"55",X"04",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"57",X"FF",X"F0",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"5F",X"FF",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"0C",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"5D",X"D5",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"57",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"5D",X"51",X"04",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"17",X"10",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"71",X"51",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"11",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"20",X"00",X"00",X"00",X"00",
		X"00",X"03",X"E0",X"08",X"00",X"10",X"00",X"00",X"00",X"03",X"F8",X"02",X"00",X"00",X"08",X"00",
		X"00",X"00",X"FE",X"80",X"80",X"00",X"00",X"00",X"08",X"10",X"3F",X"E8",X"20",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"FE",X"88",X"00",X"80",X"40",X"00",X"00",X"00",X"CF",X"E0",X"80",X"00",X"00",
		X"02",X"00",X"80",X"0F",X"FA",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"FF",X"A0",X"00",X"00",
		X"00",X"3E",X"80",X"40",X"0F",X"FA",X"AA",X"AA",X"00",X"FA",X"00",X"00",X"0F",X"CF",X"FF",X"FC",
		X"0F",X"F8",X"04",X"00",X"00",X"0F",X"FF",X"FC",X"3E",X"E0",X"00",X"02",X"00",X"00",X"03",X"80",
		X"08",X"E0",X"00",X"00",X"00",X"00",X"03",X"00",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",
		X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",
		X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",
		X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",
		X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",
		X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",
		X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",
		X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",
		X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"69",X"55",X"55",X"55",X"5D",
		X"55",X"57",X"E5",X"5A",X"55",X"55",X"55",X"55",X"55",X"57",X"F9",X"56",X"95",X"55",X"56",X"55",
		X"55",X"55",X"FE",X"95",X"A5",X"59",X"55",X"55",X"56",X"55",X"7F",X"E9",X"69",X"55",X"55",X"55",
		X"55",X"55",X"5F",X"FE",X"9A",X"55",X"55",X"55",X"55",X"55",X"55",X"DF",X"E5",X"95",X"D5",X"55",
		X"55",X"55",X"75",X"5F",X"FA",X"65",X"55",X"55",X"55",X"5F",X"95",X"55",X"FF",X"A9",X"55",X"55",
		X"65",X"7E",X"95",X"55",X"5F",X"FA",X"AA",X"AA",X"55",X"FA",X"55",X"55",X"5F",X"DF",X"FF",X"FD",
		X"5F",X"F9",X"55",X"95",X"55",X"5F",X"FF",X"FD",X"7E",X"E5",X"55",X"55",X"55",X"55",X"57",X"95",
		X"59",X"E5",X"55",X"55",X"55",X"55",X"57",X"15",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"11",X"10",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"55",X"55",X"55",X"55",X"55",X"51",X"51",X"84",
		X"55",X"55",X"55",X"55",X"55",X"55",X"14",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"04",X"55",X"55",X"55",X"55",X"55",X"55",X"14",X"80",
		X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"10",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",
		X"55",X"55",X"55",X"55",X"55",X"51",X"51",X"04",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"70",
		X"55",X"55",X"55",X"55",X"55",X"55",X"14",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"10",
		X"55",X"55",X"55",X"55",X"55",X"54",X"44",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"44",
		X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"44",X"60",
		X"55",X"55",X"55",X"55",X"55",X"45",X"51",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"14",X"90",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"56",X"D5",X"55",X"55",X"55",X"55",X"8B",X"00",
		X"54",X"D5",X"55",X"55",X"55",X"55",X"8B",X"00",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"15",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"15",X"55",X"55",X"55",X"45",
		X"00",X"10",X"40",X"45",X"55",X"55",X"75",X"75",X"00",X"00",X"04",X"15",X"55",X"75",X"55",X"15",
		X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"00",X"30",X"44",X"55",X"55",X"55",X"55",X"55",
		X"01",X"04",X"11",X"55",X"55",X"55",X"55",X"55",X"00",X"01",X"54",X"55",X"75",X"55",X"55",X"55",
		X"00",X"04",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"01",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"00",X"05",X"15",X"55",X"55",X"55",X"55",X"55",X"30",X"11",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"45",X"15",X"55",X"57",X"55",X"55",X"55",X"00",X"14",X"55",X"55",X"55",X"55",X"55",X"55",
		X"51",X"11",X"04",X"11",X"10",X"00",X"00",X"00",X"55",X"55",X"10",X"40",X"01",X"10",X"00",X"00",
		X"55",X"55",X"55",X"04",X"50",X"40",X"10",X"00",X"55",X"55",X"54",X"51",X"04",X"04",X"00",X"00",
		X"55",X"55",X"55",X"14",X"51",X"40",X"41",X"00",X"55",X"55",X"55",X"55",X"04",X"04",X"00",X"04",
		X"55",X"55",X"55",X"51",X"10",X"40",X"10",X"00",X"55",X"55",X"55",X"55",X"51",X"11",X"01",X"00",
		X"55",X"55",X"55",X"55",X"04",X"00",X"00",X"10",X"55",X"55",X"55",X"54",X"51",X"10",X"00",X"00",
		X"55",X"55",X"55",X"55",X"10",X"41",X"04",X"41",X"55",X"55",X"55",X"10",X"44",X"10",X"00",X"00",
		X"55",X"55",X"54",X"45",X"01",X"00",X"40",X"00",X"55",X"55",X"51",X"14",X"10",X"00",X"04",X"00",
		X"55",X"55",X"14",X"41",X"44",X"44",X"00",X"00",X"11",X"11",X"04",X"04",X"10",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"00",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"04",X"44",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"12",X"45",X"45",X"55",X"55",X"55",X"55",X"55",
		X"01",X"14",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"45",X"55",X"55",X"55",X"55",X"55",X"55",
		X"10",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"02",X"14",X"55",X"55",X"55",X"55",X"55",X"55",
		X"04",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"10",X"45",X"45",X"55",X"55",X"55",X"55",X"55",X"01",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"14",X"55",X"55",X"55",X"55",X"55",X"55",X"10",X"45",X"55",X"55",X"55",X"55",X"55",X"55",
		X"01",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"04",X"45",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"11",X"15",X"55",X"55",X"55",X"55",X"55",X"11",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"09",X"11",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"45",X"51",X"55",X"55",X"55",X"55",X"55",X"01",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"06",X"14",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"45",X"55",X"55",X"55",X"55",X"55",X"55",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"00",X"E2",X"55",X"55",X"55",X"55",X"57",X"95",
		X"00",X"E2",X"55",X"55",X"55",X"55",X"57",X"15",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"75",X"55",X"D5",X"5D",X"5D",X"55",X"55",X"5D",X"55",
		X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"5D",X"5D",X"75",X"75",X"55",X"57",X"55",X"5D",X"DD",X"55",X"55",X"55",X"D5",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"75",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"A9",X"55",X"45",X"55",X"55",X"55",X"55",X"56",X"A9",X"55",
		X"55",X"55",X"55",X"95",X"59",X"5A",X"99",X"55",X"55",X"55",X"55",X"65",X"5A",X"5A",X"A5",X"55",
		X"55",X"55",X"55",X"65",X"56",X"AA",X"A5",X"55",X"51",X"55",X"55",X"65",X"55",X"AA",X"99",X"55",
		X"55",X"55",X"55",X"95",X"15",X"9A",X"A6",X"55",X"51",X"55",X"56",X"55",X"55",X"96",X"A9",X"55",
		X"55",X"55",X"59",X"11",X"55",X"96",X"AA",X"55",X"45",X"55",X"65",X"55",X"55",X"9A",X"AA",X"95",
		X"55",X"55",X"95",X"41",X"55",X"5A",X"AA",X"65",X"51",X"15",X"A9",X"55",X"56",X"56",X"AA",X"95",
		X"55",X"55",X"99",X"54",X"65",X"55",X"AA",X"65",X"55",X"55",X"56",X"55",X"65",X"55",X"6A",X"95",
		X"55",X"11",X"56",X"55",X"55",X"55",X"6A",X"65",X"55",X"55",X"59",X"55",X"95",X"55",X"AA",X"95",
		X"55",X"44",X"59",X"55",X"55",X"55",X"AA",X"65",X"55",X"95",X"25",X"55",X"51",X"55",X"AA",X"95",
		X"55",X"56",X"65",X"55",X"55",X"55",X"AA",X"65",X"56",X"55",X"55",X"55",X"45",X"15",X"6A",X"95",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"A5",X"45",X"51",X"15",X"54",X"55",X"6A",X"95",
		X"65",X"55",X"55",X"55",X"61",X"55",X"AA",X"55",X"59",X"55",X"55",X"55",X"59",X"15",X"A5",X"55",
		X"59",X"14",X"55",X"55",X"56",X"56",X"99",X"55",X"59",X"55",X"55",X"55",X"56",X"5A",X"55",X"55",
		X"69",X"45",X"55",X"45",X"55",X"AA",X"66",X"55",X"65",X"11",X"54",X"55",X"55",X"6A",X"95",X"55",
		X"95",X"50",X"45",X"55",X"55",X"AA",X"99",X"55",X"55",X"45",X"55",X"51",X"56",X"5A",X"A5",X"55",
		X"55",X"54",X"45",X"55",X"55",X"56",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A5",X"55",
		X"10",X"55",X"55",X"55",X"45",X"6A",X"AF",X"FF",X"00",X"51",X"45",X"19",X"15",X"AA",X"AA",X"E5",
		X"11",X"40",X"66",X"69",X"C6",X"6A",X"AB",X"F9",X"54",X"15",X"66",X"29",X"55",X"AA",X"57",X"9D",
		X"45",X"53",X"25",X"59",X"59",X"A9",X"57",X"57",X"44",X"1A",X"51",X"69",X"66",X"AA",X"57",X"75",
		X"53",X"49",X"56",X"A9",X"5A",X"69",X"5D",X"55",X"54",X"64",X"45",X"A9",X"AA",X"A5",X"55",X"55",
		X"55",X"05",X"59",X"65",X"A9",X"95",X"55",X"95",X"56",X"05",X"1B",X"51",X"AA",X"95",X"55",X"55",
		X"55",X"41",X"65",X"55",X"AA",X"55",X"55",X"55",X"55",X"71",X"81",X"16",X"A9",X"65",X"75",X"55",
		X"54",X"55",X"81",X"55",X"6A",X"55",X"55",X"55",X"55",X"51",X"A9",X"A5",X"99",X"55",X"55",X"55",
		X"55",X"51",X"50",X"A5",X"A9",X"95",X"55",X"55",X"55",X"55",X"5A",X"92",X"A5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"51",X"55",X"55",X"55",X"54",X"00",X"00",X"00",
		X"5D",X"5D",X"55",X"55",X"51",X"01",X"04",X"00",X"54",X"55",X"5D",X"55",X"54",X"10",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"11",X"0C",X"00",
		X"55",X"55",X"55",X"55",X"55",X"44",X"10",X"40",X"55",X"55",X"55",X"5D",X"55",X"15",X"40",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"10",X"00",X"55",X"55",X"75",X"55",X"55",X"55",X"40",X"40",
		X"55",X"55",X"55",X"55",X"55",X"54",X"50",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"44",X"0C",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",
		X"55",X"55",X"55",X"D5",X"55",X"54",X"51",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"14",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"80",X"02",X"00",
		X"00",X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"08",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"08",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"04",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"02",X"00",X"80",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"E2",X"00",X"00",X"00",X"00",X"03",X"80",
		X"00",X"E2",X"00",X"00",X"00",X"00",X"03",X"00",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",
		X"3F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",X"3F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"14",X"26",X"55",X"55",
		X"55",X"55",X"54",X"56",X"50",X"55",X"95",X"55",X"55",X"55",X"19",X"15",X"61",X"55",X"A9",X"55",
		X"55",X"54",X"51",X"54",X"55",X"14",X"66",X"55",X"55",X"59",X"55",X"A1",X"14",X"55",X"69",X"95",
		X"54",X"45",X"04",X"25",X"59",X"41",X"9A",X"55",X"55",X"15",X"91",X"55",X"59",X"55",X"59",X"95",
		X"54",X"45",X"81",X"18",X"49",X"91",X"1A",X"A5",X"41",X"50",X"55",X"55",X"55",X"91",X"6B",X"55",
		X"00",X"05",X"61",X"45",X"01",X"55",X"AB",X"F5",X"51",X"55",X"59",X"59",X"5A",X"44",X"AB",X"F5",
		X"64",X"55",X"61",X"56",X"56",X"55",X"69",X"F5",X"69",X"05",X"A4",X"19",X"56",X"55",X"AA",X"A5",
		X"5A",X"51",X"65",X"49",X"5A",X"55",X"AA",X"A5",X"56",X"96",X"91",X"68",X"5A",X"75",X"AA",X"A5",
		X"56",X"92",X"54",X"A5",X"1A",X"56",X"AA",X"95",X"55",X"AA",X"56",X"A5",X"49",X"56",X"AA",X"55",
		X"55",X"6A",X"8A",X"A5",X"A9",X"5A",X"A5",X"95",X"55",X"56",X"A9",X"95",X"95",X"5A",X"9A",X"55",
		X"55",X"55",X"6A",X"45",X"A5",X"96",X"A9",X"55",X"55",X"55",X"56",X"AA",X"A2",X"9A",X"99",X"95",
		X"55",X"55",X"55",X"58",X"5B",X"AA",X"95",X"55",X"55",X"55",X"55",X"5A",X"AA",X"A9",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"56",X"18",X"46",X"55",X"55",X"55",X"55",X"94",X"44",X"46",X"48",X"95",
		X"55",X"55",X"65",X"60",X"90",X"11",X"99",X"A5",X"55",X"55",X"46",X"55",X"61",X"95",X"82",X"99",
		X"55",X"55",X"05",X"60",X"54",X"91",X"96",X"A5",X"55",X"54",X"15",X"25",X"26",X"65",X"44",X"A9",
		X"55",X"50",X"45",X"64",X"64",X"95",X"65",X"BF",X"55",X"45",X"55",X"65",X"65",X"94",X"A1",X"BF",
		X"55",X"55",X"15",X"65",X"65",X"A5",X"96",X"BF",X"55",X"55",X"54",X"A9",X"65",X"96",X"95",X"AA",
		X"55",X"55",X"95",X"95",X"65",X"95",X"99",X"AA",X"55",X"55",X"AA",X"95",X"96",X"9A",X"A4",X"AA",
		X"55",X"55",X"6A",X"6A",X"56",X"56",X"56",X"A9",X"55",X"64",X"56",X"69",X"9A",X"5A",X"9A",X"A5",
		X"55",X"12",X"45",X"5A",X"A5",X"6A",X"5A",X"A9",X"55",X"45",X"95",X"69",X"AA",X"AA",X"6A",X"A5",
		X"54",X"41",X"55",X"6A",X"4A",X"AA",X"A6",X"A5",X"60",X"55",X"A0",X"59",X"54",X"AA",X"6A",X"95",
		X"45",X"11",X"95",X"69",X"45",X"A6",X"2F",X"D5",X"64",X"45",X"85",X"25",X"55",X"91",X"6F",X"D5",
		X"59",X"16",X"A6",X"69",X"54",X"99",X"6F",X"D5",X"5A",X"16",X"65",X"6A",X"91",X"95",X"2A",X"95",
		X"56",X"62",X"94",X"69",X"55",X"A1",X"AA",X"95",X"55",X"6A",X"55",X"AA",X"16",X"96",X"AA",X"95",
		X"55",X"5A",X"55",X"A5",X"59",X"56",X"A9",X"55",X"55",X"56",X"99",X"95",X"56",X"66",X"A5",X"55",
		X"55",X"55",X"A6",X"A5",X"9A",X"4A",X"95",X"55",X"55",X"55",X"5A",X"A5",X"6A",X"6A",X"55",X"55",
		X"55",X"55",X"55",X"69",X"AA",X"6A",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"A5",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5A",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"45",X"55",X"55",X"55",X"55",X"51",X"00",X"00",X"15",X"55",X"5D",X"C5",X"51",X"54",X"10",
		X"01",X"05",X"55",X"55",X"55",X"15",X"51",X"00",X"00",X"11",X"55",X"55",X"D5",X"55",X"54",X"40",
		X"00",X"55",X"55",X"5D",X"75",X"55",X"51",X"00",X"00",X"11",X"55",X"55",X"55",X"51",X"54",X"10",
		X"00",X"05",X"55",X"55",X"D5",X"55",X"51",X"00",X"00",X"41",X"55",X"55",X"55",X"55",X"44",X"40",
		X"00",X"04",X"55",X"55",X"D5",X"55",X"51",X"00",X"00",X"01",X"15",X"5D",X"45",X"44",X"54",X"00",
		X"00",X"44",X"57",X"55",X"D5",X"55",X"55",X"00",X"00",X"01",X"55",X"75",X"55",X"15",X"55",X"40",
		X"00",X"05",X"57",X"57",X"75",X"55",X"55",X"00",X"00",X"11",X"55",X"55",X"55",X"55",X"44",X"00",
		X"00",X"01",X"55",X"55",X"D5",X"55",X"11",X"00",X"00",X"04",X"55",X"55",X"55",X"51",X"44",X"00",
		X"00",X"01",X"55",X"5D",X"45",X"15",X"50",X"40",X"00",X"04",X"55",X"55",X"55",X"55",X"54",X"00",
		X"00",X"01",X"15",X"55",X"55",X"51",X"51",X"00",X"00",X"00",X"45",X"57",X"55",X"55",X"54",X"00",
		X"00",X"01",X"15",X"55",X"55",X"55",X"50",X"10",X"00",X"00",X"41",X"55",X"55",X"55",X"44",X"00",
		X"00",X"00",X"15",X"55",X"55",X"51",X"10",X"00",X"00",X"01",X"05",X"55",X"D5",X"50",X"41",X"00",
		X"00",X"00",X"11",X"15",X"55",X"04",X"00",X"00",X"00",X"00",X"05",X"45",X"54",X"40",X"10",X"00",
		X"00",X"10",X"01",X"15",X"51",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"54",X"44",X"00",X"00",
		X"00",X"00",X"01",X"11",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"04",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"02",X"00",X"80",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"E2",X"00",X"00",X"00",X"00",X"03",X"80",
		X"00",X"E2",X"00",X"00",X"00",X"00",X"03",X"00",X"02",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"0F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"2F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",
		X"3F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",X"3F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"0B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"20",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"B8",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"00",X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"E8",X"84",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C2",X"20",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"A2",X"22",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"88",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"A2",X"20",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"E8",X"88",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"20",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"B8",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"E8",X"00",X"40",X"FB",X"FF",X"FF",X"FF",X"BF",X"F8",X"00",X"00",
		X"FB",X"FF",X"FF",X"FF",X"BF",X"B0",X"C0",X"00",X"FB",X"FF",X"FF",X"FF",X"BF",X"00",X"00",X"00",
		X"AB",X"AA",X"AA",X"AA",X"B8",X"00",X"00",X"00",X"0B",X"00",X"00",X"08",X"B0",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"08",X"B0",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"C0",X"40",X"0C",X"2A",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"30",X"0C",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"43",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"30",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"E8",X"20",X"00",
		X"00",X"00",X"00",X"03",X"03",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"C8",X"04",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"3E",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"A8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"E2",X"20",X"04",X"00",X"00",X"00",X"00",X"C3",X"E8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E2",X"00",X"C0",X"00",X"00",X"00",X"00",X"03",X"88",X"80",X"00",
		X"00",X"00",X"00",X"00",X"03",X"A2",X"08",X"00",X"00",X"00",X"00",X"00",X"33",X"E8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"03",X"FA",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"80",X"0C",
		X"00",X"00",X"00",X"00",X"03",X"E2",X"00",X"0C",X"00",X"00",X"00",X"0C",X"03",X"88",X"81",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"A2",X"20",X"00",X"00",X"00",X"00",X"00",X"0F",X"A8",X"82",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"E2",X"20",X"00",X"00",X"00",X"00",X"00",X"03",X"E8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"0C",X"00",
		X"00",X"00",X"00",X"03",X"FE",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"A2",X"08",X"10",X"00",X"00",X"00",X"30",X"0F",X"E8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"03",X"FA",X"20",X"00",X"00",X"00",X"00",X"00",X"0F",X"F8",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FA",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"80",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
