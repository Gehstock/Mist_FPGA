library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GALAXIAN_1H is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"00",X"30",X"34",X"6C",X"18",X"13",X"8F",X"8E",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"8C",X"1E",X"1F",X"63",X"70",X"1C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"03",X"00",X"60",X"E6",X"76",X"1C",X"18",X"8B",X"8F",
		X"03",X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"8E",X"88",X"18",X"1E",X"66",X"70",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"08",X"08",X"1B",X"37",X"1E",X"18",X"8B",X"8F",
		X"1F",X"1F",X"0F",X"00",X"00",X"00",X"01",X"01",X"88",X"88",X"1C",X"1C",X"67",X"63",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1C",X"1C",X"00",X"60",X"74",X"36",X"16",X"1E",X"08",X"0E",
		X"1C",X"1C",X"0F",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"18",X"1E",X"66",X"64",X"E4",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"00",X"00",X"80",X"C0",X"E0",X"58",X"38",X"20",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"3C",X"6C",X"70",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"80",X"E0",X"60",X"6C",X"3C",X"20",
		X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"68",X"C0",X"60",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"20",X"64",X"7C",X"78",X"30",X"28",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"60",X"60",X"60",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"80",X"C0",X"E8",X"78",X"30",X"2C",
		X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"30",X"60",X"30",X"70",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"30",X"60",X"60",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"50",X"60",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"50",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"40",X"60",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"40",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"D0",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"40",
		X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"60",X"C0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"00",X"08",X"1B",X"0F",X"0C",X"87",X"C7",X"C6",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"46",X"0B",X"0B",X"18",X"18",X"30",X"18",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"08",X"0C",X"1A",X"0F",X"CE",X"E6",X"E7",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"E6",X"E4",X"C6",X"0F",X"1F",X"19",X"38",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"0C",X"0C",X"18",X"0A",X"0E",X"26",X"24",
		X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"E7",X"E6",X"C4",X"0F",X"0F",X"19",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"08",X"1A",X"1E",X"0E",X"CD",X"07",X"06",
		X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"CF",X"0B",X"18",X"18",X"0C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"18",X"18",X"34",X"37",X"1F",X"18",
		X"1F",X"1F",X"10",X"10",X"00",X"00",X"00",X"00",X"8E",X"8F",X"8E",X"8F",X"13",X"1C",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"0F",X"00",X"00",X"10",X"38",X"F8",X"70",X"1E",X"1F",
		X"03",X"03",X"03",X"03",X"0F",X"00",X"00",X"00",X"89",X"8C",X"8F",X"8F",X"1E",X"1E",X"1B",X"38",
		X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"18",X"70",X"E0",X"72",X"1E",X"1C",
		X"10",X"10",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"8C",X"8E",X"8F",X"8D",X"18",X"1E",X"36",X"72",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"80",X"E0",X"3A",X"1F",X"1E",X"1E",
		X"1C",X"1C",X"1C",X"1C",X"0F",X"00",X"00",X"00",X"0D",X"0F",X"0F",X"0E",X"1E",X"16",X"3B",X"70",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"36",X"77",X"7C",X"18",X"0B",X"0E",X"8E",X"8F",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"98",X"18",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"04",X"2C",X"6F",X"3F",X"3C",X"18",X"C0",X"E0",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E8",X"CC",X"0E",X"1F",X"07",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"08",X"1C",X"3E",X"1C",X"00",X"00",X"20",
		X"04",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"20",X"E8",X"E8",X"CC",X"0E",X"1E",X"37",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1C",X"00",X"00",X"00",X"10",X"30",X"18",X"08",X"0C",
		X"1C",X"1C",X"1C",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0D",X"0E",X"0B",X"1D",X"3E",X"36",X"18",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"0C",X"18",X"18",X"1E",X"1C",X"0B",X"8F",X"8E",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"8C",X"0F",X"1B",X"38",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"03",X"00",X"00",X"1C",X"38",X"1E",X"0C",X"8D",X"8F",
		X"03",X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"8F",X"8E",X"0F",X"09",X"18",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"06",X"1E",X"1F",X"0E",X"8F",X"8F",
		X"1F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"8E",X"8E",X"0F",X"1C",X"1F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1C",X"1C",X"00",X"00",X"00",X"60",X"18",X"1F",X"0E",X"0C",
		X"1C",X"1C",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"0B",X"1C",X"1E",X"66",X"80",X"00",X"00",
		X"00",X"00",X"03",X"01",X"00",X"00",X"06",X"0F",X"00",X"00",X"D8",X"F4",X"6C",X"38",X"3C",X"38",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"00",X"00",X"06",X"03",X"00",X"00",X"D8",X"F4",X"7C",X"38",X"38",X"30",
		X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"30",X"E8",X"78",X"30",X"30",X"38",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"3C",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"06",X"0C",X"00",X"00",X"D0",X"B0",X"70",X"38",X"30",X"2C",
		X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"30",X"38",X"1C",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"00",X"00",X"00",X"18",X"78",X"70",X"3C",X"38",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"3C",X"6C",X"F8",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"00",X"F0",X"78",X"30",X"30",
		X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"70",X"F8",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"F8",X"70",X"2C",X"3C",
		X"0F",X"06",X"00",X"01",X"01",X"00",X"00",X"00",X"38",X"3C",X"74",X"F8",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"00",X"06",X"0C",X"00",X"00",X"00",X"80",X"D8",X"78",X"30",X"20",
		X"0C",X"06",X"00",X"00",X"03",X"03",X"00",X"00",X"38",X"38",X"6C",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"01",X"00",X"02",X"07",X"00",X"00",X"00",X"10",X"B0",X"E0",X"58",X"70",
		X"05",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"50",X"60",X"58",X"D0",X"80",X"00",X"00",X"00",
		X"00",X"03",X"07",X"00",X"00",X"00",X"06",X"0F",X"00",X"00",X"8C",X"D8",X"70",X"60",X"2E",X"3C",
		X"09",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"30",X"30",X"38",X"2E",X"EC",X"DC",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"6F",X"DF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"B0",
		X"3B",X"7F",X"7F",X"7F",X"3B",X"3F",X"7F",X"33",X"B0",X"30",X"60",X"60",X"C0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"33",X"7F",X"3F",X"3B",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",
		X"7F",X"7F",X"7F",X"3B",X"FF",X"DF",X"6F",X"03",X"60",X"60",X"30",X"B0",X"B0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"FF",X"F7",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",
		X"3F",X"7E",X"7E",X"37",X"FF",X"FF",X"0F",X"03",X"70",X"30",X"30",X"70",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"1C",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"37",X"7E",X"7F",X"3F",X"77",X"7F",X"3F",X"1C",X"F8",X"3C",X"1C",X"F8",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"83",X"CF",X"FF",X"7E",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",
		X"3B",X"7F",X"7F",X"3F",X"7A",X"FF",X"CF",X"83",X"70",X"30",X"30",X"70",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"33",X"7F",X"7F",X"FB",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",
		X"3F",X"7F",X"7F",X"3B",X"FF",X"7F",X"7F",X"33",X"70",X"30",X"30",X"70",X"60",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"83",X"CF",X"FF",X"77",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",
		X"3F",X"7E",X"7E",X"37",X"7F",X"FF",X"CF",X"83",X"70",X"30",X"30",X"70",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"33",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"A0",
		X"37",X"7E",X"7E",X"3F",X"F7",X"7F",X"7F",X"33",X"70",X"70",X"70",X"70",X"A0",X"C0",X"C0",X"80",
		X"00",X"03",X"07",X"07",X"03",X"01",X"42",X"A6",X"00",X"C0",X"00",X"80",X"C0",X"C0",X"60",X"50",
		X"AF",X"A6",X"42",X"01",X"03",X"07",X"07",X"03",X"D0",X"50",X"60",X"C0",X"C0",X"80",X"00",X"C0",
		X"00",X"0E",X"07",X"07",X"03",X"01",X"42",X"A6",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",X"50",
		X"AF",X"A6",X"42",X"01",X"03",X"07",X"07",X"0E",X"D0",X"50",X"60",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"7C",X"1F",X"0F",X"03",X"01",X"42",X"A6",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",X"50",
		X"AF",X"A6",X"42",X"01",X"03",X"0F",X"1F",X"7C",X"D0",X"50",X"60",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"0E",X"07",X"07",X"03",X"01",X"42",X"A6",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",X"50",
		X"AF",X"A6",X"42",X"01",X"03",X"07",X"07",X"0E",X"D0",X"50",X"60",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"0F",X"18",X"37",X"2C",X"2B",X"2A",X"00",X"00",X"F0",X"18",X"EC",X"36",X"DA",X"6A",
		X"2A",X"2B",X"2C",X"27",X"18",X"0F",X"00",X"00",X"AA",X"AA",X"6A",X"DA",X"36",X"EC",X"18",X"00",
		X"00",X"00",X"00",X"00",X"27",X"2C",X"2B",X"2A",X"00",X"00",X"00",X"00",X"E0",X"30",X"D8",X"68",
		X"2A",X"2B",X"2C",X"37",X"18",X"0F",X"00",X"00",X"A8",X"A8",X"68",X"D8",X"30",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0C",X"0B",X"0A",X"00",X"00",X"00",X"00",X"E0",X"30",X"D8",X"68",
		X"0A",X"0B",X"0C",X"07",X"00",X"00",X"00",X"00",X"A0",X"A0",X"60",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"60",X"40",X"00",X"00",X"00",X"00",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"00",X"07",X"37",X"33",X"03",X"0D",X"0C",X"00",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"0B",X"03",X"01",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"C0",X"C0",X"00",X"80",X"00",X"00",X"00",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"0E",X"0C",X"09",X"0F",X"FC",X"E4",X"CC",X"9C",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"18",X"18",X"24",X"DB",X"DB",X"24",X"18",X"18",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"60",X"03",X"03",X"1E",X"1E",X"C0",X"C0",X"60",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"28",X"10",X"28",X"64",X"64",X"74",X"38",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"05",X"00",X"00",X"00",X"02",X"A1",X"42",X"C0",X"A0",X"A0",X"90",X"90",X"A0",X"A0",X"C0",
		X"03",X"05",X"05",X"09",X"09",X"05",X"05",X"03",X"FF",X"81",X"66",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"66",X"81",X"FF",X"00",X"00",X"04",X"03",X"01",X"02",X"04",X"08",
		X"00",X"00",X"40",X"80",X"00",X"80",X"80",X"40",X"0C",X"0C",X"07",X"07",X"03",X"01",X"00",X"00",
		X"40",X"40",X"C0",X"80",X"80",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"C0",X"D8",X"10",X"02",X"1A",X"D0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"C0",X"80",X"10",X"30",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"18",X"3C",X"7E",X"E7",X"C3",X"81",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"C0",X"C0",X"FF",X"FF",X"C3",X"83",X"83",X"C3",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"FF",X"BF",X"87",X"87",X"87",X"DF",X"FF",X"C0",
		X"00",X"00",X"00",X"60",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"10",X"38",X"F8",
		X"FC",X"FC",X"F8",X"7C",X"FC",X"F8",X"40",X"00",X"00",X"00",X"00",X"24",X"3C",X"FC",X"F8",X"FE",
		X"FC",X"38",X"1C",X"0C",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"70",X"20",X"00",X"00",
		X"00",X"00",X"06",X"C7",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"06",X"00",X"00",X"00",X"18",X"3F",
		X"7F",X"FF",X"7F",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7F",X"FF",X"7F",
		X"3F",X"18",X"00",X"00",X"00",X"06",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"C7",X"02",X"00",X"00",
		X"00",X"0C",X"1F",X"3F",X"3F",X"1F",X"0C",X"00",X"80",X"00",X"00",X"00",X"21",X"00",X"00",X"00",
		X"00",X"08",X"00",X"C0",X"C0",X"60",X"60",X"60",X"60",X"60",X"C0",X"C0",X"00",X"00",X"08",X"00",
		X"00",X"0C",X"1F",X"3F",X"3F",X"1F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"42",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"01",X"00",X"40",X"20",X"00",
		X"20",X"40",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FC",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"18",X"38",X"F0",X"FC",
		X"FC",X"F8",X"F0",X"7C",X"FC",X"E4",X"40",X"00",X"00",X"00",X"00",X"08",X"18",X"F8",X"FE",X"FC",
		X"F8",X"7E",X"EC",X"60",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"20",X"00",X"00",
		X"00",X"38",X"1D",X"DF",X"FF",X"FF",X"FF",X"3F",X"1E",X"0C",X"00",X"00",X"00",X"00",X"18",X"3F",
		X"3F",X"18",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"DF",X"0F",X"06",X"00",
		X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"78",X"00",X"00",
		X"FF",X"39",X"63",X"07",X"01",X"00",X"00",X"01",X"01",X"03",X"06",X"00",X"00",X"80",X"80",X"C0",
		X"C0",X"C0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"0F",X"07",X"01",X"00",X"00",
		X"00",X"00",X"1C",X"FF",X"73",X"20",X"00",X"00",X"00",X"00",X"00",X"70",X"FD",X"DF",X"8F",X"01",
		X"1F",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C1",X"C3",X"C7",
		X"C7",X"B7",X"33",X"03",X"0D",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",
		X"01",X"00",X"10",X"40",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"36",X"64",X"6C",X"30",X"30",X"18",X"1C",X"1C",X"3C",X"3C",X"1C",
		X"00",X"00",X"00",X"00",X"14",X"2A",X"54",X"0F",X"7F",X"7F",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"01",X"00",X"00",X"00",X"02",X"06",X"CC",X"80",X"80",
		X"00",X"12",X"40",X"08",X"20",X"00",X"00",X"00",X"09",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"01",X"C3",
		X"C7",X"07",X"0F",X"0F",X"DE",X"DE",X"0E",X"06",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"00",X"00",
		X"00",X"60",X"60",X"00",X"00",X"30",X"30",X"00",X"00",X"0C",X"0C",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E1",X"E3",X"C1",X"81",X"00",X"0C",X"0C",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",
		X"00",X"00",X"00",X"00",X"12",X"36",X"64",X"6C",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",
		X"00",X"08",X"21",X"04",X"10",X"00",X"00",X"06",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"61",X"63",
		X"07",X"07",X"CF",X"CF",X"1E",X"1E",X"0E",X"C6",X"C0",X"00",X"00",X"00",X"60",X"60",X"00",X"00",
		X"00",X"00",X"60",X"60",X"00",X"00",X"30",X"30",X"00",X"18",X"18",X"00",X"03",X"03",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"07",X"07",X"07",X"07",X"07",X"87",X"87",X"07",X"87",X"87",X"07",X"07",X"07",X"07",X"07",X"03",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"01",X"01",X"00",
		X"01",X"01",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",X"FE",X"FF",X"FF",
		X"FF",X"FE",X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"67",X"67",X"07",
		X"67",X"67",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"80",X"80",X"80",X"02",X"04",X"08",X"08",X"08",
		X"08",X"10",X"10",X"10",X"20",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"3F",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"00",X"00",X"10",X"20",X"A0",X"44",X"44",X"06",
		X"40",X"A0",X"04",X"08",X"10",X"20",X"00",X"00",X"46",X"46",X"40",X"40",X"98",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"01",X"01",X"01",X"21",X"01",X"80",X"96",X"88",X"90",X"02",X"02",X"03",X"00",
		X"00",X"00",X"C0",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"88",X"00",X"22",X"00",X"00",X"00",X"10",X"00",X"04",X"00",X"00",X"00",X"30",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"00",X"00",X"00",X"01",X"06",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"86",X"64",X"B4",X"DB",X"0F",X"03",X"01",X"08",X"04",X"06",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"03",X"03",X"07",X"07",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"01",X"00",X"00",X"0C",X"0C",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",
		X"08",X"08",X"04",X"02",X"02",X"32",X"CC",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"40",X"E0",X"F0",X"F8",X"F8",X"FC",X"F8",X"00",X"00",X"10",X"20",X"A0",X"46",X"42",X"02",
		X"40",X"A0",X"0C",X"10",X"20",X"20",X"00",X"00",X"40",X"40",X"80",X"00",X"0C",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"96",X"88",X"90",X"03",X"01",X"01",X"00",
		X"00",X"03",X"04",X"C8",X"30",X"03",X"03",X"00",X"00",X"00",X"00",X"40",X"C8",X"90",X"A0",X"A0",
		X"E0",X"E0",X"C0",X"88",X"00",X"22",X"00",X"00",X"3F",X"3F",X"1F",X"0F",X"02",X"00",X"00",X"00",
		X"10",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"11",X"0B");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
