library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity LLANDER_VEC_ROM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of LLANDER_VEC_ROM_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"27",X"00",X"05",X"80",X"22",X"80",X"C6",X"80",X"22",X"00",X"C0",X"80",X"22",X"80",X"C2",
		X"00",X"20",X"80",X"C2",X"80",X"26",X"80",X"C2",X"80",X"26",X"00",X"C0",X"80",X"26",X"80",X"C6",
		X"00",X"20",X"80",X"C6",X"00",X"D0",X"00",X"36",X"40",X"04",X"C7",X"F2",X"80",X"22",X"80",X"C4",
		X"C2",X"F3",X"80",X"20",X"80",X"C2",X"C3",X"F6",X"80",X"26",X"80",X"C0",X"C6",X"F7",X"80",X"24",
		X"80",X"C6",X"00",X"D0",X"40",X"36",X"00",X"00",X"80",X"21",X"80",X"C7",X"80",X"22",X"00",X"C5",
		X"80",X"23",X"80",X"C1",X"00",X"21",X"80",X"C2",X"80",X"25",X"80",X"C3",X"80",X"26",X"00",X"C1",
		X"80",X"27",X"80",X"C5",X"00",X"25",X"80",X"C6",X"00",X"D0",X"00",X"36",X"80",X"00",X"80",X"20",
		X"80",X"C7",X"00",X"22",X"80",X"C5",X"80",X"23",X"80",X"C0",X"80",X"21",X"00",X"C2",X"80",X"24",
		X"80",X"C3",X"00",X"26",X"80",X"C1",X"80",X"27",X"80",X"C4",X"80",X"25",X"00",X"C6",X"00",X"D0",
		X"05",X"FE",X"C5",X"F9",X"80",X"23",X"00",X"C0",X"C1",X"F9",X"00",X"20",X"80",X"C3",X"C1",X"FD",
		X"80",X"27",X"00",X"C0",X"C5",X"FD",X"00",X"20",X"80",X"C7",X"00",X"D0",X"00",X"36",X"C0",X"04",
		X"80",X"21",X"00",X"C6",X"80",X"23",X"80",X"C4",X"00",X"22",X"80",X"C1",X"80",X"20",X"80",X"C3",
		X"80",X"25",X"00",X"C2",X"80",X"27",X"80",X"C0",X"00",X"26",X"80",X"C5",X"80",X"24",X"80",X"C7",
		X"00",X"D0",X"00",X"36",X"40",X"04",X"00",X"21",X"80",X"C6",X"80",X"23",X"80",X"C5",X"80",X"22",
		X"00",X"C1",X"80",X"21",X"80",X"C3",X"00",X"25",X"80",X"C2",X"80",X"27",X"80",X"C1",X"80",X"26",
		X"00",X"C5",X"80",X"25",X"80",X"C7",X"00",X"D0",X"00",X"36",X"40",X"00",X"80",X"20",X"80",X"C6",
		X"C6",X"F3",X"80",X"22",X"80",X"C0",X"C3",X"F2",X"80",X"24",X"80",X"C2",X"C2",X"F7",X"80",X"26",
		X"80",X"C4",X"C7",X"F6",X"00",X"D0",X"00",X"C4",X"C0",X"33",X"40",X"05",X"80",X"26",X"00",X"C0",
		X"80",X"26",X"00",X"00",X"80",X"26",X"00",X"C0",X"00",X"10",X"00",X"C7",X"C0",X"33",X"00",X"C0",
		X"00",X"10",X"00",X"C3",X"00",X"10",X"00",X"07",X"C6",X"F9",X"00",X"F1",X"C0",X"FD",X"60",X"46",
		X"00",X"00",X"C0",X"FD",X"00",X"F1",X"C2",X"F9",X"00",X"F9",X"80",X"25",X"00",X"C7",X"40",X"33",
		X"00",X"C0",X"80",X"25",X"00",X"C3",X"80",X"21",X"00",X"07",X"00",X"D0",X"13",X"C4",X"80",X"24",
		X"80",X"06",X"80",X"22",X"80",X"C4",X"80",X"22",X"80",X"04",X"80",X"22",X"80",X"C4",X"00",X"15",
		X"00",X"C7",X"C0",X"37",X"C0",X"C0",X"00",X"11",X"00",X"C3",X"00",X"15",X"00",X"07",X"80",X"26",
		X"80",X"C7",X"00",X"16",X"00",X"01",X"C5",X"F2",X"60",X"42",X"80",X"04",X"C0",X"F9",X"00",X"F5",
		X"C0",X"34",X"40",X"C2",X"C0",X"36",X"80",X"00",X"00",X"26",X"80",X"C6",X"40",X"33",X"C0",X"C4",
		X"00",X"25",X"80",X"C3",X"00",X"21",X"80",X"07",X"00",X"D0",X"22",X"C4",X"40",X"33",X"C0",X"06",
		X"80",X"26",X"00",X"C1",X"80",X"26",X"00",X"01",X"80",X"26",X"00",X"C1",X"00",X"15",X"00",X"C7",
		X"C0",X"33",X"80",X"C5",X"00",X"11",X"00",X"C3",X"00",X"15",X"00",X"07",X"40",X"30",X"00",X"C6",
		X"00",X"12",X"00",X"05",X"C1",X"F6",X"40",X"46",X"C0",X"00",X"C1",X"F6",X"00",X"12",X"00",X"05",
		X"C3",X"F3",X"05",X"F2",X"80",X"26",X"00",X"C6",X"40",X"33",X"40",X"C5",X"80",X"24",X"80",X"C3",
		X"80",X"20",X"80",X"07",X"00",X"D0",X"35",X"C4",X"80",X"25",X"00",X"06",X"00",X"22",X"80",X"C5",
		X"00",X"22",X"80",X"05",X"00",X"22",X"80",X"C5",X"00",X"15",X"00",X"C7",X"40",X"37",X"80",X"C2",
		X"C1",X"F1",X"05",X"F5",X"40",X"36",X"00",X"C5",X"00",X"06",X"00",X"02",X"C5",X"F1",X"40",X"42",
		X"A0",X"05",X"C5",X"F2",X"00",X"16",X"00",X"01",X"40",X"30",X"40",X"C2",X"40",X"36",X"C0",X"01",
		X"00",X"27",X"80",X"C5",X"80",X"32",X"00",X"C6",X"80",X"20",X"80",X"C3",X"80",X"24",X"80",X"07",
		X"00",X"D0",X"48",X"C4",X"01",X"FD",X"C5",X"F9",X"05",X"F9",X"C5",X"F9",X"C5",X"F5",X"C3",X"FF",
		X"C1",X"F1",X"05",X"F5",X"00",X"36",X"C0",X"C4",X"00",X"06",X"00",X"02",X"C5",X"F1",X"C0",X"33",
		X"C0",X"07",X"C5",X"F1",X"00",X"06",X"00",X"02",X"C0",X"30",X"00",X"C2",X"40",X"36",X"40",X"02",
		X"C5",X"F7",X"80",X"32",X"C0",X"C6",X"00",X"21",X"80",X"C3",X"00",X"25",X"80",X"07",X"00",X"D0",
		X"56",X"C4",X"80",X"31",X"00",X"06",X"80",X"25",X"00",X"C2",X"80",X"25",X"00",X"02",X"80",X"25",
		X"00",X"C2",X"C5",X"F5",X"40",X"32",X"00",X"C7",X"C1",X"F1",X"05",X"F5",X"C6",X"FD",X"00",X"02",
		X"00",X"06",X"C1",X"F5",X"00",X"37",X"C0",X"03",X"C2",X"F5",X"00",X"11",X"00",X"06",X"40",X"32",
		X"80",X"C0",X"00",X"12",X"00",X"07",X"80",X"27",X"80",X"C4",X"00",X"32",X"C0",X"C6",X"80",X"21",
		X"80",X"C3",X"80",X"25",X"80",X"07",X"00",X"D0",X"69",X"C4",X"00",X"25",X"80",X"02",X"00",X"21",
		X"80",X"C6",X"00",X"21",X"80",X"06",X"00",X"21",X"80",X"C6",X"00",X"17",X"00",X"C5",X"80",X"35",
		X"C0",X"C3",X"00",X"13",X"00",X"C1",X"00",X"17",X"00",X"05",X"40",X"36",X"00",X"C0",X"01",X"F0",
		X"C5",X"F8",X"00",X"41",X"60",X"06",X"C5",X"F1",X"00",X"06",X"00",X"02",X"00",X"23",X"80",X"C3",
		X"00",X"35",X"C0",X"02",X"80",X"27",X"00",X"C0",X"40",X"31",X"00",X"C7",X"00",X"22",X"80",X"C2",
		X"00",X"26",X"80",X"06",X"00",X"D0",X"7C",X"C4",X"80",X"24",X"80",X"02",X"80",X"20",X"80",X"C6",
		X"80",X"20",X"80",X"06",X"80",X"20",X"80",X"C6",X"00",X"17",X"00",X"C5",X"60",X"44",X"00",X"C2",
		X"00",X"13",X"00",X"C0",X"00",X"17",X"00",X"00",X"40",X"36",X"80",X"C0",X"01",X"F0",X"C5",X"F8",
		X"80",X"40",X"60",X"06",X"C6",X"F1",X"00",X"15",X"00",X"02",X"80",X"23",X"80",X"C2",X"80",X"34",
		X"00",X"03",X"80",X"27",X"00",X"C1",X"C0",X"30",X"80",X"C7",X"80",X"22",X"00",X"C2",X"80",X"26",
		X"00",X"C6",X"00",X"D0",X"00",X"C4",X"00",X"20",X"80",X"C6",X"00",X"17",X"00",X"C0",X"00",X"30",
		X"C0",X"C3",X"00",X"13",X"00",X"C0",X"00",X"20",X"80",X"C6",X"C0",X"34",X"80",X"06",X"C5",X"FE",
		X"05",X"F0",X"C1",X"F8",X"00",X"40",X"60",X"02",X"C1",X"F8",X"05",X"F0",X"C5",X"FA",X"05",X"F8",
		X"00",X"27",X"80",X"C1",X"00",X"30",X"40",X"C7",X"00",X"23",X"80",X"C1",X"00",X"27",X"80",X"05",
		X"00",X"D0",X"8B",X"C4",X"AE",X"C4",X"D5",X"C4",X"FB",X"C4",X"21",X"C5",X"40",X"C5",X"64",X"C5",
		X"8B",X"C5",X"B2",X"C5",X"AA",X"A2",X"40",X"00",X"00",X"70",X"00",X"00",X"E8",X"A0",X"00",X"00",
		X"40",X"A0",X"00",X"00",X"18",X"A1",X"00",X"00",X"78",X"A0",X"00",X"00",X"EA",X"00",X"AC",X"A0",
		X"80",X"00",X"E0",X"A0",X"80",X"00",X"18",X"A0",X"80",X"00",X"18",X"A0",X"80",X"00",X"80",X"A1",
		X"00",X"02",X"00",X"B0",X"80",X"20",X"80",X"06",X"00",X"13",X"00",X"C3",X"00",X"10",X"00",X"C3",
		X"00",X"17",X"00",X"C3",X"00",X"17",X"00",X"C0",X"00",X"17",X"00",X"C7",X"00",X"10",X"00",X"C7",
		X"00",X"13",X"00",X"C7",X"06",X"F7",X"C2",X"F1",X"C0",X"32",X"00",X"C0",X"C6",X"F1",X"02",X"F7",
		X"00",X"12",X"00",X"C7",X"80",X"27",X"00",X"C0",X"00",X"12",X"00",X"C3",X"80",X"22",X"80",X"05",
		X"00",X"D0",X"00",X"20",X"80",X"06",X"C1",X"F2",X"00",X"11",X"00",X"C3",X"C2",X"F5",X"00",X"17",
		X"00",X"C1",X"C5",X"F6",X"00",X"15",X"00",X"C7",X"C6",X"F1",X"C5",X"F5",X"00",X"23",X"80",X"C4",
		X"00",X"15",X"00",X"C3",X"00",X"22",X"80",X"06",X"80",X"24",X"00",X"C2",X"40",X"36",X"80",X"C0",
		X"00",X"16",X"00",X"C7",X"40",X"32",X"40",X"04",X"00",X"D0",X"00",X"20",X"80",X"06",X"C1",X"F2",
		X"00",X"11",X"00",X"C3",X"C2",X"F5",X"00",X"17",X"00",X"C1",X"C5",X"F6",X"00",X"15",X"00",X"C7",
		X"C6",X"F1",X"05",X"F7",X"00",X"13",X"00",X"C3",X"40",X"32",X"C0",X"C4",X"80",X"20",X"00",X"C6",
		X"00",X"26",X"80",X"02",X"00",X"11",X"00",X"C7",X"80",X"27",X"00",X"C1",X"00",X"13",X"00",X"C2",
		X"05",X"F9",X"00",X"D0",X"00",X"26",X"80",X"05",X"80",X"24",X"00",X"C2",X"00",X"12",X"00",X"C3",
		X"00",X"22",X"80",X"C0",X"00",X"13",X"00",X"C6",X"80",X"20",X"00",X"C6",X"00",X"16",X"00",X"C7",
		X"00",X"26",X"80",X"C4",X"80",X"21",X"80",X"C7",X"00",X"20",X"80",X"C2",X"40",X"36",X"80",X"C1",
		X"C5",X"F6",X"80",X"23",X"00",X"00",X"00",X"17",X"00",X"C5",X"C6",X"F3",X"00",X"10",X"00",X"C3",
		X"00",X"10",X"00",X"07",X"00",X"D0",X"06",X"F5",X"B0",X"F9",X"B1",X"F1",X"B1",X"F8",X"B1",X"F5",
		X"B0",X"FD",X"B5",X"F5",X"B5",X"F8",X"80",X"27",X"00",X"01",X"00",X"22",X"80",X"C0",X"CD",X"F1",
		X"80",X"24",X"00",X"C6",X"00",X"25",X"80",X"03",X"C5",X"F8",X"C3",X"F7",X"C0",X"F9",X"07",X"F1",
		X"00",X"D0",X"80",X"26",X"80",X"04",X"80",X"20",X"00",X"C2",X"00",X"13",X"00",X"C2",X"00",X"22",
		X"80",X"C4",X"00",X"12",X"00",X"C7",X"80",X"24",X"00",X"C6",X"00",X"17",X"00",X"C6",X"00",X"26",
		X"80",X"C0",X"00",X"36",X"80",X"01",X"C0",X"F9",X"80",X"31",X"40",X"C6",X"C6",X"F5",X"00",X"20",
		X"80",X"03",X"00",X"15",X"00",X"C7",X"C3",X"F6",X"00",X"13",X"00",X"C0",X"80",X"20",X"00",X"07",
		X"00",X"D0",X"00",X"26",X"80",X"05",X"C5",X"F2",X"00",X"13",X"00",X"C1",X"C2",X"F1",X"00",X"15",
		X"00",X"C3",X"C1",X"F6",X"00",X"17",X"00",X"C5",X"C6",X"F5",X"80",X"26",X"00",X"02",X"00",X"22",
		X"80",X"C4",X"C0",X"30",X"40",X"C6",X"00",X"17",X"00",X"C7",X"03",X"F1",X"00",X"16",X"00",X"C7",
		X"00",X"25",X"80",X"C3",X"00",X"13",X"00",X"C5",X"80",X"24",X"00",X"07",X"00",X"D0",X"80",X"26",
		X"00",X"00",X"C2",X"F1",X"00",X"13",X"00",X"C1",X"C5",X"F2",X"00",X"11",X"00",X"C7",X"C6",X"F5",
		X"00",X"17",X"00",X"C5",X"C1",X"F6",X"C5",X"F5",X"80",X"24",X"00",X"C3",X"00",X"13",X"00",X"C5",
		X"80",X"26",X"00",X"02",X"00",X"22",X"80",X"C4",X"80",X"30",X"40",X"C6",X"00",X"17",X"00",X"C6",
		X"00",X"10",X"00",X"03",X"00",X"D0",X"80",X"26",X"80",X"04",X"00",X"13",X"00",X"C7",X"00",X"13",
		X"00",X"C0",X"00",X"13",X"00",X"C3",X"00",X"10",X"00",X"C3",X"00",X"17",X"00",X"C3",X"00",X"17",
		X"00",X"C0",X"00",X"17",X"00",X"C7",X"03",X"F6",X"C5",X"F2",X"00",X"30",X"C0",X"C6",X"C5",X"F6",
		X"03",X"F2",X"00",X"17",X"00",X"C6",X"00",X"20",X"80",X"C3",X"00",X"13",X"00",X"C6",X"80",X"25",
		X"80",X"06",X"00",X"D0",X"F2",X"C5",X"11",X"C6",X"2D",X"C6",X"4A",X"C6",X"6B",X"C6",X"81",X"C6",
		X"A1",X"C6",X"BF",X"C6",X"DB",X"C6",X"18",X"A0",X"80",X"02",X"18",X"A0",X"60",X"03",X"38",X"A0",
		X"08",X"01",X"20",X"A0",X"30",X"03",X"68",X"A0",X"40",X"00",X"A0",X"A0",X"C8",X"03",X"E8",X"A0",
		X"00",X"00",X"C0",X"A0",X"98",X"00",X"88",X"A0",X"C8",X"00",X"70",X"A1",X"C0",X"01",X"78",X"A0",
		X"F8",X"02",X"E0",X"A0",X"80",X"01",X"F0",X"A0",X"20",X"02",X"B8",X"A0",X"30",X"02",X"40",X"A0",
		X"60",X"02",X"40",X"00",X"00",X"0A",X"40",X"00",X"80",X"0D",X"C0",X"00",X"20",X"04",X"60",X"00",
		X"C0",X"0C",X"80",X"01",X"00",X"01",X"60",X"02",X"20",X"0F",X"80",X"03",X"00",X"00",X"E0",X"02",
		X"60",X"02",X"00",X"02",X"20",X"03",X"A0",X"05",X"00",X"07",X"C0",X"01",X"E0",X"0B",X"60",X"03",
		X"00",X"06",X"A0",X"03",X"80",X"08",X"C0",X"02",X"C0",X"08",X"E0",X"00",X"80",X"09",X"00",X"80",
		X"00",X"D2",X"50",X"74",X"18",X"06",X"00",X"70",X"00",X"D2",X"A0",X"64",X"30",X"06",X"00",X"60",
		X"00",X"D2",X"40",X"55",X"60",X"06",X"00",X"40",X"E0",X"D3",X"80",X"46",X"00",X"07",X"57",X"C7",
		X"5B",X"C7",X"5F",X"C7",X"63",X"C7",X"67",X"C7",X"6A",X"C7",X"6E",X"C7",X"72",X"C7",X"00",X"C4",
		X"80",X"23",X"00",X"01",X"00",X"D0",X"13",X"C4",X"00",X"32",X"40",X"00",X"00",X"D0",X"22",X"C4",
		X"40",X"32",X"00",X"00",X"00",X"D0",X"35",X"C4",X"00",X"32",X"80",X"04",X"00",X"D0",X"48",X"C4",
		X"01",X"FA",X"00",X"D0",X"56",X"C4",X"00",X"32",X"C0",X"00",X"00",X"D0",X"69",X"C4",X"00",X"32",
		X"40",X"00",X"00",X"D0",X"7C",X"C4",X"00",X"32",X"40",X"04",X"00",X"D0",X"8E",X"C7",X"94",X"C7",
		X"9D",X"C7",X"A3",X"C7",X"A9",X"C7",X"B1",X"C7",X"B7",X"C7",X"BC",X"C7",X"C7",X"C7",X"D0",X"C7",
		X"D7",X"C7",X"DF",X"C7",X"9D",X"C7",X"DF",X"C7",X"C7",X"C7",X"B1",X"C7",X"A3",X"C7",X"DF",X"C7",
		X"BC",X"C7",X"94",X"C7",X"9D",X"C7",X"D0",X"C7",X"B1",X"C7",X"B7",X"C7",X"A5",X"F8",X"01",X"F0",
		X"A1",X"FA",X"00",X"36",X"80",X"04",X"00",X"D0",X"00",X"20",X"80",X"A6",X"00",X"17",X"00",X"A0",
		X"00",X"30",X"C0",X"A2",X"80",X"21",X"00",X"07",X"00",X"D0",X"A7",X"F0",X"00",X"23",X"80",X"A1",
		X"00",X"27",X"80",X"01",X"00",X"D0",X"00",X"20",X"80",X"A3",X"00",X"23",X"80",X"A5",X"06",X"F7",
		X"00",X"D0",X"A1",X"F8",X"00",X"13",X"00",X"A0",X"00",X"30",X"80",X"A6",X"80",X"25",X"00",X"03",
		X"00",X"D0",X"A1",X"F8",X"05",X"F0",X"A5",X"FA",X"00",X"36",X"80",X"00",X"00",X"D0",X"A0",X"F1",
		X"A1",X"F0",X"A0",X"F5",X"A5",X"F0",X"00",X"D0",X"00",X"27",X"80",X"A5",X"00",X"30",X"40",X"A3",
		X"00",X"23",X"80",X"A5",X"00",X"25",X"80",X"A6",X"00",X"11",X"00",X"A6",X"00",X"D0",X"00",X"13",
		X"00",X"A0",X"00",X"30",X"80",X"A3",X"00",X"17",X"00",X"A0",X"00",X"30",X"80",X"A7",X"00",X"D0",
		X"A5",X"F1",X"00",X"06",X"00",X"02",X"A2",X"F9",X"80",X"26",X"80",X"07",X"00",X"D0",X"A1",X"F1",
		X"00",X"06",X"00",X"06",X"C0",X"30",X"00",X"A6",X"00",X"26",X"80",X"07",X"00",X"D0",X"00",X"13",
		X"00",X"A3",X"00",X"17",X"00",X"A3",X"00",X"17",X"00",X"A7",X"00",X"13",X"00",X"A7",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"53");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
