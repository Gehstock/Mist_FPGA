library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_sprite_u is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_sprite_u is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AA",X"AA",X"AA",X"AF",X"2A",X"FF",X"06",X"F5",X"06",X"F1",X"01",X"F5",X"00",X"7C",X"00",X"7F",
		X"FF",X"FD",X"FF",X"FD",X"3F",X"FD",X"4F",X"FD",X"43",X"FD",X"03",X"FD",X"0F",X"F7",X"3F",X"F7",
		X"00",X"1F",X"00",X"07",X"00",X"07",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F7",X"FF",X"DF",X"FF",X"5F",X"7D",X"FF",X"17",X"FF",X"01",X"55",X"00",X"15",X"00",X"00",
		X"FF",X"7F",X"FF",X"5F",X"FD",X"F7",X"F7",X"F5",X"5F",X"FD",X"DF",X"F5",X"F7",X"F5",X"FD",X"D5",
		X"FF",X"C0",X"D5",X"40",X"DA",X"80",X"42",X"A0",X"02",X"A0",X"00",X"A0",X"80",X"A8",X"80",X"28",
		X"FD",X"56",X"FD",X"5A",X"F5",X"5A",X"D5",X"A5",X"56",X"6A",X"5A",X"9A",X"0A",X"A5",X"00",X"2A",
		X"80",X"0A",X"80",X"02",X"A0",X"00",X"50",X"00",X"A0",X"00",X"A0",X"00",X"54",X"00",X"AA",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"1F",X"00",X"7F",X"01",X"FF",
		X"00",X"00",X"00",X"00",X"05",X"54",X"5F",X"5D",X"FF",X"DF",X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",
		X"0A",X"AA",X"0A",X"AA",X"05",X"41",X"01",X"00",X"00",X"01",X"04",X"05",X"05",X"15",X"15",X"2A",
		X"AB",X"FD",X"AA",X"A6",X"40",X"01",X"04",X"09",X"05",X"AD",X"4A",X"BD",X"AB",X"FD",X"AF",X"FD",
		X"00",X"24",X"00",X"2A",X"00",X"AA",X"40",X"A9",X"D6",X"A6",X"F5",X"6A",X"FD",X"6A",X"FD",X"D9",
		X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"00",X"A0",X"00",X"A4",X"00",X"58",X"00",X"AA",X"02",
		X"FD",X"F6",X"FD",X"FD",X"F5",X"FD",X"5F",X"FD",X"F5",X"FD",X"FD",X"F5",X"FF",X"77",X"FF",X"5F",
		X"AA",X"0A",X"00",X"28",X"00",X"A8",X"40",X"A0",X"42",X"A0",X"52",X"A0",X"DA",X"80",X"D5",X"40",
		X"00",X"00",X"00",X"04",X"00",X"05",X"10",X"05",X"14",X"06",X"15",X"0A",X"15",X"6A",X"05",X"AA",
		X"16",X"BF",X"1A",X"BF",X"2A",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"CF",X"AF",X"43",X"BC",X"50",
		X"0A",X"AA",X"2A",X"AA",X"2A",X"AB",X"02",X"97",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"50",X"FD",X"40",X"FF",X"03",X"FF",X"FF",X"5F",X"FF",X"15",X"7D",X"00",X"55",X"00",X"00",
		X"DF",X"7F",X"DF",X"5F",X"DF",X"77",X"D5",X"F5",X"DF",X"FD",X"D7",X"FD",X"DD",X"F5",X"DF",X"75",
		X"FF",X"C0",X"D5",X"40",X"DA",X"80",X"42",X"A0",X"40",X"A8",X"40",X"2A",X"00",X"02",X"00",X"00",
		X"DF",X"56",X"DF",X"5A",X"DF",X"55",X"55",X"6A",X"55",X"55",X"56",X"AA",X"5A",X"A8",X"00",X"00",
		X"A0",X"00",X"55",X"00",X"AA",X"A0",X"AA",X"A8",X"55",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"00",X"AA",X"02",X"AA",X"01",X"5A",X"01",X"51",
		X"00",X"00",X"00",X"54",X"55",X"55",X"5F",X"5F",X"BF",X"DF",X"5F",X"DF",X"AB",X"D7",X"6A",X"F7",
		X"01",X"41",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"52",X"A9",X"41",X"5A",X"01",X"06",X"00",X"02",X"00",X"02",X"00",X"1A",X"10",X"6B",X"14",X"AF",
		X"00",X"00",X"00",X"00",X"40",X"0A",X"54",X"2A",X"F6",X"A5",X"F5",X"5A",X"FD",X"DA",X"FD",X"F5",
		X"00",X"00",X"A0",X"00",X"A8",X"00",X"A4",X"00",X"58",X"00",X"AA",X"00",X"95",X"00",X"6A",X"00",
		X"FD",X"FD",X"7D",X"FD",X"75",X"FD",X"5F",X"FD",X"55",X"FD",X"5D",X"F5",X"5F",X"77",X"DF",X"5F",
		X"AA",X"00",X"0A",X"00",X"40",X"02",X"40",X"2A",X"40",X"A8",X"42",X"A0",X"DA",X"80",X"D5",X"40",
		X"AB",X"57",X"2B",X"55",X"0B",X"55",X"03",X"5F",X"03",X"55",X"03",X"55",X"0B",X"57",X"2B",X"55",
		X"55",X"55",X"D5",X"55",X"75",X"57",X"D7",X"5D",X"75",X"F5",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"0A",X"D5",X"00",X"D5",X"00",X"35",X"00",X"B5",X"02",X"AD",X"00",X"AB",X"00",X"00",X"00",X"00",
		X"56",X"A0",X"56",X"A0",X"55",X"A8",X"55",X"6A",X"55",X"56",X"D5",X"55",X"3D",X"55",X"0F",X"FF",
		X"55",X"55",X"55",X"55",X"D5",X"7D",X"75",X"DF",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"00",X"57",X"00",X"5F",X"00",X"75",X"C0",X"D5",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",
		X"15",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"A5",X"55",X"65",X"55",X"55",X"FF",X"FF",X"00",
		X"55",X"C0",X"15",X"C0",X"05",X"C0",X"55",X"C0",X"57",X"C0",X"7F",X"00",X"C0",X"00",X"00",X"00",
		X"F5",X"55",X"0D",X"55",X"03",X"55",X"02",X"D5",X"0A",X"D7",X"0A",X"B7",X"02",X"AF",X"00",X"0F",
		X"5F",X"AA",X"75",X"C0",X"D5",X"7A",X"D5",X"5E",X"55",X"5C",X"55",X"57",X"55",X"55",X"55",X"D5",
		X"00",X"0F",X"00",X"AB",X"0A",X"AB",X"02",X"AD",X"00",X"BD",X"00",X"35",X"02",X"D5",X"2A",X"D5",
		X"55",X"F5",X"55",X"ED",X"57",X"ED",X"57",X"AD",X"57",X"AB",X"55",X"EB",X"55",X"7F",X"55",X"57",
		X"AA",X"C0",X"00",X"C0",X"AA",X"C0",X"AA",X"C0",X"00",X"C0",X"AB",X"00",X"EB",X"00",X"7B",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"57",X"F5",X"7D",
		X"7D",X"55",X"5D",X"55",X"57",X"55",X"7F",X"57",X"55",X"DC",X"5F",X"F0",X"55",X"C0",X"FF",X"FF",
		X"55",X"57",X"55",X"75",X"5F",X"5F",X"F0",X"D5",X"00",X"35",X"00",X"3F",X"00",X"00",X"FC",X"00",
		X"00",X"D5",X"03",X"55",X"03",X"57",X"03",X"5D",X"03",X"5D",X"03",X"5D",X"03",X"55",X"03",X"6A",
		X"55",X"55",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"05",X"55",
		X"03",X"5A",X"03",X"5A",X"00",X"D6",X"00",X"D5",X"00",X"35",X"00",X"0F",X"00",X"03",X"00",X"00",
		X"01",X"55",X"01",X"55",X"81",X"55",X"A9",X"55",X"69",X"55",X"55",X"55",X"F5",X"55",X"0F",X"FF",
		X"55",X"55",X"FF",X"FD",X"55",X"57",X"55",X"55",X"55",X"55",X"45",X"55",X"05",X"55",X"55",X"0A",
		X"70",X"00",X"70",X"00",X"5C",X"00",X"DF",X"00",X"D7",X"00",X"D7",X"00",X"57",X"00",X"97",X"00",
		X"54",X"0A",X"54",X"0A",X"54",X"29",X"56",X"A5",X"56",X"95",X"55",X"57",X"55",X"7C",X"FF",X"F0",
		X"5C",X"00",X"5C",X"00",X"5C",X"00",X"70",X"00",X"70",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"35",X"55",X"0D",X"55",X"03",X"55",X"02",X"D5",X"0A",X"D5",X"0A",X"95",X"02",X"A5",X"00",X"0D",
		X"5E",X"AA",X"57",X"00",X"57",X"AA",X"55",X"EA",X"55",X"7F",X"55",X"F5",X"57",X"D5",X"5D",X"55",
		X"00",X"0D",X"00",X"0B",X"00",X"2B",X"00",X"AB",X"00",X"2F",X"00",X"0D",X"00",X"F5",X"00",X"D5",
		X"75",X"55",X"55",X"55",X"55",X"57",X"55",X"5E",X"55",X"7A",X"55",X"EA",X"55",X"7F",X"55",X"57",
		X"A0",X"3F",X"30",X"F5",X"B3",X"D5",X"FF",X"55",X"55",X"D7",X"55",X"7C",X"55",X"70",X"55",X"5C",
		X"00",X"00",X"C0",X"00",X"70",X"00",X"5F",X"00",X"55",X"F0",X"D5",X"5C",X"35",X"FC",X"0D",X"5C",
		X"5D",X"57",X"F7",X"55",X"D7",X"55",X"DC",X"D5",X"F0",X"37",X"C0",X"35",X"00",X"0D",X"FF",X"FF",
		X"CD",X"7C",X"73",X"5C",X"5C",X"FC",X"DC",X"00",X"7C",X"00",X"F0",X"00",X"70",X"00",X"C0",X"00",
		X"03",X"FF",X"0D",X"55",X"3F",X"FF",X"00",X"00",X"28",X"02",X"82",X"08",X"00",X"A0",X"00",X"00",
		X"55",X"55",X"55",X"55",X"FF",X"FD",X"02",X"AD",X"8A",X"8D",X"28",X"D5",X"0F",X"55",X"F5",X"56",
		X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"35",X"54",X"35",X"50",X"35",X"55",X"0F",X"55",X"00",X"FF",
		X"55",X"5A",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"55",X"DE",X"57",X"57",X"5D",X"55",X"57",X"F5",X"5D",X"55",X"57",X"55",X"55",X"D5",X"AA",X"55",
		X"A0",X"00",X"E0",X"00",X"C0",X"00",X"70",X"00",X"70",X"00",X"7C",X"00",X"5E",X"00",X"5E",X"80",
		X"AA",X"95",X"0A",X"55",X"09",X"55",X"05",X"55",X"15",X"55",X"55",X"57",X"57",X"FC",X"FF",X"00",
		X"5E",X"00",X"5C",X"00",X"5C",X"00",X"5E",X"00",X"7A",X"00",X"EA",X"80",X"00",X"00",X"00",X"00",
		X"D5",X"55",X"35",X"55",X"0F",X"55",X"0A",X"D5",X"0A",X"B5",X"0A",X"B5",X"00",X"3D",X"00",X"03",
		X"57",X"AA",X"55",X"00",X"55",X"FE",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",
		X"00",X"03",X"00",X"0A",X"00",X"0A",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"03",
		X"57",X"FA",X"D7",X"00",X"D7",X"AA",X"D7",X"AA",X"D5",X"C0",X"D5",X"7A",X"D5",X"5F",X"55",X"55",
		X"AA",X"C0",X"00",X"C0",X"AA",X"C0",X"FF",X"C0",X"55",X"FC",X"55",X"57",X"55",X"55",X"F5",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"F0",X"FD",X"5C",X"55",X"5F",X"55",X"55",
		X"AF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"30",X"00",X"AC",X"00",X"EA",X"00",X"7F",X"FA",
		X"F5",X"7D",X"0D",X"57",X"0D",X"75",X"03",X"5F",X"00",X"D5",X"00",X"35",X"00",X"0F",X"A0",X"00",
		X"99",X"99",X"66",X"66",X"9C",X"CC",X"6C",X"CC",X"9E",X"AA",X"6E",X"55",X"9E",X"69",X"6E",X"69",
		X"99",X"99",X"66",X"66",X"CC",X"CC",X"CC",X"CC",X"AA",X"AA",X"A5",X"59",X"A6",X"99",X"A6",X"99",
		X"9E",X"A9",X"6E",X"A9",X"9E",X"A5",X"6E",X"AA",X"9C",X"CC",X"6C",X"CC",X"99",X"99",X"66",X"66",
		X"A6",X"99",X"A6",X"99",X"66",X"99",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",X"99",X"99",X"66",X"66",
		X"99",X"99",X"66",X"66",X"CC",X"CC",X"CC",X"CC",X"AA",X"AA",X"A6",X"99",X"A6",X"99",X"99",X"99",
		X"99",X"98",X"66",X"64",X"CC",X"D8",X"CC",X"E4",X"AA",X"D8",X"AA",X"E4",X"AA",X"D8",X"56",X"E4",
		X"99",X"99",X"6A",X"59",X"6A",X"59",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",X"99",X"99",X"66",X"66",
		X"A6",X"D8",X"A6",X"E4",X"56",X"D8",X"AA",X"E4",X"CC",X"D8",X"CC",X"E4",X"99",X"98",X"66",X"64",
		X"00",X"2A",X"00",X"02",X"0A",X"80",X"2A",X"A2",X"AA",X"AA",X"5A",X"82",X"56",X"80",X"55",X"45",
		X"80",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"88",X"00",X"A0",X"00",X"00",X"20",X"40",X"08",
		X"55",X"55",X"55",X"58",X"55",X"60",X"55",X"80",X"5A",X"00",X"A8",X"00",X"80",X"00",X"00",X"00",
		X"50",X"2A",X"50",X"AA",X"50",X"AA",X"50",X"68",X"11",X"50",X"15",X"40",X"05",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"02",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"00",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"00",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"0A",
		X"00",X"00",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"A0",X"0A",X"A0",X"02",X"A8",X"02",X"AA",X"00",X"AA",X"00",X"00",
		X"AA",X"80",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"AA",X"80",X"A8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"14",X"00",X"40",X"01",X"2A",X"01",X"28",X"04",X"28",
		X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"00",X"40",X"AA",X"10",X"00",X"10",X"00",X"04",
		X"04",X"2A",X"04",X"28",X"01",X"28",X"01",X"2A",X"00",X"40",X"00",X"14",X"00",X"01",X"00",X"00",
		X"A8",X"04",X"00",X"04",X"00",X"10",X"AA",X"10",X"00",X"40",X"05",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"14",X"00",X"40",X"01",X"28",X"01",X"0A",X"04",X"02",
		X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"00",X"40",X"0A",X"10",X"28",X"10",X"20",X"04",
		X"04",X"00",X"04",X"02",X"01",X"0A",X"01",X"28",X"00",X"40",X"00",X"14",X"00",X"01",X"00",X"00",
		X"80",X"04",X"20",X"04",X"28",X"10",X"0A",X"10",X"00",X"40",X"05",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"14",X"00",X"40",X"01",X"00",X"01",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"80",X"40",X"80",X"10",X"80",X"10",X"80",X"04",
		X"04",X"00",X"04",X"00",X"01",X"2A",X"01",X"2A",X"00",X"40",X"00",X"14",X"00",X"01",X"00",X"00",
		X"80",X"04",X"80",X"04",X"AA",X"10",X"AA",X"10",X"00",X"40",X"05",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"14",X"00",X"40",X"01",X"28",X"01",X"28",X"04",X"28",
		X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"00",X"40",X"0A",X"10",X"28",X"10",X"A0",X"04",
		X"04",X"2A",X"04",X"28",X"01",X"28",X"01",X"2A",X"00",X"40",X"00",X"14",X"00",X"01",X"00",X"00",
		X"A8",X"04",X"02",X"04",X"02",X"10",X"A8",X"10",X"00",X"40",X"05",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"14",X"00",X"40",X"01",X"28",X"01",X"28",X"04",X"2A",
		X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"00",X"40",X"0A",X"10",X"0A",X"10",X"AA",X"04",
		X"04",X"28",X"04",X"08",X"01",X"0A",X"01",X"02",X"00",X"40",X"00",X"14",X"00",X"01",X"00",X"00",
		X"0A",X"04",X"08",X"04",X"28",X"10",X"A0",X"10",X"80",X"40",X"05",X"00",X"50",X"00",X"00",X"00",
		X"17",X"FA",X"17",X"FE",X"17",X"FE",X"15",X"FF",X"15",X"7F",X"05",X"5E",X"05",X"57",X"01",X"55",
		X"AA",X"AB",X"AA",X"BF",X"AB",X"FF",X"AD",X"EF",X"FF",X"F5",X"FF",X"FF",X"FE",X"D5",X"7F",X"D5",
		X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"50",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"55",X"F5",X"40",X"55",X"55",X"D5",X"54",X"55",X"41",X"55",X"54",X"54",X"00",X"55",X"05",
		X"55",X"54",X"50",X"00",X"00",X"00",X"01",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"15",X"00",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"55",X"50",X"55",X"41",X"55",X"55",X"55",X"55",
		X"01",X"55",X"01",X"5F",X"05",X"5F",X"05",X"7B",X"15",X"7F",X"15",X"FE",X"15",X"FA",X"17",X"FA",
		X"73",X"D5",X"FF",X"F5",X"FE",X"F7",X"AB",X"FD",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"54",X"00",X"50",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"05",X"50",X"40",X"F5",X"55",X"4F",X"54",X"55",X"01",X"F5",X"55",X"FF",X"94",X"AF",X"F5",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"51",X"00",
		X"57",X"EA",X"17",X"FA",X"15",X"FF",X"05",X"7E",X"05",X"57",X"01",X"55",X"01",X"55",X"00",X"15",
		X"AA",X"AA",X"AA",X"BF",X"9A",X"2D",X"FF",X"FF",X"FB",X"FF",X"7F",X"F5",X"55",X"7F",X"55",X"55",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"F5",X"F5",X"55",X"3F",X"41",X"D5",X"54",X"75",X"55",X"55",X"45",X"55",X"50",X"50",X"00",
		X"55",X"50",X"51",X"40",X"54",X"00",X"00",X"00",X"01",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"15",X"40",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"40",X"55",X"55",X"55",X"50",X"55",X"55",
		X"01",X"55",X"05",X"55",X"05",X"57",X"15",X"7F",X"15",X"FF",X"15",X"FE",X"57",X"FA",X"57",X"EA",
		X"55",X"7F",X"7F",X"D5",X"FF",X"FF",X"F7",X"BC",X"2E",X"FF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"55",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"41",X"54",X"55",X"00",X"5F",X"54",X"F5",X"75",X"FD",X"D4",X"FF",X"F5",X"FF",X"FD",X"AB",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"40",X"14",X"00",X"50",X"00",X"45",X"40",X"FD",X"55",
		X"01",X"55",X"05",X"7F",X"15",X"7F",X"50",X"3F",X"55",X"55",X"58",X"14",X"58",X"14",X"5A",X"96",
		X"50",X"00",X"54",X"00",X"55",X"10",X"01",X"54",X"55",X"55",X"25",X"55",X"25",X"44",X"A5",X"04",
		X"15",X"55",X"05",X"55",X"20",X"0C",X"20",X"3F",X"20",X"3F",X"28",X"00",X"0A",X"00",X"02",X"AA",
		X"55",X"05",X"54",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"28",X"00",X"A0",X"00",
		X"01",X"DD",X"1D",X"DD",X"DE",X"AA",X"EA",X"AB",X"2A",X"AB",X"2A",X"AA",X"0A",X"4A",X"09",X"56",
		X"DD",X"DC",X"DD",X"DD",X"AA",X"A9",X"AE",X"AA",X"AE",X"AA",X"EB",X"AA",X"B0",X"A8",X"80",X"00",
		X"01",X"56",X"01",X"54",X"01",X"54",X"01",X"54",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"03",X"FF",X"03",X"FF",X"00",X"FC",X"00",X"FE",X"03",X"CE",X"0A",X"FE",X"2A",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"A9",X"80",X"A5",X"60",X"95",X"58",X"55",X"56",
		X"15",X"55",X"1F",X"FD",X"1C",X"CD",X"1F",X"FD",X"1C",X"CD",X"1F",X"FD",X"15",X"55",X"15",X"55",
		X"55",X"54",X"55",X"54",X"55",X"54",X"57",X"F4",X"57",X"B4",X"57",X"F4",X"57",X"F4",X"57",X"F4",
		X"01",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"05",X"55",
		X"55",X"40",X"55",X"50",X"55",X"D4",X"55",X"74",X"55",X"74",X"55",X"74",X"55",X"D4",X"55",X"50",
		X"81",X"55",X"AA",X"AA",X"2A",X"55",X"08",X"55",X"08",X"55",X"28",X"15",X"20",X"05",X"A0",X"01",
		X"55",X"40",X"A8",X"00",X"5D",X"00",X"5D",X"00",X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",
		X"05",X"01",X"15",X"99",X"16",X"59",X"16",X"40",X"58",X"00",X"59",X"50",X"56",X"59",X"56",X"65",
		X"40",X"50",X"66",X"54",X"65",X"94",X"00",X"94",X"01",X"65",X"05",X"65",X"65",X"95",X"59",X"95",
		X"59",X"25",X"58",X"05",X"60",X"01",X"65",X"59",X"65",X"65",X"49",X"65",X"19",X"03",X"00",X"03",
		X"59",X"25",X"50",X"29",X"40",X"09",X"65",X"59",X"59",X"59",X"59",X"65",X"C0",X"64",X"C0",X"00",
		X"00",X"00",X"00",X"05",X"00",X"55",X"01",X"5F",X"01",X"7C",X"05",X"7C",X"05",X"5F",X"15",X"55",
		X"00",X"00",X"50",X"00",X"55",X"00",X"F5",X"40",X"FD",X"40",X"FD",X"50",X"F5",X"50",X"55",X"54",
		X"15",X"0A",X"15",X"5A",X"55",X"5A",X"55",X"56",X"55",X"55",X"00",X"0A",X"00",X"22",X"00",X"14",
		X"A0",X"54",X"A5",X"54",X"A5",X"55",X"95",X"55",X"55",X"55",X"A0",X"00",X"88",X"00",X"14",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
