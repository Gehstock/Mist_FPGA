library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj_7p is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj_7p is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"00",X"00",X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"3F",X"1F",
		X"0C",X"18",X"1C",X"18",X"00",X"00",X"00",X"40",X"E0",X"C0",X"00",X"00",X"07",X"1F",X"3F",X"1F",
		X"30",X"60",X"60",X"60",X"00",X"00",X"00",X"20",X"60",X"40",X"00",X"00",X"07",X"1F",X"3F",X"1F",
		X"78",X"38",X"00",X"00",X"00",X"40",X"E0",X"C0",X"80",X"00",X"00",X"00",X"07",X"1F",X"3F",X"1F",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"1C",X"08",X"18",X"38",X"38",X"30",X"00",X"00",X"00",X"03",X"0F",X"1F",X"0F",X"0F",
		X"00",X"00",X"20",X"30",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"0F",X"0F",
		X"00",X"00",X"3C",X"00",X"00",X"40",X"E0",X"C0",X"00",X"1F",X"7F",X"3B",X"1E",X"00",X"00",X"00",
		X"7C",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"70",X"38",X"10",X"40",X"E0",X"C0",X"00",X"00",X"1F",X"7F",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0E",X"04",X"00",X"00",X"00",
		X"7D",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"20",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"20",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"FF",X"7F",
		X"78",X"00",X"00",X"00",X"00",X"C0",X"E0",X"00",X"00",X"0F",X"3F",X"1F",X"1F",X"0F",X"00",X"00",
		X"78",X"00",X"00",X"C0",X"C0",X"00",X"00",X"1F",X"7F",X"3F",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"E0",X"E0",X"C0",X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"EF",X"ED",X"2C",X"07",
		X"30",X"70",X"E0",X"E0",X"C0",X"80",X"C1",X"C3",X"03",X"07",X"07",X"07",X"0F",X"0D",X"0C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"11",X"11",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"47",X"E0",X"C0",X"C0",X"40",X"00",X"00",X"40",X"C0",X"C0",X"C1",X"0B",X"1F",
		X"0F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"EF",X"7F",X"3F",X"1F",
		X"00",X"00",X"02",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"0F",X"0F",
		X"00",X"00",X"3F",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"40",X"3F",
		X"08",X"09",X"06",X"04",X"03",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"20",X"10",X"08",X"06",
		X"5B",X"BF",X"1B",X"11",X"41",X"01",X"01",X"02",X"12",X"03",X"02",X"02",X"06",X"06",X"1A",X"0A",
		X"0A",X"09",X"09",X"06",X"01",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"20",X"10",X"08",X"06",
		X"35",X"7F",X"23",X"11",X"01",X"24",X"85",X"0A",X"0C",X"0C",X"0C",X"19",X"19",X"09",X"09",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"1E",X"7E",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"1E",X"7E",X"FE",X"FE",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"3E",X"7E",X"FE",X"FE",X"FC",X"BE",X"BE",X"3E",X"3E",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BE",X"BE",X"BE",X"BE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"BF",X"BF",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"2F",X"4F",X"17",X"22",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"60",X"C0",X"C0",X"04",X"03",X"07",X"17",X"1F",X"3F",X"3F",X"7F",X"FF",X"DD",X"5F",X"3F",
		X"20",X"60",X"C0",X"C0",X"04",X"83",X"C7",X"EF",X"7F",X"7F",X"3F",X"1F",X"0F",X"1D",X"1F",X"3F",
		X"2F",X"0F",X"1F",X"0F",X"17",X"07",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"03",X"60",X"40",X"40",X"00",X"04",X"0E",X"4E",X"FE",X"FE",X"FF",X"0B",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FE",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"10",X"20",X"20",X"00",X"80",X"40",X"00",X"70",X"7F",X"F3",X"E7",X"4F",X"0E",X"06",X"00",
		X"08",X"10",X"20",X"20",X"00",X"00",X"40",X"80",X"30",X"3F",X"33",X"73",X"71",X"21",X"00",X"00",
		X"E0",X"7F",X"61",X"C0",X"00",X"80",X"00",X"40",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"70",X"7D",X"7F",X"61",X"C0",X"00",X"80",X"00",X"40",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"FB",X"7F",X"61",X"C0",X"00",X"80",X"00",X"40",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"F9",X"7F",X"61",X"C0",X"00",X"80",X"00",X"40",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"F9",X"FF",X"61",X"C0",X"00",X"80",X"00",X"40",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1C",X"41",X"21",X"00",X"03",X"07",X"0E",X"0D",X"03",X"03",X"03",X"03",X"01",X"01",X"00",
		X"01",X"0D",X"0E",X"23",X"40",X"03",X"07",X"0E",X"0D",X"03",X"03",X"03",X"03",X"01",X"01",X"00",
		X"0E",X"1C",X"00",X"10",X"21",X"03",X"07",X"06",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"F4",X"72",X"30",X"00",X"00",X"00",X"CB",X"CB",X"7B",X"37",X"03",X"03",X"03",X"01",X"01",X"00",
		X"03",X"03",X"02",X"00",X"00",X"00",X"06",X"1D",X"3D",X"7B",X"F7",X"E7",X"67",X"26",X"02",X"01",
		X"06",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"0F",X"07",X"04",X"7E",X"37",X"0F",
		X"06",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"10",X"20",X"20",X"00",X"00",X"00",X"00",X"70",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"10",X"20",X"20",X"00",X"00",X"40",X"00",X"70",X"7F",X"37",X"00",X"00",X"00",X"00",X"00",
		X"08",X"10",X"20",X"20",X"00",X"80",X"40",X"00",X"70",X"7F",X"73",X"27",X"01",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"06",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"06",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"67",X"31",X"19",X"1C",X"0E",X"0C",X"09",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"1F",X"4E",X"64",X"31",X"19",X"1C",X"1C",X"0C",X"08",X"00",X"01",X"01",X"01",X"01",X"00",X"00",
		X"1F",X"0E",X"04",X"21",X"11",X"10",X"0C",X"0C",X"00",X"09",X"0A",X"02",X"01",X"01",X"00",X"00",
		X"0C",X"04",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"21",X"10",X"00",X"00",X"00",X"00",
		X"10",X"01",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"08",X"40",X"00",X"01",X"00",X"00",
		X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"3C",X"0C",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"8E",X"4F",X"0F",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"E8",X"DC",X"BE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"70",X"1F",X"87",X"E0",X"78",X"1F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"78",X"1F",X"87",X"E0",X"78",X"1F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"00",X"60",X"6F",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"0E",X"0E",X"10",X"11",X"E1",X"E0",X"0E",X"0E",
		X"00",X"00",X"00",X"E0",X"EE",X"0E",X"10",X"10",X"01",X"E1",X"EE",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"E1",X"E1",X"10",X"10",X"0E",X"0E",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"FF",X"FF",X"BB",X"BB",X"B7",X"7F",X"DD",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"FF",X"FF",X"BB",X"BB",X"B7",X"7F",X"DD",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7B",X"77",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"09",X"09",X"0F",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"61",X"12",X"1E",X"0B",X"79",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C1",X"C3",X"F3",X"3F",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"B8",X"FC",X"7C",X"3C",X"1F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"C3",X"C3",X"C3",X"FF",X"FF",X"00",
		X"00",X"03",X"0E",X"18",X"12",X"36",X"2A",X"2B",X"29",X"28",X"28",X"14",X"1B",X"0C",X"03",X"00",
		X"00",X"00",X"00",X"01",X"02",X"02",X"22",X"36",X"3D",X"11",X"13",X"08",X"04",X"03",X"00",X"00",
		X"00",X"03",X"0C",X"0B",X"16",X"14",X"14",X"13",X"0C",X"03",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0E",X"0A",X"15",X"16",X"15",X"15",X"0B",X"08",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"0E",X"05",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"04",X"05",X"05",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"05",X"04",X"05",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"06",X"06",X"06",X"06",X"06",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",
		X"7F",X"E0",X"1F",X"30",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"54",X"54",X"50",X"43",X"77",X"07",X"17",X"27",X"72",X"50",X"52",X"42",X"20",X"00",X"00",X"00",
		X"A4",X"A4",X"90",X"43",X"77",X"07",X"37",X"67",X"E2",X"A0",X"82",X"C2",X"00",X"00",X"00",X"00",
		X"04",X"A8",X"A8",X"50",X"43",X"37",X"07",X"37",X"27",X"72",X"68",X"62",X"32",X"18",X"00",X"00",
		X"A8",X"A8",X"92",X"42",X"72",X"26",X"57",X"E7",X"F7",X"D2",X"D0",X"40",X"71",X"03",X"04",X"08",
		X"54",X"54",X"22",X"32",X"02",X"06",X"37",X"67",X"C7",X"E2",X"F0",X"D0",X"D1",X"E3",X"74",X"38",
		X"24",X"48",X"42",X"42",X"32",X"06",X"77",X"C7",X"E7",X"F2",X"D0",X"D0",X"61",X"33",X"04",X"08",
		X"60",X"6A",X"C0",X"F0",X"E3",X"C7",X"57",X"67",X"0F",X"77",X"48",X"90",X"20",X"00",X"00",X"00",
		X"60",X"6A",X"C0",X"F0",X"E3",X"C7",X"57",X"67",X"0F",X"17",X"28",X"28",X"24",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"FF",X"63",X"C0",X"00",X"00",X"00",X"40",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"7F",X"3F",X"63",X"01",X"03",X"23",X"27",X"15",X"17",X"06",X"04",X"00",X"00",X"00",X"00",
		X"38",X"1D",X"3F",X"07",X"06",X"07",X"27",X"7F",X"7F",X"7F",X"5B",X"31",X"31",X"10",X"00",X"00",
		X"38",X"1F",X"1F",X"08",X"0B",X"4F",X"CF",X"FF",X"FF",X"BE",X"EE",X"C6",X"46",X"44",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"7F",X"7F",X"7F",X"7F",X"3B",X"30",X"33",X"27",X"20",X"26",X"20",X"26",X"2B",X"24",X"33",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3C",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"01",X"03",X"07",X"0E",X"1F",X"1E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3C",
		X"03",X"00",X"00",X"00",X"F8",X"87",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"00",X"00",X"00",X"0F",X"F8",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"00",X"00",X"00",X"01",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"88",X"62",X"32",X"0A",X"3E",X"2F",X"77",X"77",X"FA",X"D8",X"CE",X"CD",X"67",X"64",X"38",
		X"04",X"08",X"08",X"0B",X"03",X"02",X"01",X"01",X"01",X"03",X"07",X"06",X"06",X"06",X"06",X"02",
		X"05",X"09",X"08",X"03",X"03",X"03",X"1B",X"33",X"63",X"F1",X"FB",X"DB",X"CB",X"6B",X"63",X"30",
		X"04",X"08",X"08",X"0B",X"03",X"02",X"01",X"01",X"01",X"03",X"07",X"06",X"06",X"06",X"06",X"02",
		X"00",X"03",X"17",X"1F",X"00",X"05",X"05",X"01",X"0C",X"0E",X"0A",X"1E",X"34",X"0E",X"3E",X"1C",
		X"00",X"0B",X"17",X"0F",X"00",X"05",X"05",X"01",X"1C",X"7E",X"FA",X"F6",X"E0",X"40",X"00",X"00",
		X"00",X"03",X"17",X"1F",X"00",X"25",X"85",X"C1",X"FC",X"7E",X"0A",X"06",X"00",X"00",X"00",X"00",
		X"07",X"2F",X"B0",X"C8",X"66",X"23",X"0C",X"1E",X"0A",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"EA",X"FE",X"1C",X"01",X"05",X"05",X"00",X"1F",X"17",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"46",X"EA",X"FE",X"1C",X"01",X"05",X"05",X"00",X"1F",X"27",X"03",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"3F",X"3F",X"1A",X"1D",X"0F",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"3F",X"3A",X"1D",X"1F",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"3F",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"3F",X"3F",X"1A",X"1D",X"0F",X"0E",X"0E",X"0E",X"05",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"07",X"0A",X"0A",X"0F",X"07",X"02",X"0A",X"07",X"02",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"20",X"20",X"60",X"60",X"60",X"60",X"60",X"60",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"30",X"10",X"00",X"00",
		X"00",X"08",X"18",X"38",X"38",X"78",X"78",X"78",X"78",X"78",X"78",X"38",X"38",X"18",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"06",X"06",X"06",X"06",X"06",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"0B",X"0A",X"0A",X"0A",X"0A",X"0A",X"0B",X"04",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"04",X"09",X"0A",X"00",X"0A",X"09",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"08",X"13",X"16",X"14",X"00",X"14",X"16",X"13",X"08",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"05",X"07",X"02",X"07",X"05",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"19",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"04",X"04",X"05",X"0B",X"00",
		X"00",X"00",X"00",X"03",X"04",X"09",X"09",X"09",X"09",X"04",X"04",X"02",X"02",X"05",X"09",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"08",X"10",X"20",X"20",X"00",X"00",X"40",X"80",X"70",X"3F",X"33",X"73",X"71",X"21",X"00",X"00",
		X"36",X"08",X"20",X"20",X"30",X"70",X"78",X"24",X"1E",X"3F",X"38",X"13",X"07",X"07",X"05",X"03",
		X"00",X"00",X"00",X"06",X"0F",X"07",X"03",X"31",X"7A",X"B2",X"FE",X"FE",X"DF",X"5E",X"3C",X"18",
		X"00",X"03",X"5B",X"FB",X"D5",X"DC",X"F4",X"F3",X"FE",X"FC",X"7C",X"34",X"00",X"00",X"00",X"00",
		X"0F",X"19",X"1F",X"1F",X"1E",X"0F",X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"20",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"44",X"9C",X"0E",X"0E",X"04",
		X"30",X"65",X"D0",X"D0",X"F3",X"E7",X"5B",X"33",X"03",X"39",X"2C",X"48",X"90",X"00",X"00",X"00",
		X"3C",X"70",X"6C",X"78",X"20",X"1F",X"07",X"1B",X"23",X"29",X"09",X"00",X"03",X"00",X"00",X"01",
		X"01",X"00",X"00",X"03",X"00",X"08",X"2B",X"27",X"1B",X"03",X"1B",X"21",X"7C",X"30",X"1E",X"1C",
		X"00",X"00",X"00",X"10",X"92",X"4A",X"34",X"0F",X"67",X"D7",X"E7",X"E7",X"B1",X"41",X"2A",X"00",
		X"00",X"61",X"F2",X"EA",X"A4",X"25",X"0F",X"0F",X"0F",X"27",X"17",X"01",X"04",X"02",X"02",X"00",
		X"00",X"02",X"04",X"00",X"10",X"27",X"27",X"0F",X"0F",X"6F",X"C3",X"A1",X"EA",X"FA",X"39",X"10",
		X"06",X"0A",X"0E",X"1C",X"41",X"E5",X"E5",X"C0",X"1F",X"17",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1F",X"19",X"16",X"00",X"08",X"16",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"16",X"08",X"00",X"0E",X"1D",X"19",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"05",X"0B",X"0F",X"40",X"D2",X"E2",X"78",X"3E",X"07",X"05",X"03",
		X"00",X"30",X"79",X"1A",X"4B",X"73",X"25",X"08",X"62",X"D4",X"F1",X"62",X"18",X"34",X"3C",X"18",
		X"18",X"3C",X"34",X"18",X"62",X"F1",X"D4",X"62",X"08",X"25",X"33",X"2B",X"2E",X"35",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"18",X"18",X"18",X"18",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"66",X"76",X"5E",X"4E",X"46",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"7F",X"7F",X"00",X"D9",X"FB",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"00",X"7F",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"D9",X"FA",X"AA",X"AA",X"A9",X"00",X"7F",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"FB",X"AA",X"AB",X"7F",X"7F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
