library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dderby_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dderby_sp_bits_1 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"77",X"00",X"00",X"77",X"22",X"00",X"00",X"26",X"79",
		X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"69",X"00",X"00",X"22",X"79",X"00",X"00",X"72",X"99",
		X"00",X"00",X"77",X"99",X"00",X"00",X"72",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"99",
		X"00",X"00",X"26",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"72",X"99",X"00",X"00",X"77",X"99",
		X"00",X"00",X"72",X"99",X"00",X"00",X"22",X"79",X"00",X"00",X"99",X"69",X"00",X"00",X"22",X"99",
		X"00",X"00",X"26",X"79",X"00",X"00",X"77",X"22",X"00",X"00",X"99",X"77",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"77",X"00",X"22",X"77",X"77",X"00",X"96",X"22",X"66",X"00",
		X"99",X"22",X"99",X"00",X"22",X"72",X"29",X"00",X"66",X"72",X"27",X"00",X"66",X"92",X"27",X"00",
		X"66",X"92",X"27",X"00",X"66",X"92",X"27",X"00",X"66",X"92",X"27",X"00",X"66",X"92",X"67",X"00",
		X"66",X"92",X"27",X"00",X"66",X"92",X"27",X"00",X"66",X"92",X"27",X"00",X"66",X"92",X"27",X"00",
		X"66",X"92",X"27",X"00",X"66",X"72",X"27",X"00",X"22",X"72",X"29",X"00",X"99",X"22",X"99",X"00",
		X"96",X"22",X"66",X"00",X"22",X"77",X"77",X"00",X"99",X"99",X"77",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"90",X"00",X"00",X"0E",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"99",X"67",X"00",X"00",X"99",X"26",X"00",X"00",X"90",X"22",X"00",X"00",X"99",X"99",
		X"00",X"00",X"72",X"29",X"00",X"00",X"22",X"92",X"00",X"00",X"26",X"92",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"29",X"00",X"00",X"27",X"22",X"00",X"00",X"27",X"96",X"00",X"00",X"22",X"77",
		X"00",X"00",X"22",X"69",X"00",X"00",X"92",X"29",X"00",X"00",X"29",X"79",X"00",X"00",X"66",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"69",X"70",X"00",X"00",
		X"29",X"29",X"00",X"00",X"62",X"22",X"00",X"00",X"66",X"72",X"00",X"00",X"66",X"62",X"90",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"66",X"00",X"66",X"99",X"22",X"00",
		X"00",X"00",X"77",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"79",
		X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"92",X"00",X"66",X"97",X"22",X"00",X"66",X"92",X"22",X"00",X"66",X"92",X"27",X"00",
		X"66",X"72",X"27",X"00",X"22",X"22",X"27",X"00",X"92",X"22",X"70",X"00",X"99",X"29",X"70",X"00",
		X"69",X"29",X"70",X"00",X"22",X"92",X"00",X"00",X"72",X"92",X"00",X"00",X"09",X"92",X"90",X"00",
		X"00",X"29",X"99",X"00",X"00",X"62",X"09",X"00",X"00",X"76",X"99",X"00",X"00",X"97",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"76",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",
		X"00",X"00",X"09",X"22",X"00",X"00",X"99",X"72",X"00",X"00",X"90",X"27",X"00",X"00",X"07",X"22",
		X"00",X"00",X"02",X"92",X"00",X"00",X"79",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"62",X"92",
		X"00",X"00",X"26",X"29",X"00",X"00",X"22",X"26",X"00",X"00",X"92",X"97",X"00",X"00",X"99",X"69",
		X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"26",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",X"00",
		X"66",X"79",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"62",X"00",X"00",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"22",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"92",X"00",X"00",
		X"66",X"92",X"90",X"00",X"66",X"22",X"99",X"00",X"62",X"22",X"99",X"00",X"29",X"22",X"79",X"00",
		X"99",X"29",X"29",X"00",X"99",X"29",X"62",X"00",X"99",X"92",X"26",X"00",X"79",X"66",X"26",X"00",
		X"79",X"62",X"02",X"00",X"22",X"26",X"09",X"00",X"22",X"22",X"09",X"00",X"97",X"22",X"99",X"00",
		X"97",X"22",X"90",X"00",X"99",X"22",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"97",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"07",X"72",X"00",X"00",X"02",X"72",X"00",X"00",X"02",X"27",
		X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"32",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"26",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"77",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"72",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"77",X"00",X"00",
		X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"27",X"00",X"00",X"66",X"67",X"00",X"00",X"66",X"67",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"77",X"00",X"00",X"99",X"27",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"72",X"00",X"00",X"99",X"99",X"00",X"00",X"72",X"29",X"00",X"00",
		X"22",X"29",X"00",X"00",X"79",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",
		X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"29",X"79",X"00",X"00",X"29",X"00",X"00",X"00",
		X"69",X"00",X"00",X"00",X"69",X"99",X"00",X"00",X"67",X"99",X"00",X"00",X"06",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"70",X"00",X"00",X"3E",X"77",X"00",
		X"00",X"99",X"27",X"90",X"00",X"26",X"62",X"90",X"00",X"26",X"22",X"90",X"00",X"22",X"62",X"90",
		X"00",X"26",X"22",X"90",X"00",X"22",X"62",X"90",X"00",X"76",X"22",X"79",X"00",X"72",X"62",X"99",
		X"00",X"76",X"92",X"99",X"00",X"72",X"92",X"99",X"00",X"76",X"99",X"99",X"00",X"72",X"92",X"99",
		X"00",X"72",X"77",X"99",X"00",X"22",X"62",X"79",X"00",X"22",X"99",X"79",X"00",X"29",X"99",X"70",
		X"00",X"72",X"99",X"70",X"00",X"97",X"77",X"70",X"00",X"29",X"66",X"70",X"00",X"26",X"66",X"70",
		X"00",X"22",X"66",X"70",X"00",X"22",X"66",X"70",X"00",X"29",X"66",X"70",X"00",X"29",X"66",X"70",
		X"00",X"29",X"66",X"70",X"00",X"69",X"66",X"70",X"00",X"69",X"66",X"70",X"00",X"69",X"66",X"70",
		X"00",X"69",X"66",X"70",X"00",X"69",X"22",X"70",X"00",X"79",X"99",X"70",X"00",X"72",X"99",X"70",
		X"00",X"72",X"99",X"70",X"00",X"72",X"99",X"70",X"00",X"77",X"99",X"90",X"00",X"76",X"77",X"99",
		X"00",X"76",X"22",X"99",X"00",X"76",X"22",X"99",X"00",X"76",X"97",X"99",X"00",X"76",X"22",X"99",
		X"00",X"76",X"62",X"99",X"00",X"76",X"22",X"99",X"00",X"76",X"62",X"79",X"00",X"76",X"22",X"79",
		X"00",X"76",X"62",X"70",X"00",X"76",X"99",X"70",X"00",X"76",X"77",X"00",X"00",X"96",X"00",X"00",
		X"00",X"96",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9C",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",
		X"00",X"00",X"AB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"44",X"90",X"00",
		X"00",X"44",X"90",X"00",X"00",X"41",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"AD",
		X"00",X"00",X"00",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"AD",X"90",
		X"00",X"00",X"D9",X"00",X"00",X"09",X"DD",X"00",X"00",X"9D",X"DA",X"00",X"00",X"DA",X"DD",X"00",
		X"00",X"AA",X"D9",X"00",X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"0F",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"77",X"00",X"22",X"77",X"22",X"00",X"96",X"22",X"22",X"00",
		X"99",X"22",X"22",X"00",X"22",X"72",X"22",X"00",X"66",X"72",X"27",X"00",X"66",X"92",X"27",X"00",
		X"66",X"92",X"27",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",
		X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",
		X"66",X"92",X"97",X"00",X"66",X"72",X"97",X"00",X"22",X"72",X"99",X"00",X"99",X"22",X"99",X"00",
		X"96",X"22",X"96",X"00",X"22",X"77",X"67",X"00",X"99",X"99",X"77",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"69",X"70",X"00",X"00",
		X"29",X"29",X"00",X"00",X"62",X"22",X"00",X"00",X"66",X"72",X"00",X"00",X"66",X"62",X"90",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"66",X"00",X"66",X"99",X"22",X"00",
		X"66",X"99",X"22",X"00",X"66",X"97",X"22",X"00",X"66",X"92",X"22",X"00",X"66",X"92",X"97",X"00",
		X"66",X"72",X"97",X"00",X"22",X"22",X"97",X"00",X"92",X"22",X"70",X"00",X"99",X"29",X"70",X"00",
		X"99",X"29",X"70",X"00",X"22",X"92",X"00",X"00",X"72",X"92",X"00",X"00",X"09",X"99",X"90",X"00",
		X"00",X"29",X"99",X"00",X"00",X"69",X"09",X"00",X"00",X"76",X"90",X"00",X"00",X"96",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"22",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"92",X"00",X"00",
		X"66",X"92",X"00",X"00",X"66",X"22",X"90",X"00",X"62",X"22",X"99",X"00",X"29",X"22",X"79",X"00",
		X"99",X"29",X"22",X"00",X"99",X"29",X"22",X"00",X"99",X"92",X"29",X"00",X"79",X"66",X"99",X"00",
		X"79",X"62",X"09",X"00",X"22",X"99",X"09",X"00",X"22",X"99",X"09",X"00",X"97",X"99",X"99",X"00",
		X"97",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"97",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"27",X"00",X"00",X"66",X"67",X"00",X"00",X"66",X"67",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"27",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"72",X"00",X"00",X"99",X"29",X"00",X"00",X"92",X"29",X"00",X"00",
		X"22",X"22",X"00",X"00",X"79",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",
		X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"67",X"99",X"00",X"00",X"06",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"29",X"66",X"70",X"00",X"69",X"66",X"70",X"00",X"69",X"66",X"70",X"00",X"69",X"66",X"70",
		X"00",X"69",X"66",X"70",X"00",X"69",X"22",X"70",X"00",X"79",X"99",X"70",X"00",X"72",X"99",X"70",
		X"00",X"72",X"99",X"70",X"00",X"72",X"99",X"70",X"00",X"77",X"99",X"90",X"00",X"76",X"77",X"99",
		X"00",X"76",X"22",X"99",X"00",X"76",X"22",X"99",X"00",X"76",X"97",X"99",X"00",X"76",X"22",X"99",
		X"00",X"66",X"62",X"99",X"00",X"69",X"22",X"99",X"00",X"69",X"99",X"79",X"00",X"69",X"99",X"79",
		X"00",X"69",X"99",X"70",X"00",X"76",X"99",X"20",X"00",X"76",X"77",X"00",X"00",X"96",X"90",X"00",
		X"00",X"96",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"77",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"79",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"79",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"99",
		X"00",X"00",X"26",X"79",X"00",X"00",X"77",X"22",X"00",X"00",X"99",X"77",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"9D",X"92",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"77",
		X"00",X"00",X"29",X"69",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"79",X"00",X"00",X"66",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"39",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"DD",X"00",X"00",X"90",X"9D",X"00",X"00",X"07",X"D2",
		X"00",X"00",X"09",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"29",X"00",X"00",X"62",X"92",
		X"00",X"00",X"26",X"29",X"00",X"00",X"22",X"26",X"00",X"00",X"92",X"97",X"00",X"00",X"99",X"69",
		X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E2",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"77",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"72",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"07",X"9D",X"00",X"00",X"02",X"DD",X"00",X"00",X"02",X"9D",
		X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"9E",X"99",X"90",
		X"00",X"9E",X"99",X"EE",X"00",X"23",X"99",X"EE",X"00",X"26",X"99",X"33",X"00",X"22",X"9D",X"20",
		X"00",X"26",X"DD",X"20",X"00",X"22",X"9D",X"90",X"00",X"76",X"DD",X"79",X"00",X"72",X"9D",X"99",
		X"00",X"76",X"DD",X"99",X"00",X"72",X"2D",X"99",X"00",X"76",X"29",X"99",X"00",X"72",X"99",X"99",
		X"00",X"72",X"77",X"99",X"00",X"22",X"62",X"79",X"00",X"22",X"99",X"70",X"00",X"29",X"99",X"70",
		X"00",X"72",X"99",X"70",X"00",X"97",X"77",X"70",X"00",X"29",X"66",X"70",X"00",X"26",X"66",X"70",
		X"00",X"22",X"66",X"70",X"00",X"22",X"66",X"70",X"00",X"29",X"66",X"70",X"00",X"29",X"66",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"77",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"79",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"79",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"99",
		X"00",X"00",X"26",X"79",X"00",X"00",X"77",X"22",X"00",X"00",X"99",X"77",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"69",X"70",X"00",X"00",
		X"29",X"29",X"00",X"00",X"62",X"22",X"00",X"00",X"66",X"72",X"90",X"00",X"66",X"62",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"66",X"00",X"66",X"99",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"9D",X"92",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"77",
		X"00",X"00",X"29",X"69",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"79",X"00",X"00",X"66",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"DD",X"00",X"00",X"90",X"9D",X"00",X"00",X"07",X"D2",
		X"00",X"00",X"09",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"29",X"00",X"00",X"62",X"92",
		X"00",X"00",X"26",X"29",X"00",X"00",X"22",X"26",X"00",X"00",X"92",X"97",X"00",X"00",X"99",X"69",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"E2",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"77",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"72",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"0E",X"99",X"00",X"00",X"0E",X"9D",X"00",X"00",X"0E",X"DD",X"00",X"00",X"02",X"9D",
		X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"09",X"00",X"00",X"EE",X"99",X"EE",
		X"00",X"99",X"99",X"3E",X"00",X"26",X"99",X"33",X"00",X"26",X"99",X"23",X"00",X"22",X"9D",X"20",
		X"00",X"26",X"DD",X"20",X"00",X"22",X"9D",X"90",X"00",X"76",X"DD",X"70",X"00",X"72",X"9D",X"90",
		X"00",X"76",X"DD",X"90",X"00",X"72",X"2D",X"90",X"00",X"76",X"29",X"90",X"00",X"72",X"99",X"90",
		X"00",X"72",X"77",X"90",X"00",X"22",X"62",X"70",X"00",X"22",X"99",X"70",X"00",X"29",X"99",X"70",
		X"00",X"72",X"99",X"70",X"00",X"97",X"77",X"70",X"00",X"29",X"66",X"70",X"00",X"26",X"66",X"70",
		X"00",X"22",X"66",X"70",X"00",X"22",X"66",X"70",X"00",X"29",X"66",X"70",X"00",X"29",X"66",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"77",X"00",X"22",X"77",X"77",X"00",X"96",X"22",X"90",X"00",
		X"99",X"22",X"22",X"00",X"22",X"72",X"22",X"00",X"66",X"72",X"22",X"00",X"66",X"92",X"22",X"00",
		X"66",X"92",X"27",X"00",X"66",X"92",X"27",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",
		X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",X"66",X"92",X"97",X"00",
		X"66",X"92",X"97",X"00",X"66",X"72",X"97",X"00",X"22",X"72",X"99",X"00",X"99",X"22",X"99",X"00",
		X"96",X"22",X"96",X"00",X"22",X"77",X"67",X"00",X"99",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"22",X"00",X"66",X"97",X"29",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",
		X"66",X"72",X"97",X"00",X"22",X"22",X"97",X"00",X"92",X"22",X"70",X"00",X"99",X"29",X"70",X"00",
		X"99",X"29",X"70",X"00",X"22",X"92",X"00",X"00",X"72",X"92",X"00",X"00",X"09",X"99",X"90",X"00",
		X"00",X"29",X"99",X"00",X"00",X"69",X"09",X"00",X"00",X"76",X"90",X"00",X"00",X"06",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"77",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"79",
		X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"92",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"92",X"90",X"00",
		X"66",X"22",X"99",X"00",X"62",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"99",X"29",X"99",X"00",
		X"99",X"29",X"29",X"00",X"99",X"92",X"00",X"00",X"79",X"66",X"99",X"00",X"79",X"62",X"09",X"00",
		X"22",X"22",X"09",X"00",X"22",X"99",X"09",X"00",X"97",X"99",X"99",X"00",X"97",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"27",X"00",X"00",X"66",X"67",X"00",X"00",X"66",X"67",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"27",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"72",X"00",X"00",X"99",X"29",X"00",X"00",X"92",X"29",X"00",X"00",
		X"22",X"22",X"00",X"00",X"79",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"67",X"99",X"00",X"00",X"06",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"29",X"66",X"70",X"00",X"69",X"66",X"70",X"00",X"69",X"66",X"70",X"00",X"69",X"66",X"70",
		X"00",X"69",X"66",X"70",X"00",X"69",X"22",X"70",X"00",X"79",X"99",X"70",X"00",X"72",X"99",X"70",
		X"00",X"72",X"99",X"70",X"00",X"72",X"99",X"70",X"00",X"77",X"99",X"99",X"00",X"76",X"77",X"99",
		X"00",X"76",X"22",X"99",X"00",X"76",X"22",X"99",X"00",X"76",X"97",X"99",X"00",X"76",X"22",X"99",
		X"00",X"66",X"22",X"99",X"00",X"69",X"22",X"99",X"00",X"69",X"22",X"79",X"00",X"69",X"99",X"79",
		X"00",X"69",X"99",X"20",X"00",X"76",X"99",X"90",X"00",X"76",X"77",X"00",X"00",X"96",X"90",X"00",
		X"00",X"96",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"00",X"11",X"00",X"00",X"00",X"01",X"10",X"21",X"00",X"00",X"11",X"10",X"00",X"00",X"22",X"11",
		X"00",X"00",X"11",X"F0",X"00",X"99",X"12",X"90",X"00",X"99",X"12",X"90",X"00",X"00",X"99",X"11",
		X"00",X"00",X"10",X"01",X"00",X"00",X"10",X"21",X"00",X"00",X"11",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"99",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"10",
		X"00",X"00",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"22",X"00",X"00",X"10",X"0F",X"00",X"00",X"11",X"F0",X"01",X"00",X"20",X"01",X"10",
		X"00",X"20",X"00",X"11",X"00",X"2F",X"00",X"10",X"00",X"90",X"00",X"10",X"00",X"09",X"00",X"10",
		X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"99",X"00",X"00",X"01",X"90",X"00",X"11",X"01",X"00",
		X"00",X"11",X"02",X"00",X"00",X"10",X"22",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"11",X"00",
		X"00",X"09",X"00",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",
		X"00",X"09",X"91",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"29",X"99",
		X"00",X"00",X"10",X"99",X"00",X"00",X"10",X"99",X"00",X"00",X"02",X"99",X"00",X"90",X"01",X"99",
		X"00",X"90",X"01",X"99",X"00",X"09",X"00",X"99",X"00",X"11",X"09",X"99",X"00",X"01",X"00",X"99",
		X"00",X"11",X"00",X"99",X"09",X"10",X"99",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"90",X"00",X"00",
		X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"10",X"00",X"01",X"00",X"11",X"11",X"00",X"90",X"01",X"10",X"00",X"00",X"0F",X"01",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"09",X"00",X"01",X"00",X"09",X"00",X"01",X"00",
		X"99",X"00",X"10",X"00",X"90",X"09",X"91",X"00",X"99",X"00",X"10",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"11",X"99",X"99",X"11",X"11",X"99",X"99",X"10",X"01",X"99",X"99",X"00",X"99",
		X"90",X"00",X"00",X"99",X"09",X"00",X"01",X"99",X"99",X"09",X"11",X"09",X"00",X"09",X"10",X"99",
		X"00",X"11",X"00",X"00",X"91",X"10",X"10",X"00",X"09",X"01",X"99",X"00",X"99",X"09",X"01",X"00",
		X"00",X"10",X"01",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"11",X"00",X"00",X"11",X"01",X"01",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"09",X"00",
		X"99",X"99",X"99",X"00",X"09",X"99",X"11",X"10",X"00",X"99",X"21",X"10",X"00",X"99",X"11",X"00",
		X"00",X"99",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"09",X"91",X"00",X"00",X"00",X"91",X"11",
		X"00",X"11",X"11",X"01",X"00",X"10",X"10",X"91",X"00",X"00",X"11",X"01",X"00",X"11",X"10",X"00",
		X"00",X"11",X"09",X"01",X"00",X"01",X"09",X"11",X"00",X"01",X"10",X"10",X"00",X"11",X"99",X"10",
		X"00",X"19",X"99",X"00",X"00",X"99",X"09",X"09",X"00",X"99",X"90",X"99",X"00",X"99",X"90",X"99",
		X"00",X"09",X"11",X"00",X"00",X"99",X"19",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"01",
		X"00",X"91",X"01",X"00",X"00",X"99",X"10",X"00",X"09",X"00",X"01",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"01",X"00",X"00",X"10",X"00",X"00",X"99",X"00",X"11",X"01",X"00",X"F0",X"00",
		X"01",X"01",X"00",X"99",X"10",X"11",X"00",X"99",X"00",X"01",X"00",X"09",X"99",X"11",X"11",X"00",
		X"99",X"01",X"11",X"00",X"90",X"10",X"11",X"00",X"00",X"11",X"01",X"00",X"90",X"00",X"90",X"00",
		X"00",X"91",X"90",X"00",X"00",X"00",X"99",X"00",X"10",X"00",X"09",X"00",X"09",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"01",X"90",X"00",
		X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",
		X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",
		X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",X"01",X"11",X"90",X"00",
		X"01",X"11",X"90",X"00",X"01",X"19",X"90",X"00",X"01",X"19",X"90",X"00",X"01",X"90",X"90",X"00",
		X"01",X"00",X"90",X"00",X"01",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"09",X"00",X"01",X"11",X"99",
		X"00",X"14",X"14",X"90",X"00",X"91",X"41",X"90",X"00",X"09",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"99",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"F1",X"00",
		X"00",X"00",X"12",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"F1",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F9",X"00",X"00",X"99",X"99",X"09",
		X"00",X"9F",X"0F",X"F0",X"00",X"F9",X"0F",X"F0",X"00",X"09",X"FF",X"F0",X"00",X"F9",X"99",X"99",
		X"00",X"F9",X"90",X"99",X"00",X"F0",X"09",X"99",X"00",X"9F",X"00",X"FF",X"00",X"FF",X"F0",X"FF",
		X"00",X"90",X"FF",X"99",X"00",X"99",X"FF",X"99",X"00",X"99",X"F9",X"F9",X"00",X"9F",X"F9",X"0F",
		X"00",X"FF",X"09",X"FF",X"00",X"F0",X"90",X"F0",X"00",X"FF",X"99",X"F0",X"00",X"FF",X"F9",X"0F",
		X"00",X"FF",X"99",X"00",X"00",X"99",X"99",X"FF",X"00",X"99",X"00",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"F0",X"00",X"00",X"F9",X"09",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"9F",X"F9",X"00",
		X"00",X"F0",X"99",X"00",X"00",X"0F",X"0F",X"00",X"00",X"FF",X"99",X"00",X"00",X"9F",X"F9",X"00",
		X"00",X"99",X"9F",X"00",X"00",X"9F",X"9F",X"00",X"00",X"FF",X"F0",X"00",X"00",X"FF",X"0F",X"00",
		X"00",X"9F",X"F0",X"00",X"00",X"9F",X"FF",X"00",X"00",X"90",X"99",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"00",X"90",
		X"00",X"F9",X"F0",X"09",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"0F",X"00",X"09",X"00",X"9F",
		X"00",X"00",X"00",X"9F",X"00",X"00",X"90",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"0F",X"00",X"00",X"90",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"09",X"09",X"F0",X"00",X"90",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"09",X"AD",
		X"00",X"00",X"9A",X"99",X"00",X"00",X"AB",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"90",X"00",
		X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AD",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"A9",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"62",X"22",
		X"00",X"00",X"26",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"29",
		X"00",X"00",X"77",X"29",X"00",X"00",X"66",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"77",X"29",
		X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"99",X"00",X"00",X"26",X"29",
		X"00",X"00",X"62",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"90",X"00",X"99",X"99",X"90",X"00",X"22",X"99",X"99",X"00",X"99",X"22",X"29",X"00",
		X"99",X"22",X"29",X"00",X"99",X"27",X"79",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"76",X"00",
		X"66",X"99",X"76",X"00",X"66",X"99",X"76",X"00",X"66",X"99",X"76",X"00",X"66",X"99",X"96",X"00",
		X"66",X"99",X"96",X"00",X"66",X"99",X"76",X"00",X"66",X"99",X"76",X"00",X"66",X"99",X"76",X"00",
		X"66",X"99",X"76",X"00",X"66",X"99",X"99",X"00",X"99",X"27",X"79",X"00",X"99",X"22",X"29",X"00",
		X"99",X"22",X"29",X"00",X"22",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"00",X"09",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"22",X"66",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"92",
		X"00",X"09",X"22",X"29",X"00",X"09",X"26",X"29",X"00",X"00",X"72",X"69",X"00",X"00",X"27",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"99",X"00",X"00",X"26",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"79",X"99",X"00",X"00",X"67",X"29",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"99",X"00",X"00",X"66",X"22",X"90",X"00",X"66",X"97",X"99",X"00",X"66",X"99",X"99",X"00",
		X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"09",X"99",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"22",X"00",X"66",X"99",X"92",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"69",X"00",
		X"66",X"99",X"29",X"00",X"66",X"99",X"96",X"00",X"99",X"97",X"96",X"00",X"99",X"72",X"69",X"00",
		X"99",X"22",X"60",X"00",X"29",X"29",X"90",X"00",X"92",X"92",X"90",X"00",X"99",X"99",X"00",X"00",
		X"00",X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",
		X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"26",X"00",X"00",X"92",X"26",X"00",X"00",X"92",X"22",
		X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"77",X"00",X"00",X"92",X"27",
		X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",
		X"00",X"00",X"22",X"96",X"00",X"00",X"66",X"96",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"90",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"99",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"99",X"00",X"00",
		X"66",X"99",X"90",X"00",X"66",X"99",X"90",X"00",X"66",X"99",X"99",X"00",X"69",X"92",X"29",X"00",
		X"29",X"92",X"27",X"00",X"29",X"22",X"20",X"00",X"92",X"29",X"29",X"00",X"92",X"92",X"79",X"00",
		X"92",X"22",X"90",X"00",X"22",X"22",X"90",X"00",X"92",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"29",X"99",X"00",X"09",X"66",X"99",X"00",X"00",X"96",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"09",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"9E",X"22",
		X"00",X"00",X"EE",X"22",X"00",X"00",X"99",X"62",X"00",X"00",X"99",X"62",X"00",X"00",X"92",X"76",
		X"00",X"00",X"99",X"77",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"97",X"00",X"00",X"09",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"79",X"92",X"00",X"00",
		X"79",X"27",X"00",X"00",X"99",X"27",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"69",X"00",X"00",X"22",X"62",X"00",X"00",X"29",X"26",X"00",X"00",
		X"92",X"26",X"00",X"00",X"26",X"29",X"00",X"00",X"26",X"99",X"00",X"00",X"92",X"66",X"00",X"00",
		X"92",X"77",X"00",X"00",X"29",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"77",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"29",X"99",
		X"00",X"EE",X"22",X"E9",X"00",X"EE",X"22",X"E9",X"00",X"39",X"22",X"99",X"00",X"79",X"22",X"90",
		X"00",X"72",X"22",X"90",X"00",X"26",X"26",X"90",X"00",X"26",X"26",X"90",X"00",X"26",X"26",X"90",
		X"00",X"76",X"26",X"79",X"00",X"96",X"26",X"99",X"00",X"76",X"26",X"99",X"00",X"76",X"22",X"99",
		X"00",X"76",X"99",X"99",X"00",X"76",X"66",X"99",X"00",X"76",X"99",X"99",X"00",X"72",X"99",X"99",
		X"00",X"77",X"99",X"99",X"00",X"27",X"99",X"70",X"00",X"27",X"99",X"70",X"00",X"29",X"66",X"90",
		X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",
		X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",
		X"00",X"27",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"99",X"90",X"00",X"29",X"99",X"70",
		X"00",X"29",X"99",X"70",X"00",X"29",X"99",X"70",X"00",X"79",X"99",X"70",X"00",X"72",X"99",X"79",
		X"00",X"72",X"99",X"79",X"00",X"72",X"22",X"79",X"00",X"72",X"99",X"79",X"00",X"72",X"22",X"79",
		X"00",X"72",X"22",X"79",X"00",X"72",X"22",X"79",X"00",X"72",X"22",X"99",X"00",X"72",X"92",X"99",
		X"00",X"72",X"99",X"90",X"00",X"09",X"66",X"00",X"00",X"00",X"77",X"90",X"00",X"99",X"77",X"90",
		X"00",X"99",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"50",
		X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"BB",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"BB",X"00",X"00",X"09",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"0B",X"05",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"05",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"90",X"00",X"99",X"99",X"90",X"00",X"22",X"99",X"99",X"00",X"99",X"29",X"29",X"00",
		X"99",X"22",X"29",X"00",X"99",X"27",X"29",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"99",X"27",X"79",X"00",X"99",X"22",X"29",X"00",
		X"22",X"29",X"29",X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"90",X"00",X"00",X"09",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"79",X"99",X"00",X"00",X"67",X"29",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"99",X"00",X"00",X"66",X"22",X"90",X"00",X"66",X"97",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"22",X"00",X"66",X"99",X"92",X"00",X"66",X"99",X"29",X"00",X"66",X"99",X"22",X"00",
		X"66",X"99",X"22",X"00",X"66",X"99",X"77",X"00",X"99",X"97",X"79",X"00",X"99",X"72",X"99",X"00",
		X"22",X"22",X"99",X"00",X"92",X"29",X"99",X"00",X"99",X"92",X"99",X"00",X"99",X"92",X"99",X"00",
		X"00",X"29",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"99",X"00",X"00",
		X"66",X"99",X"90",X"00",X"66",X"99",X"90",X"00",X"66",X"99",X"99",X"00",X"69",X"92",X"29",X"00",
		X"29",X"92",X"27",X"00",X"29",X"22",X"20",X"00",X"92",X"29",X"29",X"00",X"92",X"92",X"79",X"00",
		X"92",X"22",X"90",X"00",X"99",X"27",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"79",X"99",X"00",
		X"99",X"79",X"99",X"00",X"09",X"79",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"79",X"92",X"00",X"00",
		X"79",X"27",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",
		X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"97",X"00",X"00",
		X"22",X"79",X"00",X"00",X"29",X"99",X"00",X"00",X"27",X"99",X"00",X"00",X"27",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"92",X"66",X"90",
		X"00",X"92",X"66",X"90",X"00",X"92",X"66",X"90",X"00",X"92",X"99",X"90",X"00",X"92",X"99",X"70",
		X"00",X"99",X"99",X"70",X"00",X"99",X"99",X"70",X"00",X"99",X"99",X"70",X"00",X"72",X"99",X"79",
		X"00",X"72",X"99",X"79",X"00",X"92",X"22",X"79",X"00",X"72",X"99",X"79",X"00",X"22",X"22",X"79",
		X"00",X"27",X"22",X"79",X"00",X"27",X"22",X"79",X"00",X"77",X"72",X"99",X"00",X"77",X"77",X"99",
		X"00",X"77",X"77",X"90",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"69",X"92",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"29",
		X"00",X"00",X"77",X"29",X"00",X"00",X"66",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"77",X"29",
		X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"66",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"92",
		X"00",X"00",X"22",X"29",X"00",X"00",X"26",X"29",X"00",X"00",X"72",X"69",X"00",X"00",X"27",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",
		X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"26",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"29",
		X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"77",X"00",X"00",X"92",X"27",
		X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"26",X"00",X"00",X"09",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"9E",X"22",
		X"00",X"00",X"3E",X"22",X"00",X"00",X"EE",X"62",X"00",X"00",X"9E",X"62",X"00",X"00",X"99",X"76",
		X"00",X"00",X"99",X"77",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"92",
		X"00",X"00",X"09",X"92",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"29",X"99",
		X"00",X"99",X"22",X"99",X"00",X"9E",X"22",X"99",X"00",X"EE",X"22",X"99",X"00",X"EE",X"22",X"90",
		X"00",X"33",X"22",X"90",X"00",X"99",X"26",X"90",X"00",X"99",X"26",X"90",X"00",X"99",X"26",X"90",
		X"00",X"99",X"26",X"99",X"00",X"99",X"26",X"99",X"00",X"79",X"26",X"99",X"00",X"79",X"22",X"99",
		X"00",X"76",X"99",X"99",X"00",X"76",X"66",X"99",X"00",X"76",X"99",X"99",X"00",X"72",X"99",X"99",
		X"00",X"77",X"99",X"99",X"00",X"27",X"99",X"70",X"00",X"27",X"99",X"70",X"00",X"29",X"66",X"90",
		X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"69",X"92",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"29",
		X"00",X"00",X"77",X"29",X"00",X"00",X"66",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"77",X"29",
		X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"79",X"99",X"00",X"00",X"67",X"29",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"99",X"90",X"00",X"66",X"22",X"99",X"00",X"66",X"97",X"99",X"00",X"66",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"90",
		X"00",X"00",X"E9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"66",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"92",
		X"00",X"00",X"22",X"29",X"00",X"00",X"26",X"29",X"00",X"00",X"72",X"69",X"00",X"00",X"27",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",
		X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"26",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"29",
		X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"77",X"00",X"00",X"92",X"27",
		X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"26",X"00",X"00",X"09",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"9E",X"22",
		X"00",X"00",X"9E",X"22",X"00",X"00",X"0E",X"62",X"00",X"00",X"9E",X"62",X"00",X"00",X"99",X"76",
		X"00",X"00",X"99",X"77",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"92",
		X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"29",X"99",
		X"00",X"99",X"22",X"99",X"00",X"9E",X"22",X"99",X"00",X"EE",X"22",X"99",X"00",X"EE",X"22",X"90",
		X"00",X"E9",X"22",X"90",X"00",X"99",X"26",X"90",X"00",X"99",X"26",X"90",X"00",X"99",X"26",X"90",
		X"00",X"99",X"26",X"90",X"00",X"99",X"26",X"90",X"00",X"79",X"26",X"90",X"00",X"79",X"22",X"90",
		X"00",X"76",X"99",X"90",X"00",X"76",X"66",X"90",X"00",X"76",X"99",X"90",X"00",X"72",X"99",X"90",
		X"00",X"77",X"99",X"90",X"00",X"27",X"99",X"70",X"00",X"27",X"99",X"70",X"00",X"29",X"66",X"90",
		X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",
		X"00",X"09",X"90",X"00",X"99",X"99",X"90",X"00",X"22",X"99",X"99",X"00",X"99",X"29",X"29",X"00",
		X"99",X"22",X"29",X"00",X"99",X"27",X"29",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"99",X"27",X"79",X"00",X"99",X"22",X"29",X"00",
		X"22",X"29",X"29",X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"22",X"00",X"66",X"99",X"92",X"00",X"66",X"99",X"29",X"00",X"66",X"99",X"22",X"00",
		X"66",X"99",X"22",X"00",X"96",X"99",X"77",X"00",X"99",X"97",X"79",X"00",X"99",X"72",X"99",X"00",
		X"22",X"22",X"99",X"00",X"92",X"29",X"99",X"00",X"99",X"92",X"99",X"00",X"99",X"92",X"99",X"00",
		X"00",X"29",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"99",
		X"00",X"00",X"09",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"99",X"90",X"00",
		X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"99",X"99",X"00",X"69",X"92",X"29",X"00",
		X"29",X"92",X"27",X"00",X"29",X"22",X"20",X"00",X"92",X"29",X"29",X"00",X"92",X"92",X"79",X"00",
		X"92",X"22",X"90",X"00",X"99",X"27",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"79",X"99",X"00",
		X"09",X"79",X"99",X"00",X"00",X"79",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"92",X"00",X"00",X"79",X"92",X"00",X"00",
		X"79",X"27",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",
		X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"97",X"00",X"00",
		X"22",X"79",X"00",X"00",X"29",X"99",X"00",X"00",X"27",X"99",X"00",X"00",X"27",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"29",X"66",X"90",X"00",X"92",X"66",X"90",
		X"00",X"92",X"66",X"90",X"00",X"92",X"66",X"90",X"00",X"92",X"99",X"90",X"00",X"92",X"99",X"70",
		X"00",X"99",X"99",X"70",X"00",X"99",X"99",X"70",X"00",X"99",X"99",X"70",X"00",X"72",X"99",X"79",
		X"00",X"72",X"99",X"79",X"00",X"92",X"22",X"79",X"00",X"72",X"99",X"79",X"00",X"22",X"22",X"79",
		X"00",X"27",X"22",X"79",X"00",X"27",X"22",X"79",X"00",X"77",X"72",X"99",X"00",X"77",X"77",X"99",
		X"00",X"77",X"77",X"90",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"02",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",
		X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",
		X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",X"02",X"22",X"90",X"00",
		X"02",X"22",X"90",X"00",X"02",X"29",X"90",X"00",X"02",X"29",X"90",X"00",X"02",X"90",X"90",X"00",
		X"02",X"00",X"90",X"00",X"02",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"09",X"00",X"02",X"22",X"99",
		X"00",X"26",X"26",X"90",X"00",X"92",X"62",X"90",X"00",X"09",X"22",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"99",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"90",X"00",X"00",X"45",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"41",
		X"00",X"00",X"54",X"44",X"00",X"00",X"54",X"99",X"00",X"00",X"15",X"11",X"00",X"00",X"55",X"41",
		X"00",X"00",X"55",X"14",X"00",X"00",X"55",X"44",X"00",X"00",X"94",X"44",X"00",X"00",X"51",X"44",
		X"00",X"00",X"59",X"94",X"00",X"00",X"51",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"51",X"44",
		X"00",X"00",X"55",X"14",X"00",X"00",X"55",X"14",X"00",X"00",X"59",X"55",X"00",X"00",X"94",X"99",
		X"00",X"00",X"91",X"11",X"00",X"00",X"95",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"99",X"99",X"99",X"00",X"55",X"55",X"11",X"00",X"55",X"51",X"55",X"00",
		X"99",X"99",X"49",X"00",X"59",X"99",X"51",X"00",X"55",X"59",X"91",X"00",X"14",X"11",X"49",X"00",
		X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",
		X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",
		X"44",X"44",X"49",X"00",X"44",X"44",X"49",X"00",X"99",X"99",X"91",X"00",X"99",X"99",X"51",X"00",
		X"59",X"99",X"55",X"00",X"59",X"55",X"51",X"00",X"99",X"99",X"99",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"15",
		X"00",X"00",X"99",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"94",X"91",X"00",X"00",X"54",X"55",
		X"00",X"00",X"15",X"44",X"00",X"00",X"45",X"44",X"00",X"00",X"55",X"14",X"00",X"00",X"55",X"41",
		X"00",X"00",X"91",X"44",X"00",X"00",X"54",X"94",X"00",X"00",X"54",X"94",X"00",X"00",X"55",X"45",
		X"00",X"00",X"95",X"49",X"00",X"00",X"49",X"49",X"00",X"00",X"14",X"19",X"00",X"00",X"11",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"19",X"90",X"00",X"00",X"15",X"59",X"00",X"00",
		X"45",X"51",X"00",X"00",X"44",X"51",X"90",X"00",X"44",X"15",X"99",X"00",X"44",X"99",X"55",X"00",
		X"44",X"15",X"11",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"15",X"00",
		X"00",X"00",X"55",X"59",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"51",X"00",X"00",X"00",X"45",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"59",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",
		X"54",X"44",X"99",X"00",X"59",X"44",X"99",X"00",X"99",X"44",X"55",X"00",X"19",X"44",X"94",X"00",
		X"91",X"54",X"91",X"00",X"91",X"95",X"55",X"00",X"09",X"99",X"59",X"00",X"00",X"59",X"19",X"00",
		X"00",X"55",X"59",X"00",X"00",X"51",X"59",X"00",X"00",X"59",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"35",X"00",X"00",X"00",X"31",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"09",X"15",
		X"00",X"00",X"99",X"11",X"00",X"00",X"94",X"41",X"00",X"00",X"51",X"44",X"00",X"00",X"49",X"44",
		X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"44",X"00",X"00",X"55",X"54",X"00",X"00",X"45",X"95",
		X"00",X"00",X"45",X"51",X"00",X"00",X"44",X"49",X"00",X"00",X"14",X"99",X"00",X"00",X"51",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"45",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"19",X"00",X"00",
		X"44",X"45",X"90",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"45",X"00",
		X"14",X"44",X"44",X"00",X"54",X"44",X"55",X"00",X"95",X"44",X"55",X"00",X"99",X"44",X"59",X"00",
		X"99",X"44",X"90",X"00",X"59",X"44",X"90",X"00",X"55",X"49",X"90",X"00",X"15",X"99",X"00",X"00",
		X"91",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"09",X"95",X"00",X"00",X"09",X"91",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"95",X"00",X"00",X"09",X"54",X"00",X"00",X"09",X"49",
		X"00",X"00",X"09",X"45",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"51",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"41",X"99",X"00",X"00",
		X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"51",X"00",X"00",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"91",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"11",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"41",X"00",X"00",
		X"14",X"44",X"00",X"00",X"54",X"44",X"00",X"00",X"91",X"99",X"00",X"00",X"54",X"99",X"90",X"00",
		X"95",X"99",X"90",X"00",X"94",X"09",X"90",X"00",X"49",X"59",X"90",X"00",X"19",X"54",X"00",X"00",
		X"99",X"59",X"00",X"00",X"49",X"99",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"EE",X"11",X"59",X"00",X"EE",X"99",X"59",
		X"00",X"33",X"55",X"59",X"00",X"14",X"15",X"90",X"00",X"14",X"99",X"00",X"00",X"14",X"11",X"90",
		X"00",X"14",X"11",X"90",X"00",X"41",X"14",X"90",X"00",X"45",X"41",X"90",X"00",X"15",X"11",X"90",
		X"00",X"45",X"14",X"90",X"00",X"45",X"11",X"90",X"00",X"45",X"11",X"90",X"00",X"45",X"99",X"50",
		X"00",X"49",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"15",X"99",X"00",X"00",X"59",X"99",X"00",
		X"00",X"15",X"11",X"00",X"00",X"55",X"44",X"00",X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"15",X"44",X"00",X"00",X"14",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"19",X"44",X"90",X"00",X"59",X"44",X"90",
		X"00",X"19",X"44",X"90",X"00",X"59",X"44",X"90",X"00",X"19",X"44",X"90",X"00",X"59",X"44",X"90",
		X"00",X"19",X"44",X"90",X"00",X"59",X"11",X"90",X"00",X"19",X"99",X"90",X"00",X"51",X"99",X"00",
		X"00",X"19",X"55",X"00",X"00",X"55",X"15",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"55",X"90",
		X"00",X"59",X"99",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"09",X"90",X"99",X"00",X"99",X"00",X"39",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"39",X"00",
		X"99",X"00",X"99",X"00",X"99",X"00",X"39",X"00",X"99",X"00",X"39",X"00",X"99",X"00",X"93",X"00",
		X"99",X"90",X"99",X"00",X"09",X"99",X"39",X"00",X"09",X"99",X"99",X"00",X"09",X"39",X"99",X"00",
		X"00",X"93",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"50",
		X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"50",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"50",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"93",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"9A",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"50",
		X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"50",
		X"00",X"90",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"99",X"99",X"99",X"00",X"55",X"55",X"11",X"00",X"15",X"51",X"55",X"00",
		X"99",X"99",X"49",X"00",X"59",X"99",X"59",X"00",X"55",X"59",X"99",X"00",X"14",X"11",X"99",X"00",
		X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"91",X"00",X"99",X"99",X"95",X"00",X"99",X"99",X"99",X"00",
		X"59",X"99",X"99",X"00",X"51",X"51",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"19",X"90",X"00",X"00",X"15",X"59",X"00",X"00",
		X"45",X"51",X"90",X"00",X"44",X"51",X"99",X"00",X"44",X"15",X"99",X"00",X"44",X"99",X"55",X"00",
		X"44",X"15",X"11",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"45",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"49",X"99",X"00",
		X"54",X"54",X"99",X"00",X"59",X"45",X"99",X"00",X"99",X"54",X"55",X"00",X"19",X"45",X"94",X"00",
		X"91",X"54",X"91",X"00",X"91",X"95",X"55",X"00",X"09",X"99",X"59",X"00",X"00",X"59",X"19",X"00",
		X"00",X"55",X"59",X"00",X"00",X"51",X"59",X"00",X"00",X"59",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"90",X"00",X"44",X"19",X"90",X"00",
		X"44",X"45",X"90",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"59",X"00",X"44",X"55",X"45",X"00",
		X"14",X"99",X"44",X"00",X"54",X"99",X"55",X"00",X"95",X"99",X"55",X"00",X"99",X"99",X"59",X"00",
		X"99",X"99",X"90",X"00",X"59",X"99",X"90",X"00",X"55",X"99",X"90",X"00",X"15",X"95",X"00",X"00",
		X"91",X"55",X"00",X"00",X"95",X"99",X"00",X"00",X"09",X"95",X"00",X"00",X"09",X"91",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"91",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"11",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"91",X"00",X"00",
		X"11",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"91",X"99",X"00",X"00",X"55",X"55",X"90",X"00",
		X"49",X"95",X"90",X"00",X"49",X"99",X"90",X"00",X"49",X"59",X"90",X"00",X"15",X"54",X"00",X"00",
		X"95",X"59",X"00",X"00",X"49",X"99",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"15",X"44",X"00",X"00",X"14",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"19",X"44",X"99",X"00",X"59",X"54",X"99",
		X"00",X"19",X"55",X"99",X"00",X"59",X"99",X"99",X"00",X"19",X"59",X"99",X"00",X"59",X"99",X"99",
		X"00",X"11",X"99",X"99",X"00",X"54",X"99",X"99",X"00",X"11",X"99",X"99",X"00",X"55",X"95",X"00",
		X"00",X"15",X"99",X"00",X"00",X"55",X"55",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"55",X"90",
		X"00",X"59",X"99",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"45",X"99",X"00",X"00",X"E5",X"11",X"00",X"00",X"E3",X"41",
		X"00",X"00",X"E3",X"44",X"00",X"00",X"53",X"55",X"00",X"00",X"15",X"55",X"00",X"00",X"55",X"51",
		X"00",X"00",X"55",X"54",X"00",X"00",X"59",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"59",X"54",
		X"00",X"00",X"59",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"59",X"54",
		X"00",X"00",X"99",X"54",X"00",X"00",X"55",X"54",X"00",X"00",X"E5",X"55",X"00",X"00",X"E3",X"99",
		X"00",X"00",X"E3",X"11",X"00",X"00",X"93",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"15",
		X"00",X"00",X"99",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"94",X"51",X"00",X"00",X"54",X"55",
		X"00",X"00",X"1D",X"99",X"00",X"00",X"4D",X"99",X"00",X"00",X"DD",X"D9",X"00",X"00",X"D5",X"D5",
		X"00",X"00",X"D9",X"91",X"00",X"00",X"59",X"91",X"00",X"00",X"59",X"51",X"00",X"00",X"35",X"15",
		X"00",X"00",X"35",X"19",X"00",X"00",X"49",X"19",X"00",X"00",X"14",X"19",X"00",X"00",X"11",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"31",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"09",X"55",
		X"00",X"00",X"99",X"95",X"00",X"00",X"94",X"99",X"00",X"00",X"5D",X"D9",X"00",X"00",X"49",X"DD",
		X"00",X"00",X"95",X"9D",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"59",X"00",X"00",X"45",X"95",
		X"00",X"00",X"45",X"51",X"00",X"00",X"44",X"19",X"00",X"00",X"14",X"99",X"00",X"00",X"51",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"41",X"99",X"00",X"00",
		X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"51",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"1D",X"00",X"00",X"00",X"DD",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"9D",
		X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"EE",X"1D",X"00",X"00",X"EE",X"DD",X"59",
		X"00",X"33",X"99",X"39",X"00",X"14",X"9D",X"90",X"00",X"14",X"DD",X"00",X"00",X"14",X"9D",X"99",
		X"00",X"14",X"9D",X"99",X"00",X"41",X"DD",X"99",X"00",X"45",X"DD",X"99",X"00",X"15",X"9D",X"99",
		X"00",X"45",X"99",X"99",X"00",X"45",X"99",X"99",X"00",X"45",X"11",X"99",X"00",X"41",X"99",X"90",
		X"00",X"49",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"15",X"99",X"00",X"00",X"59",X"99",X"00",
		X"00",X"15",X"11",X"00",X"00",X"55",X"44",X"00",X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"35",X"99",X"00",X"00",X"35",X"11",X"00",X"00",X"35",X"41",
		X"00",X"00",X"34",X"44",X"00",X"00",X"34",X"55",X"00",X"00",X"15",X"55",X"00",X"00",X"55",X"51",
		X"00",X"00",X"55",X"54",X"00",X"00",X"59",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"59",X"54",
		X"00",X"00",X"59",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"59",X"54",
		X"00",X"00",X"99",X"54",X"00",X"00",X"35",X"54",X"00",X"00",X"35",X"55",X"00",X"00",X"34",X"99",
		X"00",X"00",X"91",X"11",X"00",X"00",X"95",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"19",X"90",X"00",X"00",X"15",X"59",X"00",X"00",
		X"45",X"51",X"00",X"00",X"44",X"51",X"90",X"00",X"44",X"15",X"99",X"00",X"44",X"99",X"55",X"00",
		X"44",X"15",X"11",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"45",X"00",X"44",X"44",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"15",
		X"00",X"00",X"99",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"94",X"51",X"00",X"00",X"54",X"55",
		X"00",X"00",X"1D",X"99",X"00",X"00",X"4D",X"99",X"00",X"00",X"DD",X"D9",X"00",X"00",X"D5",X"D5",
		X"00",X"00",X"D9",X"91",X"00",X"00",X"59",X"91",X"00",X"00",X"59",X"51",X"00",X"00",X"35",X"15",
		X"00",X"00",X"35",X"19",X"00",X"00",X"49",X"19",X"00",X"00",X"14",X"19",X"00",X"00",X"11",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"31",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"09",X"55",
		X"00",X"00",X"99",X"95",X"00",X"00",X"94",X"99",X"00",X"00",X"5D",X"D9",X"00",X"00",X"49",X"DD",
		X"00",X"00",X"95",X"9D",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"59",X"00",X"00",X"45",X"95",
		X"00",X"00",X"45",X"51",X"00",X"00",X"44",X"19",X"00",X"00",X"14",X"99",X"00",X"00",X"51",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"41",X"99",X"00",X"00",
		X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"51",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"1D",X"00",X"00",X"00",X"DD",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"9D",
		X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"EE",X"1D",X"00",X"00",X"EE",X"DD",X"59",
		X"00",X"E4",X"99",X"59",X"00",X"33",X"9D",X"90",X"00",X"14",X"DD",X"00",X"00",X"14",X"9D",X"50",
		X"00",X"14",X"9D",X"50",X"00",X"41",X"DD",X"50",X"00",X"45",X"DD",X"50",X"00",X"15",X"9D",X"50",
		X"00",X"45",X"99",X"50",X"00",X"45",X"99",X"50",X"00",X"45",X"11",X"50",X"00",X"41",X"99",X"50",
		X"00",X"49",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"15",X"99",X"00",X"00",X"59",X"99",X"00",
		X"00",X"15",X"11",X"00",X"00",X"55",X"44",X"00",X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"99",X"99",X"99",X"00",X"55",X"55",X"11",X"00",X"15",X"51",X"55",X"00",
		X"99",X"99",X"49",X"00",X"59",X"99",X"59",X"00",X"55",X"59",X"99",X"00",X"14",X"11",X"99",X"00",
		X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"91",X"00",X"99",X"99",X"95",X"00",X"99",X"99",X"99",X"00",
		X"59",X"99",X"99",X"00",X"51",X"51",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"49",X"99",X"00",
		X"54",X"54",X"99",X"00",X"59",X"45",X"99",X"00",X"99",X"54",X"55",X"00",X"19",X"45",X"94",X"00",
		X"91",X"54",X"91",X"00",X"91",X"95",X"55",X"00",X"09",X"99",X"59",X"00",X"09",X"59",X"19",X"00",
		X"00",X"55",X"59",X"00",X"00",X"51",X"59",X"00",X"00",X"59",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"59",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"51",X"00",X"00",X"99",X"45",
		X"00",X"00",X"99",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"19",X"00",X"00",
		X"44",X"45",X"90",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"59",X"00",X"44",X"55",X"45",X"00",
		X"14",X"99",X"44",X"00",X"54",X"99",X"55",X"00",X"95",X"99",X"55",X"00",X"99",X"99",X"59",X"00",
		X"99",X"99",X"90",X"00",X"59",X"99",X"90",X"00",X"55",X"99",X"90",X"00",X"15",X"95",X"00",X"00",
		X"91",X"55",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"91",X"00",X"00",
		X"99",X"55",X"00",X"00",X"09",X"59",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"91",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"11",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"91",X"00",X"00",
		X"11",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"91",X"99",X"00",X"00",X"55",X"55",X"90",X"00",
		X"49",X"95",X"90",X"00",X"49",X"99",X"90",X"00",X"49",X"59",X"90",X"00",X"15",X"54",X"00",X"00",
		X"95",X"59",X"00",X"00",X"49",X"99",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"15",X"44",X"00",X"00",X"14",X"44",X"00",
		X"00",X"19",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"19",X"44",X"90",X"00",X"59",X"54",X"90",
		X"00",X"19",X"55",X"90",X"00",X"59",X"99",X"90",X"00",X"19",X"59",X"90",X"00",X"59",X"99",X"90",
		X"00",X"11",X"99",X"90",X"00",X"54",X"99",X"90",X"00",X"11",X"99",X"90",X"00",X"55",X"95",X"00",
		X"00",X"15",X"99",X"00",X"00",X"55",X"55",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"55",X"90",
		X"00",X"59",X"99",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"09",X"09",X"00",X"99",X"09",X"09",X"00",X"22",X"09",X"09",X"00",X"22",X"09",X"09",
		X"00",X"92",X"09",X"09",X"00",X"92",X"09",X"09",X"00",X"92",X"09",X"09",X"00",X"92",X"09",X"09",
		X"00",X"92",X"09",X"09",X"00",X"92",X"99",X"99",X"00",X"92",X"99",X"99",X"00",X"22",X"22",X"22",
		X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"09",X"92",X"92",X"92",X"09",X"29",X"29",X"29",X"99",X"29",X"29",X"29",
		X"92",X"29",X"29",X"29",X"32",X"29",X"29",X"29",X"39",X"29",X"29",X"29",X"99",X"29",X"29",X"29",
		X"09",X"29",X"29",X"29",X"09",X"29",X"29",X"29",X"09",X"29",X"29",X"29",X"09",X"29",X"29",X"29",
		X"09",X"29",X"29",X"29",X"09",X"29",X"29",X"29",X"99",X"29",X"29",X"29",X"92",X"92",X"92",X"92",
		X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"09",X"09",X"09",X"92",X"99",X"99",X"99",X"92",X"92",X"92",X"92",X"92",X"22",X"22",X"22",
		X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",
		X"99",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"99",X"22",X"22",X"22",
		X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"99",X"92",X"92",X"92",X"99",X"99",X"99",X"99",
		X"00",X"09",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"99",X"99",X"99",X"99",X"22",X"92",X"92",X"92",X"29",X"29",X"29",X"92",X"29",X"29",X"29",
		X"99",X"29",X"29",X"29",X"00",X"99",X"29",X"29",X"00",X"22",X"29",X"29",X"09",X"22",X"29",X"29",
		X"09",X"99",X"29",X"29",X"99",X"00",X"29",X"29",X"92",X"00",X"29",X"29",X"92",X"99",X"29",X"29",
		X"92",X"29",X"29",X"29",X"92",X"29",X"29",X"29",X"92",X"29",X"29",X"29",X"92",X"92",X"92",X"92",
		X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"90",
		X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"AA",X"99",X"00",X"A9",X"99",X"99",X"00",X"9A",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"99",
		X"00",X"99",X"00",X"99",X"00",X"A9",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"90",
		X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"93",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"50",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"95",X"99",X"00",X"00",X"15",X"11",X"00",X"00",X"31",X"44",
		X"00",X"00",X"31",X"59",X"00",X"00",X"34",X"91",X"00",X"00",X"31",X"15",X"00",X"00",X"15",X"49",
		X"00",X"00",X"99",X"49",X"00",X"00",X"95",X"49",X"00",X"00",X"11",X"49",X"00",X"00",X"15",X"49",
		X"00",X"00",X"95",X"49",X"00",X"00",X"49",X"49",X"00",X"00",X"51",X"49",X"00",X"00",X"95",X"49",
		X"00",X"00",X"59",X"49",X"00",X"00",X"31",X"45",X"00",X"00",X"31",X"55",X"00",X"00",X"31",X"95",
		X"00",X"00",X"31",X"15",X"00",X"00",X"15",X"11",X"00",X"00",X"55",X"15",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"99",X"99",X"00",X"99",X"91",X"11",X"00",X"15",X"15",X"44",X"00",
		X"99",X"55",X"44",X"00",X"99",X"14",X"99",X"00",X"99",X"44",X"55",X"00",X"44",X"41",X"55",X"00",
		X"44",X"19",X"55",X"00",X"44",X"19",X"51",X"00",X"44",X"59",X"51",X"00",X"44",X"99",X"51",X"00",
		X"44",X"59",X"99",X"00",X"44",X"99",X"51",X"00",X"44",X"59",X"51",X"00",X"44",X"19",X"51",X"00",
		X"44",X"19",X"51",X"00",X"44",X"41",X"15",X"00",X"99",X"44",X"55",X"00",X"99",X"14",X"99",X"00",
		X"99",X"55",X"44",X"00",X"51",X"44",X"44",X"00",X"99",X"51",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"05",X"99",X"00",X"00",X"95",X"59",
		X"00",X"00",X"55",X"41",X"00",X"00",X"59",X"44",X"00",X"00",X"95",X"44",X"00",X"00",X"55",X"51",
		X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"11",X"00",X"00",X"59",X"14",X"00",X"00",X"95",X"14",
		X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"51",X"00",X"00",X"91",X"44",
		X"00",X"00",X"E3",X"14",X"00",X"00",X"E3",X"44",X"00",X"00",X"31",X"11",X"00",X"00",X"14",X"45",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"90",X"00",X"00",
		X"19",X"59",X"00",X"00",X"44",X"11",X"00",X"00",X"44",X"44",X"95",X"00",X"44",X"99",X"99",X"00",
		X"44",X"99",X"41",X"00",X"44",X"11",X"44",X"00",X"44",X"44",X"54",X"00",X"44",X"44",X"95",X"00",
		X"00",X"00",X"54",X"49",X"00",X"00",X"55",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"05",X"59",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"95",X"00",X"44",X"45",X"95",X"00",X"44",X"49",X"95",X"00",X"44",X"59",X"55",X"00",
		X"14",X"99",X"51",X"00",X"99",X"99",X"55",X"00",X"99",X"99",X"51",X"00",X"99",X"99",X"95",X"00",
		X"19",X"19",X"15",X"00",X"95",X"44",X"15",X"00",X"59",X"14",X"59",X"00",X"00",X"55",X"59",X"00",
		X"00",X"49",X"91",X"00",X"00",X"44",X"94",X"00",X"00",X"54",X"14",X"00",X"00",X"99",X"41",X"00",
		X"00",X"59",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",
		X"00",X"00",X"00",X"34",X"00",X"00",X"00",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"99",X"91",
		X"00",X"00",X"95",X"59",X"00",X"00",X"59",X"11",X"00",X"00",X"99",X"44",X"00",X"00",X"59",X"44",
		X"00",X"00",X"E5",X"44",X"00",X"00",X"E3",X"44",X"00",X"00",X"31",X"54",X"00",X"00",X"14",X"45",
		X"00",X"00",X"14",X"44",X"00",X"00",X"14",X"14",X"00",X"00",X"54",X"49",X"00",X"00",X"95",X"59",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"14",X"50",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"95",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"51",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"95",X"90",X"00",X"44",X"99",X"55",X"00",X"44",X"91",X"49",X"00",X"44",X"54",X"44",X"00",
		X"91",X"44",X"44",X"00",X"91",X"44",X"49",X"00",X"91",X"44",X"55",X"00",X"91",X"44",X"54",X"00",
		X"91",X"44",X"45",X"00",X"45",X"45",X"55",X"00",X"14",X"95",X"59",X"00",X"54",X"55",X"90",X"00",
		X"95",X"51",X"00",X"00",X"99",X"15",X"00",X"00",X"09",X"55",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"09",X"94",
		X"00",X"00",X"59",X"51",X"00",X"00",X"55",X"59",X"00",X"00",X"59",X"51",X"00",X"00",X"09",X"54",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"14",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"50",X"00",X"00",X"44",X"19",X"00",X"00",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"54",X"00",X"00",X"44",X"94",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"41",X"00",X"00",X"44",X"44",X"00",X"00",
		X"49",X"14",X"00",X"00",X"59",X"45",X"00",X"00",X"99",X"45",X"00",X"00",X"99",X"45",X"00",X"00",
		X"54",X"49",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"55",X"00",X"00",X"54",X"51",X"00",X"00",
		X"95",X"15",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"59",X"00",X"00",X"15",X"54",X"00",X"00",
		X"49",X"55",X"00",X"00",X"49",X"55",X"00",X"00",X"95",X"50",X"00",X"00",X"95",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"5E",X"55",X"90",
		X"00",X"EE",X"99",X"55",X"00",X"9E",X"59",X"95",X"00",X"13",X"45",X"95",X"00",X"14",X"51",X"95",
		X"00",X"14",X"11",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"41",X"41",X"95",
		X"00",X"44",X"44",X"95",X"00",X"44",X"14",X"95",X"00",X"44",X"44",X"95",X"00",X"14",X"41",X"95",
		X"00",X"45",X"44",X"95",X"00",X"49",X"95",X"95",X"00",X"49",X"99",X"95",X"00",X"49",X"99",X"95",
		X"00",X"99",X"99",X"95",X"00",X"94",X"99",X"95",X"00",X"19",X"44",X"90",X"00",X"55",X"41",X"90",
		X"00",X"19",X"41",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",
		X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",
		X"00",X"15",X"44",X"50",X"00",X"14",X"44",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",
		X"00",X"19",X"14",X"95",X"00",X"51",X"99",X"95",X"00",X"55",X"99",X"95",X"00",X"55",X"99",X"95",
		X"00",X"15",X"11",X"95",X"00",X"19",X"44",X"95",X"00",X"15",X"44",X"95",X"00",X"49",X"44",X"95",
		X"00",X"45",X"44",X"95",X"00",X"45",X"55",X"95",X"00",X"45",X"55",X"95",X"00",X"45",X"15",X"95",
		X"00",X"45",X"55",X"55",X"00",X"99",X"55",X"50",X"00",X"95",X"91",X"95",X"00",X"95",X"55",X"95",
		X"00",X"99",X"99",X"90",X"00",X"05",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"9A",X"90",X"00",X"00",X"A9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"93",X"99",X"00",
		X"00",X"93",X"90",X"00",X"00",X"33",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"50",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"50",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"50",X"00",X"99",X"05",X"00",X"00",X"09",X"50",X"50",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"99",X"99",X"00",X"99",X"91",X"59",X"00",X"15",X"15",X"45",X"00",
		X"99",X"55",X"54",X"00",X"99",X"14",X"99",X"00",X"99",X"44",X"99",X"00",X"44",X"41",X"99",X"00",
		X"44",X"19",X"99",X"00",X"44",X"19",X"99",X"00",X"44",X"59",X"99",X"00",X"44",X"99",X"99",X"00",
		X"44",X"59",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"59",X"99",X"00",X"44",X"19",X"99",X"00",
		X"44",X"19",X"99",X"00",X"44",X"41",X"95",X"00",X"99",X"44",X"55",X"00",X"99",X"14",X"99",X"00",
		X"99",X"55",X"49",X"00",X"51",X"44",X"99",X"00",X"99",X"51",X"19",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"90",X"00",X"00",
		X"19",X"59",X"00",X"00",X"44",X"11",X"90",X"00",X"44",X"44",X"95",X"00",X"44",X"99",X"99",X"00",
		X"44",X"99",X"41",X"00",X"44",X"11",X"44",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"95",X"00",
		X"44",X"44",X"95",X"00",X"44",X"45",X"95",X"00",X"44",X"49",X"99",X"00",X"44",X"59",X"99",X"00",
		X"14",X"99",X"59",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"19",X"19",X"99",X"00",X"95",X"44",X"99",X"00",X"59",X"14",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"49",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"59",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"55",X"90",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",
		X"44",X"95",X"99",X"00",X"44",X"99",X"55",X"00",X"44",X"91",X"49",X"00",X"44",X"54",X"44",X"00",
		X"91",X"44",X"54",X"00",X"91",X"44",X"45",X"00",X"91",X"45",X"55",X"00",X"91",X"55",X"59",X"00",
		X"91",X"55",X"99",X"00",X"45",X"55",X"55",X"00",X"14",X"99",X"50",X"00",X"54",X"99",X"90",X"00",
		X"95",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"54",X"00",X"00",X"44",X"94",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"41",X"00",X"00",X"44",X"44",X"00",X"00",
		X"49",X"14",X"00",X"00",X"59",X"45",X"00",X"00",X"99",X"45",X"00",X"00",X"99",X"45",X"00",X"00",
		X"54",X"54",X"00",X"00",X"14",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",
		X"95",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"50",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",
		X"00",X"15",X"44",X"50",X"00",X"14",X"44",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",
		X"00",X"19",X"14",X"95",X"00",X"51",X"99",X"95",X"00",X"55",X"99",X"95",X"00",X"55",X"99",X"95",
		X"00",X"15",X"11",X"95",X"00",X"19",X"44",X"95",X"00",X"15",X"45",X"95",X"00",X"49",X"54",X"95",
		X"00",X"49",X"55",X"95",X"00",X"15",X"99",X"95",X"00",X"95",X"95",X"95",X"00",X"15",X"99",X"95",
		X"00",X"95",X"99",X"55",X"00",X"99",X"99",X"50",X"00",X"99",X"99",X"95",X"00",X"95",X"55",X"95",
		X"00",X"99",X"09",X"90",X"00",X"05",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"95",X"99",X"00",X"00",X"35",X"11",X"00",X"00",X"35",X"44",
		X"00",X"00",X"35",X"59",X"00",X"00",X"34",X"91",X"00",X"00",X"11",X"15",X"00",X"00",X"15",X"49",
		X"00",X"00",X"99",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"D9",X"49",X"00",X"00",X"D9",X"49",
		X"00",X"00",X"99",X"49",X"00",X"00",X"D9",X"49",X"00",X"00",X"59",X"49",X"00",X"00",X"95",X"49",
		X"00",X"00",X"59",X"49",X"00",X"00",X"31",X"45",X"00",X"00",X"31",X"55",X"00",X"00",X"31",X"95",
		X"00",X"00",X"31",X"15",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"15",X"00",X"00",X"99",X"99",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"05",X"99",X"00",X"00",X"95",X"59",
		X"00",X"00",X"05",X"41",X"00",X"00",X"59",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"55",X"51",
		X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"95",X"D9",
		X"00",X"00",X"9D",X"DD",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"94",
		X"00",X"00",X"EE",X"94",X"00",X"00",X"E3",X"94",X"00",X"00",X"E3",X"11",X"00",X"00",X"34",X"45",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",
		X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"34",X"00",X"00",X"09",X"44",X"00",X"00",X"99",X"91",
		X"00",X"00",X"95",X"99",X"00",X"00",X"59",X"D9",X"00",X"00",X"99",X"9D",X"00",X"00",X"59",X"DD",
		X"00",X"00",X"EE",X"D9",X"00",X"00",X"EE",X"99",X"00",X"00",X"E3",X"99",X"00",X"00",X"34",X"95",
		X"00",X"00",X"14",X"94",X"00",X"00",X"54",X"14",X"00",X"00",X"55",X"49",X"00",X"00",X"95",X"59",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"50",X"00",X"00",X"44",X"19",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"09",X"99",
		X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"DD",X"00",X"00",X"59",X"DD",X"00",X"00",X"09",X"DD",
		X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"59",X"55",X"90",
		X"00",X"5E",X"99",X"50",X"00",X"9E",X"DD",X"90",X"00",X"13",X"93",X"50",X"00",X"54",X"D9",X"59",
		X"00",X"14",X"9D",X"95",X"00",X"54",X"9D",X"99",X"00",X"44",X"D9",X"95",X"00",X"51",X"99",X"99",
		X"00",X"44",X"9D",X"95",X"00",X"44",X"99",X"99",X"00",X"44",X"99",X"99",X"00",X"14",X"99",X"95",
		X"00",X"45",X"11",X"95",X"00",X"49",X"95",X"95",X"00",X"41",X"99",X"95",X"00",X"49",X"99",X"95",
		X"00",X"99",X"99",X"90",X"00",X"94",X"99",X"95",X"00",X"19",X"44",X"90",X"00",X"55",X"41",X"90",
		X"00",X"19",X"41",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"95",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"44",
		X"00",X"00",X"35",X"59",X"00",X"00",X"E3",X"91",X"00",X"00",X"31",X"15",X"00",X"00",X"15",X"49",
		X"00",X"00",X"99",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"D9",X"49",X"00",X"00",X"D9",X"49",
		X"00",X"00",X"99",X"49",X"00",X"00",X"D9",X"49",X"00",X"00",X"59",X"49",X"00",X"00",X"95",X"49",
		X"00",X"00",X"59",X"49",X"00",X"00",X"E3",X"45",X"00",X"00",X"E3",X"55",X"00",X"00",X"31",X"95",
		X"00",X"00",X"51",X"15",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"15",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"90",X"00",X"00",
		X"19",X"59",X"00",X"00",X"44",X"11",X"00",X"00",X"44",X"44",X"90",X"00",X"44",X"99",X"99",X"00",
		X"44",X"99",X"41",X"00",X"44",X"11",X"44",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"95",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"05",X"99",X"00",X"00",X"95",X"59",
		X"00",X"00",X"05",X"41",X"00",X"00",X"59",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"55",X"51",
		X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"95",X"D9",
		X"00",X"00",X"9D",X"DD",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"94",
		X"00",X"00",X"EE",X"94",X"00",X"00",X"EE",X"94",X"00",X"00",X"E3",X"11",X"00",X"00",X"33",X"45",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",
		X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"33",X"00",X"00",X"09",X"44",X"00",X"00",X"99",X"91",
		X"00",X"00",X"95",X"99",X"00",X"00",X"59",X"D9",X"00",X"00",X"99",X"9D",X"00",X"00",X"59",X"DD",
		X"00",X"00",X"EE",X"D9",X"00",X"00",X"E3",X"99",X"00",X"00",X"E3",X"99",X"00",X"00",X"54",X"95",
		X"00",X"00",X"14",X"94",X"00",X"00",X"54",X"14",X"00",X"00",X"55",X"49",X"00",X"00",X"95",X"59",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"50",X"00",X"00",X"44",X"19",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"09",X"99",
		X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"DD",X"00",X"00",X"59",X"DD",X"00",X"00",X"09",X"DD",
		X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"99",X"9D",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"59",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"59",X"55",X"90",
		X"00",X"5E",X"99",X"50",X"00",X"9E",X"DD",X"90",X"00",X"13",X"95",X"50",X"00",X"54",X"D9",X"59",
		X"00",X"11",X"9D",X"95",X"00",X"54",X"9D",X"99",X"00",X"44",X"D9",X"95",X"00",X"51",X"99",X"99",
		X"00",X"44",X"9D",X"95",X"00",X"44",X"99",X"99",X"00",X"44",X"99",X"99",X"00",X"14",X"99",X"95",
		X"00",X"45",X"11",X"95",X"00",X"49",X"95",X"95",X"00",X"41",X"99",X"95",X"00",X"49",X"99",X"95",
		X"00",X"99",X"99",X"90",X"00",X"94",X"99",X"95",X"00",X"19",X"44",X"90",X"00",X"55",X"41",X"90",
		X"00",X"19",X"41",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"99",X"91",X"59",X"00",X"15",X"15",X"45",X"00",
		X"99",X"55",X"54",X"00",X"99",X"14",X"99",X"00",X"99",X"44",X"99",X"00",X"44",X"41",X"99",X"00",
		X"44",X"19",X"99",X"00",X"44",X"19",X"99",X"00",X"44",X"59",X"99",X"00",X"44",X"99",X"99",X"00",
		X"44",X"59",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"59",X"99",X"00",X"44",X"19",X"99",X"00",
		X"44",X"19",X"99",X"00",X"44",X"41",X"95",X"00",X"99",X"44",X"55",X"00",X"99",X"14",X"99",X"00",
		X"99",X"55",X"49",X"00",X"51",X"44",X"99",X"00",X"99",X"51",X"19",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"95",X"00",X"44",X"45",X"95",X"00",X"44",X"49",X"99",X"00",X"44",X"59",X"99",X"00",
		X"14",X"99",X"59",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"19",X"19",X"99",X"00",X"95",X"44",X"99",X"00",X"59",X"14",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"49",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"95",X"00",X"00",X"09",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"49",X"00",X"00",X"55",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",
		X"00",X"00",X"99",X"15",X"00",X"00",X"09",X"51",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"90",X"00",
		X"44",X"95",X"99",X"00",X"44",X"99",X"55",X"00",X"44",X"91",X"49",X"00",X"44",X"54",X"44",X"00",
		X"91",X"44",X"54",X"00",X"91",X"44",X"45",X"00",X"91",X"45",X"55",X"00",X"91",X"55",X"59",X"00",
		X"91",X"55",X"99",X"00",X"45",X"55",X"55",X"00",X"14",X"99",X"50",X"00",X"54",X"99",X"90",X"00",
		X"95",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"95",X"00",X"00",X"09",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"54",X"00",X"00",X"44",X"94",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"41",X"00",X"00",X"44",X"44",X"00",X"00",
		X"49",X"14",X"00",X"00",X"59",X"45",X"00",X"00",X"99",X"45",X"00",X"00",X"99",X"45",X"00",X"00",
		X"54",X"54",X"00",X"00",X"14",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",
		X"95",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"50",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",X"00",X"59",X"44",X"50",
		X"00",X"15",X"44",X"50",X"00",X"14",X"44",X"50",X"00",X"59",X"44",X"50",X"00",X"19",X"44",X"50",
		X"00",X"19",X"14",X"95",X"00",X"51",X"99",X"95",X"00",X"55",X"99",X"95",X"00",X"55",X"99",X"95",
		X"00",X"15",X"11",X"95",X"00",X"19",X"44",X"95",X"00",X"15",X"45",X"95",X"00",X"49",X"54",X"95",
		X"00",X"49",X"55",X"95",X"00",X"15",X"99",X"95",X"00",X"95",X"95",X"95",X"00",X"15",X"99",X"95",
		X"00",X"95",X"99",X"55",X"00",X"99",X"99",X"50",X"00",X"99",X"99",X"95",X"00",X"95",X"55",X"95",
		X"00",X"99",X"09",X"90",X"00",X"05",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"0C",X"C0",X"00",
		X"00",X"0C",X"0C",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"99",X"00",X"00",X"C0",X"99",X"00",X"00",X"C0",X"99",X"0C",X"00",X"00",X"99",X"C0",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"50",X"CC",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"C0",
		X"00",X"C0",X"99",X"C0",X"00",X"00",X"99",X"0C",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"CC",X"05",X"00",X"00",X"C0",X"50",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"75",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"74",
		X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"74",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"71",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"11",
		X"75",X"77",X"70",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",
		X"47",X"77",X"77",X"70",X"11",X"77",X"77",X"00",X"21",X"77",X"77",X"00",X"31",X"77",X"77",X"70",
		X"31",X"77",X"77",X"77",X"32",X"77",X"77",X"77",X"32",X"77",X"77",X"77",X"32",X"77",X"77",X"77",
		X"22",X"77",X"77",X"77",X"22",X"77",X"77",X"77",X"32",X"77",X"77",X"77",X"21",X"77",X"77",X"77",
		X"17",X"77",X"77",X"77",X"47",X"77",X"77",X"77",X"74",X"74",X"77",X"77",X"41",X"14",X"77",X"77",
		X"44",X"11",X"77",X"77",X"44",X"21",X"77",X"77",X"44",X"11",X"77",X"77",X"44",X"11",X"77",X"77",
		X"74",X"11",X"77",X"77",X"77",X"14",X"77",X"77",X"77",X"17",X"77",X"77",X"47",X"47",X"77",X"77",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"71",
		X"00",X"00",X"00",X"71",X"00",X"00",X"00",X"74",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"BB",X"BB",X"99",X"00",X"CB",X"AA",X"99",X"00",X"BB",X"9A",X"94",X"00",X"BB",X"A9",X"99",
		X"00",X"BB",X"AA",X"99",X"00",X"BB",X"AA",X"99",X"00",X"BB",X"AA",X"79",X"00",X"BB",X"AA",X"79",
		X"77",X"47",X"77",X"77",X"41",X"77",X"77",X"77",X"22",X"17",X"77",X"77",X"12",X"47",X"77",X"77",
		X"44",X"47",X"77",X"77",X"F6",X"47",X"77",X"77",X"11",X"77",X"77",X"77",X"21",X"77",X"77",X"77",
		X"41",X"77",X"77",X"77",X"22",X"77",X"77",X"77",X"33",X"74",X"77",X"77",X"33",X"74",X"77",X"77",
		X"22",X"44",X"A7",X"77",X"21",X"44",X"A9",X"77",X"44",X"44",X"7B",X"77",X"11",X"41",X"47",X"77",
		X"11",X"11",X"14",X"77",X"21",X"11",X"14",X"77",X"22",X"11",X"24",X"77",X"22",X"21",X"14",X"47",
		X"22",X"12",X"19",X"99",X"22",X"21",X"19",X"99",X"22",X"22",X"49",X"99",X"23",X"22",X"9A",X"99",
		X"22",X"11",X"AB",X"99",X"22",X"32",X"AB",X"99",X"22",X"22",X"AC",X"99",X"22",X"22",X"CC",X"A9",
		X"22",X"22",X"CB",X"A9",X"22",X"22",X"AB",X"A9",X"22",X"22",X"B9",X"AA",X"22",X"22",X"97",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"99",X"BB",X"A9",X"79",X"9B",X"9A",X"99",X"79",X"BB",X"9B",X"AA",X"97",X"BB",X"AA",X"AA",X"99",
		X"BB",X"AA",X"AA",X"97",X"BB",X"9A",X"A9",X"99",X"BB",X"99",X"AA",X"99",X"AB",X"9B",X"AA",X"99",
		X"BB",X"BA",X"AA",X"99",X"BB",X"9A",X"AA",X"99",X"BB",X"AA",X"AA",X"99",X"B9",X"AA",X"AA",X"A9",
		X"B9",X"9A",X"AA",X"99",X"BB",X"9A",X"A9",X"99",X"BB",X"A9",X"99",X"99",X"9B",X"99",X"99",X"99",
		X"99",X"9A",X"99",X"99",X"7A",X"AA",X"A9",X"99",X"97",X"AB",X"AA",X"97",X"99",X"BB",X"A9",X"99",
		X"77",X"BA",X"A9",X"77",X"47",X"AA",X"A9",X"97",X"44",X"BA",X"AA",X"79",X"44",X"A9",X"AA",X"97",
		X"47",X"B9",X"AA",X"77",X"41",X"B9",X"AA",X"77",X"47",X"BA",X"AA",X"77",X"17",X"BA",X"AA",X"97",
		X"70",X"CB",X"AA",X"77",X"70",X"DC",X"AA",X"79",X"00",X"CC",X"AA",X"97",X"00",X"BB",X"AA",X"79",
		X"22",X"12",X"99",X"AB",X"22",X"22",X"99",X"BB",X"22",X"22",X"9A",X"BB",X"22",X"24",X"9A",X"7A",
		X"22",X"49",X"9A",X"AA",X"22",X"9B",X"B9",X"AA",X"22",X"AB",X"AA",X"AA",X"22",X"BB",X"AA",X"BC",
		X"22",X"BB",X"AA",X"BB",X"22",X"BA",X"AA",X"BB",X"22",X"AA",X"BA",X"BB",X"22",X"AA",X"BB",X"AB",
		X"22",X"BA",X"BB",X"BA",X"22",X"BA",X"BA",X"A7",X"23",X"AA",X"BB",X"AA",X"13",X"AA",X"BB",X"AA",
		X"22",X"AA",X"AA",X"9A",X"12",X"AA",X"AB",X"99",X"22",X"AA",X"AA",X"99",X"12",X"AA",X"AA",X"97",
		X"14",X"AA",X"AA",X"97",X"1A",X"AA",X"AA",X"97",X"1B",X"AA",X"AA",X"77",X"1A",X"BA",X"AA",X"77",
		X"1A",X"AA",X"AA",X"77",X"4B",X"BB",X"A9",X"77",X"BB",X"AB",X"A9",X"77",X"BB",X"BB",X"A9",X"77",
		X"BB",X"BB",X"A9",X"77",X"BB",X"BB",X"AA",X"77",X"AB",X"BB",X"BA",X"77",X"AB",X"BB",X"AA",X"77",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"02",X"21",X"00",X"00",X"22",X"11",
		X"00",X"00",X"22",X"14",X"00",X"00",X"22",X"11",X"00",X"00",X"22",X"41",X"00",X"00",X"22",X"10",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"10",
		X"00",X"00",X"22",X"10",X"00",X"00",X"23",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"21",X"00",X"00",X"22",X"12",X"00",X"00",X"12",X"11",X"00",X"00",X"12",X"21",
		X"00",X"00",X"12",X"21",X"00",X"00",X"02",X"21",X"00",X"00",X"01",X"21",X"00",X"00",X"00",X"21",
		X"00",X"BB",X"AA",X"79",X"00",X"AB",X"AA",X"97",X"00",X"AA",X"AA",X"79",X"00",X"AA",X"A9",X"97",
		X"00",X"AA",X"AA",X"79",X"00",X"AA",X"A9",X"99",X"00",X"AA",X"99",X"99",X"00",X"9A",X"99",X"AA",
		X"00",X"99",X"99",X"A9",X"00",X"99",X"99",X"AA",X"00",X"99",X"99",X"AA",X"00",X"AA",X"A9",X"9A",
		X"00",X"9A",X"AA",X"AA",X"00",X"99",X"AA",X"A9",X"00",X"44",X"9A",X"99",X"00",X"17",X"99",X"9A",
		X"00",X"41",X"99",X"99",X"00",X"24",X"B9",X"9A",X"00",X"21",X"BB",X"9A",X"00",X"21",X"79",X"B9",
		X"00",X"22",X"47",X"B9",X"00",X"21",X"11",X"B9",X"00",X"22",X"21",X"BB",X"00",X"21",X"12",X"B9",
		X"00",X"21",X"21",X"AA",X"00",X"12",X"22",X"79",X"00",X"02",X"22",X"77",X"00",X"02",X"22",X"77",
		X"00",X"02",X"2B",X"79",X"00",X"02",X"BB",X"9B",X"00",X"02",X"BB",X"9C",X"00",X"02",X"14",X"9C",
		X"AB",X"CC",X"AA",X"74",X"AA",X"CB",X"79",X"77",X"BA",X"CC",X"77",X"77",X"BB",X"CC",X"97",X"77",
		X"BA",X"DC",X"77",X"77",X"BA",X"DC",X"79",X"77",X"AB",X"CC",X"99",X"77",X"A9",X"CC",X"99",X"77",
		X"A9",X"BC",X"A9",X"77",X"AA",X"CB",X"A9",X"77",X"AA",X"BB",X"99",X"74",X"AA",X"BB",X"99",X"77",
		X"AA",X"AB",X"97",X"74",X"9A",X"AA",X"77",X"77",X"99",X"AA",X"77",X"74",X"B9",X"99",X"97",X"44",
		X"99",X"99",X"79",X"44",X"99",X"79",X"77",X"44",X"9A",X"97",X"77",X"44",X"BB",X"99",X"77",X"41",
		X"BA",X"97",X"77",X"41",X"AA",X"B7",X"79",X"42",X"AA",X"99",X"79",X"41",X"AB",X"77",X"79",X"42",
		X"99",X"77",X"99",X"41",X"99",X"B7",X"70",X"12",X"77",X"77",X"90",X"11",X"47",X"77",X"00",X"12",
		X"11",X"14",X"90",X"11",X"C2",X"14",X"90",X"12",X"22",X"44",X"00",X"11",X"22",X"44",X"00",X"11",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"22",X"17",X"00",X"02",X"22",X"12",X"00",X"00",X"22",X"11",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"40",X"00",X"22",X"22",X"20",X"00",X"22",X"22",
		X"20",X"00",X"22",X"22",X"24",X"00",X"22",X"22",X"12",X"00",X"22",X"22",X"22",X"00",X"22",X"22",
		X"11",X"00",X"12",X"22",X"21",X"00",X"21",X"22",X"12",X"22",X"42",X"22",X"21",X"11",X"44",X"12",
		X"12",X"22",X"14",X"12",X"21",X"12",X"21",X"11",X"22",X"12",X"22",X"11",X"22",X"21",X"11",X"11",
		X"22",X"21",X"11",X"11",X"22",X"12",X"17",X"74",X"22",X"12",X"14",X"45",X"11",X"11",X"14",X"4E",
		X"41",X"21",X"21",X"EE",X"00",X"21",X"14",X"E5",X"00",X"22",X"12",X"55",X"00",X"11",X"42",X"55",
		X"22",X"11",X"00",X"11",X"22",X"12",X"00",X"11",X"22",X"22",X"00",X"41",X"22",X"22",X"20",X"01",
		X"22",X"21",X"E7",X"01",X"22",X"22",X"EE",X"04",X"22",X"22",X"7E",X"00",X"23",X"22",X"77",X"00",
		X"23",X"22",X"77",X"00",X"23",X"22",X"75",X"00",X"32",X"11",X"77",X"00",X"22",X"21",X"77",X"00",
		X"23",X"11",X"57",X"00",X"32",X"17",X"57",X"00",X"22",X"7E",X"75",X"00",X"22",X"7E",X"57",X"00",
		X"22",X"E5",X"55",X"00",X"22",X"55",X"55",X"50",X"22",X"55",X"55",X"E5",X"22",X"E5",X"55",X"55",
		X"22",X"E5",X"55",X"5E",X"2E",X"E5",X"55",X"55",X"EE",X"E5",X"55",X"55",X"E5",X"E5",X"55",X"5E",
		X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"E5",X"5E",X"55",X"55",
		X"E5",X"EE",X"55",X"75",X"E5",X"5E",X"55",X"55",X"55",X"5E",X"55",X"75",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"41",X"42",X"57",X"00",X"77",X"71",X"57",X"00",X"77",X"71",X"55",X"00",X"77",X"74",X"55",
		X"00",X"77",X"77",X"55",X"00",X"57",X"77",X"75",X"00",X"55",X"57",X"57",X"00",X"EE",X"75",X"57",
		X"00",X"EE",X"57",X"75",X"00",X"E5",X"55",X"57",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"57",
		X"04",X"55",X"55",X"57",X"41",X"E5",X"55",X"74",X"42",X"57",X"E5",X"55",X"22",X"21",X"EE",X"55",
		X"22",X"21",X"EE",X"E5",X"33",X"21",X"5E",X"54",X"32",X"22",X"EE",X"54",X"22",X"11",X"EE",X"57",
		X"22",X"22",X"5E",X"75",X"22",X"21",X"7E",X"77",X"22",X"12",X"17",X"57",X"22",X"22",X"12",X"75",
		X"22",X"12",X"22",X"77",X"22",X"22",X"21",X"77",X"22",X"22",X"11",X"77",X"22",X"21",X"11",X"74",
		X"21",X"22",X"11",X"47",X"12",X"22",X"17",X"74",X"22",X"22",X"11",X"44",X"12",X"11",X"17",X"44",
		X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"57",X"77",X"55",X"55",X"55",
		X"55",X"55",X"55",X"57",X"57",X"55",X"55",X"55",X"77",X"55",X"55",X"55",X"57",X"55",X"55",X"55",
		X"75",X"55",X"E5",X"55",X"57",X"55",X"E5",X"55",X"75",X"55",X"55",X"55",X"75",X"55",X"55",X"55",
		X"75",X"55",X"EE",X"55",X"75",X"55",X"55",X"55",X"7E",X"55",X"55",X"55",X"75",X"55",X"77",X"55",
		X"5E",X"55",X"11",X"55",X"75",X"75",X"11",X"55",X"5E",X"27",X"22",X"05",X"75",X"21",X"23",X"00",
		X"5E",X"22",X"32",X"14",X"4E",X"22",X"32",X"14",X"57",X"22",X"23",X"14",X"41",X"22",X"23",X"14",
		X"41",X"22",X"22",X"11",X"41",X"22",X"22",X"14",X"41",X"22",X"23",X"11",X"41",X"22",X"22",X"14",
		X"41",X"22",X"32",X"11",X"44",X"22",X"23",X"14",X"41",X"22",X"32",X"11",X"41",X"22",X"22",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"07",X"40",X"00",X"C4",X"07",X"44",X"44",X"CC",
		X"04",X"CC",X"CD",X"CC",X"04",X"CD",X"CC",X"CC",X"04",X"CB",X"AC",X"FC",X"00",X"CC",X"DD",X"FC",
		X"00",X"CF",X"DD",X"FC",X"00",X"CF",X"DD",X"FC",X"00",X"CF",X"DD",X"CC",X"00",X"C6",X"DD",X"CC",
		X"00",X"C6",X"DD",X"CC",X"00",X"CD",X"DD",X"C4",X"00",X"CD",X"DD",X"C0",X"00",X"CD",X"DD",X"C0",
		X"00",X"CD",X"DD",X"70",X"00",X"CD",X"DD",X"00",X"00",X"CC",X"DC",X"00",X"00",X"CC",X"DC",X"00",
		X"00",X"CC",X"DC",X"00",X"00",X"CC",X"DC",X"00",X"00",X"CC",X"D7",X"00",X"00",X"4C",X"4D",X"00",
		X"00",X"44",X"4C",X"00",X"00",X"C4",X"CF",X"00",X"00",X"7D",X"FA",X"00",X"00",X"77",X"47",X"00",
		X"00",X"07",X"C7",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"C7",X"00",X"00",X"0C",X"CC",X"00",X"00",X"CD",X"CC",X"00",X"00",X"CD",X"DC",X"00",
		X"00",X"CD",X"DC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"76",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"67",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"57",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"BB",X"A9",X"79",X"9B",X"9A",X"99",X"79",X"BB",X"9B",X"AA",X"97",X"BB",X"AA",X"AA",X"99",
		X"BB",X"AA",X"AA",X"97",X"BB",X"9A",X"A9",X"99",X"BB",X"99",X"AA",X"99",X"AB",X"9B",X"AA",X"99",
		X"BB",X"BA",X"AA",X"99",X"BB",X"9A",X"AA",X"99",X"BB",X"AA",X"AA",X"99",X"B9",X"AA",X"AA",X"A9",
		X"B9",X"9A",X"AA",X"99",X"BB",X"9A",X"A9",X"99",X"BB",X"A9",X"99",X"99",X"9B",X"99",X"99",X"99",
		X"99",X"9A",X"99",X"99",X"7A",X"AA",X"A9",X"99",X"97",X"AB",X"AA",X"97",X"99",X"BB",X"A9",X"99",
		X"77",X"BA",X"A9",X"77",X"47",X"AB",X"A9",X"97",X"44",X"BB",X"AA",X"79",X"44",X"BB",X"AA",X"97",
		X"47",X"BB",X"AA",X"77",X"41",X"9A",X"AA",X"77",X"47",X"B9",X"AA",X"77",X"17",X"BB",X"AA",X"97",
		X"70",X"CB",X"AA",X"77",X"70",X"DC",X"AA",X"79",X"00",X"CC",X"AA",X"97",X"00",X"BB",X"AA",X"79",
		X"AB",X"CC",X"AA",X"74",X"AA",X"CB",X"A9",X"77",X"BA",X"CC",X"AA",X"77",X"BB",X"CC",X"B4",X"77",
		X"BA",X"DC",X"44",X"77",X"BA",X"DC",X"49",X"77",X"AB",X"CC",X"99",X"77",X"A9",X"CC",X"99",X"77",
		X"A9",X"BC",X"A9",X"77",X"AA",X"CB",X"A9",X"77",X"AA",X"BB",X"99",X"74",X"AA",X"BB",X"99",X"77",
		X"AA",X"AB",X"97",X"74",X"9A",X"AA",X"77",X"77",X"99",X"AA",X"77",X"74",X"B9",X"99",X"97",X"44",
		X"99",X"99",X"79",X"44",X"99",X"79",X"77",X"44",X"9A",X"97",X"77",X"44",X"BB",X"99",X"77",X"41",
		X"BA",X"97",X"77",X"41",X"AA",X"B7",X"79",X"42",X"AA",X"99",X"79",X"41",X"AB",X"77",X"79",X"42",
		X"99",X"77",X"99",X"41",X"99",X"B7",X"70",X"12",X"77",X"77",X"90",X"11",X"47",X"77",X"00",X"12",
		X"11",X"14",X"90",X"11",X"C2",X"14",X"90",X"12",X"22",X"44",X"00",X"11",X"22",X"44",X"00",X"11",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",
		X"00",X"07",X"77",X"77",X"00",X"07",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"14",X"77",
		X"00",X"77",X"14",X"77",X"00",X"77",X"21",X"77",X"00",X"07",X"21",X"77",X"00",X"07",X"24",X"77",
		X"00",X"07",X"77",X"77",X"00",X"07",X"16",X"77",X"00",X"04",X"21",X"77",X"00",X"00",X"13",X"77",
		X"00",X"00",X"13",X"77",X"00",X"07",X"42",X"77",X"00",X"07",X"41",X"77",X"00",X"07",X"24",X"77",
		X"00",X"07",X"44",X"77",X"00",X"00",X"12",X"77",X"00",X"00",X"12",X"77",X"00",X"00",X"21",X"77",
		X"00",X"00",X"14",X"77",X"00",X"00",X"47",X"A7",X"00",X"00",X"11",X"A7",X"00",X"00",X"21",X"9A",
		X"00",X"00",X"22",X"CA",X"00",X"9C",X"22",X"9B",X"00",X"BB",X"22",X"CB",X"09",X"AB",X"22",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"02",
		X"99",X"A9",X"22",X"97",X"BB",X"A9",X"22",X"79",X"BB",X"A9",X"22",X"99",X"BB",X"A9",X"22",X"AB",
		X"BB",X"AA",X"22",X"AB",X"BB",X"AA",X"22",X"BB",X"BA",X"A9",X"23",X"BB",X"B9",X"99",X"22",X"BB",
		X"9A",X"99",X"22",X"AB",X"9A",X"A9",X"24",X"AA",X"77",X"A9",X"1A",X"AA",X"47",X"AA",X"1A",X"AA",
		X"47",X"AA",X"1A",X"A9",X"40",X"AA",X"BA",X"A9",X"70",X"AA",X"BA",X"A9",X"00",X"AA",X"AA",X"A9",
		X"00",X"AA",X"AA",X"A9",X"00",X"AA",X"AA",X"A9",X"00",X"AA",X"AA",X"A9",X"00",X"99",X"9A",X"A9",
		X"00",X"99",X"99",X"A9",X"00",X"9A",X"9A",X"99",X"00",X"A9",X"99",X"97",X"00",X"99",X"99",X"77",
		X"00",X"9A",X"99",X"77",X"00",X"B9",X"9B",X"77",X"00",X"44",X"BA",X"77",X"00",X"24",X"AB",X"77",
		X"00",X"21",X"99",X"70",X"00",X"21",X"77",X"70",X"00",X"2B",X"12",X"70",X"00",X"B4",X"22",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"50",X"00",X"22",X"22",X"E5",X"00",X"23",X"22",X"7E",
		X"00",X"23",X"22",X"77",X"40",X"22",X"33",X"77",X"20",X"22",X"22",X"57",X"10",X"22",X"23",X"77",
		X"14",X"12",X"11",X"57",X"11",X"47",X"77",X"55",X"12",X"17",X"55",X"55",X"22",X"21",X"5E",X"55",
		X"22",X"12",X"55",X"55",X"22",X"14",X"57",X"55",X"41",X"27",X"E5",X"55",X"00",X"14",X"55",X"55",
		X"00",X"44",X"55",X"55",X"00",X"74",X"55",X"55",X"00",X"77",X"57",X"55",X"0E",X"55",X"75",X"55",
		X"00",X"55",X"75",X"E5",X"00",X"55",X"7E",X"55",X"01",X"55",X"7E",X"E5",X"12",X"EE",X"75",X"55",
		X"23",X"EE",X"55",X"77",X"32",X"EE",X"55",X"22",X"22",X"5E",X"57",X"32",X"22",X"47",X"52",X"22",
		X"22",X"24",X"42",X"22",X"22",X"11",X"42",X"22",X"22",X"14",X"41",X"32",X"21",X"17",X"41",X"32",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"F0",X"0D",X"00",X"00",X"F0",X"0D",
		X"06",X"FF",X"F0",X"0D",X"06",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",
		X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"FF",X"F0",X"00",
		X"66",X"FF",X"F0",X"00",X"06",X"00",X"F0",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"DD",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"DD",
		X"0D",X"DD",X"00",X"00",X"D0",X"DD",X"00",X"00",X"D0",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"0D",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"DD",X"00",X"00",X"D0",X"DD",X"00",X"00",X"D0",X"0D",X"00",X"00",
		X"D0",X"0D",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"0D",X"0D",X"0D",X"00",
		X"0D",X"0D",X"00",X"00",X"D0",X"0D",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"13",X"30",X"30",
		X"00",X"13",X"33",X"33",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",
		X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",
		X"00",X"13",X"33",X"33",X"00",X"11",X"30",X"30",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"11",X"11",X"13",
		X"00",X"31",X"33",X"11",X"00",X"31",X"33",X"31",X"00",X"31",X"33",X"31",X"00",X"31",X"11",X"31",
		X"00",X"11",X"31",X"31",X"00",X"13",X"31",X"31",X"00",X"33",X"31",X"31",X"00",X"33",X"31",X"31",
		X"00",X"33",X"11",X"11",X"00",X"11",X"13",X"13",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"11",X"13",X"13",
		X"00",X"31",X"11",X"11",X"00",X"33",X"31",X"31",X"00",X"33",X"31",X"31",X"00",X"11",X"31",X"31",
		X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",
		X"00",X"11",X"11",X"11",X"00",X"13",X"13",X"13",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"11",X"11",X"13",
		X"00",X"11",X"33",X"11",X"00",X"33",X"33",X"31",X"00",X"03",X"33",X"31",X"00",X"31",X"11",X"31",
		X"00",X"11",X"31",X"31",X"00",X"13",X"31",X"31",X"00",X"30",X"31",X"31",X"00",X"30",X"31",X"31",
		X"00",X"30",X"11",X"11",X"00",X"30",X"13",X"13",X"00",X"30",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"31",X"31",X"31",
		X"00",X"11",X"11",X"11",X"00",X"13",X"13",X"13",X"03",X"13",X"13",X"13",X"03",X"13",X"13",X"13",
		X"03",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",
		X"03",X"11",X"11",X"11",X"03",X"31",X"31",X"31",X"03",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"03",X"00",X"31",X"11",X"33",
		X"00",X"11",X"11",X"31",X"03",X"13",X"11",X"11",X"03",X"33",X"11",X"11",X"03",X"30",X"11",X"11",
		X"00",X"00",X"33",X"11",X"00",X"03",X"00",X"11",X"00",X"33",X"33",X"11",X"00",X"31",X"13",X"11",
		X"03",X"11",X"11",X"31",X"03",X"11",X"31",X"33",X"03",X"33",X"33",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"03",X"00",X"11",X"33",X"33",
		X"00",X"11",X"31",X"31",X"00",X"11",X"11",X"11",X"03",X"11",X"11",X"11",X"03",X"11",X"11",X"11",
		X"03",X"33",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"33",X"11",X"11",X"00",X"13",X"11",X"11",
		X"03",X"11",X"31",X"31",X"03",X"31",X"33",X"33",X"03",X"33",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"30",X"30",
		X"00",X"23",X"33",X"33",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",
		X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",
		X"00",X"23",X"33",X"33",X"00",X"22",X"30",X"30",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"22",X"22",X"23",
		X"00",X"32",X"33",X"22",X"00",X"32",X"33",X"32",X"00",X"32",X"33",X"32",X"00",X"32",X"22",X"32",
		X"00",X"22",X"32",X"32",X"00",X"23",X"32",X"32",X"00",X"33",X"32",X"32",X"00",X"33",X"32",X"32",
		X"00",X"33",X"22",X"22",X"00",X"22",X"23",X"23",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"22",X"23",X"23",
		X"00",X"32",X"22",X"22",X"00",X"33",X"32",X"32",X"00",X"33",X"32",X"32",X"00",X"22",X"32",X"32",
		X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",
		X"00",X"22",X"22",X"22",X"00",X"23",X"23",X"23",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"22",X"22",X"23",
		X"00",X"22",X"33",X"22",X"00",X"33",X"33",X"32",X"00",X"03",X"33",X"32",X"00",X"32",X"22",X"32",
		X"00",X"22",X"32",X"32",X"00",X"23",X"32",X"32",X"00",X"30",X"32",X"32",X"00",X"30",X"32",X"32",
		X"00",X"30",X"22",X"22",X"00",X"30",X"23",X"23",X"00",X"30",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"32",X"32",X"32",
		X"00",X"22",X"22",X"22",X"00",X"23",X"23",X"23",X"03",X"23",X"23",X"23",X"03",X"23",X"23",X"23",
		X"03",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",
		X"03",X"22",X"22",X"22",X"03",X"32",X"32",X"32",X"03",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"03",X"00",X"32",X"22",X"33",
		X"00",X"22",X"22",X"32",X"03",X"23",X"22",X"22",X"03",X"33",X"22",X"22",X"03",X"30",X"22",X"22",
		X"00",X"00",X"33",X"22",X"00",X"03",X"00",X"22",X"00",X"33",X"33",X"22",X"00",X"32",X"23",X"22",
		X"03",X"22",X"22",X"32",X"03",X"22",X"32",X"33",X"03",X"33",X"33",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"03",X"00",X"22",X"33",X"33",
		X"00",X"22",X"32",X"32",X"00",X"22",X"22",X"22",X"03",X"22",X"22",X"22",X"03",X"22",X"22",X"22",
		X"03",X"33",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"33",X"22",X"22",X"00",X"23",X"22",X"22",
		X"03",X"22",X"32",X"32",X"03",X"32",X"33",X"33",X"03",X"33",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
