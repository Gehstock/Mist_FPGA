library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_spr_bit4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_spr_bit4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"7F",X"93",X"93",X"93",X"93",X"93",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FE",X"92",X"92",X"82",X"82",X"93",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"11",X"31",X"E1",X"E3",X"E2",X"E2",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"7F",X"FF",X"FF",X"27",X"27",X"27",X"27",X"27",X"26",X"26",
		X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FE",X"FF",X"FF",X"26",X"26",X"22",X"02",X"12",X"13",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"60",X"73",X"33",X"33",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"70",X"F8",X"FC",X"FC",X"FE",X"FE",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"0C",X"1E",X"1E",X"1E",X"1E",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"14",X"04",X"06",X"1C",X"04",X"00",X"09",X"07",X"0E",X"02",X"04",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"06",X"4C",X"06",X"07",X"8F",X"DF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"20",X"00",X"04",X"00",X"00",X"20",X"01",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"04",X"00",X"00",
		X"80",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"80",X"08",X"00",X"00",X"02",X"40",X"00",X"00",
		X"00",X"00",X"02",X"03",X"01",X"00",X"01",X"00",X"00",X"04",X"0F",X"1D",X"39",X"23",X"42",X"02",
		X"3C",X"04",X"44",X"68",X"F0",X"F0",X"70",X"D0",X"10",X"33",X"CF",X"F9",X"FC",X"FE",X"F2",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"C3",X"C2",X"C2",X"C2",X"C2",X"C2",X"40",X"C0",X"C0",X"60",X"70",X"70",X"30",X"30",X"60",X"60",
		X"00",X"03",X"07",X"0F",X"0F",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"3F",X"3F",
		X"00",X"E0",X"E0",X"F0",X"F0",X"70",X"70",X"70",X"30",X"00",X"00",X"40",X"C0",X"F8",X"FC",X"FE",
		X"38",X"3F",X"1F",X"0F",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"E0",X"F0",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"04",X"04",
		X"60",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"01",X"03",X"07",X"07",X"03",X"03",X"07",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"E4",X"F8",X"E2",X"FC",X"F8",X"E4",X"B8",X"48",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"0B",X"0B",X"17",X"07",X"07",X"05",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"F0",X"E8",X"F6",X"F8",X"C0",X"A0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"05",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"05",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"60",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"0D",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"60",X"C0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"08",X"1D",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"60",X"F0",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"00",X"00",X"00",X"00",X"10",X"38",X"0D",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"18",X"18",X"30",X"78",X"FC",X"F0",X"E0",
		X"00",X"06",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"70",X"3F",X"0F",X"03",
		X"00",X"00",X"08",X"08",X"04",X"04",X"04",X"0C",X"0C",X"18",X"1C",X"3E",X"FE",X"FC",X"F0",X"C0",
		X"08",X"00",X"08",X"18",X"18",X"10",X"00",X"80",X"C0",X"C0",X"60",X"60",X"30",X"3F",X"5F",X"07",
		X"04",X"04",X"02",X"02",X"02",X"02",X"06",X"07",X"0F",X"0F",X"1E",X"7E",X"FC",X"FC",X"F8",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"0B",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"D0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0C",X"13",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"30",X"C8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"15",X"27",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"28",X"E4",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"29",X"01",X"8F",X"CF",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"24",X"20",X"F0",X"F5",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"15",X"55",X"D5",X"3B",X"3F",X"7F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"10",X"12",X"13",X"54",X"FC",X"FF",X"FF",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"08",X"04",X"03",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"15",X"55",X"D5",X"35",X"2B",X"22",X"3F",X"7F",X"7F",X"EF",
		X"00",X"00",X"80",X"C0",X"F0",X"F8",X"50",X"54",X"5A",X"08",X"28",X"AC",X"FC",X"FE",X"FE",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"10",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"04",X"00",X"00",X"00",X"01",X"21",X"3B",X"1F",
		X"03",X"07",X"0F",X"15",X"15",X"95",X"95",X"B5",X"A5",X"21",X"73",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"E0",X"F0",X"F8",X"A8",X"AA",X"8D",X"84",X"94",X"56",X"76",X"76",X"FF",X"FF",X"FF",X"FF",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"00",X"00",X"00",X"80",X"84",X"CC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"02",X"06",X"0C",X"1C",X"34",X"00",X"01",X"03",X"03",X"03",X"C7",X"FF",X"1F",
		X"7F",X"49",X"49",X"49",X"49",X"49",X"C9",X"93",X"92",X"C6",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"FE",X"96",X"96",X"82",X"92",X"9A",X"09",X"49",X"79",X"79",X"FF",X"FF",X"FF",X"FF",X"F3",X"01",
		X"00",X"00",X"00",X"40",X"20",X"00",X"08",X"3C",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E1",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0F",X"0F",X"03",X"00",
		X"38",X"79",X"01",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"FF",X"FF",X"3E",
		X"93",X"93",X"13",X"32",X"22",X"86",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"11",X"59",X"49",X"49",X"78",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"71",X"82",
		X"0C",X"3E",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F1",X"FF",X"FF",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"E0",X"C0",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",X"F0",X"3F",X"0F",X"01",
		X"02",X"06",X"04",X"04",X"0E",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"FF",X"FF",X"F3",
		X"66",X"46",X"44",X"44",X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"E7",
		X"99",X"89",X"C8",X"78",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"0C",
		X"00",X"80",X"80",X"80",X"80",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FF",X"FF",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"87",X"FC",X"F0",X"08",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FC",X"FC",X"FC",X"7C",X"7C",X"3E",X"3E",X"3E",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"01",X"10",X"04",X"00",X"00",X"00",X"00",X"18",X"07",X"01",X"2D",X"59",
		X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"40",X"A8",X"F0",X"68",X"E8",X"AC",X"94",X"38",X"EB",
		X"00",X"00",X"00",X"00",X"08",X"02",X"01",X"02",X"14",X"12",X"46",X"19",X"A7",X"22",X"67",X"3A",
		X"00",X"00",X"08",X"20",X"40",X"90",X"20",X"E0",X"50",X"C8",X"9C",X"F4",X"50",X"6A",X"B6",X"D4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"5A",X"95",X"36",X"AD",X"B5",
		X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"01",X"0A",X"07",X"05",X"0D",X"02",X"04",X"46",X"03",
		X"00",X"00",X"00",X"00",X"10",X"80",X"08",X"A0",X"C4",X"E2",X"EC",X"A1",X"91",X"7A",X"EF",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"C0",X"20",X"30",X"82",X"20",X"20",X"3D",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"12",X"14",X"26",X"6A",X"79",X"D3",X"FA",
		X"00",X"00",X"08",X"05",X"00",X"03",X"05",X"02",X"07",X"05",X"0B",X"02",X"82",X"03",X"01",X"87",
		X"00",X"00",X"00",X"E1",X"40",X"28",X"DA",X"B4",X"9A",X"27",X"98",X"C4",X"69",X"60",X"B1",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"A8",X"12",X"08",X"65",X"12",X"86",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"13",X"0E",X"3C",X"0B",X"ED",
		X"00",X"00",X"00",X"00",X"14",X"0B",X"09",X"16",X"03",X"01",X"83",X"01",X"00",X"C0",X"80",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"08",X"C2",X"81",X"B1",X"EA",X"94",X"48",X"B7",X"F3",X"31",X"AD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"42",X"4A",X"30",X"41",X"A2",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"02",X"04",X"20",X"0A",X"35",X"AD",X"1E",X"7E",
		X"08",X"02",X"00",X"02",X"09",X"07",X"03",X"05",X"83",X"02",X"81",X"C0",X"C2",X"61",X"E1",X"50",
		X"00",X"00",X"10",X"08",X"A3",X"E5",X"30",X"5A",X"CB",X"5D",X"7B",X"BF",X"ED",X"27",X"7D",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"10",X"C0",X"A8",X"20",X"60",X"A4",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0A",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"20",X"B8",X"6C",X"38",X"0D",X"02",X"09",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1D",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"80",X"00",X"00",X"50",X"0D",X"1A",X"0F",X"03",X"09",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"22",X"6F",X"15",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"14",X"38",X"78",X"7D",X"1E",X"86",X"1A",X"6C",
		X"02",X"01",X"23",X"11",X"1B",X"0B",X"01",X"01",X"02",X"03",X"01",X"04",X"01",X"02",X"20",X"0C",
		X"F5",X"5F",X"BF",X"F4",X"7E",X"DF",X"76",X"ED",X"FE",X"DA",X"64",X"F0",X"E1",X"DC",X"3B",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",
		X"00",X"20",X"00",X"00",X"08",X"00",X"00",X"82",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"02",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"04",X"0C",X"1F",X"00",X"07",X"07",X"07",
		X"38",X"1C",X"0C",X"18",X"F4",X"FE",X"DA",X"FB",X"F9",X"F0",X"01",X"81",X"81",X"C1",X"C1",X"E3",
		X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"04",X"05",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"3F",X"1F",X"0F",X"07",X"07",X"0A",X"07",X"00",X"00",X"00",X"08",X"0C",X"4F",X"47",X"47",X"63",
		X"FE",X"7E",X"7B",X"71",X"70",X"70",X"F0",X"30",X"30",X"38",X"18",X"18",X"38",X"B8",X"98",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"DF",X"FC",X"FF",X"79",X"7E",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"60",X"80",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"FF",X"FF",X"7E",X"0D",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"60",X"90",X"60",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"05",X"0D",X"0F",X"0F",X"07",X"03",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"A0",X"A0",X"40",X"40",X"E0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"05",X"02",X"0A",X"05",X"07",X"03",X"07",X"07",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"40",X"50",X"A0",X"E0",X"C0",X"80",X"80",X"80",X"00",
		X"01",X"03",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"1F",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"70",X"10",X"78",X"FC",X"FE",X"FF",X"FF",X"C7",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"01",X"00",X"00",X"01",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"1E",X"E8",X"C0",X"B0",X"60",X"C0",X"80",X"00",X"00",
		X"80",X"E0",X"F0",X"F0",X"F8",X"38",X"3C",X"1C",X"8E",X"8E",X"C7",X"F3",X"79",X"7F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0E",X"08",X"1E",X"3F",X"7F",X"FF",X"FF",X"E3",X"87",
		X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"78",X"17",X"03",X"0D",X"06",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"80",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"01",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"3E",X"78",X"58",X"D8",X"B0",X"B0",X"E0",X"C0",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"70",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"87",X"0F",X"1F",X"1F",X"3F",X"3F",X"3E",X"1E",X"9C",X"F0",X"38",X"03",X"07",X"07",X"03",X"01",
		X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"38",X"08",X"08",X"04",X"04",X"80",X"C0",X"C0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"15",X"1E",X"1A",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"3F",X"3E",X"3E",X"1E",X"1C",
		X"FF",X"FF",X"FC",X"FC",X"FB",X"67",X"1F",X"BE",X"FC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"40",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"05",X"06",X"0F",X"0F",X"1F",X"1F",X"1F",X"3E",X"3C",X"30",X"60",X"40",
		X"00",X"10",X"2C",X"78",X"78",X"70",X"18",X"1E",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"FF",X"7F",X"1E",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"76",X"66",X"7C",X"F0",X"FC",X"FF",X"7E",X"3D",X"1B",X"0B",X"05",X"0C",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"EC",X"F6",X"F7",X"FB",X"FB",X"7D",X"7F",
		X"00",X"00",X"00",X"28",X"14",X"1C",X"0E",X"0E",X"06",X"04",X"0C",X"5C",X"B8",X"D0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"18",X"18",X"50",X"D0",X"D0",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"06",X"00",X"37",X"6F",X"EF",X"DF",X"BF",X"B8",X"7C",
		X"7C",X"FC",X"EC",X"E0",X"F0",X"CF",X"3F",X"FF",X"7E",X"BC",X"D0",X"C0",X"BC",X"3C",X"7C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"28",X"38",X"70",X"70",X"60",X"20",X"30",X"3A",X"1D",X"09",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"C3",X"67",X"71",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"41",X"A8",X"7B",X"E7",X"1E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"3F",X"FF",X"F6",X"81",X"03",X"02",X"06",X"03",X"03",X"00",X"00",X"00",X"00",X"01",X"03",
		X"C0",X"80",X"77",X"F9",X"FE",X"FF",X"EF",X"1F",X"1F",X"3F",X"3F",X"3F",X"0C",X"E3",X"F3",X"FF",
		X"00",X"00",X"80",X"C0",X"E0",X"70",X"F0",X"F8",X"F8",X"E8",X"E8",X"C2",X"1E",X"FE",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",X"60",X"50",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"FC",X"3F",X"E7",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3E",X"FC",
		X"07",X"07",X"C3",X"C1",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"FF",X"FF",X"FF",X"3F",
		X"E4",X"E0",X"F0",X"F2",X"F6",X"F6",X"66",X"06",X"0F",X"1E",X"FE",X"FE",X"8E",X"C2",X"E2",X"E2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"60",X"60",X"C0",X"70",X"30",X"00",X"00",X"10",X"18",X"18",X"08",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"F8",X"7C",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0E",X"0C",X"00",X"00",X"00",X"00",X"F0",X"F8",X"7F",X"1F",X"1F",X"07",X"03",X"10",X"1C",
		X"03",X"09",X"0F",X"11",X"0D",X"1D",X"79",X"F1",X"21",X"C1",X"F1",X"FC",X"FD",X"FE",X"FE",X"3E",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"88",X"C8",X"F0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"E0",X"E0",X"30",X"38",X"2C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"D0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"0E",X"06",X"03",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"70",X"38",X"3D",X"1E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"DC",X"6C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"38",X"38",X"0C",X"1C",X"1A",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6C",X"CC",X"CE",X"1E",X"1E",X"1E",X"9E",X"BE",X"BE",X"3E",X"3E",X"3C",X"7C",X"5C",X"5C",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"87",X"2F",X"7F",X"BF",X"DF",X"DF",X"DE",X"DE",X"DC",X"9C",X"3A",X"32",X"63",X"C1",X"81",
		X"F8",X"38",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"38",X"30",X"30",X"70",X"70",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",
		X"07",X"0F",X"1F",X"1F",X"13",X"1B",X"3E",X"31",X"43",X"3B",X"77",X"77",X"E0",X"CF",X"9F",X"DF",
		X"F8",X"F8",X"78",X"70",X"F0",X"E0",X"8E",X"3F",X"BF",X"BC",X"B8",X"60",X"1A",X"79",X"7B",X"72",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"3C",X"04",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",
		X"18",X"18",X"18",X"98",X"98",X"98",X"98",X"98",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"02",X"03",X"03",X"03",X"00",X"01",X"03",X"03",X"07",X"07",X"0C",X"0B",X"0B",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"C0",X"E0",X"F8",X"FC",X"1F",X"E7",X"E9",X"C8",X"D8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0E",X"18",X"11",
		X"00",X"00",X"00",X"03",X"06",X"0C",X"0F",X"0F",X"08",X"1D",X"7D",X"FD",X"98",X"03",X"1B",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"F8",X"F0",X"06",X"7B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FD",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"05",X"24",X"02",X"00",X"01",X"10",X"04",X"19",X"00",X"21",X"00",
		X"68",X"60",X"32",X"8B",X"71",X"09",X"E6",X"07",X"14",X"00",X"02",X"40",X"08",X"31",X"64",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"60",X"C0",X"40",X"04",X"DA",X"7F",X"FD",X"FE",
		X"02",X"02",X"07",X"01",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"02",X"86",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"87",X"DE",X"87",X"31",X"0C",X"C5",X"63",X"03",X"11",X"1C",X"0B",X"03",X"00",X"02",X"03",
		X"3D",X"8C",X"E1",X"D0",X"C2",X"B3",X"F9",X"A0",X"C2",X"F1",X"78",X"7C",X"28",X"72",X"32",X"B1",
		X"8B",X"42",X"87",X"D1",X"E2",X"A4",X"C0",X"E2",X"58",X"F4",X"DE",X"6C",X"CC",X"08",X"59",X"EC",
		X"DF",X"EF",X"FE",X"AE",X"7F",X"FB",X"7F",X"5F",X"C7",X"67",X"B3",X"E5",X"E7",X"73",X"5B",X"3D",
		X"27",X"31",X"59",X"7C",X"36",X"8D",X"CF",X"DF",X"9F",X"87",X"4B",X"EE",X"EF",X"B7",X"FE",X"FD",
		X"26",X"97",X"9A",X"EE",X"FA",X"EC",X"50",X"D0",X"C0",X"94",X"8E",X"87",X"1B",X"2F",X"7F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"8C",X"8C",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"3B",X"3B",X"2C",X"24",X"62",X"42",X"41",X"81",X"00",X"04",X"0A",X"05",X"06",X"00",X"00",
		X"C0",X"A0",X"70",X"F0",X"EE",X"FF",X"FF",X"7E",X"5C",X"9C",X"88",X"49",X"09",X"0D",X"0F",X"1E",
		X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"7C",X"7E",X"7E",X"7C",X"38",X"00",
		X"01",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"01",X"00",X"07",X"0F",X"1F",X"3E",X"38",X"00",X"00",
		X"1F",X"07",X"01",X"04",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"38",X"B8",X"FC",X"FC",X"FE",X"FE",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",
		X"03",X"05",X"0E",X"0F",X"77",X"FF",X"FF",X"7A",X"38",X"39",X"11",X"02",X"30",X"70",X"F4",X"F4",
		X"D8",X"DC",X"DC",X"34",X"24",X"46",X"42",X"82",X"81",X"00",X"20",X"50",X"A0",X"60",X"00",X"00",
		X"80",X"F7",X"CF",X"BF",X"7F",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"40",X"FE",X"7E",X"3E",X"3E",X"1C",X"00",
		X"07",X"07",X"0C",X"08",X"18",X"19",X"3F",X"3F",X"7F",X"7F",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",
		X"90",X"30",X"60",X"60",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"54",X"2C",X"40",X"04",X"04",X"06",X"05",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1F",X"3D",X"7D",X"DB",X"D8",X"87",X"37",X"2F",X"2F",X"3F",X"7E",X"7F",X"C0",
		X"00",X"E0",X"F0",X"FC",X"FE",X"FF",X"FF",X"CF",X"27",X"D3",X"D9",X"B0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"70",X"78",X"AC",X"84",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"3C",X"06",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"18",X"9C",X"C8",X"C8",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"FF",X"FF",X"FE",X"F0",X"70",X"00",X"38",X"DC",X"DC",X"EE",X"F7",X"FB",X"FF",X"FF",
		X"30",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0E",X"1E",X"35",X"21",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FE",X"E7",X"8B",X"1B",X"09",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"0D",X"1B",X"1A",X"1E",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"F0",X"E6",X"4F",X"1F",X"3F",X"3F",X"7F",X"7C",X"F0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"7E",X"30",X"0F",X"8F",X"9F",X"3F",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"70",X"30",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"71",X"01",X"03",X"06",X"0C",X"F0",X"C0",X"80",X"00",
		X"71",X"71",X"E3",X"63",X"63",X"61",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"20",X"70",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"04",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"06",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"AB",X"7B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"39",X"3F",X"1E",X"14",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"1F",X"3C",X"20",X"40",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F1",X"C0",X"03",X"06",X"0C",X"CC",X"E8",X"D8",X"70",X"60",X"40",X"00",X"00",X"00",X"00",
		X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"30",X"38",X"1C",X"17",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"68",
		X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"C0",X"F8",X"3E",X"1F",X"0D",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"70",X"3C",X"1E",X"0F",X"03",X"31",X"F8",X"FC",X"7C",X"3C",X"1E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"00",X"00",X"78",X"9C",
		X"F7",X"3F",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"3F",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FF",X"3F",X"03",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0D",X"1E",X"1F",X"1B",X"09",
		X"06",X"86",X"86",X"C4",X"44",X"E0",X"60",X"62",X"32",X"B3",X"FB",X"DB",X"1B",X"1B",X"13",X"83",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"00",X"00",X"87",X"FF",X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"70",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"01",X"04",X"03",X"04",X"01",
		X"B8",X"00",X"6C",X"06",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"05",
		X"00",X"0C",X"0C",X"0C",X"18",X"18",X"98",X"B8",X"B0",X"70",X"60",X"60",X"C0",X"80",X"80",X"80",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"1F",X"39",X"F0",X"C0",X"00",X"00",
		X"78",X"B0",X"A1",X"C3",X"E2",X"F0",X"F0",X"FB",X"FB",X"FD",X"7C",X"7E",X"7E",X"3E",X"3E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"0F",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"60",X"FC",X"1F",X"03",X"00",X"00",
		X"38",X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"1F",X"1F",X"EB",X"F1",X"FC",X"FF",X"CF",
		X"00",X"00",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"F0",X"F0",X"F0",X"F0",X"30",X"10",X"10",X"30",X"20",X"20",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"BC",X"80",X"00",X"01",X"06",X"3E",X"30",X"60",
		X"78",X"7E",X"FF",X"FF",X"FC",X"60",X"00",X"01",X"03",X"07",X"07",X"CC",X"F0",X"C0",X"F0",X"01",
		X"00",X"00",X"00",X"80",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"60",X"20",X"10",X"10",X"18",
		X"02",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"01",
		X"70",X"30",X"30",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"11",X"13",X"03",X"03",X"07",X"07",X"04",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"90",X"01",X"81",X"82",X"64",X"33",X"06",X"C4",X"E4",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"98",X"88",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"01",
		X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",
		X"02",X"03",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9B",X"17",X"3F",X"7F",X"68",X"C0",X"80",X"00",X"01",X"03",X"07",X"67",X"FF",X"70",X"60",X"00",
		X"F2",X"E2",X"C2",X"16",X"18",X"18",X"0C",X"74",X"F0",X"F1",X"F0",X"E0",X"80",X"80",X"00",X"00",
		X"C0",X"40",X"60",X"20",X"30",X"10",X"10",X"08",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"06",X"07",X"07",X"07",X"03",X"01",
		X"40",X"40",X"40",X"60",X"70",X"70",X"70",X"70",X"30",X"20",X"60",X"E0",X"E0",X"E0",X"C0",X"80",
		X"06",X"04",X"04",X"14",X"24",X"18",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"07",X"0F",X"18",X"20",X"00",X"00",X"00",X"00",X"73",X"7F",X"73",X"60",X"40",X"60",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"90",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7D",X"7F",X"DF",X"FF",X"BF",X"33",X"19",X"43",X"C0",X"60",X"1F",X"07",X"0C",X"00",X"00",X"00",
		X"7F",X"FB",X"FC",X"FF",X"FF",X"FF",X"FE",X"FF",X"73",X"C4",X"00",X"88",X"F0",X"00",X"00",X"00",
		X"10",X"08",X"40",X"62",X"E9",X"CF",X"BC",X"F8",X"E0",X"7C",X"86",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"E0",X"68",X"C4",X"80",X"10",X"68",X"A1",X"04",X"38",X"00",X"00",X"00",X"00",
		X"30",X"20",X"00",X"80",X"00",X"40",X"00",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"10",X"30",X"00",X"02",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"02",X"07",X"01",X"19",
		X"C4",X"6C",X"E6",X"B2",X"93",X"48",X"6C",X"3E",X"96",X"50",X"86",X"CB",X"67",X"43",X"15",X"D7",
		X"8F",X"E7",X"83",X"58",X"49",X"00",X"00",X"9C",X"6E",X"3C",X"34",X"59",X"1D",X"3F",X"B6",X"8E",
		X"00",X"30",X"30",X"30",X"10",X"20",X"28",X"40",X"10",X"14",X"58",X"38",X"3C",X"3E",X"4A",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"01",X"01",X"03",X"02",X"01",X"01",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"28",X"91",X"10",X"22",X"2F",X"15",X"92",X"81",X"C9",X"5E",X"93",X"0C",X"46",X"31",X"00",
		X"1A",X"3F",X"7A",X"7E",X"1F",X"86",X"1B",X"6C",X"70",X"E2",X"F7",X"FC",X"C9",X"3E",X"0C",X"00",
		X"3B",X"38",X"7E",X"4F",X"65",X"B0",X"E2",X"E7",X"71",X"20",X"00",X"00",X"00",X"40",X"33",X"00",
		X"FE",X"5A",X"64",X"B0",X"E1",X"DC",X"3B",X"7F",X"B8",X"FF",X"78",X"03",X"07",X"1C",X"E0",X"00",
		X"2F",X"5F",X"3E",X"54",X"3D",X"DB",X"7E",X"FC",X"E0",X"F8",X"F1",X"8E",X"1C",X"36",X"81",X"00",
		X"BA",X"60",X"30",X"6A",X"C2",X"04",X"18",X"70",X"80",X"02",X"30",X"18",X"34",X"41",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
