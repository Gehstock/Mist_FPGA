library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"31",X"00",X"81",X"C3",X"43",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"D1",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"70",X"00",X"3C",X"71",X"00",X"3C",X"9E",X"00",X"3C",X"CB",X"00",X"3B",X"F8",X"00",X"3D",
		X"25",X"01",X"78",X"80",X"01",X"7D",X"A1",X"01",X"64",X"D7",X"01",X"64",X"FB",X"01",X"5F",X"19",
		X"02",X"73",X"40",X"02",X"74",X"77",X"02",X"74",X"B1",X"02",X"79",X"EB",X"02",X"7E",X"0C",X"03",
		X"21",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"10",X"10",X"10",X"18",X"03",X"03",X"02",
		X"03",X"03",X"03",X"1F",X"00",X"20",X"01",X"1B",X"1F",X"04",X"06",X"FF",X"03",X"81",X"0B",X"06",
		X"00",X"23",X"81",X"0B",X"07",X"00",X"25",X"81",X"01",X"03",X"03",X"81",X"F1",X"10",X"19",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1D",X"10",X"10",X"10",X"18",X"03",X"03",X"02",X"03",X"03",X"03",
		X"1F",X"00",X"20",X"01",X"1B",X"10",X"04",X"06",X"FF",X"03",X"81",X"0B",X"06",X"00",X"23",X"81",
		X"0B",X"07",X"00",X"25",X"81",X"01",X"03",X"03",X"81",X"F1",X"10",X"19",X"06",X"06",X"05",X"05",
		X"07",X"00",X"1D",X"10",X"10",X"10",X"18",X"02",X"02",X"02",X"03",X"03",X"03",X"1F",X"00",X"20",
		X"01",X"1B",X"1F",X"04",X"06",X"FF",X"03",X"81",X"0B",X"06",X"00",X"23",X"81",X"0B",X"07",X"00",
		X"25",X"81",X"01",X"03",X"03",X"81",X"F1",X"10",X"19",X"01",X"01",X"01",X"01",X"01",X"00",X"1D",
		X"10",X"10",X"10",X"18",X"03",X"03",X"02",X"03",X"03",X"03",X"1F",X"00",X"10",X"01",X"1B",X"09",
		X"04",X"06",X"FF",X"03",X"81",X"0B",X"06",X"00",X"23",X"81",X"0B",X"07",X"00",X"25",X"81",X"01",
		X"03",X"03",X"81",X"F1",X"10",X"19",X"C8",X"C8",X"64",X"01",X"00",X"FA",X"1D",X"0F",X"0F",X"0F",
		X"18",X"02",X"02",X"02",X"03",X"03",X"03",X"1B",X"1F",X"04",X"06",X"0A",X"03",X"81",X"01",X"01",
		X"0B",X"03",X"00",X"23",X"81",X"0B",X"04",X"00",X"25",X"81",X"0B",X"10",X"00",X"27",X"81",X"03",
		X"03",X"81",X"EC",X"06",X"0D",X"05",X"81",X"06",X"1E",X"03",X"81",X"01",X"0B",X"0A",X"00",X"23",
		X"81",X"0B",X"0A",X"00",X"25",X"81",X"0B",X"40",X"00",X"27",X"81",X"03",X"03",X"81",X"EC",X"0A",
		X"FF",X"2B",X"81",X"0A",X"FF",X"2C",X"81",X"0A",X"FF",X"2D",X"81",X"03",X"05",X"81",X"D8",X"10",
		X"1D",X"0C",X"05",X"09",X"18",X"03",X"03",X"03",X"03",X"03",X"03",X"19",X"00",X"01",X"50",X"01",
		X"90",X"01",X"06",X"28",X"05",X"81",X"0B",X"F9",X"FF",X"23",X"81",X"01",X"03",X"05",X"81",X"F6",
		X"10",X"1D",X"0D",X"0D",X"00",X"18",X"02",X"02",X"02",X"03",X"03",X"03",X"06",X"0F",X"05",X"81",
		X"19",X"37",X"00",X"30",X"00",X"00",X"00",X"06",X"14",X"03",X"81",X"01",X"0B",X"10",X"00",X"23",
		X"81",X"0B",X"12",X"00",X"25",X"81",X"03",X"03",X"81",X"F1",X"0A",X"FF",X"2B",X"81",X"0A",X"FF",
		X"2C",X"81",X"03",X"05",X"81",X"DA",X"10",X"1D",X"10",X"F0",X"F0",X"1F",X"80",X"00",X"01",X"18",
		X"03",X"03",X"03",X"03",X"03",X"03",X"19",X"01",X"00",X"00",X"00",X"00",X"00",X"06",X"20",X"05",
		X"81",X"0B",X"02",X"00",X"23",X"81",X"01",X"03",X"05",X"81",X"F6",X"1D",X"10",X"F0",X"A0",X"1F",
		X"80",X"01",X"01",X"19",X"08",X"00",X"00",X"00",X"00",X"00",X"06",X"10",X"05",X"81",X"0B",X"20",
		X"00",X"23",X"81",X"01",X"03",X"05",X"81",X"F6",X"10",X"19",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"02",X"03",X"03",X"03",X"03",X"03",X"1D",X"10",X"50",X"50",X"1B",X"1F",X"07",X"1F",X"C0",
		X"04",X"0C",X"06",X"1E",X"03",X"81",X"17",X"0A",X"FF",X"29",X"81",X"03",X"03",X"81",X"F7",X"10",
		X"19",X"30",X"00",X"F0",X"00",X"00",X"00",X"1D",X"0F",X"0F",X"00",X"18",X"03",X"03",X"03",X"03",
		X"03",X"03",X"06",X"0D",X"05",X"81",X"06",X"14",X"03",X"81",X"01",X"01",X"0B",X"01",X"00",X"23",
		X"81",X"0B",X"FF",X"FF",X"25",X"81",X"03",X"03",X"81",X"F1",X"0A",X"FF",X"2B",X"81",X"0A",X"FF",
		X"2C",X"81",X"03",X"05",X"81",X"E0",X"10",X"19",X"F0",X"00",X"90",X"00",X"90",X"00",X"1D",X"0F",
		X"0F",X"F0",X"18",X"03",X"03",X"03",X"03",X"03",X"03",X"1B",X"1F",X"07",X"06",X"0D",X"05",X"81",
		X"06",X"14",X"03",X"81",X"01",X"01",X"0B",X"02",X"00",X"23",X"81",X"0B",X"02",X"00",X"25",X"81",
		X"03",X"03",X"81",X"F1",X"0A",X"01",X"2B",X"81",X"0A",X"FF",X"2C",X"81",X"03",X"05",X"81",X"E0",
		X"10",X"19",X"F0",X"00",X"90",X"00",X"90",X"00",X"1D",X"0F",X"0F",X"F0",X"18",X"03",X"03",X"03",
		X"03",X"03",X"03",X"1B",X"1F",X"07",X"06",X"0D",X"05",X"81",X"06",X"14",X"03",X"81",X"01",X"01",
		X"0B",X"FE",X"FF",X"23",X"81",X"0B",X"FE",X"FF",X"25",X"81",X"03",X"03",X"81",X"F1",X"0A",X"01",
		X"2B",X"81",X"0A",X"FF",X"2C",X"81",X"03",X"05",X"81",X"E0",X"10",X"1D",X"0F",X"0F",X"0F",X"18",
		X"03",X"03",X"03",X"03",X"03",X"03",X"19",X"F0",X"02",X"50",X"03",X"90",X"08",X"06",X"28",X"05",
		X"81",X"0B",X"F7",X"FF",X"23",X"81",X"17",X"03",X"05",X"81",X"F6",X"10",X"19",X"F0",X"00",X"90",
		X"00",X"90",X"00",X"1D",X"0F",X"0F",X"F0",X"18",X"02",X"02",X"02",X"03",X"03",X"03",X"06",X"0D",
		X"05",X"81",X"06",X"14",X"03",X"81",X"01",X"01",X"0B",X"FE",X"FF",X"23",X"81",X"0B",X"FE",X"FF",
		X"25",X"81",X"03",X"03",X"81",X"F1",X"0A",X"01",X"2B",X"81",X"0A",X"FF",X"2C",X"81",X"03",X"05",
		X"81",X"E0",X"10",X"0E",X"10",X"CD",X"70",X"06",X"0E",X"40",X"CD",X"70",X"06",X"CD",X"FE",X"03",
		X"21",X"00",X"80",X"01",X"00",X"04",X"36",X"00",X"23",X"0D",X"20",X"FA",X"10",X"F8",X"3E",X"3F",
		X"32",X"2A",X"81",X"32",X"38",X"81",X"CD",X"0C",X"04",X"01",X"00",X"00",X"ED",X"56",X"FB",X"ED",
		X"5B",X"01",X"81",X"7A",X"B3",X"28",X"16",X"F3",X"31",X"00",X"81",X"CD",X"70",X"06",X"CD",X"51",
		X"06",X"ED",X"4B",X"01",X"81",X"11",X"00",X"00",X"ED",X"53",X"01",X"81",X"FB",X"0A",X"03",X"26",
		X"00",X"87",X"6F",X"11",X"9C",X"03",X"19",X"7E",X"23",X"66",X"6F",X"E9",X"D3",X"04",X"E5",X"04",
		X"05",X"05",X"11",X"05",X"1E",X"05",X"28",X"05",X"34",X"05",X"41",X"05",X"53",X"05",X"5D",X"05",
		X"69",X"05",X"78",X"05",X"92",X"05",X"A3",X"05",X"B9",X"05",X"CD",X"05",X"D3",X"05",X"F3",X"05",
		X"06",X"06",X"15",X"06",X"3A",X"06",X"46",X"06",X"4A",X"06",X"F5",X"04",X"36",X"04",X"45",X"04",
		X"4E",X"04",X"82",X"04",X"87",X"04",X"A5",X"04",X"AA",X"04",X"B9",X"04",X"BE",X"04",X"E3",X"05",
		X"21",X"44",X"81",X"06",X"06",X"11",X"00",X"00",X"CB",X"23",X"CB",X"12",X"CB",X"23",X"CB",X"12",
		X"7E",X"E6",X"03",X"B3",X"5F",X"2B",X"10",X"F0",X"21",X"00",X"90",X"19",X"77",X"C9",X"3E",X"03",
		X"21",X"3F",X"81",X"06",X"06",X"77",X"10",X"FD",X"CD",X"E0",X"03",X"C9",X"11",X"23",X"81",X"0E",
		X"10",X"CD",X"1D",X"04",X"11",X"31",X"81",X"0E",X"40",X"CD",X"1D",X"04",X"C9",X"2E",X"00",X"06",
		X"0E",X"7D",X"FE",X"0B",X"1A",X"13",X"38",X"06",X"CD",X"C8",X"06",X"BC",X"28",X"04",X"67",X"CD",
		X"B9",X"06",X"2C",X"10",X"EC",X"C9",X"21",X"3F",X"81",X"1E",X"06",X"0A",X"77",X"23",X"03",X"1D",
		X"20",X"F9",X"C3",X"6F",X"03",X"DD",X"21",X"2A",X"81",X"21",X"23",X"81",X"18",X"07",X"DD",X"21",
		X"38",X"81",X"21",X"31",X"81",X"CD",X"73",X"04",X"28",X"04",X"DD",X"CB",X"00",X"86",X"CD",X"73",
		X"04",X"28",X"04",X"DD",X"CB",X"00",X"8E",X"CD",X"73",X"04",X"28",X"04",X"DD",X"CB",X"00",X"96",
		X"C3",X"6F",X"03",X"EB",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"EB",X"73",X"23",X"72",X"23",X"7A",
		X"B3",X"C9",X"21",X"29",X"81",X"18",X"03",X"21",X"37",X"81",X"0A",X"03",X"77",X"23",X"0A",X"03",
		X"CB",X"47",X"28",X"02",X"CB",X"9E",X"CB",X"4F",X"28",X"02",X"CB",X"A6",X"CB",X"57",X"28",X"02",
		X"CB",X"AE",X"C3",X"6F",X"03",X"21",X"2B",X"81",X"18",X"03",X"21",X"39",X"81",X"16",X"03",X"0A",
		X"77",X"03",X"23",X"15",X"20",X"F9",X"C3",X"6F",X"03",X"21",X"2E",X"81",X"18",X"03",X"21",X"3C",
		X"81",X"EB",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"EB",X"73",X"23",X"72",X"23",X"0A",X"03",X"77",
		X"C3",X"6F",X"03",X"AF",X"32",X"00",X"81",X"01",X"00",X"00",X"ED",X"4B",X"01",X"81",X"78",X"B1",
		X"C2",X"6F",X"03",X"18",X"F5",X"C5",X"CD",X"E0",X"03",X"CD",X"0C",X"04",X"3E",X"13",X"3D",X"20",
		X"FD",X"C1",X"C3",X"6F",X"03",X"C5",X"CD",X"0C",X"04",X"CD",X"E0",X"03",X"3E",X"CF",X"3D",X"20",
		X"FD",X"C1",X"C3",X"6F",X"03",X"0A",X"03",X"6F",X"87",X"9F",X"67",X"09",X"44",X"4D",X"C3",X"6F",
		X"03",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"35",X"20",X"EB",X"03",X"C3",X"6F",X"03",X"0A",X"03",
		X"6F",X"0A",X"03",X"67",X"5E",X"C3",X"37",X"05",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"23",
		X"56",X"C3",X"47",X"05",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"73",X"C3",X"6F",
		X"03",X"0A",X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"73",X"23",X"72",
		X"C3",X"6F",X"03",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"C3",X"6C",X"05",X"0A",X"03",X"6F",
		X"0A",X"03",X"67",X"5E",X"23",X"56",X"C3",X"7E",X"05",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",
		X"03",X"67",X"7E",X"83",X"77",X"C3",X"6F",X"03",X"0A",X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",
		X"6F",X"0A",X"03",X"67",X"E5",X"7E",X"23",X"66",X"6F",X"19",X"EB",X"E1",X"73",X"23",X"72",X"C3",
		X"6F",X"03",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"CB",X"2E",X"1D",X"20",X"FB",
		X"C3",X"6F",X"03",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"23",X"CB",X"2E",X"2B",
		X"CB",X"1E",X"23",X"1D",X"20",X"F7",X"C3",X"6F",X"03",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",
		X"03",X"67",X"0A",X"77",X"23",X"03",X"1D",X"C2",X"C2",X"05",X"C3",X"6F",X"03",X"0A",X"03",X"87",
		X"C3",X"BB",X"05",X"CD",X"70",X"06",X"CD",X"51",X"06",X"01",X"70",X"00",X"AF",X"32",X"00",X"81",
		X"C3",X"6F",X"03",X"CD",X"70",X"06",X"CD",X"51",X"06",X"01",X"00",X"00",X"AF",X"32",X"00",X"81",
		X"C3",X"6F",X"03",X"0A",X"03",X"57",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"7E",
		X"B2",X"A3",X"77",X"C3",X"6F",X"03",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"7E",
		X"B3",X"77",X"C3",X"6F",X"03",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"35",X"20",X"09",X"23",X"7E",
		X"B7",X"20",X"03",X"C3",X"6F",X"03",X"35",X"0B",X"0B",X"0B",X"C5",X"CD",X"E0",X"03",X"CD",X"0C",
		X"04",X"3E",X"13",X"3D",X"20",X"FD",X"C1",X"C3",X"6F",X"03",X"0A",X"03",X"6F",X"0A",X"03",X"67",
		X"C5",X"44",X"4D",X"C3",X"6F",X"03",X"C1",X"C3",X"6F",X"03",X"DD",X"36",X"02",X"00",X"C3",X"6F",
		X"03",X"C5",X"21",X"23",X"81",X"06",X"0E",X"AF",X"77",X"23",X"10",X"FC",X"21",X"31",X"81",X"06",
		X"0E",X"AF",X"77",X"23",X"10",X"FC",X"3E",X"3F",X"32",X"2A",X"81",X"32",X"38",X"81",X"C1",X"C9",
		X"CD",X"8C",X"06",X"0E",X"10",X"2E",X"08",X"26",X"00",X"CD",X"B9",X"06",X"2E",X"09",X"26",X"00",
		X"CD",X"B9",X"06",X"2E",X"0A",X"26",X"00",X"CD",X"B9",X"06",X"18",X"17",X"0E",X"40",X"2E",X"08",
		X"26",X"00",X"CD",X"B9",X"06",X"2E",X"09",X"26",X"00",X"CD",X"B9",X"06",X"2E",X"0A",X"26",X"00",
		X"CD",X"B9",X"06",X"06",X"0D",X"ED",X"41",X"CB",X"21",X"16",X"00",X"78",X"FE",X"07",X"20",X"02",
		X"16",X"3F",X"ED",X"51",X"CB",X"39",X"10",X"ED",X"C9",X"ED",X"69",X"CB",X"21",X"ED",X"61",X"CB",
		X"39",X"C9",X"0E",X"10",X"18",X"02",X"0E",X"40",X"ED",X"69",X"CB",X"21",X"ED",X"60",X"CB",X"39",
		X"C9",X"F5",X"C5",X"D5",X"E5",X"CD",X"0A",X"07",X"6C",X"7D",X"FE",X"1F",X"38",X"02",X"2E",X"00",
		X"26",X"00",X"54",X"5D",X"19",X"19",X"11",X"40",X"00",X"19",X"EB",X"1A",X"21",X"00",X"81",X"BE",
		X"30",X"03",X"C3",X"02",X"07",X"32",X"00",X"81",X"13",X"1A",X"32",X"01",X"81",X"13",X"1A",X"32",
		X"02",X"81",X"E1",X"D1",X"C1",X"F1",X"ED",X"56",X"FB",X"C9",X"3E",X"0E",X"D3",X"40",X"DB",X"80",
		X"67",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
