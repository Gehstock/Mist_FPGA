library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"A3",X"80",X"A1",X"15",X"0F",X"EE",X"A6",X"A8",X"8F",X"A7",X"7D",X"D7",X"A2",X"7D",X"F6",X"8C",
		X"D6",X"8B",X"20",X"8C",X"DD",X"63",X"2A",X"6E",X"CD",X"23",X"B1",X"75",X"34",X"AB",X"C9",X"86",
		X"A1",X"30",X"79",X"7D",X"6B",X"A9",X"E6",X"6C",X"06",X"C8",X"6D",X"97",X"E0",X"69",X"7D",X"96",
		X"AA",X"89",X"DD",X"9E",X"A9",X"AF",X"C9",X"1A",X"24",X"28",X"07",X"E0",X"DD",X"5E",X"AA",X"1D",
		X"A0",X"8C",X"7D",X"D7",X"22",X"69",X"7D",X"96",X"21",X"88",X"7D",X"94",X"23",X"69",X"7D",X"96",
		X"BF",X"8A",X"C9",X"75",X"F6",X"AB",X"39",X"FC",X"68",X"E3",X"8F",X"A5",X"D2",X"B7",X"E6",X"C8",
		X"37",X"C8",X"46",X"C8",X"5A",X"B7",X"46",X"C8",X"37",X"C8",X"46",X"C8",X"66",X"C8",X"7D",X"6B",
		X"A9",X"CE",X"CC",X"F1",X"68",X"65",X"0A",X"C8",X"C9",X"75",X"36",X"AA",X"2A",X"75",X"36",X"A9",
		X"27",X"69",X"B2",X"84",X"28",X"CE",X"37",X"E8",X"7D",X"56",X"22",X"15",X"A0",X"8C",X"7D",X"D7",
		X"AA",X"61",X"DD",X"9E",X"A9",X"88",X"DD",X"9C",X"AB",X"61",X"DD",X"5E",X"AB",X"91",X"03",X"C8",
		X"4B",X"2F",X"05",X"15",X"E0",X"E6",X"E0",X"34",X"E0",X"E6",X"E0",X"15",X"E0",X"E6",X"E0",X"34",
		X"68",X"E6",X"68",X"4E",X"68",X"65",X"5A",X"C8",X"CD",X"72",X"B7",X"61",X"CD",X"6E",X"68",X"65",
		X"37",X"C8",X"6D",X"C7",X"E1",X"69",X"6D",X"E2",X"06",X"7D",X"96",X"BF",X"A2",X"69",X"8E",X"89",
		X"B8",X"8A",X"2E",X"88",X"DD",X"5E",X"2C",X"A7",X"08",X"87",X"2F",X"87",X"3E",X"88",X"FF",X"89",
		X"87",X"C9",X"B9",X"66",X"83",X"E6",X"83",X"F6",X"83",X"76",X"83",X"56",X"7D",X"D7",X"B0",X"FD",
		X"CD",X"E7",X"A1",X"F1",X"5D",X"75",X"CB",X"98",X"7E",X"08",X"29",X"14",X"73",X"F1",X"CD",X"B8",
		X"E1",X"5D",X"65",X"C7",X"01",X"59",X"7D",X"DD",X"63",X"18",X"F6",X"20",X"A1",X"BC",X"DB",X"59",
		X"CD",X"18",X"69",X"3D",X"3D",X"20",X"D8",X"C9",X"DD",X"CB",X"38",X"46",X"A0",X"01",X"AC",X"DD",
		X"63",X"18",X"66",X"A0",X"A1",X"2C",X"61",X"08",X"A1",X"14",X"B4",X"09",X"A0",X"08",X"A0",X"08",
		X"29",X"1C",X"3C",X"05",X"28",X"00",X"28",X"00",X"20",X"1C",X"3C",X"01",X"28",X"00",X"28",X"00",
		X"80",X"14",X"B4",X"0D",X"A0",X"08",X"A0",X"08",X"A1",X"88",X"B2",X"0A",X"A0",X"08",X"A0",X"08",
		X"29",X"20",X"3A",X"06",X"28",X"00",X"28",X"1B",X"29",X"20",X"3A",X"02",X"28",X"00",X"28",X"1B",
		X"A1",X"88",X"B2",X"0E",X"A0",X"08",X"A0",X"DD",X"89",X"08",X"2D",X"CD",X"AC",X"49",X"75",X"21",
		X"20",X"8D",X"CD",X"84",X"69",X"DD",X"21",X"40",X"8D",X"CD",X"0C",X"41",X"DD",X"21",X"60",X"8D",
		X"65",X"2C",X"E1",X"C9",X"75",X"EE",X"A0",X"DD",X"4E",X"09",X"75",X"F6",X"37",X"07",X"60",X"D6",
		X"2A",X"48",X"B2",X"84",X"8D",X"39",X"9B",X"41",X"4B",X"8F",X"A5",X"A3",X"69",X"AC",X"69",X"B2",
		X"E1",X"B0",X"E1",X"B6",X"B0",X"90",X"68",X"DD",X"9E",X"17",X"A3",X"C9",X"96",X"F8",X"B0",X"48",
		X"B8",X"F5",X"B6",X"18",X"91",X"48",X"B8",X"EF",X"B6",X"D8",X"91",X"48",X"B8",X"E9",X"DD",X"21",
		X"88",X"25",X"19",X"63",X"E1",X"DD",X"D6",X"17",X"6B",X"27",X"05",X"50",X"93",X"71",X"E1",X"B5",
		X"6B",X"E9",X"6C",X"29",X"6D",X"59",X"33",X"68",X"33",X"DD",X"45",X"D5",X"41",X"DD",X"21",X"80",
		X"2D",X"CD",X"50",X"96",X"F5",X"36",X"30",X"08",X"F5",X"36",X"31",X"08",X"75",X"F6",X"A4",X"39",
		X"BA",X"43",X"CD",X"8F",X"A5",X"20",X"75",X"CD",X"F0",X"43",X"DD",X"F6",X"2C",X"39",X"01",X"43",
		X"6D",X"2F",X"05",X"00",X"22",X"5E",X"D0",X"7A",X"BC",X"CA",X"76",X"08",X"5A",X"1C",X"E2",X"6D",
		X"F0",X"CB",X"CD",X"21",X"6B",X"7D",X"CB",X"B8",X"66",X"E4",X"D1",X"CA",X"CD",X"FE",X"6A",X"65",
		X"50",X"CB",X"F0",X"A7",X"8F",X"A7",X"CF",X"51",X"4E",X"8A",X"8F",X"A7",X"8F",X"67",X"7D",X"56",
		X"2C",X"7D",X"45",X"75",X"41",X"75",X"77",X"8C",X"DD",X"D9",X"28",X"75",X"70",X"89",X"CD",X"7B",
		X"E3",X"7D",X"96",X"AF",X"A0",X"16",X"D0",X"7D",X"6B",X"B8",X"C6",X"00",X"A2",X"16",X"D4",X"7D",
		X"77",X"8A",X"CD",X"23",X"B1",X"75",X"34",X"BF",X"2E",X"8D",X"CD",X"27",X"B8",X"61",X"CD",X"67",
		X"E2",X"F8",X"B2",X"48",X"2D",X"B8",X"6B",X"5F",X"75",X"D7",X"31",X"69",X"B6",X"98",X"36",X"00",
		X"39",X"1C",X"96",X"08",X"AD",X"75",X"36",X"BF",X"2A",X"7D",X"45",X"75",X"41",X"75",X"36",X"BF",
		X"A0",X"69",X"7D",X"96",X"37",X"8D",X"75",X"CD",X"7D",X"C9",X"7D",X"96",X"37",X"88",X"8E",X"8B",
		X"CD",X"27",X"B8",X"61",X"DD",X"9E",X"BF",X"8C",X"D5",X"63",X"B8",X"C6",X"A0",X"8D",X"D5",X"9E",
		X"37",X"88",X"69",X"6D",X"50",X"CB",X"75",X"CD",X"7D",X"C9",X"7D",X"96",X"37",X"88",X"4D",X"A6",
		X"2A",X"65",X"87",X"B8",X"49",X"65",X"4E",X"CA",X"CB",X"6E",X"CB",X"DE",X"C8",X"89",X"98",X"2D",
		X"95",X"81",X"7D",X"2D",X"95",X"69",X"81",X"48",X"2C",X"B6",X"A5",X"6B",X"F6",X"00",X"22",X"83",
		X"23",X"8B",X"23",X"8B",X"23",X"95",X"20",X"53",X"C9",X"9E",X"08",X"ED",X"23",X"9E",X"A9",X"8B",
		X"D1",X"83",X"D0",X"83",X"83",X"96",X"A1",X"6D",X"4F",X"CA",X"41",X"F8",X"96",X"48",X"69",X"6D",
		X"AA",X"90",X"58",X"2F",X"77",X"8B",X"77",X"9F",X"C9",X"C8",X"E1",X"6D",X"FB",X"10",X"8D",X"65",
		X"39",X"85",X"60",X"D5",X"9C",X"10",X"E5",X"FB",X"9A",X"25",X"65",X"31",X"05",X"C8",X"F5",X"34",
		X"B8",X"C5",X"FB",X"B4",X"8D",X"CD",X"99",X"2D",X"C8",X"C9",X"22",X"43",X"37",X"43",X"ED",X"43",
		X"C2",X"4B",X"0D",X"CD",X"47",X"81",X"96",X"12",X"B6",X"C8",X"F5",X"CB",X"30",X"EE",X"96",X"16",
		X"96",X"C8",X"D5",X"CB",X"B8",X"A6",X"C9",X"2C",X"2C",X"CD",X"E7",X"29",X"B6",X"18",X"96",X"C8",
		X"F5",X"CB",X"30",X"EE",X"96",X"14",X"B6",X"C8",X"F5",X"CB",X"30",X"AE",X"61",X"AD",X"65",X"C7",
		X"A1",X"B6",X"B9",X"96",X"C8",X"D5",X"CB",X"18",X"46",X"B6",X"BD",X"96",X"C8",X"D5",X"CB",X"18",
		X"8E",X"C9",X"04",X"AC",X"65",X"C7",X"01",X"B6",X"30",X"96",X"60",X"D5",X"63",X"10",X"CE",X"B6",
		X"BC",X"96",X"C8",X"D5",X"CB",X"18",X"06",X"C9",X"CD",X"78",X"B6",X"DD",X"F6",X"04",X"39",X"85",
		X"E3",X"CD",X"2F",X"85",X"61",X"25",X"E3",X"3A",X"E3",X"3F",X"E3",X"34",X"E3",X"F0",X"7E",X"0A",
		X"6F",X"C9",X"F0",X"4E",X"2A",X"6F",X"C9",X"F1",X"5E",X"02",X"EF",X"C9",X"F1",X"4E",X"2A",X"EF",
		X"61",X"07",X"11",X"1F",X"11",X"13",X"11",X"16",X"11",X"C5",X"4B",X"08",X"28",X"CD",X"A0",X"81",
		X"CD",X"00",X"A1",X"CD",X"BE",X"29",X"CD",X"00",X"A1",X"CD",X"28",X"29",X"C9",X"DD",X"34",X"07",
		X"75",X"F6",X"A7",X"DD",X"B6",X"0E",X"70",X"DD",X"9E",X"0F",X"A0",X"CD",X"CD",X"4B",X"89",X"73",
		X"6B",X"45",X"DD",X"F6",X"2C",X"39",X"4E",X"33",X"4B",X"8F",X"A5",X"DD",X"F6",X"05",X"DD",X"45",
		X"E9",X"CD",X"F4",X"99",X"61",X"DD",X"D6",X"08",X"EE",X"07",X"F6",X"00",X"68",X"DD",X"D6",X"09",
		X"46",X"0F",X"48",X"CD",X"31",X"44",X"CD",X"78",X"B6",X"DD",X"F6",X"04",X"39",X"85",X"6B",X"CD",
		X"2F",X"A5",X"7D",X"56",X"A4",X"B1",X"89",X"CB",X"6D",X"2F",X"05",X"68",X"76",X"D0",X"B0",X"8B",
		X"D6",X"08",X"D8",X"75",X"34",X"BF",X"CD",X"F0",X"B6",X"75",X"F6",X"8C",X"39",X"0D",X"6B",X"65",
		X"2F",X"A5",X"B6",X"88",X"92",X"8A",X"28",X"4D",X"CB",X"88",X"28",X"16",X"34",X"6D",X"A0",X"A7",
		X"C9",X"7D",X"21",X"88",X"8D",X"65",X"EE",X"CC",X"D5",X"89",X"20",X"2D",X"CD",X"EE",X"6C",X"7D",
		X"81",X"C8",X"2D",X"6D",X"66",X"CC",X"75",X"81",X"C0",X"2D",X"6D",X"EE",X"E4",X"69",X"75",X"56",
		X"BF",X"AF",X"C8",X"7E",X"2E",X"F0",X"DD",X"5E",X"2C",X"91",X"FF",X"CC",X"4B",X"2F",X"A5",X"C7",
		X"E4",X"2E",X"E4",X"20",X"E4",X"6F",X"E4",X"6D",X"50",X"B6",X"D8",X"71",X"6D",X"2F",X"16",X"52",
		X"90",X"08",X"AC",X"1C",X"90",X"08",X"A8",X"1D",X"B5",X"38",X"A0",X"8B",X"B5",X"38",X"48",X"5B",
		X"31",X"00",X"A3",X"15",X"31",X"E8",X"7D",X"94",X"27",X"5D",X"96",X"BF",X"21",X"69",X"6D",X"F0",
		X"B6",X"D0",X"F9",X"65",X"8F",X"B6",X"F2",X"38",X"A0",X"45",X"B5",X"38",X"A0",X"41",X"B4",X"1C",
		X"30",X"00",X"7C",X"14",X"30",X"00",X"78",X"69",X"6D",X"F0",X"16",X"F0",X"F9",X"6D",X"2F",X"B6",
		X"F3",X"39",X"A0",X"AC",X"B4",X"39",X"A0",X"A8",X"B5",X"1D",X"91",X"08",X"2B",X"1D",X"91",X"E0",
		X"F2",X"18",X"A0",X"8B",X"B5",X"18",X"48",X"7D",X"94",X"AF",X"75",X"96",X"37",X"A9",X"69",X"6D",
		X"F0",X"B6",X"78",X"51",X"CD",X"2F",X"B6",X"5B",X"91",X"08",X"45",X"1D",X"91",X"08",X"41",X"1C",
		X"B4",X"19",X"A0",X"7C",X"B4",X"19",X"A0",X"78",X"69",X"6D",X"0D",X"B2",X"75",X"81",X"A0",X"2D",
		X"D5",X"5E",X"BF",X"7E",X"AA",X"88",X"2C",X"7D",X"36",X"A8",X"28",X"7D",X"21",X"80",X"8D",X"7D",
		X"D6",X"17",X"F6",X"02",X"88",X"0C",X"F5",X"36",X"20",X"08",X"F5",X"21",X"E0",X"25",X"F5",X"F6",
		X"BF",X"D6",X"AA",X"20",X"2C",X"D5",X"36",X"08",X"28",X"D5",X"21",X"60",X"8D",X"D5",X"F6",X"1F",
		X"F6",X"02",X"88",X"0C",X"F5",X"36",X"20",X"08",X"61",X"CD",X"50",X"96",X"E5",X"6B",X"A0",X"20",
		X"DD",X"CB",X"B8",X"66",X"4A",X"BC",X"6D",X"DD",X"F6",X"19",X"CB",X"F7",X"A0",X"11",X"46",X"7F",
		X"2F",X"3E",X"A0",X"FF",X"89",X"6A",X"2D",X"B9",X"D9",X"23",X"D8",X"DD",X"9E",X"11",X"A0",X"B6",
		X"A9",X"32",X"2A",X"88",X"CD",X"FE",X"A6",X"DD",X"34",X"1F",X"2E",X"04",X"CD",X"AF",X"B8",X"DD",
		X"D6",X"07",X"AF",X"C8",X"0E",X"0D",X"65",X"6F",X"30",X"39",X"80",X"08",X"96",X"02",X"F5",X"21",
		X"28",X"8D",X"D5",X"96",X"BF",X"A0",X"38",X"D5",X"B9",X"D5",X"96",X"1F",X"A0",X"09",X"D5",X"B9",
		X"F5",X"96",X"37",X"A0",X"A2",X"D5",X"11",X"DD",X"4E",X"07",X"F5",X"70",X"32",X"D5",X"9C",X"17",
		X"D5",X"21",X"20",X"8D",X"D5",X"96",X"BF",X"20",X"2F",X"D5",X"36",X"1A",X"28",X"D5",X"34",X"1F",
		X"F5",X"B9",X"F5",X"96",X"37",X"20",X"A7",X"D5",X"9E",X"12",X"A0",X"D5",X"9C",X"17",X"F5",X"B9",
		X"D5",X"96",X"BF",X"48",X"D5",X"36",X"BA",X"00",X"D5",X"34",X"BF",X"C9",X"DD",X"F6",X"B8",X"46",
		X"27",X"0F",X"1E",X"08",X"57",X"21",X"98",X"25",X"11",X"71",X"8B",X"70",X"96",X"01",X"9A",X"0A",
		X"88",X"CD",X"81",X"2F",X"DD",X"36",X"28",X"00",X"DD",X"36",X"29",X"00",X"CD",X"CE",X"33",X"DD",
		X"9C",X"17",X"65",X"E3",X"E5",X"CD",X"62",X"4E",X"6B",X"52",X"E5",X"DD",X"63",X"1E",X"56",X"48",
		X"C5",X"EB",X"10",X"8D",X"CD",X"D8",X"EB",X"C5",X"EB",X"B2",X"8D",X"CD",X"D8",X"4B",X"C5",X"EB",
		X"9C",X"2D",X"6D",X"78",X"63",X"7D",X"96",X"9F",X"A0",X"6D",X"B2",X"CE",X"48",X"7D",X"96",X"9F",
		X"D7",X"61",X"C5",X"43",X"10",X"2D",X"C5",X"53",X"12",X"2D",X"CD",X"A2",X"6E",X"60",X"C5",X"53",
		X"9C",X"2D",X"6D",X"A2",X"E6",X"68",X"65",X"63",X"9A",X"2D",X"86",X"88",X"F0",X"EE",X"A2",X"BA",
		X"D8",X"7E",X"2D",X"F0",X"5E",X"8A",X"A0",X"89",X"24",X"59",X"4E",X"8A",X"1B",X"70",X"D6",X"8D",
		X"58",X"FE",X"A2",X"00",X"A1",X"84",X"B6",X"89",X"1C",X"69",X"7D",X"6B",X"B6",X"F6",X"48",X"6D",
		X"1E",X"E8",X"A0",X"8C",X"CD",X"C3",X"E8",X"E0",X"DD",X"9E",X"3F",X"88",X"2E",X"8B",X"CD",X"29",
		X"30",X"36",X"81",X"6D",X"52",X"A6",X"8E",X"C8",X"4D",X"50",X"46",X"8B",X"99",X"3E",X"E7",X"6D",
		X"8F",X"A5",X"B6",X"8A",X"CD",X"59",X"A0",X"E1",X"4D",X"58",X"B5",X"EE",X"2F",X"1C",X"CD",X"76",
		X"E7",X"E9",X"4D",X"60",X"6D",X"9F",X"60",X"16",X"A2",X"6D",X"F9",X"A0",X"49",X"B0",X"79",X"6D",
		X"17",X"91",X"CD",X"38",X"AF",X"89",X"E4",X"CF",X"CD",X"A6",X"AF",X"89",X"F1",X"CF",X"DD",X"63",
		X"B6",X"F6",X"A0",X"8B",X"81",X"28",X"E7",X"6D",X"DC",X"A1",X"81",X"D1",X"E7",X"6D",X"DC",X"A1",
		X"21",X"09",X"6F",X"65",X"54",X"A1",X"B6",X"A2",X"CD",X"59",X"A0",X"86",X"2F",X"65",X"4F",X"B8",
		X"8E",X"C4",X"81",X"60",X"A3",X"7D",X"6B",X"9E",X"56",X"00",X"A5",X"A6",X"92",X"81",X"DC",X"89",
		X"4D",X"ED",X"F0",X"EE",X"2B",X"64",X"EF",X"CF",X"39",X"AA",X"28",X"65",X"87",X"A0",X"41",X"91",
		X"22",X"88",X"27",X"4D",X"DA",X"CD",X"6D",X"C8",X"03",X"86",X"B2",X"06",X"22",X"82",X"A0",X"28",
		X"CD",X"DC",X"A4",X"1E",X"2A",X"65",X"59",X"A0",X"41",X"E1",X"4D",X"ED",X"E8",X"65",X"3F",X"E8",
		X"E9",X"49",X"18",X"64",X"0E",X"F7",X"65",X"6F",X"30",X"2E",X"20",X"CD",X"EF",X"10",X"96",X"48",
		X"CD",X"D1",X"A0",X"CD",X"92",X"0F",X"DD",X"36",X"3E",X"FF",X"B6",X"09",X"CD",X"FE",X"6F",X"CD",
		X"42",X"86",X"75",X"45",X"75",X"21",X"A0",X"25",X"65",X"38",X"E7",X"DD",X"89",X"88",X"2D",X"CD",
		X"18",X"47",X"DD",X"21",X"68",X"8D",X"CD",X"90",X"6F",X"DD",X"21",X"60",X"8D",X"CD",X"18",X"47",
		X"75",X"21",X"A8",X"25",X"65",X"66",X"93",X"B6",X"80",X"CD",X"F9",X"80",X"75",X"41",X"61",X"CB",
		X"78",X"A0",X"3C",X"4D",X"AE",X"24",X"B6",X"0B",X"32",X"02",X"88",X"CD",X"9E",X"28",X"B5",X"A0",
		X"A4",X"6F",X"65",X"8E",X"05",X"49",X"61",X"4D",X"06",X"80",X"10",X"E2",X"21",X"18",X"B0",X"02",
		X"2D",X"0A",X"39",X"18",X"6A",X"4F",X"EE",X"55",X"5B",X"0B",X"3A",X"10",X"31",X"30",X"30",X"30",
		X"98",X"06",X"B3",X"11",X"F0",X"5C",X"F3",X"B2",X"23",X"1A",X"B0",X"88",X"95",X"98",X"90",X"B8",
		X"CD",X"CE",X"33",X"B6",X"2A",X"DD",X"96",X"1F",X"48",X"DD",X"36",X"1F",X"2B",X"C9",X"5A",X"47",
		X"48",X"4F",X"8E",X"4F",X"1C",X"4F",X"E5",X"EB",X"98",X"25",X"65",X"70",X"63",X"C5",X"43",X"BA",
		X"8D",X"CD",X"4A",X"4B",X"C5",X"EB",X"14",X"8D",X"CD",X"C2",X"EB",X"C9",X"C5",X"EB",X"10",X"8D",
		X"65",X"6A",X"63",X"C5",X"43",X"BA",X"2D",X"CD",X"78",X"43",X"E5",X"EB",X"9C",X"25",X"65",X"6A",
		X"EB",X"C9",X"C5",X"EB",X"10",X"8D",X"CD",X"C2",X"EB",X"C5",X"EB",X"B2",X"8D",X"CD",X"4A",X"4B",
		X"E5",X"EB",X"9C",X"25",X"65",X"70",X"63",X"C9",X"E5",X"EB",X"98",X"25",X"65",X"70",X"63",X"C5",
		X"EB",X"B2",X"8D",X"CD",X"D8",X"4B",X"C5",X"EB",X"14",X"8D",X"CD",X"D8",X"EB",X"C9",X"21",X"62",
		X"AC",X"B1",X"C3",X"0C",X"8E",X"BA",X"4D",X"A1",X"35",X"88",X"D7",X"4D",X"10",X"83",X"83",X"83",
		X"3B",X"93",X"3B",X"E1",X"38",X"50",X"C9",X"89",X"01",X"0F",X"39",X"80",X"28",X"86",X"AE",X"59",
		X"46",X"8F",X"4E",X"9E",X"D7",X"8F",X"65",X"F2",X"D7",X"8F",X"65",X"F2",X"AC",X"B0",X"D8",X"81",
		X"6A",X"0C",X"2E",X"AF",X"F1",X"EE",X"2F",X"E6",X"3E",X"DF",X"23",X"DF",X"23",X"04",X"38",X"54",
		X"81",X"8A",X"AC",X"A6",X"26",X"51",X"46",X"8F",X"4E",X"9E",X"D7",X"83",X"D7",X"83",X"AC",X"B0",
		X"54",X"89",X"97",X"0F",X"2E",X"AF",X"F1",X"EE",X"2F",X"E6",X"3E",X"DF",X"A3",X"DF",X"A3",X"04",
		X"98",X"54",X"69",X"81",X"98",X"2D",X"F6",X"83",X"83",X"1E",X"48",X"83",X"83",X"1E",X"48",X"6D",
		X"58",X"E8",X"21",X"11",X"8D",X"91",X"2A",X"88",X"F6",X"11",X"B5",X"1D",X"96",X"E0",X"B9",X"1D",
		X"B5",X"1E",X"48",X"12",X"98",X"2D",X"76",X"89",X"A0",X"8E",X"76",X"B9",X"A0",X"8A",X"27",X"69",
		X"DD",X"9E",X"3E",X"77",X"87",X"61",X"21",X"11",X"8D",X"5E",X"23",X"8B",X"96",X"E0",X"23",X"8B",
		X"36",X"E8",X"6D",X"4B",X"60",X"81",X"98",X"2D",X"99",X"8A",X"A0",X"56",X"B9",X"15",X"B5",X"1E",
		X"48",X"11",X"B5",X"1D",X"96",X"E0",X"B2",X"11",X"8D",X"7E",X"2A",X"08",X"5B",X"7E",X"BE",X"08",
		X"6F",X"0F",X"69",X"81",X"98",X"2D",X"8E",X"8A",X"4D",X"6D",X"7D",X"E8",X"49",X"B0",X"59",X"69",
		X"21",X"10",X"8D",X"86",X"2A",X"E5",X"CD",X"73",X"E8",X"E1",X"38",X"71",X"C9",X"ED",X"FE",X"8B",
		X"DE",X"83",X"F3",X"1E",X"B0",X"AA",X"83",X"83",X"98",X"71",X"41",X"D3",X"83",X"D2",X"83",X"69",
		X"F6",X"DB",X"FF",X"8B",X"F6",X"DA",X"7F",X"8B",X"F3",X"10",X"C5",X"ED",X"FE",X"8B",X"7E",X"8B",
		X"D2",X"23",X"B6",X"B0",X"21",X"23",X"18",X"F1",X"E9",X"73",X"8B",X"72",X"8B",X"C9",X"83",X"F6",
		X"73",X"FF",X"23",X"F6",X"72",X"7F",X"23",X"B8",X"C5",X"DD",X"21",X"C0",X"8C",X"2E",X"2D",X"4D",
		X"75",X"CB",X"A0",X"D6",X"6C",X"98",X"61",X"39",X"A6",X"08",X"75",X"B9",X"69",X"38",X"D8",X"C9",
		X"DD",X"F6",X"2D",X"39",X"B1",X"49",X"4B",X"8F",X"A5",X"58",X"33",X"4D",X"E9",X"67",X"E9",X"72",
		X"61",X"1F",X"62",X"8A",X"62",X"DF",X"62",X"2A",X"62",X"6E",X"62",X"ED",X"62",X"DD",X"63",X"08",
		X"76",X"A0",X"AD",X"21",X"49",X"8D",X"F6",X"DD",X"77",X"04",X"35",X"2E",X"2C",X"CD",X"4F",X"18",
		X"75",X"34",X"A5",X"21",X"77",X"24",X"9D",X"DD",X"D6",X"08",X"FE",X"0A",X"75",X"77",X"A0",X"DD",
		X"34",X"05",X"B2",X"24",X"88",X"46",X"BF",X"48",X"DD",X"35",X"28",X"DD",X"F6",X"00",X"46",X"07",
		X"68",X"DD",X"D6",X"09",X"95",X"A0",X"E1",X"DD",X"DF",X"09",X"75",X"35",X"A5",X"6F",X"96",X"00",
		X"18",X"DD",X"CB",X"00",X"76",X"A0",X"2E",X"D6",X"2E",X"B0",X"2A",X"B6",X"A8",X"0F",X"0F",X"4E",
		X"C0",X"55",X"75",X"EE",X"A2",X"DD",X"4E",X"0B",X"E5",X"6B",X"A0",X"20",X"65",X"C7",X"01",X"B6",
		X"BC",X"96",X"A0",X"0A",X"B6",X"09",X"32",X"02",X"88",X"51",X"CD",X"00",X"A7",X"C9",X"51",X"DD",
		X"9E",X"08",X"A0",X"DD",X"9E",X"0D",X"A0",X"C9",X"75",X"CB",X"A0",X"DE",X"88",X"88",X"75",X"EE",
		X"2A",X"DD",X"6E",X"03",X"CD",X"A9",X"6B",X"DD",X"CB",X"00",X"E6",X"39",X"2B",X"00",X"DD",X"45",
		X"6C",X"A7",X"00",X"DD",X"E9",X"DD",X"9E",X"08",X"A0",X"DD",X"9E",X"0D",X"A0",X"C9",X"89",X"68",
		X"8D",X"F6",X"6F",X"B6",X"AC",X"18",X"CB",X"B7",X"4E",X"08",X"EF",X"DD",X"F6",X"04",X"18",X"C5",
		X"CC",X"A9",X"86",X"88",X"E7",X"82",X"A0",X"28",X"7D",X"D4",X"A1",X"7D",X"D5",X"8C",X"B6",X"9F",
		X"CD",X"B4",X"A1",X"75",X"34",X"8D",X"C9",X"75",X"F6",X"88",X"56",X"AF",X"DD",X"DF",X"28",X"75",
		X"94",X"8D",X"B2",X"84",X"28",X"CE",X"27",X"E8",X"7D",X"E6",X"A3",X"7D",X"EE",X"8A",X"7D",X"6B",
		X"28",X"CE",X"A0",X"8F",X"B6",X"98",X"CD",X"4C",X"EB",X"10",X"2D",X"1E",X"AC",X"65",X"4C",X"EB",
		X"7D",X"95",X"A0",X"7D",X"F6",X"88",X"46",X"AF",X"48",X"7D",X"C6",X"89",X"7D",X"46",X"A4",X"82",
		X"28",X"28",X"B6",X"80",X"CD",X"B4",X"A1",X"75",X"CB",X"88",X"E6",X"88",X"3A",X"75",X"6E",X"8B",
		X"7D",X"66",X"A2",X"6D",X"09",X"CB",X"7D",X"96",X"A0",X"88",X"7D",X"96",X"A5",X"88",X"69",X"7D",
		X"34",X"8D",X"DD",X"9E",X"29",X"8D",X"C9",X"75",X"F6",X"88",X"56",X"8B",X"DD",X"DF",X"28",X"75",
		X"94",X"8D",X"B2",X"84",X"28",X"CE",X"37",X"E8",X"7D",X"95",X"A0",X"7D",X"F6",X"88",X"46",X"8F",
		X"48",X"75",X"F6",X"89",X"B5",X"08",X"A3",X"75",X"77",X"89",X"DD",X"9D",X"2D",X"C7",X"B6",X"8C",
		X"18",X"AF",X"0F",X"EE",X"A8",X"7D",X"EE",X"8A",X"7D",X"E6",X"A3",X"4D",X"CB",X"88",X"28",X"DD",
		X"B6",X"98",X"DD",X"63",X"29",X"CE",X"A0",X"8A",X"B6",X"AC",X"32",X"8A",X"88",X"F9",X"CD",X"88",
		X"07",X"69",X"7D",X"94",X"A5",X"69",X"7D",X"56",X"A0",X"DE",X"20",X"7D",X"D7",X"88",X"7D",X"94",
		X"2D",X"75",X"EE",X"8A",X"DD",X"C6",X"2B",X"6D",X"6B",X"88",X"88",X"1E",X"38",X"9A",X"2A",X"28",
		X"B6",X"38",X"6D",X"88",X"07",X"12",X"84",X"28",X"46",X"B7",X"48",X"7D",X"95",X"88",X"7D",X"56",
		X"28",X"EE",X"AF",X"E0",X"DD",X"46",X"2A",X"75",X"6E",X"8B",X"CD",X"21",X"6B",X"91",X"32",X"88",
		X"65",X"A7",X"00",X"DD",X"9E",X"08",X"A0",X"DD",X"9E",X"0D",X"A0",X"C9",X"75",X"21",X"88",X"25",
		X"DD",X"CB",X"3F",X"7E",X"C8",X"B2",X"24",X"88",X"6F",X"46",X"B7",X"48",X"CB",X"70",X"A0",X"06",
		X"96",X"01",X"65",X"84",X"63",X"C9",X"96",X"04",X"65",X"84",X"63",X"C9",X"75",X"EE",X"B0",X"DD",
		X"6E",X"11",X"CD",X"C4",X"EB",X"DD",X"EE",X"12",X"DD",X"6E",X"3B",X"CD",X"4C",X"4B",X"DD",X"EE",
		X"B4",X"DD",X"4E",X"1D",X"65",X"6C",X"63",X"C9",X"75",X"21",X"E8",X"25",X"75",X"CB",X"37",X"D6",
		X"C8",X"DD",X"CB",X"1F",X"66",X"CC",X"FC",X"4B",X"CD",X"69",X"EB",X"C9",X"DD",X"F6",X"BF",X"56",
		X"26",X"DD",X"DF",X"17",X"75",X"CB",X"37",X"EE",X"61",X"B2",X"84",X"20",X"EE",X"07",X"68",X"DD",
		X"35",X"1F",X"DD",X"F6",X"BF",X"46",X"AF",X"48",X"DD",X"CB",X"BF",X"A6",X"DD",X"F6",X"BE",X"B5",
		X"80",X"0F",X"75",X"77",X"36",X"CD",X"3B",X"43",X"61",X"DD",X"9E",X"17",X"A0",X"B2",X"9E",X"25",
		X"07",X"C8",X"DD",X"36",X"BF",X"80",X"DD",X"36",X"BE",X"08",X"C9",X"DD",X"6E",X"00",X"21",X"C2",
		X"2D",X"4D",X"ED",X"EE",X"8B",X"6E",X"D0",X"09",X"80",X"19",X"92",X"0B",X"2D",X"DD",X"63",X"16",
		X"6E",X"CC",X"4C",X"4B",X"DD",X"CB",X"BE",X"46",X"4C",X"D8",X"EB",X"41",X"49",X"23",X"23",X"38",
		X"C8",X"C9",X"96",X"04",X"65",X"74",X"63",X"77",X"04",X"CD",X"7C",X"43",X"DF",X"2C",X"65",X"74",
		X"EB",X"77",X"AD",X"CD",X"DC",X"4B",X"77",X"C9",X"B6",X"09",X"B8",X"E8",X"55",X"CD",X"E7",X"29",
		X"19",X"08",X"A4",X"B9",X"F9",X"C9",X"75",X"21",X"A8",X"25",X"75",X"F6",X"37",X"07",X"60",X"D6",
		X"2E",X"58",X"CD",X"78",X"B6",X"60",X"E1",X"DD",X"21",X"00",X"8D",X"CD",X"BC",X"4C",X"B0",X"2E",
		X"7D",X"81",X"80",X"2D",X"6D",X"BC",X"64",X"10",X"85",X"7D",X"81",X"C8",X"2D",X"6D",X"34",X"EC",
		X"B0",X"BC",X"DD",X"89",X"60",X"2D",X"CD",X"BC",X"EC",X"18",X"3B",X"61",X"DD",X"5E",X"BF",X"7E",
		X"A4",X"F8",X"6D",X"F0",X"16",X"F0",X"F9",X"6D",X"39",X"A5",X"97",X"68",X"B7",X"69",X"7D",X"81",
		X"08",X"2D",X"DD",X"9E",X"BF",X"88",X"DD",X"9E",X"BE",X"77",X"B6",X"BA",X"2F",X"87",X"DD",X"DF",
		X"A2",X"6D",X"0B",X"B1",X"6D",X"3E",X"00",X"15",X"68",X"E7",X"B6",X"AB",X"92",X"8A",X"28",X"26",
		X"A4",X"65",X"26",X"A5",X"C9",X"75",X"21",X"08",X"8D",X"75",X"F6",X"BF",X"07",X"60",X"D6",X"8E",
		X"58",X"6D",X"50",X"B6",X"C0",X"41",X"7D",X"81",X"A0",X"2D",X"6D",X"0B",X"64",X"7D",X"81",X"80",
		X"8D",X"65",X"0B",X"EC",X"DD",X"89",X"68",X"2D",X"CD",X"0B",X"EC",X"75",X"21",X"C0",X"8D",X"65",
		X"AB",X"EC",X"69",X"7D",X"F6",X"BF",X"76",X"8C",X"A0",X"8B",X"76",X"8D",X"48",X"6D",X"50",X"B6",
		X"78",X"51",X"CD",X"39",X"A5",X"E0",X"DD",X"9E",X"A9",X"88",X"DD",X"9E",X"BF",X"8E",X"C9",X"77",
		X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",
		X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",
		X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",
		X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",
		X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",X"5F",X"77",
		X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",X"D7",X"77",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"91",X"11",X"B0",X"92",X"B2",X"11",X"B2",X"91",X"80",X"62",X"C9",X"F0",X"C9",X"66",X"80",
		X"20",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"31",X"80",X"EA",X"C9",X"78",X"C9",X"EE",X"80",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"80",X"99",X"11",X"90",X"92",X"92",X"11",X"92",X"91",X"88",X"62",X"49",X"F0",X"49",X"66",X"88",
		X"20",X"31",X"B1",X"38",X"32",X"3A",X"B1",X"3A",X"31",X"20",X"EA",X"41",X"78",X"41",X"EE",X"20",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"4E",X"EF",X"42",X"7D",X"4F",X"20",X"4B",X"EF",X"44",X"6D",X"52",X"69",X"20",X"20",X"3A",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"66",X"67",X"6A",X"7D",X"67",X"A8",X"63",X"67",X"6C",X"6D",X"7A",X"69",X"A8",X"A8",X"B2",
		X"1A",X"EE",X"47",X"6A",X"D5",X"EF",X"88",X"EB",X"47",X"6C",X"C5",X"7A",X"C1",X"20",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"54",X"7B",X"55",X"7C",X"4F",X"ED",X"55",X"20",X"49",X"7F",X"41",X"EE",X"45",X"20",X"3A",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"7C",X"7B",X"7D",X"7C",X"67",X"65",X"7D",X"A8",X"61",X"7F",X"69",X"66",X"6D",X"A8",X"B2",
		X"1A",X"7C",X"D3",X"7D",X"D4",X"EF",X"45",X"7D",X"88",X"E9",X"D7",X"69",X"46",X"6D",X"88",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"41",X"EB",X"49",X"7A",X"41",X"20",X"4E",X"69",X"4B",X"69",X"4B",X"7D",X"4D",X"69",X"3A",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"69",X"63",X"61",X"7A",X"69",X"A8",X"66",X"69",X"63",X"69",X"63",X"7D",X"65",X"69",X"B2",
		X"1A",X"69",X"43",X"E9",X"D2",X"69",X"88",X"EE",X"C1",X"EB",X"C1",X"EB",X"D5",X"ED",X"C1",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"53",X"E8",X"49",X"EE",X"4A",X"E9",X"20",X"6D",X"47",X"E9",X"20",X"20",X"20",X"20",X"3A",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"B2",X"7B",X"60",X"61",X"66",X"62",X"61",X"A8",X"6D",X"6F",X"61",X"A8",X"A8",X"A8",X"A8",X"B2",
		X"1A",X"7B",X"40",X"E9",X"46",X"EA",X"41",X"20",X"C5",X"6F",X"41",X"20",X"88",X"20",X"88",X"B2",
		X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"8F",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",
		X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"A3",X"A0",X"B7",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"62",X"88",X"28",X"88",X"28",X"45",X"1A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"88",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"B2",X"A2",X"A0",X"B7",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"61",X"D0",X"28",X"88",X"28",X"0E",X"8F",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"06",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"A1",X"A0",X"B7",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"28",X"E7",X"28",X"88",X"28",X"E2",X"19",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"B1",X"A0",X"16",X"C8",X"67",X"88",X"A0",X"88",
		X"28",X"88",X"28",X"E6",X"28",X"88",X"28",X"E2",X"8A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"B0",X"87",X"15",X"C8",X"66",X"DD",X"F0",X"88",
		X"28",X"88",X"28",X"B7",X"28",X"88",X"28",X"E1",X"8A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",
		X"18",X"35",X"A2",X"8A",X"A2",X"8A",X"A2",X"41",X"27",X"86",X"A0",X"C8",X"65",X"DC",X"F0",X"88",
		X"28",X"88",X"28",X"E5",X"28",X"88",X"28",X"E2",X"8A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",
		X"A4",X"0C",X"EB",X"61",X"69",X"61",X"78",X"E8",X"26",X"8D",X"A0",X"49",X"64",X"5B",X"F0",X"08",
		X"28",X"00",X"28",X"6C",X"28",X"00",X"28",X"69",X"18",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",
		X"A4",X"0C",X"A4",X"0C",X"6D",X"7C",X"FF",X"77",X"CC",X"8C",X"A0",X"49",X"63",X"08",X"66",X"08",
		X"28",X"00",X"28",X"6C",X"74",X"00",X"28",X"85",X"8F",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"A5",
		X"9F",X"BF",X"9F",X"60",X"A1",X"09",X"EA",X"B4",X"25",X"08",X"A0",X"49",X"A0",X"08",X"66",X"08",
		X"28",X"00",X"28",X"6B",X"73",X"00",X"28",X"E5",X"8E",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"00",
		X"A1",X"09",X"A1",X"09",X"EA",X"B4",X"A3",X"64",X"24",X"8B",X"14",X"4D",X"62",X"08",X"66",X"08",
		X"28",X"00",X"28",X"6A",X"2A",X"00",X"28",X"84",X"8D",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"00",
		X"A1",X"09",X"EA",X"B4",X"A3",X"0B",X"6C",X"76",X"23",X"8A",X"13",X"4C",X"61",X"08",X"64",X"08",
		X"28",X"00",X"28",X"69",X"2A",X"7A",X"28",X"83",X"8C",X"02",X"2A",X"02",X"2A",X"02",X"04",X"00",
		X"9E",X"B4",X"A3",X"0B",X"A3",X"64",X"FE",X"75",X"22",X"89",X"12",X"4B",X"60",X"08",X"F7",X"08",
		X"28",X"00",X"28",X"69",X"2A",X"79",X"28",X"01",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"03",X"00",
		X"A3",X"0B",X"A3",X"0B",X"6C",X"08",X"FD",X"7A",X"CB",X"88",X"11",X"4A",X"E7",X"08",X"F6",X"08",
		X"28",X"00",X"28",X"68",X"2A",X"78",X"28",X"82",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"02",X"00",
		X"A3",X"0B",X"E9",X"6F",X"A0",X"68",X"FB",X"09",X"CA",X"17",X"A0",X"49",X"E6",X"58",X"A0",X"08",
		X"28",X"5D",X"28",X"68",X"2A",X"02",X"F5",X"81",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"28",X"00",
		X"9D",X"33",X"A0",X"88",X"E8",X"8B",X"FA",X"59",X"7B",X"BE",X"10",X"C9",X"E6",X"EE",X"A0",X"88",
		X"28",X"FC",X"28",X"C7",X"72",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",X"28",X"88",
		X"A0",X"88",X"A0",X"48",X"A3",X"5B",X"A1",X"58",X"7A",X"BD",X"97",X"C9",X"A0",X"DA",X"A0",X"88",
		X"28",X"FC",X"28",X"C6",X"E1",X"D7",X"2A",X"8A",X"2A",X"8A",X"2A",X"3B",X"9D",X"01",X"28",X"88",
		X"A0",X"88",X"E8",X"8B",X"A3",X"5A",X"F9",X"8C",X"79",X"8A",X"96",X"C9",X"A0",X"D9",X"A0",X"88",
		X"28",X"C9",X"28",X"C5",X"71",X"D6",X"2A",X"8A",X"2A",X"8A",X"2A",X"3A",X"9C",X"00",X"28",X"88",
		X"9C",X"10",X"A3",X"8B",X"1A",X"89",X"F8",X"7C",X"A2",X"BC",X"95",X"C9",X"A0",X"EC",X"A0",X"88",
		X"28",X"FF",X"28",X"C4",X"28",X"D5",X"F4",X"8A",X"2A",X"8A",X"2A",X"39",X"28",X"3F",X"28",X"88",
		X"A3",X"8B",X"A3",X"32",X"A1",X"59",X"A4",X"7B",X"A2",X"BB",X"94",X"C9",X"A0",X"EC",X"A0",X"88",
		X"28",X"FE",X"28",X"C4",X"28",X"88",X"F3",X"08",X"2A",X"8A",X"98",X"88",X"28",X"3E",X"28",X"88",
		X"A3",X"8B",X"1A",X"89",X"A1",X"58",X"A4",X"7A",X"21",X"BA",X"93",X"C9",X"A0",X"EC",X"A0",X"88",
		X"28",X"D8",X"28",X"FC",X"28",X"88",X"28",X"F7",X"8B",X"8A",X"3B",X"88",X"28",X"88",X"28",X"88",
		X"A3",X"32",X"A1",X"89",X"6B",X"8C",X"A4",X"79",X"20",X"B9",X"A0",X"C9",X"A0",X"EE",X"A0",X"88",
		X"FD",X"88",X"FD",X"C9",X"28",X"88",X"28",X"EC",X"8A",X"8A",X"3B",X"88",X"28",X"88",X"28",X"88",
		X"9B",X"89",X"A1",X"4E",X"6A",X"8C",X"6F",X"8A",X"A7",X"B8",X"92",X"C9",X"A0",X"EE",X"A0",X"88",
		X"FC",X"88",X"60",X"C3",X"28",X"88",X"28",X"E0",X"8A",X"8A",X"1F",X"88",X"28",X"88",X"28",X"88",
		X"A1",X"09",X"A1",X"6D",X"A4",X"0C",X"6E",X"0A",X"A2",X"1F",X"91",X"49",X"A0",X"58",X"A0",X"08",
		X"FB",X"00",X"28",X"00",X"28",X"00",X"28",X"7E",X"8A",X"02",X"1F",X"00",X"28",X"00",X"28",X"00",
		X"A1",X"09",X"1F",X"0C",X"A4",X"67",X"A2",X"0A",X"A6",X"08",X"90",X"48",X"A0",X"08",X"A0",X"08",
		X"FA",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"89",X"02",X"1E",X"00",X"28",X"00",X"28",X"00",
		X"08",X"A6",X"A4",X"0C",X"A4",X"66",X"A2",X"0A",X"A5",X"1E",X"07",X"48",X"A0",X"08",X"A0",X"08",
		X"F9",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"88",X"94",X"69",X"00",X"28",X"00",X"28",X"00",
		X"A4",X"0C",X"A4",X"0C",X"EC",X"0A",X"A2",X"0A",X"A2",X"1D",X"06",X"97",X"A0",X"08",X"A0",X"08",
		X"F8",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"EC",X"93",X"1D",X"00",X"28",X"00",X"28",X"00",
		X"A4",X"0C",X"A4",X"6C",X"A2",X"0A",X"A2",X"0A",X"A2",X"1C",X"05",X"97",X"A0",X"08",X"A0",X"08",
		X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"0F",X"00",X"28",X"00",X"28",X"00",X"28",X"00",
		X"A4",X"B1",X"1E",X"0A",X"A2",X"0A",X"A2",X"0A",X"A2",X"1B",X"04",X"97",X"A0",X"08",X"A0",X"08",
		X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",
		X"A0",X"08",X"A2",X"0A",X"A2",X"A5",X"A4",X"0C",X"A4",X"0C",X"0C",X"09",X"A1",X"A3",X"A3",X"0B",
		X"2B",X"00",X"28",X"00",X"82",X"03",X"2B",X"A9",X"29",X"01",X"29",X"A8",X"2C",X"04",X"28",X"00",
		X"A0",X"08",X"A2",X"0A",X"A2",X"0A",X"0D",X"0C",X"A4",X"0C",X"9A",X"09",X"A1",X"A3",X"A3",X"0B",
		X"11",X"00",X"28",X"00",X"10",X"03",X"2B",X"AF",X"29",X"01",X"29",X"AE",X"2C",X"04",X"28",X"00",
		X"0A",X"22",X"0A",X"22",X"0A",X"22",X"0E",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"28",X"88",X"00",X"6A",X"90",X"33",X"93",X"18",X"8B",X"34",X"CB",X"20",X"82",X"26",
		X"3A",X"39",X"39",X"3D",X"39",X"08",X"1B",X"28",X"0A",X"28",X"0A",X"39",X"39",X"28",X"7A",X"88",
		X"99",X"39",X"99",X"39",X"99",X"39",X"99",X"A9",X"9B",X"31",X"93",X"33",X"93",X"33",X"93",X"33",
		X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",
		X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",
		X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"5B",X"33",X"08",X"26",
		X"AA",X"20",X"8A",X"28",X"90",X"68",X"93",X"A9",X"08",X"7A",X"99",X"39",X"99",X"88",X"88",X"A8",
		X"0A",X"3D",X"39",X"29",X"18",X"33",X"1B",X"33",X"3B",X"31",X"1B",X"33",X"1B",X"33",X"1B",X"33",
		X"97",X"3B",X"82",X"22",X"82",X"22",X"18",X"3A",X"81",X"3A",X"99",X"39",X"99",X"39",X"99",X"39",
		X"39",X"A9",X"3B",X"31",X"1B",X"AB",X"18",X"2B",X"28",X"22",X"0A",X"22",X"1E",X"33",X"1B",X"08",
		X"88",X"2C",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"C8",X"28",
		X"28",X"26",X"21",X"33",X"1B",X"33",X"1B",X"33",X"5B",X"33",X"23",X"39",X"3D",X"A9",X"98",X"22",
		X"99",X"31",X"93",X"33",X"08",X"60",X"82",X"22",X"08",X"20",X"82",X"22",X"82",X"3A",X"D9",X"10",
		X"3B",X"31",X"28",X"33",X"19",X"2B",X"0C",X"39",X"3B",X"AA",X"79",X"39",X"39",X"10",X"1B",X"33",
		X"18",X"33",X"8B",X"A8",X"82",X"22",X"82",X"22",X"18",X"33",X"93",X"33",X"93",X"08",X"93",X"33",
		X"1B",X"B3",X"1B",X"B3",X"1B",X"38",X"39",X"01",X"A0",X"20",X"1B",X"B3",X"2F",X"31",X"88",X"B2",
		X"88",X"88",X"88",X"88",X"AA",X"88",X"88",X"0B",X"93",X"0B",X"28",X"AA",X"9A",X"99",X"99",X"B0",
		X"A0",X"20",X"28",X"20",X"39",X"31",X"39",X"20",X"1B",X"35",X"39",X"B3",X"39",X"A2",X"0A",X"A6",
		X"C2",X"AA",X"82",X"AA",X"82",X"AA",X"81",X"BC",X"9B",X"99",X"81",X"AA",X"AA",X"A8",X"9D",X"99",
		X"39",X"31",X"39",X"31",X"39",X"31",X"39",X"31",X"39",X"31",X"39",X"31",X"39",X"31",X"39",X"31",
		X"99",X"09",X"8A",X"88",X"88",X"88",X"88",X"C8",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",
		X"A0",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",
		X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",
		X"A0",X"31",X"1B",X"31",X"09",X"93",X"A0",X"93",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"0A",X"22",X"0A",X"22",X"0A",X"22",X"0A",X"22",X"0A",X"22",X"0A",X"22",X"0A",X"22",X"0E",X"2A",
		X"88",X"28",X"88",X"28",X"A8",X"10",X"88",X"28",X"88",X"68",X"10",X"33",X"93",X"33",X"D3",X"2B",
		X"1B",X"33",X"1B",X"33",X"1B",X"08",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",
		X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",
		X"1B",X"33",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"5B",X"18",X"39",X"10",X"1B",X"37",X"1B",X"33",
		X"AB",X"39",X"D9",X"33",X"93",X"33",X"93",X"88",X"99",X"39",X"99",X"39",X"99",X"39",X"99",X"39",
		X"39",X"39",X"39",X"3B",X"39",X"33",X"1B",X"37",X"1B",X"33",X"1B",X"33",X"1B",X"33",X"A8",X"28",
		X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"A8",
		X"88",X"22",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"A9",X"3B",X"39",X"39",X"39",
		X"00",X"3A",X"91",X"68",X"A8",X"18",X"99",X"39",X"99",X"39",X"99",X"A9",X"10",X"33",X"93",X"33",
		X"1B",X"AB",X"19",X"33",X"1B",X"33",X"A8",X"28",X"28",X"2A",X"68",X"30",X"20",X"00",X"0A",X"22",
		X"82",X"22",X"88",X"22",X"82",X"22",X"AA",X"21",X"88",X"68",X"81",X"39",X"91",X"33",X"97",X"39",
		X"39",X"A9",X"3B",X"22",X"0A",X"62",X"1A",X"39",X"39",X"39",X"39",X"39",X"3D",X"39",X"1D",X"2B",
		X"88",X"26",X"9A",X"22",X"C2",X"22",X"82",X"AA",X"88",X"2C",X"88",X"22",X"82",X"22",X"82",X"22",
		X"0A",X"2E",X"28",X"28",X"28",X"20",X"A0",X"39",X"59",X"28",X"28",X"10",X"1B",X"33",X"1B",X"33",
		X"93",X"37",X"93",X"33",X"97",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",X"93",X"33",
		X"1B",X"B3",X"1B",X"B7",X"1B",X"B3",X"1B",X"B3",X"1B",X"B3",X"23",X"31",X"5B",X"F3",X"1B",X"B3",
		X"93",X"BB",X"93",X"BB",X"93",X"BB",X"93",X"BB",X"93",X"BB",X"93",X"BB",X"93",X"BB",X"93",X"90",
		X"39",X"31",X"79",X"31",X"0A",X"62",X"1B",X"33",X"1F",X"B3",X"1B",X"B3",X"1B",X"B3",X"1B",X"B3",
		X"93",X"90",X"8A",X"A8",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"28",X"AA",X"88",X"BB",
		X"1B",X"31",X"0A",X"A6",X"22",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",X"A0",X"08",X"0A",X"20",
		X"88",X"88",X"10",X"88",X"88",X"C8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"28",X"20",X"28",X"20",X"28",X"20",X"3A",X"31",X"39",X"35",X"39",X"93",X"A0",X"93",X"A0",X"93",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",X"5F",X"F7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"F7",X"2F",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8E",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",
		X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2E",X"8B",X"8E",X"8B",X"2B",X"8B",X"2B",X"8B",
		X"A3",X"8B",X"A3",X"8E",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"2D",X"A3",X"8B",X"A3",X"8B",
		X"2B",X"8B",X"2B",X"8E",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2E",X"8B",X"2B",X"8B",X"2B",X"8B",
		X"A3",X"8B",X"A6",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8E",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",
		X"2E",X"8B",X"2B",X"8B",X"7E",X"8B",X"2E",X"2E",X"2B",X"8B",X"2B",X"8E",X"2B",X"8B",X"2B",X"8E",
		X"A3",X"8B",X"A6",X"8B",X"A6",X"8B",X"A3",X"8E",X"F5",X"2F",X"A6",X"8E",X"A6",X"8E",X"A6",X"89",
		X"2E",X"89",X"29",X"89",X"7C",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"2F",X"DB",X"29",X"89",
		X"A7",X"89",X"A7",X"8F",X"A7",X"8F",X"2E",X"8F",X"77",X"8A",X"A7",X"8A",X"A2",X"8F",X"2D",X"8A",
		X"2A",X"8A",X"2A",X"8F",X"2A",X"8A",X"2A",X"8A",X"2F",X"8A",X"2A",X"8A",X"8C",X"8A",X"2A",X"8F",
		X"A2",X"8A",X"A2",X"8A",X"A7",X"8A",X"A2",X"8A",X"A2",X"8F",X"A2",X"8A",X"A2",X"FE",X"A2",X"8F",
		X"2A",X"8A",X"2A",X"8A",X"2F",X"8A",X"2A",X"8A",X"2A",X"8F",X"8A",X"8A",X"2A",X"8A",X"2F",X"8A",
		X"A2",X"8A",X"A2",X"8A",X"A7",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A7",X"8A",X"A2",X"2B",
		X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2F",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",
		X"2C",X"8A",X"A2",X"8A",X"A7",X"8A",X"A2",X"8A",X"A2",X"2D",X"A2",X"8A",X"A2",X"8A",X"2E",X"8A",
		X"2A",X"8A",X"2A",X"DA",X"8F",X"89",X"48",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"2F",X"4F",X"A7",X"0A",X"A2",X"0F",X"A2",X"0A",X"A7",X"0A",X"A2",X"0F",X"A2",X"0A",X"A7",X"0A",
		X"2A",X"07",X"2A",X"07",X"2A",X"07",X"2A",X"46",X"2F",X"02",X"2F",X"02",X"2F",X"01",X"2E",X"03",
		X"2C",X"0B",X"A6",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0E",X"A3",X"0B",X"A3",X"0B",X"A3",X"4D",
		X"2E",X"03",X"2B",X"03",X"2B",X"06",X"2B",X"03",X"2B",X"03",X"2B",X"06",X"2B",X"03",X"2B",X"03",
		X"A6",X"0B",X"2F",X"0E",X"A3",X"0E",X"A3",X"0E",X"E4",X"09",X"A1",X"0F",X"A7",X"0A",X"A7",X"0A",
		X"8E",X"02",X"2F",X"02",X"2A",X"02",X"2F",X"02",X"2A",X"02",X"2A",X"07",X"8C",X"02",X"2A",X"02",
		X"A7",X"47",X"A2",X"0A",X"A7",X"0A",X"A2",X"0A",X"A7",X"0A",X"A2",X"0F",X"A2",X"0F",X"A2",X"0A",
		X"2A",X"07",X"2A",X"8B",X"2F",X"02",X"2A",X"07",X"2A",X"07",X"2A",X"02",X"2F",X"02",X"2F",X"02",
		X"A7",X"0A",X"A2",X"0F",X"A2",X"0A",X"A7",X"0A",X"A2",X"0A",X"A7",X"0A",X"2A",X"0A",X"A7",X"0A",
		X"2F",X"4E",X"2A",X"02",X"2F",X"02",X"2A",X"07",X"2A",X"02",X"2F",X"02",X"2A",X"07",X"2A",X"07",
		X"A2",X"0F",X"A2",X"0F",X"A2",X"0F",X"2B",X"0A",X"A7",X"0A",X"A7",X"0A",X"A7",X"0A",X"A7",X"24",
		X"2F",X"07",X"2F",X"07",X"ED",X"07",X"2F",X"07",X"2F",X"8D",X"2F",X"07",X"2F",X"07",X"2F",X"41",
		X"A1",X"0F",X"A7",X"26",X"A7",X"0F",X"A1",X"0F",X"A1",X"0F",X"A7",X"09",X"A7",X"09",X"A1",X"0F",
		X"29",X"07",X"29",X"01",X"29",X"07",X"29",X"01",X"29",X"01",X"29",X"01",X"29",X"01",X"29",X"01",
		X"A1",X"09",X"A1",X"09",X"A1",X"09",X"A1",X"09",X"E0",X"09",X"A1",X"09",X"A1",X"09",X"A6",X"09",
		X"29",X"8D",X"29",X"01",X"2E",X"01",X"2E",X"01",X"2E",X"01",X"E4",X"06",X"2E",X"06",X"2E",X"06",
		X"A6",X"8B",X"A6",X"2C",X"A3",X"8B",X"A3",X"8E",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",
		X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"68",X"88",X"29",X"88",X"29",X"88",X"29",X"48",
		X"2F",X"CF",X"A1",X"89",X"A1",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",
		X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8A",X"2A",X"8F",X"2F",X"8A",X"2A",X"8A",X"2A",X"8A",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",
		X"2A",X"8A",X"2A",X"8F",X"2F",X"8A",X"2A",X"8F",X"2A",X"8A",X"2F",X"CE",X"2A",X"8A",X"2A",X"8A",
		X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A7",X"8F",X"A7",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",
		X"2A",X"8A",X"2A",X"8A",X"2A",X"8F",X"2A",X"8A",X"2A",X"8F",X"2F",X"8F",X"6D",X"8F",X"2F",X"8F",
		X"A2",X"8F",X"A7",X"8F",X"A2",X"8F",X"A7",X"8A",X"A2",X"8F",X"E4",X"8F",X"A7",X"8F",X"A7",X"8F",
		X"2F",X"8F",X"2F",X"CB",X"2F",X"8F",X"29",X"89",X"2F",X"89",X"29",X"8F",X"29",X"89",X"29",X"89",
		X"A3",X"8E",X"A1",X"89",X"E2",X"8E",X"A6",X"8E",X"A6",X"8E",X"A6",X"8E",X"A6",X"8E",X"A6",X"8E",
		X"2E",X"8E",X"2E",X"8E",X"2E",X"C9",X"2E",X"8E",X"2E",X"8E",X"2E",X"8E",X"2E",X"8E",X"2E",X"8E",
		X"A6",X"8E",X"A6",X"8E",X"A6",X"8E",X"A3",X"8B",X"A1",X"8B",X"A3",X"89",X"A3",X"8B",X"A1",X"8B",
		X"2B",X"89",X"2B",X"8B",X"29",X"8B",X"2B",X"89",X"2B",X"8B",X"29",X"8B",X"2B",X"89",X"E5",X"8B",
		X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"C9",X"E8",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"88",X"29",X"88",X"29",X"88",X"29",X"88",X"29",X"88",X"29",X"88",X"29",X"88",X"29",X"88",
		X"2F",X"4F",X"A2",X"0F",X"A2",X"0A",X"A2",X"0A",X"A7",X"0A",X"A2",X"0A",X"A2",X"0A",X"A7",X"0A",
		X"2A",X"02",X"2A",X"07",X"2A",X"02",X"2A",X"02",X"2F",X"02",X"2A",X"02",X"2A",X"07",X"2A",X"02",
		X"A2",X"0A",X"A7",X"0A",X"A2",X"0A",X"2E",X"4E",X"A7",X"0A",X"A2",X"0F",X"A2",X"0A",X"A2",X"0F",
		X"2A",X"02",X"2A",X"07",X"2A",X"02",X"2F",X"02",X"2A",X"07",X"2A",X"02",X"2F",X"02",X"2A",X"07",
		X"A2",X"0A",X"2D",X"4D",X"A7",X"0A",X"A2",X"0F",X"A2",X"0A",X"A7",X"0A",X"A7",X"0A",X"A2",X"0F",
		X"2A",X"07",X"2A",X"07",X"2A",X"07",X"8C",X"44",X"2F",X"02",X"2F",X"07",X"29",X"06",X"2E",X"03",
		X"A3",X"0E",X"A3",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0B",X"A3",X"0B",X"A3",X"0B",X"A3",X"0B",
		X"2B",X"8B",X"E7",X"06",X"2B",X"03",X"2B",X"03",X"2B",X"03",X"2B",X"03",X"2E",X"03",X"2B",X"03",
		X"A3",X"0B",X"A3",X"0B",X"A3",X"0E",X"A3",X"0B",X"A3",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0B",
		X"2B",X"06",X"2B",X"03",X"2B",X"03",X"2B",X"06",X"2B",X"03",X"2B",X"03",X"2E",X"03",X"2B",X"03",
		X"A3",X"0B",X"A6",X"0B",X"A3",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0B",X"A3",X"0B",X"A3",X"0B",
		X"2E",X"03",X"2B",X"03",X"2B",X"03",X"2E",X"03",X"2B",X"03",X"2B",X"03",X"2B",X"03",X"2E",X"03",
		X"A3",X"0B",X"A3",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0B",X"A3",X"0B",X"A3",X"0E",X"A3",X"0B",
		X"2B",X"03",X"2E",X"03",X"2B",X"03",X"2B",X"06",X"2B",X"03",X"2B",X"03",X"8A",X"6E",X"2E",X"03",
		X"A3",X"0B",X"A3",X"0E",X"A3",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0B",X"A3",X"0E",X"A3",X"0B",
		X"2B",X"03",X"2B",X"03",X"2E",X"03",X"2B",X"03",X"2B",X"06",X"2B",X"03",X"2B",X"03",X"2E",X"03",
		X"A3",X"8B",X"A6",X"8B",X"A3",X"CA",X"E8",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",
		X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",X"29",X"89",
		X"2F",X"5F",X"A3",X"0B",X"A3",X"0E",X"A3",X"0B",X"A3",X"0B",X"A3",X"0E",X"A3",X"0B",X"A3",X"0B",
		X"2B",X"06",X"2B",X"03",X"2B",X"03",X"2B",X"03",X"2E",X"03",X"2B",X"03",X"2E",X"03",X"2B",X"03",
		X"A6",X"0B",X"A6",X"0B",X"2E",X"5E",X"A6",X"0B",X"A6",X"0B",X"A6",X"0B",X"A6",X"0E",X"A6",X"0E",
		X"2B",X"06",X"8D",X"55",X"2E",X"03",X"2E",X"03",X"2E",X"03",X"2E",X"06",X"2B",X"06",X"2B",X"03",
		X"A6",X"0B",X"A3",X"0E",X"A3",X"0B",X"2C",X"5C",X"A6",X"0B",X"A3",X"0E",X"A3",X"0B",X"A3",X"0E",
		X"2B",X"03",X"2E",X"03",X"2E",X"03",X"2E",X"03",X"2E",X"06",X"8B",X"53",X"2E",X"01",X"2E",X"01",
		X"A6",X"0E",X"A6",X"0E",X"A1",X"0E",X"A1",X"09",X"A6",X"09",X"A1",X"09",X"2A",X"5A",X"A6",X"09",
		X"29",X"01",X"2E",X"01",X"29",X"01",X"2E",X"01",X"29",X"01",X"2E",X"06",X"89",X"5E",X"2E",X"06",
		X"A6",X"0B",X"A6",X"0B",X"A3",X"0B",X"A6",X"0B",X"A3",X"0E",X"20",X"00",X"F1",X"0E",X"A6",X"09",
		X"29",X"01",X"2F",X"01",X"29",X"07",X"2F",X"07",X"2F",X"87",X"FD",X"07",X"2A",X"07",X"2A",X"07",
		X"A2",X"0A",X"A2",X"0F",X"A2",X"0A",X"A2",X"0A",X"A2",X"0A",X"A2",X"0A",X"A7",X"0A",X"A2",X"0A",
		X"2A",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",
		X"A2",X"0F",X"A2",X"0A",X"A2",X"0A",X"A2",X"0A",X"A2",X"0A",X"A7",X"0A",X"A2",X"0A",X"A2",X"0A",
		X"2A",X"02",X"2A",X"02",X"2F",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"79",X"C0",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"2F",X"CF",X"A1",X"8F",X"A7",X"89",X"A7",X"89",X"A7",X"2F",X"E6",X"8F",X"A7",X"8F",X"A7",X"8F",
		X"29",X"8F",X"2F",X"2F",X"6D",X"8F",X"2F",X"8F",X"2F",X"8F",X"2F",X"89",X"2F",X"2F",X"6C",X"8F",
		X"A7",X"8F",X"A7",X"8F",X"A2",X"8F",X"A7",X"8F",X"2F",X"CB",X"A7",X"8F",X"A2",X"8F",X"A7",X"8F",
		X"2F",X"8F",X"2F",X"8F",X"2A",X"8F",X"2F",X"8F",X"2F",X"8A",X"2F",X"8A",X"2F",X"8F",X"8F",X"CA",
		X"A7",X"8F",X"A7",X"8A",X"A7",X"8F",X"A7",X"8F",X"A7",X"8A",X"A7",X"8F",X"A7",X"8F",X"A7",X"8F",
		X"2F",X"8F",X"2F",X"2F",X"69",X"8F",X"2F",X"8F",X"2F",X"8F",X"2F",X"8F",X"2F",X"8F",X"2F",X"8F",
		X"A7",X"8F",X"A7",X"8F",X"A7",X"8F",X"A7",X"8F",X"A7",X"8F",X"A7",X"8F",X"A7",X"8F",X"A7",X"89",
		X"2F",X"8F",X"2F",X"89",X"2F",X"8F",X"2F",X"8F",X"29",X"8F",X"29",X"8F",X"29",X"8F",X"29",X"8F",
		X"A1",X"89",X"A1",X"89",X"A1",X"2F",X"E0",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"89",X"A1",X"8E",
		X"29",X"89",X"2E",X"89",X"29",X"8E",X"29",X"8E",X"29",X"8E",X"2E",X"89",X"2E",X"8E",X"29",X"8E",
		X"A6",X"8E",X"A6",X"8E",X"A6",X"8E",X"A6",X"2D",X"44",X"8E",X"A6",X"8B",X"A6",X"8E",X"A6",X"8E",
		X"2E",X"8B",X"2E",X"8B",X"2E",X"8B",X"2E",X"8B",X"2B",X"8E",X"2B",X"8B",X"2B",X"8B",X"2E",X"8B",
		X"A3",X"8B",X"A3",X"8E",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",
		X"2B",X"8E",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",
		X"A3",X"8B",X"A3",X"8B",X"A6",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",X"A3",X"8B",
		X"2B",X"8E",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",X"2B",X"8B",
		X"E8",X"0B",X"A3",X"0B",X"A3",X"0B",X"A1",X"09",X"E0",X"68",X"A1",X"09",X"A1",X"09",X"A1",X"09",
		X"29",X"C0",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",X"A0",X"09",
		X"28",X"01",X"28",X"01",X"28",X"01",X"28",X"01",X"66",X"01",X"06",X"01",X"C3",X"01",X"C2",X"C0",
		X"40",X"70",X"28",X"74",X"28",X"7D",X"08",X"72",X"08",X"77",X"08",X"74",X"D7",X"70",X"08",X"75",
		X"80",X"F0",X"A0",X"F6",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"40",X"70",X"20",X"74",X"08",X"7D",X"00",X"72",X"00",X"77",X"48",X"74",X"D7",X"70",X"38",X"76",
		X"80",X"F1",X"80",X"F7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"40",X"70",X"68",X"74",X"28",X"7E",X"48",X"72",X"48",X"77",X"28",X"75",X"D7",X"70",X"00",X"76",
		X"80",X"F2",X"A0",X"F7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"48",X"71",X"30",X"72",X"78",X"72",X"68",X"73",X"18",X"73",X"40",X"71",X"D7",X"70",
		X"7F",X"D7",X"80",X"71",X"C0",X"77",X"C0",X"71",X"88",X"73",X"E0",X"73",X"F8",X"71",X"E8",X"71",
		X"D7",X"70",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"80",X"71",X"C0",X"71",X"88",X"73",X"E0",X"73",X"F8",X"71",X"C0",X"77",X"E8",X"71",
		X"D7",X"70",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"00",X"D6",X"05",X"56",X"00",X"D1",X"01",X"22",X"02",X"24",X"02",X"25",X"02",
		X"8F",X"2A",X"09",X"2A",X"0B",X"2A",X"98",X"2A",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D2",
		X"D7",X"2A",X"D6",X"22",X"D1",X"2A",X"DE",X"29",X"A1",X"2C",X"AF",X"2A",X"AD",X"2A",X"AC",X"2A",
		X"88",X"2A",X"8A",X"2A",X"8C",X"2A",X"8D",X"2A",X"88",X"2A",X"8A",X"2A",X"8C",X"2A",X"8D",X"2C",
		X"BD",X"2C",X"D2",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"28",X"D6",X"27",X"D1",X"29",X"28",X"28",X"29",X"28",X"2A",X"28",X"2B",X"28",X"2C",X"28",
		X"85",X"28",X"86",X"28",X"87",X"28",X"00",X"28",X"01",X"28",X"02",X"28",X"03",X"28",X"90",X"28",
		X"39",X"28",X"3A",X"28",X"3B",X"28",X"3C",X"28",X"3D",X"28",X"3E",X"28",X"3F",X"28",X"30",X"28",
		X"11",X"28",X"12",X"28",X"13",X"28",X"88",X"28",X"89",X"28",X"8A",X"28",X"8B",X"28",X"8C",X"28",
		X"AD",X"28",X"AE",X"28",X"AF",X"28",X"A0",X"28",X"A1",X"28",X"A2",X"28",X"A3",X"28",X"B8",X"28",
		X"99",X"28",X"9A",X"28",X"9B",X"28",X"9C",X"28",X"9D",X"28",X"9E",X"28",X"9F",X"28",X"18",X"28",
		X"B1",X"28",X"B2",X"28",X"B3",X"28",X"D2",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2F",X"D6",X"27",X"DE",X"28",X"D1",X"2A",X"A8",X"28",X"AC",X"28",X"AF",X"28",X"AC",X"28",
		X"88",X"28",X"8C",X"28",X"8F",X"28",X"7D",X"2A",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2D",X"D6",X"27",X"D1",X"29",X"DE",X"28",X"28",X"2C",X"B8",X"2C",X"D5",X"B8",X"D2",X"D7",
		X"7F",X"2B",X"7E",X"AA",X"FE",X"28",X"79",X"28",X"90",X"2A",X"91",X"2A",X"90",X"2A",X"7D",X"2B",
		X"AB",X"00",X"AA",X"00",X"A9",X"00",X"A8",X"00",X"2F",X"00",X"2E",X"00",X"2D",X"00",X"2C",X"00",
		X"83",X"28",X"82",X"28",X"81",X"28",X"80",X"28",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"2D",X"7E",X"AF",X"79",X"28",X"80",X"AF",X"90",X"A8",X"7F",X"2C",X"7E",X"A8",X"98",X"2C",
		X"D6",X"04",X"30",X"08",X"D6",X"00",X"D2",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"2D",X"7E",X"AF",X"79",X"28",X"98",X"A8",X"7E",X"2C",X"7E",X"A8",X"88",X"2C",X"7E",X"2C",
		X"20",X"08",X"D6",X"00",X"D2",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"00",X"D6",X"04",X"D1",X"01",X"56",X"00",X"28",X"04",X"2C",X"04",X"2F",X"04",X"38",X"04",
		X"94",X"2C",X"97",X"2C",X"88",X"2C",X"8C",X"2C",X"8F",X"2C",X"98",X"2C",X"7D",X"2B",X"7A",X"28",
		X"D7",X"01",X"D6",X"04",X"D1",X"01",X"56",X"00",X"2C",X"04",X"2F",X"04",X"38",X"04",X"3C",X"04",
		X"97",X"2C",X"88",X"2C",X"8C",X"2C",X"8F",X"2C",X"98",X"2C",X"9C",X"2C",X"7D",X"2B",X"7A",X"28",
		X"D7",X"06",X"D6",X"04",X"D1",X"01",X"56",X"00",X"2F",X"04",X"38",X"04",X"3C",X"04",X"3F",X"04",
		X"88",X"2C",X"8C",X"2C",X"8F",X"2C",X"98",X"2C",X"9C",X"2C",X"9F",X"2C",X"7D",X"2B",X"7A",X"28",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2D",X"D6",X"2F",X"D1",X"28",X"38",X"2E",X"D0",X"2C",X"38",X"2E",X"68",X"2C",X"D0",X"2C",
		X"C0",X"A8",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"29",X"D6",X"27",X"DE",X"28",X"D1",X"28",X"28",X"28",X"D6",X"26",X"28",X"28",X"D6",X"25",
		X"80",X"28",X"7E",X"AC",X"80",X"28",X"7E",X"AB",X"80",X"28",X"7E",X"AA",X"80",X"28",X"7E",X"A9",
		X"28",X"2D",X"D6",X"20",X"28",X"28",X"D6",X"2F",X"28",X"28",X"D6",X"2E",X"28",X"28",X"D6",X"2D",
		X"80",X"28",X"7E",X"2C",X"80",X"28",X"7E",X"2B",X"80",X"28",X"7E",X"2A",X"80",X"28",X"7E",X"29",
		X"28",X"28",X"D6",X"28",X"D5",X"29",X"D2",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"2A",X"7E",X"AF",X"FE",X"28",X"79",X"28",X"42",X"2C",X"43",X"28",X"D0",X"28",X"D1",X"28",
		X"7A",X"28",X"7B",X"28",X"7C",X"28",X"7D",X"28",X"7E",X"28",X"7F",X"28",X"70",X"28",X"71",X"28",
		X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2D",X"D6",X"28",X"DE",X"28",X"D1",X"28",X"D6",X"27",X"38",X"28",X"D6",X"25",X"23",X"28",
		X"7E",X"AD",X"02",X"28",X"7F",X"2D",X"01",X"28",X"7E",X"A8",X"00",X"28",X"7E",X"2F",X"87",X"28",
		X"D6",X"2E",X"2E",X"28",X"D6",X"2D",X"2D",X"28",X"D6",X"2C",X"2C",X"28",X"D6",X"2B",X"2B",X"28",
		X"7E",X"2A",X"82",X"28",X"7E",X"29",X"81",X"28",X"7E",X"28",X"7D",X"29",X"7A",X"D7",X"7F",X"D7",
		X"D7",X"07",X"D6",X"04",X"56",X"01",X"D1",X"05",X"38",X"02",X"20",X"02",X"38",X"02",X"38",X"02",
		X"88",X"2A",X"90",X"2A",X"88",X"2A",X"88",X"2A",X"90",X"2A",X"7D",X"2B",X"7A",X"2A",X"98",X"2A",
		X"D7",X"01",X"D6",X"04",X"56",X"01",X"D1",X"05",X"3C",X"02",X"24",X"02",X"3C",X"02",X"3C",X"02",
		X"8C",X"2A",X"94",X"2A",X"8C",X"2A",X"8C",X"2A",X"94",X"2A",X"7D",X"2B",X"7A",X"2A",X"9D",X"2A",
		X"D7",X"02",X"D6",X"04",X"56",X"01",X"D1",X"05",X"3F",X"02",X"27",X"02",X"3F",X"02",X"3F",X"02",
		X"8F",X"2A",X"97",X"2A",X"8F",X"2A",X"8F",X"2A",X"97",X"2A",X"7D",X"2B",X"7A",X"D7",X"80",X"23",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"06",X"D6",X"06",X"56",X"01",X"D1",X"05",X"3F",X"02",X"24",X"02",X"3F",X"02",X"3E",X"02",
		X"8B",X"2A",X"96",X"2A",X"95",X"2A",X"8A",X"2A",X"95",X"2A",X"88",X"2A",X"8A",X"2A",X"8B",X"2A",
		X"24",X"08",X"D2",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"06",X"D6",X"06",X"56",X"01",X"D1",X"05",X"28",X"02",X"D0",X"02",X"28",X"02",X"28",X"02",
		X"78",X"2A",X"80",X"2A",X"80",X"2A",X"78",X"2A",X"80",X"2A",X"94",X"2A",X"95",X"2A",X"96",X"2A",
		X"3F",X"08",X"D2",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2E",X"D6",X"2E",X"DE",X"29",X"D1",X"2D",X"3F",X"2A",X"AC",X"2A",X"3F",X"2A",X"3E",X"2A",
		X"8B",X"2A",X"96",X"2A",X"95",X"2A",X"8A",X"2A",X"95",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",
		X"28",X"20",X"D2",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2A",X"D6",X"2C",X"DE",X"29",X"D1",X"2B",X"33",X"2C",X"33",X"2C",X"A8",X"2C",X"AA",X"2C",
		X"8A",X"2C",X"88",X"2C",X"13",X"2C",X"11",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",
		X"33",X"2E",X"31",X"2A",X"31",X"2E",X"33",X"2C",X"33",X"2C",X"A8",X"2C",X"AA",X"2C",X"AA",X"2C",
		X"88",X"2C",X"13",X"2C",X"11",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",X"11",X"2E",
		X"3F",X"2A",X"3F",X"2E",X"31",X"2C",X"31",X"2C",X"33",X"2C",X"3F",X"2C",X"31",X"2C",X"33",X"2A",
		X"88",X"2A",X"13",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2A",X"88",X"2A",X"13",X"2C",X"11",X"2C",
		X"3F",X"2C",X"31",X"2C",X"3A",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"A8",X"2C",X"AA",X"2C",
		X"8A",X"2C",X"88",X"2C",X"13",X"2C",X"11",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",
		X"B9",X"06",X"3F",X"02",X"3F",X"06",X"56",X"00",X"D0",X"04",X"D2",X"00",X"28",X"00",X"28",X"00",
		X"7F",X"28",X"7E",X"2C",X"FE",X"29",X"79",X"2B",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",
		X"BB",X"04",X"B9",X"04",X"3F",X"04",X"3A",X"04",X"AB",X"04",X"AB",X"04",X"3A",X"04",X"3F",X"04",
		X"97",X"2E",X"96",X"2A",X"96",X"2E",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",X"13",X"2C",
		X"B9",X"04",X"3F",X"04",X"3A",X"04",X"AB",X"04",X"AB",X"04",X"3A",X"04",X"3F",X"04",X"3E",X"06",
		X"97",X"2A",X"97",X"2E",X"96",X"2C",X"92",X"2C",X"97",X"2C",X"03",X"2C",X"92",X"2C",X"97",X"2A",
		X"B9",X"02",X"3F",X"04",X"3F",X"04",X"3E",X"04",X"3F",X"02",X"B9",X"02",X"BB",X"04",X"3E",X"04",
		X"94",X"2C",X"91",X"2C",X"92",X"2C",X"97",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",
		X"BB",X"04",X"B9",X"04",X"3F",X"04",X"3A",X"04",X"AB",X"04",X"AB",X"04",X"3A",X"04",X"3F",X"04",
		X"96",X"2E",X"97",X"2A",X"97",X"2E",X"FE",X"28",X"78",X"2C",X"7A",X"28",X"80",X"28",X"80",X"28",
		X"D7",X"03",X"D6",X"04",X"56",X"01",X"D1",X"03",X"BB",X"04",X"BB",X"04",X"20",X"04",X"22",X"04",
		X"8A",X"2C",X"88",X"2C",X"13",X"2C",X"11",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",
		X"BB",X"06",X"B9",X"02",X"B9",X"06",X"BB",X"04",X"BB",X"04",X"20",X"04",X"22",X"04",X"22",X"04",
		X"88",X"2C",X"13",X"2C",X"11",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",X"11",X"2E",
		X"3F",X"02",X"3F",X"06",X"B9",X"04",X"B9",X"04",X"BB",X"04",X"3F",X"04",X"B9",X"04",X"BB",X"02",
		X"88",X"2A",X"13",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2A",X"88",X"2A",X"13",X"2C",X"11",X"2C",
		X"3F",X"2C",X"31",X"2C",X"3A",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"A8",X"2C",X"AA",X"2C",
		X"8A",X"2C",X"88",X"2C",X"13",X"2C",X"11",X"2C",X"97",X"2C",X"97",X"2C",X"11",X"2C",X"13",X"2C",
		X"31",X"2E",X"3F",X"2A",X"3F",X"2E",X"DE",X"28",X"D0",X"2C",X"D2",X"28",X"28",X"28",X"28",X"28",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2A",X"D6",X"22",X"DE",X"28",X"D1",X"28",X"A8",X"29",X"AA",X"29",X"AC",X"29",X"AD",X"29",
		X"8F",X"29",X"09",X"29",X"0B",X"29",X"98",X"2A",X"7D",X"2B",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2E",X"D6",X"20",X"DE",X"29",X"D1",X"2A",X"38",X"2C",X"31",X"2C",X"38",X"2C",X"3C",X"2C",
		X"95",X"2E",X"95",X"2A",X"94",X"2C",X"92",X"2C",X"7D",X"2B",X"90",X"2C",X"90",X"2C",X"7A",X"D7",
		X"D7",X"2D",X"D6",X"20",X"DE",X"29",X"D1",X"2A",X"A8",X"2C",X"B8",X"2C",X"A8",X"2C",X"AF",X"2C",
		X"09",X"A8",X"8F",X"2C",X"8D",X"2C",X"7D",X"2B",X"98",X"2C",X"98",X"2C",X"7A",X"D7",X"7F",X"D7",
		X"D7",X"2D",X"D6",X"20",X"DE",X"29",X"D1",X"2A",X"A8",X"2C",X"B8",X"2C",X"A8",X"2C",X"AF",X"2C",
		X"09",X"A8",X"8F",X"2C",X"8D",X"2C",X"7D",X"2B",X"98",X"2C",X"98",X"2C",X"7A",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"03",X"D6",X"06",X"56",X"01",X"B1",X"02",X"37",X"02",X"B1",X"02",X"34",X"02",X"30",X"02",
		X"9C",X"2A",X"09",X"2C",X"19",X"2A",X"9F",X"2A",X"19",X"2A",X"9C",X"2A",X"98",X"2A",X"9C",X"2A",
		X"A1",X"04",X"B1",X"02",X"B3",X"02",X"68",X"02",X"B3",X"01",X"68",X"01",X"68",X"02",X"B1",X"02",
		X"1B",X"2A",X"19",X"29",X"1B",X"29",X"1B",X"2A",X"9F",X"2A",X"19",X"2A",X"9D",X"2A",X"98",X"2A",
		X"35",X"02",X"B1",X"02",X"D0",X"02",X"D5",X"02",X"57",X"01",X"34",X"02",X"32",X"02",X"34",X"02",
		X"98",X"2A",X"8F",X"2A",X"98",X"2A",X"8C",X"2C",X"7D",X"2A",X"FF",X"28",X"9C",X"2A",X"9E",X"2A",
		X"37",X"02",X"36",X"01",X"37",X"02",X"37",X"01",X"34",X"02",X"36",X"02",X"34",X"01",X"36",X"02",
		X"9E",X"29",X"9A",X"2A",X"9C",X"2A",X"0B",X"2A",X"8F",X"2A",X"0B",X"2A",X"9C",X"2A",X"78",X"2A",
		X"55",X"FF",X"D2",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"29",X"D6",X"2C",X"DE",X"29",X"3C",X"2A",X"AC",X"2A",X"31",X"2A",X"AC",X"2A",X"3C",X"2A",
		X"8C",X"2A",X"11",X"2A",X"8C",X"2A",X"94",X"2A",X"8C",X"2A",X"11",X"2A",X"8C",X"2A",X"94",X"2A",
		X"AC",X"2A",X"31",X"2A",X"AC",X"2A",X"3C",X"2A",X"AC",X"2A",X"31",X"2A",X"AC",X"2A",X"3C",X"2A",
		X"8C",X"2A",X"97",X"2A",X"8A",X"2A",X"92",X"2A",X"8A",X"2A",X"95",X"2A",X"88",X"2A",X"90",X"2A",
		X"A8",X"2A",X"3D",X"2A",X"A8",X"2A",X"D5",X"2A",X"DF",X"29",X"3F",X"2A",X"AF",X"2A",X"A8",X"2A",
		X"8F",X"2A",X"97",X"2A",X"8F",X"2A",X"88",X"2A",X"8F",X"2A",X"7D",X"2A",X"FF",X"28",X"97",X"2A",
		X"AF",X"2A",X"A8",X"2A",X"AF",X"2A",X"3F",X"2A",X"AF",X"2A",X"AA",X"2A",X"A1",X"2A",X"31",X"2A",
		X"09",X"2A",X"8C",X"2A",X"0B",X"2A",X"13",X"2A",X"0B",X"2A",X"8C",X"2A",X"78",X"2A",X"FD",X"D7",
		X"D2",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"06",X"D6",X"04",X"56",X"01",X"2C",X"02",X"20",X"02",X"A9",X"02",X"20",X"02",X"2C",X"02",
		X"88",X"2A",X"01",X"2A",X"88",X"2A",X"84",X"2A",X"88",X"2A",X"01",X"2A",X"88",X"2A",X"84",X"2A",
		X"20",X"02",X"A9",X"02",X"20",X"02",X"2C",X"02",X"20",X"02",X"A9",X"02",X"20",X"02",X"2C",X"02",
		X"88",X"2A",X"87",X"2A",X"13",X"2A",X"82",X"2A",X"13",X"2A",X"85",X"2A",X"11",X"2A",X"80",X"2A",
		X"B9",X"02",X"2D",X"02",X"B9",X"02",X"D5",X"02",X"57",X"01",X"2F",X"02",X"24",X"02",X"38",X"02",
		X"8C",X"2A",X"87",X"2A",X"8C",X"2A",X"90",X"2A",X"8C",X"2A",X"7D",X"2A",X"FF",X"28",X"87",X"2A",
		X"24",X"02",X"38",X"02",X"24",X"02",X"2F",X"02",X"24",X"02",X"3A",X"02",X"26",X"02",X"A9",X"02",
		X"8E",X"2A",X"94",X"2A",X"8F",X"2A",X"03",X"2A",X"8F",X"2A",X"94",X"2A",X"78",X"2A",X"FD",X"D7",
		X"D2",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"2A",X"D6",X"20",X"D1",X"2A",X"DE",X"29",X"38",X"2C",X"38",X"2C",X"3C",X"2C",X"3F",X"2C",
		X"78",X"2C",X"94",X"2C",X"97",X"38",X"88",X"2C",X"88",X"2C",X"8C",X"2C",X"8F",X"2C",X"78",X"2C",
		X"AC",X"2C",X"AF",X"38",X"D2",X"2C",X"B8",X"2C",X"BC",X"2C",X"BF",X"2C",X"D0",X"2C",X"BC",X"2C",
		X"9F",X"38",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"29",X"D6",X"20",X"D1",X"2A",X"DE",X"29",X"3C",X"2C",X"3C",X"2C",X"3F",X"2C",X"A8",X"2C",
		X"78",X"2C",X"97",X"2C",X"88",X"38",X"7D",X"2A",X"7A",X"B8",X"7D",X"2A",X"7A",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"06",X"D6",X"08",X"D1",X"02",X"56",X"01",X"3F",X"04",X"3F",X"04",X"20",X"04",X"24",X"04",
		X"78",X"2C",X"88",X"2C",X"8C",X"38",X"7D",X"2A",X"7A",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"03",X"D6",X"08",X"56",X"01",X"D1",X"03",X"6D",X"04",X"6D",X"04",X"6D",X"04",X"78",X"08",
		X"D0",X"2A",X"D0",X"2A",X"D0",X"2C",X"D0",X"2C",X"C5",X"2C",X"C5",X"2C",X"C5",X"2C",X"D0",X"A8",
		X"78",X"02",X"78",X"02",X"78",X"04",X"78",X"04",X"6F",X"04",X"6F",X"04",X"6F",X"04",X"7A",X"08",
		X"D2",X"2A",X"D2",X"2A",X"D2",X"2C",X"D2",X"2C",X"C7",X"2C",X"C7",X"2C",X"C7",X"2C",X"D2",X"A8",
		X"7A",X"02",X"7A",X"02",X"7A",X"04",X"7A",X"04",X"D5",X"04",X"6D",X"04",X"6D",X"04",X"D2",X"00",
		X"80",X"28",X"7F",X"D7",X"80",X"28",X"7F",X"D7",X"80",X"D7",X"7F",X"28",X"80",X"D7",X"7F",X"28",
		X"28",X"FF",X"D7",X"00",X"28",X"FF",X"D7",X"00",X"28",X"FF",X"D7",X"00",X"28",X"FF",X"D7",X"00",
		X"80",X"D7",X"7F",X"28",X"80",X"D7",X"7F",X"28",X"80",X"D7",X"7F",X"28",X"80",X"D7",X"7F",X"28",
		X"D7",X"2A",X"D6",X"20",X"DE",X"29",X"D1",X"2B",X"2D",X"2C",X"2D",X"2A",X"2D",X"2A",X"D0",X"2C",
		X"80",X"2C",X"78",X"2C",X"82",X"2C",X"78",X"2C",X"84",X"2C",X"85",X"2C",X"85",X"2A",X"85",X"2A",
		X"D0",X"2C",X"28",X"2C",X"D0",X"2C",X"2A",X"2C",X"D0",X"2C",X"2C",X"2C",X"2F",X"2C",X"2F",X"2A",
		X"87",X"2A",X"78",X"2C",X"82",X"2C",X"78",X"2C",X"84",X"2C",X"78",X"2C",X"85",X"2C",X"87",X"2C",
		X"2F",X"2A",X"2F",X"2A",X"D0",X"2C",X"2A",X"2C",X"D0",X"2C",X"2C",X"2C",X"D0",X"2C",X"2F",X"2C",
		X"7D",X"2C",X"85",X"2C",X"85",X"2C",X"7A",X"28",X"7F",X"D7",X"80",X"28",X"7F",X"D7",X"80",X"28",
		X"D7",X"D7",X"28",X"28",X"D7",X"D7",X"28",X"28",X"D7",X"D7",X"28",X"28",X"D7",X"D7",X"28",X"28",
		X"7F",X"D7",X"80",X"28",X"7F",X"D7",X"80",X"28",X"7F",X"D7",X"80",X"28",X"7F",X"D7",X"80",X"28",
		X"D7",X"2E",X"D6",X"20",X"DE",X"29",X"D1",X"2E",X"2D",X"2A",X"28",X"2A",X"2A",X"2C",X"2D",X"2A",
		X"80",X"2A",X"82",X"2C",X"85",X"2A",X"80",X"2A",X"82",X"2A",X"85",X"2C",X"80",X"2A",X"82",X"2C",
		X"2F",X"2A",X"2A",X"2A",X"2C",X"2C",X"2F",X"2A",X"2A",X"2A",X"2C",X"2C",X"2F",X"2A",X"2A",X"2A",
		X"84",X"2A",X"87",X"2C",X"82",X"2A",X"84",X"2C",X"7D",X"2C",X"85",X"2A",X"85",X"2A",X"7A",X"28",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",X"7F",X"D7",
		X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"7C",X"28",X"80",X"28",X"80",X"28",X"80",X"28",X"12",X"28",X"7D",X"28",X"9C",X"28",X"D9",X"28");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
