library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_8N is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_8N is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"15",X"AA",X"54",X"AA",X"51",X"A8",X"54",X"A2",X"45",X"AA",X"50",X"8A",X"44",X"A2",X"55",
		X"2A",X"50",X"A2",X"40",X"AA",X"50",X"28",X"00",X"AA",X"54",X"AA",X"45",X"A8",X"54",X"AA",X"00",
		X"A2",X"50",X"AA",X"01",X"AA",X"41",X"0A",X"41",X"A0",X"40",X"2A",X"01",X"0A",X"10",X"AA",X"41",
		X"A8",X"00",X"A8",X"41",X"AA",X"55",X"20",X"00",X"8A",X"55",X"AA",X"40",X"AA",X"00",X"00",X"00",
		X"BF",X"FF",X"FF",X"7F",X"BF",X"7F",X"FF",X"7F",X"FD",X"FC",X"FE",X"F0",X"E9",X"E2",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"BF",X"5F",X"C8",X"82",X"D0",X"FB",X"FE",X"D1",X"E0",X"D2",
		X"FF",X"7E",X"BD",X"FE",X"FE",X"7F",X"BF",X"7F",X"E4",X"08",X"45",X"31",X"40",X"9A",X"F4",X"40",
		X"FF",X"7E",X"FC",X"F8",X"FD",X"7E",X"FF",X"7F",X"B5",X"04",X"90",X"B0",X"49",X"02",X"04",X"FE",
		X"C7",X"97",X"A3",X"43",X"13",X"51",X"B1",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"89",X"8C",X"2C",X"26",X"06",X"47",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FC",X"FA",X"D1",X"E3",X"F8",X"F9",X"FC",X"EE",
		X"BF",X"7F",X"BF",X"7F",X"BF",X"7F",X"FF",X"7F",X"FD",X"E8",X"E0",X"F9",X"F2",X"FA",X"FE",X"F8",
		X"01",X"06",X"83",X"47",X"6F",X"7F",X"3E",X"E5",X"80",X"00",X"00",X"C0",X"E0",X"26",X"19",X"0C",
		X"C8",X"A0",X"42",X"00",X"20",X"AC",X"0F",X"01",X"06",X"41",X"00",X"1B",X"26",X"08",X"18",X"C0",
		X"0A",X"0F",X"1A",X"15",X"20",X"03",X"01",X"44",X"04",X"0B",X"1C",X"0C",X"04",X"60",X"C0",X"20",
		X"D0",X"10",X"32",X"5C",X"0C",X"05",X"02",X"0A",X"11",X"26",X"47",X"4E",X"92",X"05",X"02",X"00",
		X"AA",X"15",X"AA",X"54",X"AA",X"51",X"A8",X"54",X"A2",X"45",X"AA",X"50",X"8A",X"44",X"A2",X"55",
		X"2A",X"50",X"A2",X"40",X"AA",X"00",X"28",X"15",X"AA",X"54",X"AA",X"45",X"A8",X"54",X"A2",X"00",
		X"AA",X"44",X"AA",X"45",X"2A",X"15",X"AA",X"11",X"AA",X"55",X"AA",X"40",X"AA",X"15",X"AA",X"51",
		X"AA",X"44",X"A2",X"15",X"8A",X"01",X"AA",X"14",X"AA",X"40",X"AA",X"55",X"AA",X"51",X"AA",X"51",
		X"88",X"72",X"78",X"32",X"B9",X"1B",X"D3",X"07",X"03",X"17",X"9E",X"FC",X"FE",X"F8",X"FF",X"FC",
		X"8F",X"6F",X"BF",X"5F",X"BF",X"7F",X"BF",X"7F",X"FC",X"F8",X"F8",X"F0",X"FE",X"F8",X"F0",X"F8",
		X"01",X"03",X"01",X"00",X"01",X"03",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"01",X"03",X"07",X"01",X"01",X"09",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"00",X"00",X"3F",X"3F",X"BF",X"BF",X"7F",X"3F",
		X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"3F",X"BF",X"BF",X"7F",X"3F",X"3F",X"BF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"3F",X"7F",X"3F",X"3F",X"BF",X"BF",X"7F",X"3F",X"3F",
		X"1F",X"1F",X"1E",X"1F",X"1E",X"17",X"17",X"16",X"BF",X"80",X"EF",X"EF",X"EF",X"E0",X"80",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"1F",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"FF",X"FF",X"FF",X"BF",X"DF",X"FF",X"0F",X"00",
		X"04",X"17",X"16",X"1F",X"17",X"1F",X"1E",X"16",X"40",X"E0",X"E7",X"E3",X"EF",X"EF",X"E0",X"C0",
		X"00",X"1E",X"16",X"17",X"17",X"17",X"1F",X"13",X"40",X"C0",X"E0",X"EF",X"EF",X"EF",X"6F",X"3F",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"3D",X"3F",X"FF",X"FF",X"FF",X"F7",X"EF",X"FF",
		X"07",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"3F",X"BF",X"BF",X"7F",X"3F",X"3F",X"BF",X"BF",
		X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"7F",X"3F",X"3F",X"BF",X"BF",X"7F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"BF",X"BF",X"7F",X"3F",X"3F",X"BF",X"BF",X"7F",
		X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"3F",X"3F",X"BF",X"BF",X"7F",X"3F",X"3F",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",
		X"7C",X"44",X"FC",X"C4",X"FF",X"FF",X"E7",X"FF",X"BF",X"7F",X"00",X"BF",X"BF",X"BF",X"FF",X"FF",
		X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"FF",X"C0",X"80",X"BF",X"BF",X"BF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"37",X"0F",
		X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"FF",X"C0",X"80",X"BF",X"BF",X"BF",X"FF",X"FF",
		X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"FF",X"C0",X"80",X"BF",X"BF",X"BF",X"FF",X"FF",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"1F",X"1F",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"03",X"03",X"00",X"00",
		X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"FF",X"C0",X"80",X"BF",X"BF",X"BF",X"FF",X"FF",
		X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"E7",X"FF",X"FF",X"C0",X"80",X"BF",X"BF",X"BF",X"80",X"00",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"07",X"03",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"08",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"24",X"90",X"84",X"11",X"80",X"10",X"02",X"00",X"BF",X"06",X"00",X"2A",X"C2",X"3B",X"08",X"03",
		X"20",X"86",X"11",X"21",X"02",X"00",X"B0",X"05",X"01",X"0A",X"00",X"03",X"40",X"10",X"02",X"63",
		X"FF",X"12",X"08",X"00",X"10",X"02",X"80",X"10",X"FF",X"8C",X"04",X"A6",X"00",X"40",X"84",X"25",
		X"C0",X"60",X"1C",X"17",X"11",X"10",X"00",X"A4",X"84",X"00",X"C0",X"84",X"C4",X"74",X"94",X"A7",
		X"DF",X"10",X"50",X"14",X"00",X"10",X"10",X"80",X"D7",X"10",X"00",X"18",X"20",X"10",X"91",X"50",
		X"34",X"11",X"00",X"12",X"10",X"10",X"80",X"10",X"10",X"14",X"40",X"30",X"00",X"14",X"00",X"91",
		X"FF",X"10",X"12",X"10",X"15",X"90",X"10",X"22",X"28",X"00",X"08",X"40",X"00",X"00",X"00",X"04",
		X"11",X"10",X"48",X"12",X"10",X"14",X"10",X"30",X"00",X"20",X"04",X"A0",X"10",X"00",X"00",X"28",
		X"00",X"82",X"04",X"0A",X"20",X"80",X"00",X"00",X"28",X"42",X"6A",X"08",X"A4",X"02",X"92",X"41",
		X"20",X"0A",X"82",X"00",X"20",X"01",X"00",X"21",X"10",X"2A",X"A9",X"00",X"52",X"12",X"09",X"0D",
		X"88",X"44",X"68",X"10",X"48",X"0C",X"0A",X"0A",X"84",X"04",X"90",X"01",X"04",X"84",X"80",X"44",
		X"80",X"08",X"44",X"00",X"08",X"52",X"08",X"C0",X"82",X"C0",X"A4",X"00",X"2C",X"04",X"02",X"05",
		X"D1",X"70",X"1C",X"03",X"02",X"08",X"10",X"90",X"40",X"00",X"44",X"40",X"C0",X"70",X"0C",X"47",
		X"20",X"80",X"10",X"54",X"03",X"10",X"08",X"10",X"81",X"44",X"00",X"40",X"00",X"40",X"C8",X"00",
		X"90",X"10",X"22",X"10",X"90",X"90",X"24",X"30",X"00",X"04",X"00",X"01",X"20",X"00",X"00",X"00",
		X"D0",X"70",X"1C",X"37",X"81",X"10",X"18",X"50",X"04",X"90",X"00",X"00",X"C4",X"01",X"00",X"60",
		X"00",X"80",X"20",X"00",X"14",X"80",X"00",X"00",X"90",X"00",X"45",X"20",X"42",X"84",X"09",X"81",
		X"00",X"82",X"00",X"00",X"20",X"00",X"22",X"80",X"10",X"04",X"02",X"02",X"00",X"10",X"03",X"04",
		X"46",X"88",X"40",X"40",X"08",X"48",X"04",X"00",X"08",X"94",X"01",X"04",X"80",X"85",X"44",X"80",
		X"C8",X"89",X"08",X"00",X"4A",X"00",X"49",X"08",X"AC",X"10",X"0C",X"86",X"84",X"00",X"44",X"8C",
		X"90",X"40",X"30",X"10",X"18",X"44",X"12",X"11",X"A0",X"21",X"00",X"20",X"20",X"20",X"20",X"02",
		X"08",X"10",X"00",X"18",X"91",X"00",X"84",X"10",X"80",X"60",X"20",X"10",X"20",X"24",X"0A",X"21",
		X"10",X"18",X"91",X"00",X"08",X"01",X"25",X"00",X"20",X"05",X"4A",X"5F",X"3B",X"3F",X"DF",X"FF",
		X"01",X"04",X"0D",X"87",X"03",X"0C",X"03",X"01",X"7F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"90",X"00",X"00",X"00",X"11",X"40",X"00",X"24",X"02",X"52",X"01",X"10",X"09",X"04",X"02",
		X"04",X"00",X"80",X"80",X"84",X"00",X"10",X"40",X"88",X"00",X"42",X"04",X"04",X"01",X"26",X"40",
		X"A0",X"80",X"40",X"00",X"21",X"08",X"05",X"08",X"86",X"00",X"04",X"88",X"00",X"85",X"04",X"00",
		X"22",X"20",X"00",X"22",X"00",X"42",X"00",X"43",X"88",X"04",X"04",X"20",X"80",X"04",X"03",X"01",
		X"20",X"90",X"50",X"21",X"08",X"10",X"08",X"08",X"20",X"20",X"42",X"20",X"00",X"20",X"40",X"18",
		X"14",X"10",X"22",X"01",X"10",X"00",X"54",X"00",X"20",X"22",X"A2",X"00",X"80",X"A0",X"68",X"A1",
		X"86",X"0B",X"04",X"93",X"01",X"04",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"41",X"87",X"01",X"53",X"14",X"0C",X"87",X"23",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"00",X"00",X"10",X"00",X"00",X"A0",X"04",X"02",X"00",X"80",X"02",X"09",X"10",X"00",X"03",
		X"00",X"00",X"02",X"20",X"80",X"00",X"01",X"40",X"00",X"00",X"28",X"02",X"00",X"08",X"04",X"02",
		X"05",X"20",X"04",X"02",X"10",X"04",X"10",X"00",X"40",X"01",X"84",X"D0",X"0C",X"10",X"84",X"08",
		X"08",X"06",X"80",X"34",X"00",X"00",X"44",X"88",X"22",X"24",X"04",X"01",X"C2",X"54",X"90",X"21",
		X"90",X"98",X"00",X"14",X"42",X"01",X"14",X"00",X"29",X"90",X"28",X"28",X"46",X"12",X"22",X"A5",
		X"00",X"90",X"50",X"05",X"10",X"12",X"08",X"90",X"10",X"20",X"26",X"00",X"21",X"44",X"00",X"60",
		X"14",X"03",X"83",X"00",X"51",X"0F",X"27",X"88",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"43",X"11",X"8C",X"07",X"0B",X"03",X"84",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"20",X"12",X"00",X"03",X"2C",X"80",X"08",X"01",
		X"00",X"04",X"00",X"08",X"40",X"00",X"00",X"80",X"02",X"00",X"10",X"04",X"00",X"00",X"40",X"09",
		X"02",X"88",X"43",X"00",X"2A",X"00",X"10",X"91",X"24",X"12",X"14",X"20",X"04",X"08",X"85",X"14",
		X"00",X"02",X"40",X"08",X"00",X"01",X"84",X"10",X"40",X"11",X"82",X"0A",X"84",X"22",X"05",X"D0",
		X"50",X"82",X"14",X"00",X"50",X"51",X"20",X"08",X"A4",X"20",X"40",X"00",X"A0",X"04",X"30",X"20",
		X"10",X"00",X"14",X"40",X"00",X"10",X"50",X"40",X"28",X"84",X"04",X"00",X"A3",X"20",X"45",X"88",
		X"91",X"A5",X"00",X"10",X"A0",X"25",X"00",X"13",X"FF",X"3F",X"FF",X"FF",X"9F",X"3F",X"7F",X"BF",
		X"81",X"12",X"A1",X"00",X"51",X"09",X"52",X"22",X"1F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"BF",
		X"00",X"84",X"00",X"00",X"00",X"02",X"80",X"00",X"21",X"00",X"04",X"22",X"01",X"00",X"00",X"41",
		X"00",X"20",X"00",X"08",X"00",X"82",X"00",X"00",X"08",X"01",X"02",X"00",X"08",X"01",X"10",X"04",
		X"80",X"44",X"08",X"00",X"00",X"50",X"42",X"01",X"02",X"10",X"80",X"44",X"00",X"04",X"50",X"01",
		X"08",X"00",X"00",X"84",X"00",X"00",X"00",X"40",X"00",X"02",X"A0",X"00",X"00",X"55",X"00",X"81",
		X"42",X"90",X"01",X"08",X"50",X"20",X"02",X"22",X"26",X"00",X"20",X"95",X"08",X"A2",X"04",X"28",
		X"00",X"90",X"02",X"04",X"10",X"80",X"08",X"04",X"42",X"19",X"22",X"04",X"B5",X"00",X"01",X"2A",
		X"82",X"22",X"40",X"01",X"A7",X"09",X"80",X"42",X"FF",X"7F",X"7F",X"FF",X"FF",X"BF",X"FF",X"7F",
		X"03",X"01",X"08",X"50",X"40",X"00",X"13",X"81",X"3F",X"FF",X"FF",X"7F",X"7F",X"FF",X"9F",X"3F",
		X"EA",X"D5",X"EA",X"D4",X"EA",X"F1",X"E8",X"D4",X"A2",X"45",X"AA",X"50",X"8A",X"44",X"A2",X"55",
		X"EA",X"D0",X"E2",X"C0",X"EA",X"E0",X"E8",X"D5",X"AA",X"54",X"AA",X"41",X"A8",X"54",X"A2",X"00",
		X"AA",X"C4",X"EA",X"C5",X"EA",X"95",X"AA",X"91",X"AA",X"55",X"AA",X"40",X"AA",X"15",X"AA",X"51",
		X"EA",X"C4",X"82",X"D5",X"8A",X"81",X"CA",X"D4",X"AA",X"40",X"AA",X"55",X"AA",X"51",X"AA",X"51",
		X"AA",X"D0",X"EA",X"E1",X"AA",X"E5",X"EA",X"C1",X"A8",X"40",X"2A",X"11",X"AA",X"14",X"AA",X"41",
		X"A8",X"D0",X"AA",X"C1",X"EA",X"D5",X"AA",X"C4",X"AA",X"55",X"AA",X"44",X"AA",X"21",X"CA",X"20",
		X"AA",X"95",X"EA",X"D4",X"AA",X"D1",X"E8",X"D4",X"A2",X"45",X"AA",X"50",X"8A",X"44",X"A2",X"55",
		X"AA",X"D0",X"E2",X"C0",X"EA",X"D0",X"EA",X"E0",X"AA",X"54",X"AA",X"45",X"A8",X"54",X"AA",X"00",
		X"AF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FC",X"FF",X"FE",X"F8",X"FE",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FE",X"FF",X"FE",X"FE",X"FC",X"FF",X"FE",
		X"03",X"1F",X"0F",X"13",X"0F",X"07",X"0F",X"3F",X"FC",X"F8",X"FE",X"FF",X"FE",X"FE",X"FF",X"FE",
		X"5F",X"1F",X"1F",X"BF",X"7F",X"BF",X"5F",X"BF",X"FC",X"FF",X"FA",X"FD",X"FE",X"FC",X"FE",X"FF",
		X"3F",X"7F",X"BF",X"1F",X"4F",X"3F",X"1F",X"3F",X"FE",X"FC",X"FE",X"FF",X"FE",X"FE",X"FF",X"FE",
		X"CF",X"7F",X"1F",X"BF",X"7F",X"BF",X"7F",X"BF",X"FD",X"F8",X"F2",X"FC",X"FA",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FD",X"FF",X"FE",X"F8",X"FE",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FE",X"FF",X"FE",X"FE",X"FC",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"E4",X"F8",X"FC",X"F0",X"F8",X"E8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"F8",X"C4",X"F0",X"FC",X"F0",X"FF",X"FE",
		X"00",X"00",X"00",X"02",X"03",X"0B",X"07",X"05",X"00",X"00",X"00",X"40",X"80",X"C0",X"E0",X"F0",
		X"03",X"07",X"0A",X"03",X"06",X"01",X"02",X"00",X"E0",X"F0",X"F0",X"E0",X"C0",X"40",X"80",X"00",
		X"00",X"00",X"00",X"00",X"02",X"0C",X"26",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2F",X"1F",X"3F",X"17",X"0F",X"17",X"0A",X"14",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"7F",X"7B",X"63",X"6B",X"63",X"7F",X"7F",X"01",X"7F",X"7B",X"63",X"6B",X"63",X"7F",X"7F",
		X"01",X"7F",X"7B",X"63",X"6B",X"63",X"7F",X"7F",X"01",X"7F",X"7B",X"63",X"6B",X"63",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"10",X"50",X"50",X"50",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"D0",X"D0",X"D0",X"50",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"FA",X"FA",X"FE",X"F7",X"F7",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FD",X"F7",X"F7",X"F6",X"F6",X"F6",
		X"EE",X"EB",X"EB",X"FB",X"FF",X"FB",X"EB",X"EF",X"DF",X"FF",X"DF",X"DF",X"5F",X"7F",X"6F",X"7F",
		X"EF",X"EF",X"EB",X"EA",X"FA",X"FA",X"FE",X"FF",X"5F",X"7F",X"EF",X"EF",X"AF",X"EF",X"DF",X"F7",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",
		X"00",X"00",X"00",X"06",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"99",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"06",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"99",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"99",X"00",X"66",
		X"00",X"99",X"00",X"66",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"66",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"EE",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"EE",X"FF",
		X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",
		X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",
		X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"7F",X"7F",X"3F",X"3F",X"1F",X"00",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"92",X"92",X"92",X"92",X"92",X"92",X"00",X"00",X"49",X"49",X"49",X"49",X"49",X"49",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"49",X"49",X"49",X"49",X"49",X"49",X"49",X"49",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"00",X"1F",X"06",X"0C",X"1F",X"00",X"1F",X"14",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"1F",X"04",X"AE",X"BF",X"AA",X"BF",X"BF",X"BF",
		X"AA",X"AA",X"AA",X"FF",X"7F",X"3F",X"1F",X"00",X"BF",X"AA",X"BA",X"FF",X"FF",X"FF",X"FF",X"00",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"49",X"49",X"49",X"49",X"49",X"49",X"49",X"49",
		X"92",X"92",X"92",X"92",X"92",X"92",X"00",X"00",X"49",X"49",X"49",X"49",X"49",X"49",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"B8",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B8",X"00",X"03",X"00",X"B8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"3B",X"00",X"00",X"00",
		X"0F",X"0F",X"7E",X"7E",X"7E",X"7F",X"7E",X"7E",X"3B",X"00",X"00",X"00",X"3B",X"00",X"00",X"00",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"3B",X"00",X"00",X"00",X"3B",X"00",X"00",X"00",
		X"7F",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"00",X"3B",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B8",X"00",X"03",X"00",X"B8",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"B8",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",
		X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",
		X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",
		X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",
		X"00",X"66",X"3F",X"19",X"0F",X"06",X"03",X"01",X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"66",X"3F",X"19",X"0F",X"06",X"03",X"00",
		X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",
		X"FF",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"00",X"FF",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"00",
		X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",
		X"CC",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"80",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",X"00",X"66",X"FF",X"99",X"FF",X"66",X"FF",X"99",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"08",X"08",X"08",X"0F",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"0F",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"0F",X"08",X"08",X"08",
		X"C0",X"80",X"C0",X"80",X"C0",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"C0",X"80",X"C0",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"10",X"70",X"E0",X"C0",X"C0",X"80",X"00",X"80",
		X"7F",X"7D",X"3E",X"7C",X"7E",X"FF",X"74",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"01",X"01",X"03",X"01",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"03",X"01",X"03",X"03",X"01",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"52",X"FC",X"FF",X"FF",X"FF",X"FF",X"01",X"0B",X"47",X"EF",X"C7",X"F7",X"FB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"F7",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"06",X"0C",X"40",X"80",X"C0",X"C0",X"00",X"20",X"20",X"60",
		X"30",X"41",X"47",X"4B",X"5F",X"47",X"4F",X"5B",X"64",X"FA",X"FE",X"FE",X"FF",X"FF",X"FF",X"DF",
		X"E3",X"C5",X"C3",X"C3",X"83",X"C1",X"C3",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CB",X"C3",X"C1",X"C3",X"C3",X"CB",X"81",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"FF",X"00",X"00",X"00",X"3E",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"3C",X"FB",X"F7",X"F6",X"F4",X"45",X"69",X"75",X"E8",X"05",X"54",X"E2",X"C4",
		X"00",X"00",X"00",X"00",X"02",X"23",X"3A",X"33",X"00",X"00",X"06",X"03",X"01",X"01",X"01",X"41",
		X"33",X"21",X"F8",X"BC",X"FF",X"DE",X"F8",X"C0",X"41",X"49",X"B9",X"F8",X"F1",X"73",X"7B",X"7F",
		X"49",X"39",X"30",X"10",X"00",X"00",X"00",X"03",X"CF",X"8F",X"87",X"83",X"81",X"01",X"01",X"03",
		X"1F",X"33",X"71",X"F8",X"F9",X"F8",X"F8",X"F8",X"FF",X"F1",X"C0",X"80",X"C0",X"E0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1D",X"01",X"07",X"17",X"77",X"F7",X"D5",X"55",X"55",
		X"7D",X"C0",X"80",X"7F",X"FE",X"FE",X"FA",X"FC",X"50",X"00",X"00",X"01",X"03",X"05",X"08",X"08",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"FE",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F8",
		X"03",X"07",X"07",X"06",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0B",X"19",X"19",X"1D",X"10",X"39",X"F9",X"F8",X"F9",X"FD",X"FD",X"FC",
		X"E0",X"E0",X"01",X"01",X"01",X"01",X"00",X"00",X"84",X"82",X"02",X"82",X"C2",X"82",X"A2",X"C0",
		X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"F1",X"FD",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"C4",X"61",X"71",X"61",X"43",X"42",X"61",X"00",X"7F",X"F5",X"FB",X"AB",X"DF",X"DF",X"1F",X"1D",
		X"28",X"25",X"24",X"0C",X"24",X"4C",X"34",X"24",X"3F",X"15",X"5F",X"2F",X"37",X"3F",X"1F",X"5D",
		X"F8",X"E0",X"F3",X"F0",X"F8",X"F0",X"D0",X"F8",X"C0",X"D0",X"C8",X"E0",X"48",X"48",X"C0",X"64",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"FF",X"FF",X"FC",X"40",X"E0",X"71",X"7F",X"FF",X"D3",X"01",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"18",X"30",X"20",X"7C",X"03",X"0F",
		X"00",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"70",X"00",X"00",X"00",X"00",X"00",X"C0",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"10",
		X"7F",X"3D",X"9D",X"CD",X"CD",X"05",X"C1",X"C1",X"F0",X"F8",X"FC",X"7E",X"3E",X"0E",X"0F",X"0F",
		X"C1",X"C9",X"C1",X"C0",X"40",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"03",
		X"18",X"19",X"1D",X"8F",X"BF",X"9D",X"98",X"BC",X"FE",X"FF",X"FD",X"F9",X"F9",X"F9",X"F1",X"F9",
		X"9D",X"9F",X"8F",X"9F",X"BF",X"1F",X"0F",X"1F",X"F9",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"C0",X"C0",X"C0",X"F8",X"FC",X"FC",X"7F",X"7C",X"35",X"3D",X"18",X"37",X"2E",X"0B",
		X"FC",X"E7",X"8F",X"CF",X"DF",X"FF",X"FF",X"FE",X"13",X"15",X"EF",X"DD",X"EF",X"FF",X"9F",X"1F",
		X"C0",X"80",X"80",X"87",X"8F",X"C7",X"C1",X"A0",X"01",X"01",X"00",X"70",X"30",X"B8",X"B0",X"F8",
		X"80",X"B0",X"D8",X"CC",X"8C",X"C2",X"80",X"C0",X"38",X"38",X"1C",X"18",X"00",X"00",X"00",X"00",
		X"C5",X"C7",X"CD",X"C3",X"DF",X"DF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"F2",X"E2",X"F2",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"82",X"86",X"84",X"80",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"08",X"08",X"00",X"11",X"11",X"11",X"00",X"01",
		X"00",X"04",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"30",X"14",X"00",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"80",X"07",X"07",X"07",X"07",X"0F",X"8F",X"8F",X"9F",
		X"81",X"87",X"1F",X"7F",X"00",X"00",X"00",X"00",X"E7",X"8F",X"7F",X"FF",X"1F",X"03",X"04",X"1A",
		X"67",X"B3",X"94",X"88",X"CB",X"C1",X"80",X"C0",X"FF",X"FD",X"FF",X"FF",X"FF",X"F9",X"CF",X"09",
		X"C0",X"80",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"87",X"04",X"00",X"80",X"E8",X"EC",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FD",X"32",X"83",X"C1",X"18",X"98",X"18",X"1C",X"1E",X"1E",
		X"00",X"C0",X"F2",X"7E",X"BE",X"B8",X"30",X"30",X"1E",X"1F",X"0C",X"58",X"CC",X"C0",X"81",X"01",
		X"C9",X"D9",X"DD",X"DC",X"EE",X"D7",X"C0",X"D0",X"60",X"60",X"B0",X"78",X"C0",X"C0",X"06",X"0C",
		X"C0",X"F8",X"E0",X"E8",X"E0",X"E0",X"C8",X"E8",X"06",X"06",X"70",X"1C",X"1C",X"0C",X"0C",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"E9",X"E1",X"F5",X"EA",X"F4",X"E0",X"D4",X"E0",
		X"FD",X"F8",X"F0",X"F0",X"F0",X"C0",X"C0",X"C0",X"E8",X"D0",X"E4",X"D0",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"C6",X"0C",X"00",X"02",X"0A",X"2A",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"52",X"52",X"56",X"D6",X"D3",X"6E",X"EE",X"EE",X"EE",X"AA",X"AA",X"AA",X"AA",
		X"F3",X"F7",X"F7",X"1F",X"03",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"1E",X"00",
		X"16",X"00",X"10",X"11",X"17",X"1F",X"0F",X"0F",X"00",X"06",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"07",X"07",X"03",X"02",X"05",X"02",X"2D",X"95",X"F0",X"FB",X"95",X"B5",X"EA",X"A5",X"52",X"25",
		X"20",X"10",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",X"03",X"07",X"03",X"03",X"03",X"05",X"01",X"03",
		X"3E",X"07",X"A1",X"58",X"D4",X"AA",X"92",X"6D",X"00",X"00",X"04",X"01",X"01",X"03",X"02",X"00",
		X"83",X"81",X"01",X"00",X"89",X"82",X"8B",X"8B",X"66",X"66",X"26",X"23",X"41",X"E3",X"C0",X"40",
		X"8F",X"0D",X"8A",X"97",X"1D",X"0C",X"84",X"84",X"41",X"61",X"60",X"E3",X"31",X"B1",X"93",X"4D",
		X"60",X"70",X"78",X"7C",X"44",X"64",X"40",X"E2",X"0C",X"0E",X"06",X"0A",X"0E",X"06",X"02",X"06",
		X"E1",X"C1",X"C1",X"E1",X"FD",X"80",X"81",X"81",X"16",X"0E",X"0C",X"88",X"18",X"08",X"0C",X"04",
		X"08",X"11",X"11",X"03",X"23",X"01",X"01",X"02",X"00",X"80",X"08",X"00",X"02",X"00",X"00",X"00",
		X"06",X"06",X"04",X"06",X"04",X"0C",X"08",X"10",X"02",X"00",X"10",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"05",X"0D",X"0B",X"3C",X"35",
		X"00",X"00",X"02",X"04",X"06",X"1F",X"3A",X"2F",X"DD",X"D7",X"DD",X"9B",X"DF",X"76",X"5D",X"35",
		X"7A",X"EF",X"BB",X"5A",X"F3",X"BB",X"6E",X"FF",X"C0",X"80",X"E0",X"E0",X"B0",X"A8",X"9C",X"BE",
		X"DB",X"7B",X"7B",X"56",X"FB",X"5F",X"9D",X"DB",X"BD",X"EB",X"7B",X"FA",X"F7",X"BB",X"3B",X"96",
		X"84",X"84",X"86",X"42",X"02",X"20",X"20",X"3C",X"CF",X"EF",X"F7",X"67",X"FF",X"78",X"78",X"7C",
		X"0C",X"8E",X"46",X"C4",X"44",X"E2",X"B0",X"68",X"FE",X"7F",X"2F",X"09",X"08",X"00",X"00",X"00",
		X"80",X"80",X"80",X"00",X"78",X"18",X"98",X"98",X"07",X"07",X"07",X"03",X"01",X"03",X"07",X"1E",
		X"0C",X"06",X"97",X"7B",X"3F",X"0F",X"1F",X"00",X"1C",X"30",X"78",X"3C",X"B6",X"D9",X"D8",X"7C",
		X"80",X"00",X"A0",X"80",X"40",X"A0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"40",X"20",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"03",X"09",X"0F",X"2A",
		X"00",X"00",X"02",X"02",X"0A",X"1A",X"2A",X"29",X"2B",X"A1",X"EB",X"BB",X"AB",X"8D",X"AA",X"AA",
		X"AD",X"7A",X"AD",X"DD",X"B4",X"3B",X"BF",X"AB",X"AF",X"ED",X"EA",X"7F",X"EA",X"67",X"DA",X"6D",
		X"DB",X"BE",X"BB",X"7D",X"AB",X"BB",X"BB",X"75",X"7F",X"F3",X"BA",X"6B",X"6F",X"6E",X"BB",X"7E",
		X"6E",X"FA",X"9E",X"FA",X"EC",X"5C",X"DA",X"BA",X"8B",X"0B",X"0A",X"C4",X"60",X"66",X"67",X"27",
		X"BA",X"6C",X"DE",X"76",X"DD",X"DF",X"D3",X"BD",X"21",X"01",X"21",X"03",X"03",X"03",X"00",X"00",
		X"01",X"41",X"20",X"37",X"11",X"18",X"08",X"08",X"BC",X"EC",X"E7",X"E0",X"E0",X"C0",X"F8",X"F0",
		X"0F",X"0C",X"07",X"03",X"83",X"83",X"03",X"03",X"60",X"60",X"78",X"62",X"FA",X"F2",X"C2",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"0A",
		X"00",X"00",X"01",X"02",X"03",X"01",X"01",X"40",X"2E",X"33",X"FA",X"38",X"9E",X"EE",X"AB",X"2A",
		X"AE",X"A2",X"AA",X"8A",X"8A",X"A9",X"AA",X"6E",X"AA",X"CA",X"AA",X"AA",X"A8",X"AA",X"AB",X"A2",
		X"AA",X"BA",X"F2",X"EA",X"AA",X"AE",X"A9",X"8A",X"EA",X"AF",X"4A",X"3A",X"B8",X"AA",X"AA",X"A2",
		X"F3",X"AF",X"FF",X"F7",X"7D",X"DE",X"D6",X"DF",X"0C",X"2E",X"2E",X"26",X"86",X"82",X"92",X"91",
		X"BD",X"6D",X"F9",X"DB",X"FF",X"77",X"DF",X"5D",X"1B",X"D6",X"D3",X"81",X"A9",X"69",X"48",X"E8",
		X"0F",X"1F",X"3F",X"1F",X"1F",X"7F",X"FF",X"FF",X"7A",X"7C",X"7E",X"7C",X"78",X"60",X"BC",X"BE",
		X"FF",X"6F",X"3F",X"3F",X"0B",X"0F",X"0F",X"23",X"9E",X"9E",X"82",X"C6",X"80",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"24",X"26",X"03",X"C1",X"C1",X"A5",X"25",X"25",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"39",X"2A",X"32",X"36",X"2B",X"3A",X"35",X"31",
		X"10",X"20",X"A0",X"80",X"20",X"22",X"22",X"23",X"7A",X"76",X"7A",X"71",X"72",X"3A",X"1E",X"0E",
		X"F5",X"BE",X"AC",X"FD",X"DB",X"7D",X"FD",X"AD",X"D8",X"E8",X"EE",X"A7",X"FE",X"6B",X"DF",X"FD",
		X"BF",X"77",X"BD",X"9D",X"BF",X"F7",X"6F",X"BD",X"6F",X"CE",X"EF",X"6F",X"E9",X"FC",X"BD",X"ED",
		X"20",X"A0",X"AF",X"BF",X"FC",X"F6",X"FA",X"EF",X"80",X"80",X"80",X"80",X"80",X"C0",X"40",X"40",
		X"F5",X"FE",X"F5",X"FA",X"FD",X"FE",X"F5",X"FB",X"40",X"C0",X"3C",X"D7",X"4A",X"10",X"A8",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"0A",X"08",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"3A",X"32",X"12",X"02",X"00",X"00",X"00",
		X"04",X"04",X"84",X"82",X"A2",X"A6",X"A4",X"24",X"48",X"40",X"48",X"48",X"42",X"42",X"20",X"20",
		X"04",X"25",X"21",X"05",X"14",X"44",X"50",X"54",X"21",X"21",X"22",X"02",X"02",X"82",X"80",X"80",
		X"22",X"12",X"22",X"26",X"24",X"AC",X"A8",X"A1",X"0A",X"0E",X"1E",X"05",X"0A",X"0C",X"0F",X"0E",
		X"81",X"A0",X"B0",X"A4",X"A2",X"21",X"22",X"04",X"06",X"87",X"A3",X"82",X"0B",X"02",X"0E",X"8E",
		X"FF",X"FE",X"FB",X"FD",X"FF",X"FF",X"FD",X"FF",X"AA",X"E8",X"54",X"A4",X"78",X"C2",X"28",X"D4",
		X"FE",X"FB",X"FF",X"FD",X"FF",X"FF",X"FB",X"FE",X"B0",X"C8",X"32",X"60",X"D4",X"68",X"D0",X"A8",
		X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"94",X"94",X"11",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"28",X"29",X"29",X"21",X"00",X"08",X"08",X"2A",X"A6",X"86",X"86",X"1E",X"39",X"3A",X"3E",X"BF",
		X"3B",X"3B",X"3E",X"3B",X"3E",X"36",X"3E",X"1E",X"AE",X"E6",X"A6",X"EA",X"8B",X"BF",X"E9",X"AB",
		X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AB",X"EC",X"82",X"2A",X"3A",X"0B",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AE",X"E2",X"8A",X"2A",X"A9",X"A8",X"AA",X"AA",X"9A",X"AC",X"E8",X"EC",X"A4",X"A8",X"A8",X"28",
		X"9A",X"EE",X"EA",X"AA",X"6A",X"0B",X"02",X"06",X"B9",X"A2",X"AB",X"AA",X"47",X"A7",X"A7",X"AD",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"AB",X"B7",X"27",X"1A",X"07",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DB",X"7D",X"D5",X"FD",X"B6",X"65",X"DE",X"DD",X"DE",X"F7",X"77",X"E4",X"B7",X"B3",X"B6",X"D7",
		X"55",X"7D",X"1D",X"17",X"0D",X"03",X"02",X"00",X"BF",X"F7",X"4F",X"9D",X"D7",X"D7",X"77",X"D9",
		X"A6",X"B6",X"94",X"97",X"37",X"B7",X"1F",X"3B",X"3B",X"27",X"AD",X"16",X"8D",X"9D",X"C7",X"F2",
		X"5A",X"36",X"22",X"20",X"30",X"78",X"F0",X"20",X"F9",X"C8",X"1C",X"2A",X"1F",X"1B",X"FD",X"3D",
		X"E2",X"76",X"66",X"67",X"33",X"A3",X"67",X"F3",X"38",X"1E",X"AC",X"0C",X"0D",X"19",X"31",X"1D",
		X"F7",X"63",X"37",X"33",X"5B",X"9B",X"1F",X"97",X"1A",X"03",X"B1",X"AB",X"11",X"A5",X"33",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"30",X"30",X"3B",X"1B",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F7",X"FD",X"01",X"27",X"00",X"40",X"30",X"3B",X"ED",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"60",X"3C",X"A7",X"83",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",
		X"01",X"00",X"03",X"87",X"0F",X"3F",X"FF",X"FF",X"F0",X"FC",X"01",X"00",X"80",X"80",X"80",X"80",
		X"04",X"03",X"3E",X"FE",X"FE",X"3E",X"00",X"00",X"80",X"FF",X"20",X"00",X"00",X"FF",X"8C",X"8F",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"8F",X"8F",X"FF",X"FF",X"07",X"07",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"C4",X"04",X"0F",
		X"FE",X"FF",X"07",X"07",X"03",X"00",X"00",X"00",X"7F",X"FF",X"FD",X"FD",X"FD",X"0D",X"01",X"07",
		X"FF",X"FF",X"0F",X"07",X"07",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"01",X"FF",X"3F",
		X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3F",X"1B",X"14",X"10",X"10",X"30",
		X"20",X"FF",X"20",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"3F",X"07",X"00",X"00",X"00",X"FC",X"FC",X"FD",X"FD",X"E3",X"C3",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"FD",X"F7",X"F7",X"FD",X"01",X"00",X"FC",X"FC",X"FC",X"FD",X"E1",X"E1",X"C3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"3F",X"A7",X"BF",X"A7",X"B8",X"22",
		X"00",X"07",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"02",X"FE",X"FD",X"FB",X"F7",X"EF",X"DC",X"BC",
		X"FF",X"3F",X"07",X"80",X"C0",X"E0",X"01",X"F9",X"80",X"80",X"80",X"FE",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"03",X"09",
		X"00",X"00",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"07",X"07",X"07",X"07",X"07",X"F8",X"88",X"88",
		X"FC",X"86",X"87",X"FF",X"87",X"87",X"FF",X"FF",X"F8",X"F8",X"60",X"60",X"3F",X"80",X"FF",X"FF",
		X"00",X"FF",X"F8",X"F0",X"F8",X"FF",X"FF",X"55",X"00",X"FF",X"F8",X"F0",X"F8",X"FF",X"FF",X"50",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"80",X"80",X"50",X"50",X"50",X"50",X"50",X"51",X"01",X"01",
		X"00",X"FF",X"FF",X"F8",X"F0",X"F8",X"FF",X"03",X"04",X"F8",X"EF",X"EF",X"FB",X"FB",X"EF",X"EF",
		X"73",X"73",X"F3",X"F3",X"F3",X"F2",X"F2",X"F2",X"FB",X"F8",X"CF",X"CF",X"CF",X"7F",X"7F",X"7F",
		X"5F",X"1F",X"5E",X"1F",X"5F",X"1F",X"5E",X"1F",X"EF",X"FC",X"2C",X"FC",X"EF",X"FC",X"2C",X"FC",
		X"5F",X"1F",X"1F",X"18",X"1F",X"1E",X"1F",X"01",X"EF",X"FF",X"FF",X"FF",X"83",X"7C",X"8E",X"84",
		X"FF",X"08",X"08",X"08",X"F8",X"08",X"08",X"08",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"18",X"F8",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0F",X"03",X"10",X"78",X"3C",X"8E",X"E3",
		X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FE",X"FF",X"7F",X"1F",X"0F",X"03",X"00",
		X"FF",X"FE",X"FD",X"FB",X"33",X"19",X"0C",X"06",X"7F",X"F9",X"F9",X"FF",X"F3",X"F3",X"FF",X"79",
		X"83",X"41",X"20",X"80",X"E0",X"F8",X"FC",X"FE",X"39",X"9F",X"CC",X"64",X"33",X"19",X"0C",X"06",
		X"CF",X"D8",X"D8",X"9F",X"B0",X"B0",X"9F",X"D8",X"8D",X"0D",X"0D",X"8D",X"0D",X"0D",X"8D",X"0D",
		X"D8",X"CF",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"0D",X"8D",X"0B",X"87",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"87",X"87",X"FF",X"87",X"87",X"FF",X"FF",X"FF",X"C3",X"C3",X"FF",X"C3",X"C3",X"FF",
		X"FF",X"FF",X"FF",X"87",X"87",X"FF",X"87",X"87",X"FF",X"FF",X"FF",X"C3",X"C2",X"FC",X"C0",X"C0",
		X"FF",X"FF",X"E1",X"E1",X"FE",X"E0",X"E0",X"F0",X"ED",X"CD",X"8D",X"0D",X"0D",X"0D",X"0F",X"0F",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"0F",X"0D",X"0C",X"0C",X"0E",X"0E",X"0E",X"0E",
		X"F3",X"F3",X"F3",X"9F",X"9F",X"9F",X"FF",X"FF",X"FE",X"FD",X"FB",X"F7",X"EF",X"DF",X"BF",X"3C",
		X"FF",X"1F",X"9F",X"9F",X"E3",X"F3",X"73",X"72",X"9F",X"CF",X"E7",X"F3",X"F9",X"FC",X"FE",X"7F",
		X"01",X"01",X"FF",X"FF",X"87",X"FF",X"FF",X"FF",X"80",X"81",X"B3",X"A3",X"83",X"A3",X"A3",X"83",
		X"FF",X"FF",X"87",X"FF",X"FF",X"01",X"01",X"01",X"A3",X"A3",X"81",X"A0",X"B3",X"81",X"80",X"FC",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"7F",X"3F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",
		X"1E",X"1E",X"1E",X"1E",X"1F",X"1F",X"1E",X"1E",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"FF",X"07",X"00",X"00",X"00",X"00",X"3E",X"FE",X"FE",X"FE",X"7E",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"03",X"00",X"00",
		X"FF",X"7B",X"7B",X"00",X"00",X"00",X"00",X"7B",X"82",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"F0",X"07",X"3F",X"FC",X"FC",X"FF",X"3F",X"07",X"1F",X"E0",X"F7",X"00",X"00",X"F7",X"F7",X"E0",
		X"00",X"F2",X"E7",X"0F",X"1F",X"0D",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"01",X"E7",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"00",X"1F",X"00",X"00",X"3F",X"7F",X"FF",
		X"F1",X"03",X"F3",X"F7",X"87",X"87",X"87",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"00",X"00",X"FF",X"C0",X"C0",X"00",X"4F",X"4F",X"0F",X"00",X"FF",X"83",X"83",X"00",X"9F",X"9F",
		X"0F",X"8F",X"8F",X"8F",X"8F",X"00",X"00",X"F1",X"9F",X"9F",X"9F",X"9F",X"9F",X"00",X"00",X"E3",
		X"B2",X"52",X"53",X"43",X"63",X"33",X"33",X"13",X"7F",X"7F",X"CF",X"CF",X"CF",X"FB",X"FB",X"EF",
		X"13",X"23",X"23",X"23",X"23",X"03",X"03",X"C3",X"EF",X"FB",X"FB",X"EF",X"EF",X"F8",X"C4",X"84",
		X"1F",X"1F",X"1F",X"18",X"1F",X"1F",X"1F",X"5F",X"8E",X"86",X"FF",X"FF",X"FF",X"FF",X"EF",X"FC",
		X"1E",X"5F",X"1F",X"5F",X"1E",X"5F",X"00",X"7F",X"2C",X"FC",X"EF",X"FC",X"2C",X"FC",X"01",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"02",X"07",X"E0",X"E0",X"E0",X"C0",X"C0",X"CA",X"DF",X"FF",
		X"0B",X"07",X"0F",X"3F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DE",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"73",X"71",X"70",X"00",X"00",X"00",X"00",X"00",X"F8",X"F1",X"F1",X"78",X"3C",X"3E",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"F3",X"F3",X"81",X"F1",X"00",X"00",X"FF",X"02",X"E7",X"E7",X"02",X"E3",X"00",X"00",X"FF",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C2",X"C1",X"07",X"C7",X"03",X"02",X"FF",X"0F",X"7D",X"FD",X"FD",X"FD",X"FD",X"1D",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"C0",X"C0",X"C0",X"C1",X"C2",X"C3",X"3F",X"3F",X"07",X"0F",X"3F",X"CF",X"FF",X"FF",
		X"0F",X"07",X"1F",X"0F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"3F",X"2F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"1B",X"07",X"07",X"03",X"05",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"03",X"03",X"07",X"0F",X"07",X"0F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"1F",X"2F",X"1F",X"3F",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"1F",X"2F",X"0F",X"17",X"1F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0B",X"07",X"03",X"05",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"67",X"02",
		X"FE",X"FF",X"FA",X"FF",X"EE",X"FD",X"FB",X"FD",X"AF",X"77",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"BF",X"7F",X"5F",X"17",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"07",X"03",X"05",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"D7",X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"C5",X"A0",X"00",X"FF",X"FF",X"FF",X"3F",X"9F",X"3F",X"0F",X"06",
		X"DF",X"BF",X"EF",X"FF",X"AB",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F7",X"F3",X"D7",X"DB",X"77",X"77",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EF",X"FF",X"EF",X"F7",X"EF",X"F7",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"E9",X"F7",X"F9",X"F3",X"FF",X"EF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"BF",X"DF",X"BF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"FF",X"5F",X"FF",X"FF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"F7",X"FF",X"F7",X"DF",X"F7",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
