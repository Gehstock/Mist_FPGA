library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"88",X"90",X"B9",X"FF",X"FC",X"23",X"77",X"18",X"99",X"89",X"98",X"98",X"9C",X"FB",X"01",
		X"11",X"12",X"11",X"21",X"12",X"22",X"27",X"78",X"E9",X"08",X"00",X"00",X"00",X"54",X"99",X"9A",
		X"F8",X"80",X"00",X"00",X"00",X"15",X"1C",X"A8",X"00",X"08",X"00",X"00",X"15",X"78",X"9A",X"D8",
		X"80",X"00",X"00",X"00",X"17",X"18",X"AD",X"98",X"00",X"01",X"00",X"01",X"54",X"0A",X"CC",X"88",
		X"00",X"10",X"01",X"02",X"72",X"8A",X"E9",X"90",X"00",X"10",X"00",X"13",X"61",X"9C",X"BA",X"80",
		X"01",X"01",X"01",X"24",X"52",X"BD",X"B9",X"80",X"10",X"10",X"11",X"24",X"40",X"BE",X"B9",X"00",
		X"11",X"10",X"02",X"35",X"39",X"EC",X"B8",X"81",X"11",X"21",X"12",X"35",X"1A",X"FC",X"A8",X"81",
		X"12",X"21",X"13",X"34",X"8C",X"FB",X"A8",X"82",X"22",X"33",X"23",X"32",X"AF",X"EB",X"A9",X"01",
		X"32",X"33",X"43",X"31",X"9F",X"CB",X"A9",X"81",X"23",X"33",X"43",X"42",X"8D",X"CC",X"A9",X"81",
		X"12",X"22",X"42",X"32",X"9C",X"EB",X"B9",X"80",X"22",X"33",X"35",X"32",X"8C",X"EB",X"BA",X"80",
		X"22",X"32",X"44",X"32",X"8B",X"DC",X"BB",X"88",X"12",X"24",X"33",X"42",X"0A",X"CD",X"BA",X"98",
		X"11",X"23",X"43",X"33",X"0B",X"DD",X"BB",X"88",X"11",X"42",X"33",X"41",X"0A",X"DC",X"AB",X"80",
		X"02",X"33",X"44",X"21",X"89",X"DC",X"AA",X"91",X"13",X"34",X"32",X"20",X"9C",X"EB",X"C9",X"82",
		X"13",X"35",X"12",X"19",X"AD",X"CB",X"BA",X"01",X"35",X"34",X"22",X"18",X"AF",X"BA",X"C9",X"01",
		X"32",X"43",X"32",X"18",X"AD",X"CC",X"A9",X"91",X"24",X"42",X"32",X"10",X"AC",X"DB",X"CA",X"80",
		X"13",X"43",X"42",X"10",X"9C",X"CB",X"D9",X"90",X"03",X"24",X"33",X"21",X"8B",X"DD",X"B9",X"A8",
		X"12",X"34",X"42",X"31",X"0A",X"CC",X"BC",X"A0",X"00",X"25",X"23",X"31",X"88",X"CC",X"BC",X"9A",
		X"02",X"13",X"53",X"23",X"0A",X"AB",X"DB",X"A8",X"08",X"22",X"43",X"32",X"08",X"AB",X"B9",X"C9",
		X"00",X"22",X"22",X"30",X"19",X"9B",X"A9",X"0B",X"02",X"01",X"31",X"10",X"0A",X"9A",X"A8",X"A8",
		X"02",X"01",X"31",X"19",X"0A",X"9B",X"0C",X"08",X"12",X"02",X"21",X"10",X"8A",X"9B",X"8B",X"08",
		X"38",X"22",X"30",X"18",X"89",X"BA",X"9B",X"80",X"38",X"22",X"20",X"28",X"8A",X"AB",X"8C",X"89",
		X"11",X"31",X"22",X"10",X"89",X"9B",X"9B",X"89",X"10",X"31",X"31",X"20",X"89",X"9A",X"9A",X"0B",
		X"02",X"01",X"21",X"28",X"08",X"8A",X"AA",X"08",X"A2",X"08",X"21",X"20",X"08",X"8A",X"9A",X"0B",
		X"08",X"08",X"08",X"0A",X"28",X"08",X"08",X"0A",X"01",X"98",X"28",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"28",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"91",X"0A",X"2A",X"2A",X"2A",X"28",X"91",X"90",X"1C",X"48",X"A0",X"10",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"89",X"18",X"09",X"10",X"80",X"80",X"89",X"10",X"91",X"80",
		X"8A",X"85",X"B1",X"00",X"A2",X"A2",X"A2",X"B3",X"B3",X"89",X"18",X"00",X"A2",X"80",X"A0",X"80",
		X"82",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"80",X"90",X"80",X"91",X"80",X"80",
		X"02",X"80",X"80",X"00",X"23",X"77",X"FF",X"F7",X"A3",X"98",X"1A",X"18",X"10",X"AA",X"2C",X"83",
		X"8C",X"13",X"B6",X"0A",X"A4",X"00",X"08",X"3A",X"B0",X"0C",X"21",X"B0",X"90",X"00",X"C0",X"40",
		X"1C",X"85",X"8A",X"0A",X"2A",X"AC",X"45",X"A8",X"01",X"AA",X"22",X"2A",X"92",X"12",X"F2",X"81",
		X"1A",X"7F",X"29",X"80",X"F1",X"24",X"A4",X"0A",X"BC",X"31",X"9B",X"13",X"E4",X"A8",X"95",X"88",
		X"08",X"10",X"0D",X"01",X"01",X"92",X"99",X"92",X"A0",X"89",X"49",X"0C",X"29",X"93",X"91",X"C8",
		X"A8",X"08",X"C3",X"21",X"C9",X"04",X"B7",X"C4",X"00",X"18",X"1A",X"89",X"20",X"C2",X"3C",X"9A",
		X"60",X"81",X"D3",X"82",X"F9",X"38",X"09",X"02",X"A0",X"0B",X"89",X"72",X"8C",X"5D",X"59",X"19",
		X"9C",X"93",X"0C",X"7B",X"20",X"A0",X"01",X"18",X"81",X"91",X"98",X"18",X"01",X"D9",X"5D",X"02",
		X"90",X"81",X"82",X"1A",X"BA",X"79",X"00",X"81",X"D1",X"00",X"1A",X"18",X"A4",X"1A",X"09",X"AA",
		X"29",X"18",X"01",X"BC",X"59",X"92",X"0F",X"6A",X"08",X"00",X"00",X"0A",X"21",X"A9",X"68",X"90",
		X"89",X"4A",X"38",X"1D",X"4A",X"1A",X"5A",X"6D",X"3B",X"10",X"A0",X"80",X"91",X"88",X"80",X"18",
		X"B5",X"1F",X"6A",X"81",X"09",X"81",X"09",X"80",X"2B",X"1A",X"29",X"08",X"19",X"B1",X"5C",X"13",
		X"B1",X"81",X"2A",X"2F",X"28",X"0A",X"59",X"1B",X"4F",X"28",X"90",X"93",X"13",X"F9",X"1A",X"30",
		X"87",X"B8",X"18",X"A1",X"09",X"95",X"B1",X"1B",X"B7",X"82",X"C0",X"3C",X"10",X"90",X"02",X"A0",
		X"29",X"02",X"B2",X"97",X"C8",X"01",X"3D",X"12",X"8A",X"83",X"F1",X"8B",X"40",X"9A",X"C3",X"93",
		X"99",X"6B",X"01",X"80",X"A3",X"B3",X"08",X"19",X"00",X"88",X"79",X"2A",X"01",X"0C",X"4A",X"81",
		X"09",X"04",X"9D",X"3F",X"39",X"80",X"09",X"39",X"C4",X"1D",X"20",X"89",X"1A",X"F5",X"99",X"48",
		X"98",X"0A",X"94",X"90",X"08",X"93",X"99",X"93",X"C3",X"09",X"A2",X"4F",X"3F",X"78",X"B0",X"20",
		X"A0",X"8A",X"34",X"B1",X"2A",X"1F",X"39",X"81",X"09",X"19",X"84",X"D2",X"80",X"B6",X"AD",X"5A",
		X"18",X"08",X"80",X"8B",X"49",X"10",X"A2",X"0B",X"54",X"E1",X"A8",X"10",X"84",X"B0",X"08",X"2B",
		X"3C",X"3A",X"09",X"33",X"D4",X"CA",X"23",X"DB",X"70",X"F4",X"89",X"01",X"89",X"81",X"90",X"0F",
		X"69",X"1B",X"20",X"7E",X"19",X"91",X"20",X"A3",X"E3",X"9A",X"24",X"1F",X"03",X"A9",X"1A",X"04",
		X"1A",X"B0",X"98",X"12",X"93",X"7A",X"D2",X"91",X"93",X"92",X"B0",X"10",X"A9",X"4E",X"10",X"10",
		X"98",X"91",X"02",X"C1",X"80",X"0B",X"17",X"9A",X"4D",X"11",X"88",X"09",X"00",X"08",X"18",X"9A",
		X"03",X"1D",X"13",X"A8",X"1C",X"1A",X"15",X"99",X"12",X"91",X"CA",X"13",X"A7",X"C1",X"00",X"B0",
		X"22",X"AE",X"20",X"08",X"81",X"A2",X"88",X"F4",X"1B",X"2F",X"30",X"98",X"00",X"91",X"88",X"02",
		X"89",X"1B",X"10",X"1B",X"23",X"83",X"F9",X"08",X"46",X"D8",X"19",X"89",X"17",X"D1",X"92",X"00",
		X"B3",X"8B",X"39",X"93",X"19",X"A8",X"01",X"2F",X"39",X"A1",X"2D",X"38",X"09",X"81",X"8B",X"22",
		X"19",X"79",X"B0",X"13",X"F7",X"0F",X"7C",X"29",X"81",X"80",X"88",X"00",X"88",X"18",X"90",X"81",
		X"88",X"00",X"91",X"88",X"8A",X"47",X"9A",X"B6",X"A0",X"92",X"09",X"2A",X"08",X"88",X"21",X"98",
		X"0F",X"38",X"20",X"AB",X"12",X"09",X"09",X"21",X"1A",X"C2",X"9D",X"59",X"88",X"3A",X"08",X"0D",
		X"21",X"19",X"20",X"8B",X"3C",X"1F",X"1F",X"7F",X"7F",X"02",X"82",X"91",X"C2",X"89",X"94",X"C2",
		X"90",X"00",X"C9",X"78",X"B5",X"A1",X"2B",X"2A",X"3C",X"40",X"F4",X"C2",X"09",X"82",X"98",X"8A",
		X"6A",X"19",X"28",X"A3",X"9A",X"05",X"B1",X"3D",X"18",X"A1",X"83",X"B8",X"2B",X"14",X"C8",X"2B",
		X"7A",X"81",X"81",X"A2",X"09",X"02",X"B7",X"A8",X"81",X"81",X"D3",X"09",X"2A",X"08",X"88",X"3A",
		X"20",X"C8",X"49",X"9A",X"04",X"BF",X"40",X"09",X"14",X"AA",X"C1",X"23",X"A0",X"A3",X"9E",X"1F",
		X"10",X"90",X"81",X"B7",X"90",X"29",X"08",X"10",X"88",X"81",X"8B",X"4B",X"12",X"B9",X"22",X"7C",
		X"08",X"88",X"2C",X"81",X"80",X"1B",X"40",X"B8",X"4D",X"4A",X"1E",X"39",X"81",X"1C",X"2A",X"93",
		X"9C",X"79",X"81",X"91",X"81",X"89",X"09",X"58",X"82",X"88",X"0A",X"80",X"09",X"81",X"A3",X"B0",
		X"E2",X"80",X"27",X"99",X"31",X"F0",X"91",X"8B",X"11",X"11",X"88",X"AB",X"7A",X"01",X"B1",X"2D",
		X"1B",X"89",X"32",X"F3",X"2C",X"02",X"92",X"93",X"40",X"9C",X"19",X"92",X"AA",X"4B",X"38",X"88",
		X"0F",X"7A",X"04",X"AB",X"21",X"7E",X"21",X"3E",X"A2",X"AA",X"F6",X"98",X"39",X"10",X"0A",X"09",
		X"90",X"02",X"AA",X"02",X"59",X"B8",X"38",X"B1",X"2F",X"5D",X"48",X"98",X"3C",X"3B",X"10",X"0B",
		X"29",X"22",X"8E",X"48",X"B2",X"1D",X"10",X"88",X"19",X"00",X"88",X"81",X"90",X"28",X"A1",X"80",
		X"8B",X"F3",X"38",X"1F",X"10",X"97",X"98",X"87",X"F0",X"10",X"88",X"83",X"85",X"F1",X"29",X"9A",
		X"01",X"91",X"B5",X"0A",X"82",X"B3",X"88",X"68",X"A0",X"29",X"A9",X"08",X"8A",X"48",X"96",X"A9",
		X"28",X"81",X"B1",X"3A",X"C5",X"8E",X"4A",X"10",X"0A",X"39",X"89",X"10",X"82",X"A8",X"90",X"7B",
		X"57",X"F5",X"B8",X"90",X"49",X"39",X"AE",X"22",X"09",X"B8",X"25",X"1C",X"99",X"32",X"8C",X"13",
		X"E0",X"10",X"88",X"91",X"28",X"C0",X"20",X"8B",X"40",X"C1",X"81",X"0B",X"82",X"01",X"8D",X"06",
		X"99",X"08",X"10",X"B1",X"39",X"B2",X"3B",X"02",X"F2",X"19",X"99",X"48",X"8A",X"1A",X"7B",X"18",
		X"3B",X"0A",X"15",X"BC",X"69",X"0A",X"38",X"90",X"90",X"49",X"99",X"31",X"BB",X"21",X"12",X"F0",
		X"5A",X"88",X"82",X"80",X"B1",X"29",X"89",X"13",X"BF",X"05",X"90",X"91",X"23",X"BF",X"84",X"8D",
		X"11",X"00",X"A0",X"08",X"A0",X"78",X"89",X"02",X"9E",X"18",X"10",X"A1",X"12",X"B9",X"17",X"C1",
		X"09",X"18",X"85",X"B8",X"A1",X"03",X"AC",X"70",X"A1",X"88",X"1C",X"01",X"8A",X"06",X"8A",X"1A",
		X"13",X"B9",X"5B",X"02",X"9A",X"01",X"C5",X"88",X"39",X"91",X"1A",X"D9",X"30",X"5A",X"91",X"3A",
		X"F2",X"19",X"83",X"3D",X"B2",X"D3",X"1B",X"48",X"A1",X"2A",X"A8",X"20",X"99",X"5C",X"B5",X"4D",
		X"88",X"87",X"99",X"29",X"80",X"1A",X"10",X"98",X"2A",X"95",X"A8",X"7B",X"92",X"1C",X"29",X"A6",
		X"19",X"90",X"91",X"98",X"0B",X"80",X"7F",X"36",X"F3",X"97",X"D1",X"0A",X"08",X"23",X"F0",X"29",
		X"2D",X"12",X"D4",X"B1",X"0A",X"2A",X"29",X"3B",X"21",X"A9",X"92",X"09",X"12",X"C1",X"19",X"8B",
		X"79",X"83",X"E3",X"A8",X"81",X"1A",X"02",X"0C",X"2C",X"03",X"D3",X"90",X"38",X"0A",X"0B",X"11",
		X"C2",X"8C",X"7A",X"12",X"E1",X"80",X"18",X"08",X"09",X"00",X"97",X"D2",X"90",X"11",X"C9",X"5B",
		X"28",X"81",X"A0",X"1A",X"4B",X"00",X"09",X"29",X"80",X"18",X"92",X"88",X"90",X"7F",X"3A",X"18",
		X"00",X"8A",X"21",X"B9",X"69",X"A0",X"22",X"81",X"F7",X"F8",X"21",X"28",X"B8",X"0B",X"7A",X"91",
		X"09",X"4A",X"C6",X"A1",X"00",X"88",X"91",X"81",X"B2",X"1B",X"28",X"09",X"08",X"82",X"B1",X"88",
		X"4C",X"68",X"E1",X"83",X"0A",X"90",X"91",X"1A",X"13",X"9A",X"1B",X"7D",X"3A",X"03",X"9A",X"10",
		X"C1",X"09",X"13",X"3F",X"21",X"AA",X"A2",X"27",X"AA",X"93",X"A3",X"C0",X"13",X"3F",X"81",X"8A",
		X"07",X"8A",X"09",X"12",X"B8",X"3C",X"2A",X"38",X"D3",X"1B",X"D2",X"31",X"91",X"AF",X"49",X"88",
		X"18",X"10",X"8F",X"20",X"19",X"A1",X"92",X"09",X"01",X"88",X"8B",X"42",X"C4",X"F2",X"09",X"19",
		X"19",X"28",X"B2",X"90",X"48",X"A1",X"AD",X"7E",X"28",X"00",X"81",X"99",X"29",X"1A",X"19",X"07",
		X"BA",X"49",X"93",X"98",X"7F",X"3C",X"84",X"0C",X"6B",X"5B",X"1A",X"28",X"91",X"88",X"2C",X"A7",
		X"A0",X"29",X"08",X"2A",X"A5",X"C2",X"1A",X"83",X"A0",X"B4",X"0C",X"28",X"0A",X"3C",X"21",X"B2",
		X"89",X"01",X"0B",X"A7",X"A1",X"29",X"E1",X"10",X"C4",X"90",X"2A",X"08",X"89",X"29",X"08",X"59",
		X"88",X"80",X"2E",X"4C",X"3B",X"4B",X"02",X"91",X"1A",X"4C",X"81",X"90",X"B3",X"A4",X"0B",X"14",
		X"F2",X"0A",X"01",X"80",X"98",X"2A",X"18",X"1C",X"5A",X"2A",X"01",X"1C",X"00",X"1A",X"C7",X"A0",
		X"91",X"29",X"89",X"10",X"01",X"08",X"10",X"3C",X"03",X"F2",X"2B",X"B4",X"4B",X"88",X"B3",X"80",
		X"80",X"14",X"9F",X"80",X"10",X"C6",X"A1",X"99",X"18",X"2A",X"3B",X"80",X"20",X"B0",X"29",X"19",
		X"98",X"10",X"3D",X"20",X"7F",X"3A",X"19",X"4B",X"00",X"92",X"90",X"09",X"08",X"08",X"89",X"82",
		X"C0",X"18",X"20",X"C3",X"A8",X"12",X"A8",X"92",X"A4",X"83",X"B0",X"80",X"8A",X"29",X"10",X"81",
		X"C8",X"4B",X"12",X"8A",X"2C",X"13",X"88",X"B3",X"98",X"6C",X"10",X"3E",X"10",X"98",X"83",X"9B",
		X"13",X"D2",X"09",X"90",X"09",X"31",X"C3",X"B3",X"80",X"8B",X"3A",X"02",X"81",X"C2",X"08",X"08",
		X"91",X"08",X"00",X"88",X"08",X"00",X"8A",X"2A",X"01",X"2C",X"83",X"B3",X"2F",X"00",X"10",X"08",
		X"88",X"91",X"98",X"2B",X"4A",X"12",X"C9",X"82",X"38",X"C1",X"81",X"90",X"92",X"0A",X"00",X"80",
		X"80",X"82",X"A2",X"A8",X"29",X"10",X"80",X"81",X"91",X"90",X"80",X"82",X"C7",X"C1",X"09",X"19",
		X"80",X"80",X"02",X"B1",X"82",X"11",X"BA",X"68",X"0A",X"89",X"82",X"80",X"A2",X"A8",X"C2",X"3B",
		X"19",X"01",X"05",X"F2",X"91",X"89",X"12",X"C1",X"90",X"18",X"11",X"91",X"89",X"08",X"01",X"88",
		X"81",X"99",X"18",X"A4",X"B3",X"99",X"1A",X"02",X"80",X"A2",X"A2",X"B8",X"11",X"88",X"18",X"90",
		X"A2",X"88",X"3B",X"92",X"17",X"9A",X"C4",X"A0",X"F7",X"90",X"1B",X"18",X"80",X"91",X"80",X"80",
		X"91",X"21",X"98",X"2A",X"80",X"89",X"37",X"9F",X"01",X"3C",X"80",X"01",X"98",X"81",X"08",X"98",
		X"23",X"F2",X"C4",X"A2",X"80",X"0B",X"09",X"3A",X"1B",X"A4",X"1B",X"3B",X"4A",X"09",X"21",X"89",
		X"10",X"80",X"C4",X"88",X"48",X"DB",X"83",X"F7",X"0C",X"21",X"C0",X"02",X"B1",X"3B",X"00",X"90",
		X"19",X"19",X"08",X"80",X"2B",X"2B",X"11",X"10",X"B8",X"27",X"FB",X"77",X"FA",X"97",X"3A",X"98",
		X"9B",X"53",X"8E",X"A2",X"33",X"BA",X"B0",X"25",X"2B",X"C9",X"32",X"2C",X"A9",X"22",X"3A",X"BB",
		X"84",X"41",X"BC",X"82",X"30",X"BB",X"00",X"35",X"AA",X"B1",X"36",X"99",X"B0",X"13",X"1A",X"BA",
		X"13",X"79",X"B9",X"21",X"22",X"F9",X"18",X"20",X"0B",X"81",X"01",X"3E",X"88",X"03",X"0A",X"A1",
		X"91",X"69",X"C0",X"11",X"00",X"C1",X"1A",X"92",X"3F",X"2B",X"58",X"8A",X"10",X"91",X"1B",X"13",
		X"A9",X"3B",X"A3",X"B0",X"70",X"9B",X"08",X"78",X"0B",X"81",X"00",X"09",X"08",X"A2",X"79",X"B9",
		X"19",X"71",X"F1",X"1A",X"08",X"2A",X"91",X"28",X"A0",X"14",X"C0",X"93",X"89",X"82",X"C8",X"0F",
		X"AF",X"35",X"13",X"10",X"DA",X"C8",X"10",X"09",X"00",X"11",X"8A",X"A2",X"04",X"84",X"8B",X"81",
		X"31",X"C9",X"94",X"A1",X"80",X"D1",X"08",X"10",X"08",X"01",X"87",X"77",X"FF",X"C3",X"53",X"E8",
		X"01",X"00",X"1C",X"80",X"14",X"8B",X"B0",X"22",X"19",X"BC",X"03",X"40",X"C9",X"81",X"21",X"BA",
		X"12",X"11",X"9D",X"80",X"35",X"9B",X"98",X"14",X"19",X"CA",X"22",X"18",X"81",X"A0",X"99",X"2A",
		X"B7",X"39",X"BC",X"13",X"39",X"0C",X"A0",X"16",X"8A",X"A2",X"93",X"1A",X"9B",X"03",X"78",X"9D",
		X"01",X"18",X"98",X"92",X"01",X"0B",X"00",X"93",X"90",X"F5",X"A0",X"2B",X"01",X"2D",X"28",X"12",
		X"E9",X"11",X"19",X"2A",X"8A",X"90",X"78",X"B8",X"06",X"8A",X"92",X"12",X"D9",X"32",X"C9",X"86",
		X"9A",X"A2",X"28",X"0B",X"30",X"B8",X"07",X"89",X"A2",X"08",X"B8",X"58",X"8B",X"03",X"1A",X"B3",
		X"0C",X"08",X"21",X"B8",X"B3",X"78",X"88",X"81",X"90",X"88",X"08",X"92",X"3A",X"D2",X"01",X"88",
		X"BB",X"45",X"A2",X"9B",X"90",X"38",X"08",X"A9",X"21",X"0A",X"09",X"00",X"24",X"F1",X"89",X"07",
		X"D3",X"8A",X"18",X"08",X"80",X"00",X"89",X"90",X"12",X"80",X"A8",X"00",X"10",X"19",X"91",X"03",
		X"A9",X"80",X"80",X"80",X"8B",X"81",X"29",X"A0",X"14",X"88",X"B2",X"8A",X"03",X"99",X"93",X"8A",
		X"80",X"93",X"29",X"80",X"A8",X"21",X"88",X"B2",X"00",X"A2",X"81",X"90",X"81",X"99",X"93",X"80",
		X"89",X"82",X"0A",X"1B",X"01",X"A4",X"A8",X"03",X"90",X"A9",X"12",X"89",X"88",X"02",X"A0",X"82",
		X"A9",X"87",X"5F",X"11",X"B2",X"90",X"08",X"08",X"08",X"08",X"08",X"A5",X"B8",X"3B",X"3B",X"03",
		X"0D",X"02",X"A2",X"0A",X"28",X"B8",X"78",X"F4",X"B3",X"9A",X"5B",X"10",X"80",X"80",X"00",X"89",
		X"19",X"81",X"90",X"19",X"10",X"80",X"A8",X"09",X"70",X"F4",X"A8",X"18",X"08",X"09",X"18",X"08",
		X"09",X"11",X"80",X"88",X"99",X"11",X"08",X"0A",X"2A",X"20",X"A8",X"80",X"28",X"91",X"99",X"38",
		X"0A",X"01",X"91",X"89",X"2A",X"01",X"98",X"01",X"08",X"19",X"0A",X"80",X"28",X"09",X"18",X"91",
		X"0A",X"28",X"08",X"98",X"28",X"08",X"08",X"93",X"9C",X"04",X"88",X"80",X"80",X"8A",X"03",X"8A",
		X"90",X"48",X"C2",X"B7",X"99",X"82",X"0A",X"01",X"0B",X"39",X"00",X"89",X"10",X"A0",X"83",X"90",
		X"A2",X"8A",X"00",X"19",X"93",X"A2",X"A2",X"A0",X"10",X"80",X"80",X"89",X"91",X"A7",X"B3",X"1F",
		X"28",X"09",X"80",X"28",X"A3",X"8B",X"95",X"A1",X"98",X"10",X"80",X"C2",X"82",X"A2",X"88",X"90",
		X"82",X"B0",X"29",X"82",X"80",X"89",X"10",X"80",X"80",X"A2",X"80",X"89",X"19",X"10",X"C1",X"83",
		X"B3",X"08",X"C1",X"20",X"80",X"80",X"8A",X"20",X"A0",X"10",X"80",X"89",X"10",X"8A",X"02",X"80",
		X"80",X"80",X"A0",X"89",X"40",X"D2",X"1A",X"10",X"80",X"80",X"80",X"A0",X"82",X"89",X"18",X"00",
		X"80",X"89",X"19",X"01",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"82",X"80",X"89",X"10",X"B1",
		X"92",X"90",X"80",X"82",X"A0",X"89",X"30",X"08",X"08",X"08",X"80",X"82",X"80",X"A0",X"89",X"91",
		X"80",X"10",X"A2",X"A1",X"00",X"80",X"80",X"89",X"80",X"90",X"7F",X"FE",X"13",X"62",X"32",X"F9",
		X"98",X"09",X"99",X"11",X"19",X"89",X"01",X"52",X"8A",X"80",X"31",X"09",X"A8",X"03",X"8C",X"B8",
		X"23",X"19",X"EA",X"02",X"48",X"BB",X"91",X"32",X"DB",X"84",X"82",X"39",X"A2",X"B5",X"AC",X"81",
		X"52",X"8B",X"C0",X"12",X"38",X"AB",X"B2",X"08",X"D9",X"27",X"02",X"99",X"98",X"20",X"1A",X"88",
		X"00",X"88",X"0A",X"88",X"38",X"08",X"91",X"19",X"B8",X"2D",X"20",X"33",X"89",X"29",X"19",X"BA",
		X"88",X"01",X"30",X"89",X"91",X"0A",X"89",X"01",X"08",X"2A",X"01",X"18",X"08",X"00",X"28",X"9A",
		X"99",X"38",X"A2",X"08",X"08",X"A3",X"C1",X"09",X"5B",X"0A",X"01",X"88",X"3A",X"10",X"08",X"0A",
		X"88",X"00",X"08",X"91",X"10",X"08",X"19",X"08",X"08",X"08",X"18",X"08",X"8A",X"28",X"98",X"80",
		X"28",X"08",X"08",X"91",X"90",X"18",X"08",X"08",X"98",X"08",X"08",X"08",X"09",X"19",X"00",X"08",
		X"28",X"08",X"08",X"91",X"08",X"08",X"08",X"08",X"19",X"08",X"0A",X"08",X"08",X"28",X"08",X"08",
		X"08",X"08",X"08",X"08",X"0A",X"01",X"99",X"00",X"7F",X"F7",X"71",X"FA",X"33",X"8E",X"93",X"19",
		X"88",X"88",X"02",X"29",X"E8",X"32",X"9A",X"01",X"88",X"03",X"AE",X"84",X"2A",X"99",X"81",X"20",
		X"8B",X"98",X"42",X"8C",X"99",X"35",X"9A",X"A3",X"B4",X"4A",X"AA",X"13",X"28",X"E0",X"80",X"30",
		X"8C",X"90",X"61",X"BA",X"83",X"01",X"B8",X"00",X"21",X"0F",X"10",X"0A",X"11",X"91",X"B8",X"33",
		X"CA",X"10",X"5A",X"8B",X"42",X"8C",X"B2",X"79",X"89",X"13",X"C3",X"C1",X"90",X"02",X"1D",X"90",
		X"58",X"9A",X"94",X"18",X"B0",X"02",X"A1",X"4A",X"BB",X"63",X"9A",X"A0",X"20",X"1A",X"0C",X"05",
		X"93",X"B8",X"B0",X"31",X"2F",X"82",X"19",X"89",X"10",X"F2",X"28",X"AB",X"21",X"39",X"B8",X"05",
		X"A0",X"A1",X"10",X"B5",X"98",X"B3",X"28",X"8B",X"02",X"19",X"B1",X"19",X"28",X"80",X"80",X"A2",
		X"A2",X"80",X"C1",X"48",X"B9",X"03",X"08",X"C3",X"08",X"98",X"0A",X"21",X"19",X"9A",X"14",X"89",
		X"B3",X"08",X"0A",X"28",X"08",X"08",X"8A",X"18",X"2A",X"01",X"A2",X"18",X"B0",X"08",X"28",X"0A",
		X"1A",X"3A",X"08",X"80",X"21",X"98",X"99",X"49",X"2C",X"08",X"21",X"89",X"B1",X"21",X"98",X"99",
		X"02",X"0A",X"88",X"38",X"08",X"9A",X"40",X"1A",X"9A",X"21",X"3B",X"A9",X"14",X"0B",X"90",X"39",
		X"08",X"0C",X"12",X"08",X"A0",X"93",X"0C",X"30",X"A2",X"90",X"81",X"91",X"08",X"91",X"19",X"08",
		X"08",X"91",X"0A",X"08",X"28",X"08",X"99",X"12",X"09",X"99",X"38",X"0B",X"11",X"08",X"08",X"00",
		X"B8",X"30",X"8A",X"08",X"28",X"08",X"98",X"08",X"28",X"98",X"01",X"08",X"91",X"0A",X"01",X"08",
		X"98",X"01",X"98",X"28",X"08",X"08",X"90",X"10",X"88",X"08",X"08",X"08",X"98",X"82",X"08",X"0B",
		X"10",X"3A",X"90",X"82",X"09",X"89",X"28",X"78",X"FB",X"2C",X"25",X"24",X"90",X"09",X"9D",X"8D",
		X"91",X"00",X"83",X"90",X"02",X"00",X"A3",X"32",X"A9",X"A2",X"05",X"09",X"DB",X"04",X"2A",X"99",
		X"32",X"0B",X"A9",X"08",X"2A",X"BC",X"91",X"18",X"38",X"08",X"60",X"99",X"A0",X"13",X"09",X"80",
		X"10",X"98",X"89",X"82",X"80",X"C0",X"B3",X"81",X"02",X"01",X"80",X"90",X"09",X"10",X"A0",X"A0",
		X"91",X"88",X"90",X"03",X"0A",X"89",X"00",X"8B",X"33",X"89",X"12",X"81",X"99",X"80",X"A2",X"A6",
		X"F0",X"2A",X"3A",X"83",X"90",X"71",X"3F",X"B2",X"80",X"9B",X"18",X"42",X"A9",X"80",X"11",X"81",
		X"2A",X"A6",X"19",X"C8",X"23",X"9B",X"81",X"08",X"21",X"DA",X"02",X"29",X"9B",X"A2",X"00",X"0C",
		X"83",X"12",X"0A",X"80",X"28",X"49",X"A8",X"03",X"99",X"88",X"08",X"1B",X"89",X"00",X"18",X"0A",
		X"58",X"00",X"0A",X"00",X"00",X"88",X"8A",X"08",X"08",X"90",X"81",X"2A",X"09",X"18",X"2A",X"01",
		X"90",X"10",X"FF",X"57",X"8B",X"A1",X"21",X"B9",X"00",X"02",X"0C",X"A1",X"33",X"9B",X"A2",X"21",
		X"11",X"CD",X"13",X"2B",X"B9",X"41",X"81",X"8F",X"A4",X"28",X"B9",X"11",X"08",X"18",X"BD",X"51",
		X"8B",X"0A",X"26",X"8A",X"90",X"05",X"89",X"98",X"82",X"01",X"AB",X"05",X"1B",X"99",X"02",X"08",
		X"08",X"08",X"19",X"91",X"0A",X"92",X"1A",X"08",X"88",X"33",X"FF",X"63",X"8D",X"B2",X"31",X"BB",
		X"10",X"11",X"8B",X"99",X"62",X"8B",X"91",X"21",X"90",X"9A",X"02",X"4B",X"B8",X"12",X"01",X"AF",
		X"84",X"29",X"A9",X"01",X"11",X"88",X"C1",X"30",X"90",X"A9",X"34",X"9C",X"90",X"14",X"9B",X"08",
		X"08",X"28",X"0C",X"04",X"09",X"0F",X"F7",X"10",X"BB",X"22",X"2B",X"B0",X"02",X"18",X"AB",X"86",
		X"18",X"9B",X"21",X"28",X"89",X"B0",X"24",X"9D",X"82",X"01",X"2B",X"B8",X"34",X"A9",X"B8",X"31",
		X"90",X"A8",X"83",X"80",X"A0",X"A2",X"10",X"A9",X"03",X"FC",X"71",X"1B",X"C2",X"12",X"AB",X"80",
		X"30",X"8C",X"80",X"33",X"99",X"B1",X"21",X"29",X"AC",X"12",X"4A",X"9A",X"28",X"10",X"9A",X"82",
		X"28",X"9A",X"88",X"11",X"08",X"8F",X"B7",X"31",X"CC",X"12",X"18",X"C8",X"01",X"11",X"BA",X"83",
		X"40",X"9B",X"02",X"29",X"93",X"F8",X"12",X"89",X"A1",X"21",X"0A",X"CA",X"33",X"10",X"B9",X"38",
		X"92",X"AA",X"F4",X"50",X"9D",X"82",X"18",X"A8",X"00",X"12",X"AA",X"B3",X"32",X"AA",X"2B",X"38",
		X"19",X"A9",X"13",X"09",X"99",X"11",X"18",X"88",X"B3",X"2E",X"B7",X"11",X"BD",X"83",X"18",X"09",
		X"24",X"01",X"AA",X"9B",X"BB",X"8B",X"0B",X"22",X"10",X"A2",X"34",X"08",X"00",X"82",X"10",X"C8",
		X"03",X"1B",X"98",X"82",X"A8",X"18",X"A8",X"21",X"98",X"B2",X"80",X"88",X"81",X"83",X"98",X"92",
		X"89",X"19",X"01",X"80",X"89",X"1A",X"20",X"80",X"B0",X"02",X"A9",X"18",X"81",X"01",X"91",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"89",X"96",X"B1",X"18",X"B3",X"B3",X"80",X"89",X"10",X"80",
		X"A2",X"A2",X"B1",X"10",X"80",X"80",X"81",X"9F",X"32",X"B9",X"02",X"09",X"10",X"19",X"88",X"A0",
		X"2F",X"58",X"A0",X"80",X"A2",X"22",X"19",X"08",X"3A",X"0B",X"0A",X"0C",X"08",X"B8",X"18",X"3B",
		X"08",X"85",X"11",X"B9",X"08",X"30",X"12",X"A8",X"81",X"80",X"81",X"90",X"98",X"80",X"81",X"92",
		X"D2",X"91",X"08",X"08",X"98",X"08",X"08",X"08",X"08",X"08",X"08",X"28",X"0A",X"08",X"28",X"08",
		X"91",X"08",X"08",X"08",X"19",X"08",X"08",X"08",X"08",X"08",X"91",X"91",X"08",X"0A",X"01",X"80",
		X"08",X"0A",X"2A",X"28",X"08",X"98",X"2A",X"28",X"0A",X"28",X"0A",X"01",X"91",X"08",X"08",X"0A",
		X"28",X"08",X"98",X"01",X"91",X"08",X"08",X"08",X"0A",X"2A",X"28",X"08",X"90",X"18",X"08",X"08",
		X"90",X"18",X"08",X"08",X"08",X"0A",X"28",X"B1",X"08",X"2A",X"28",X"98",X"01",X"08",X"08",X"08",
		X"08",X"08",X"0A",X"08",X"08",X"09",X"08",X"00",X"08",X"08",X"28",X"08",X"10",X"08",X"28",X"08",
		X"0A",X"09",X"8A",X"89",X"08",X"08",X"08",X"00",X"08",X"19",X"19",X"88",X"07",X"FF",X"7D",X"1F",
		X"6C",X"13",X"84",X"89",X"98",X"C9",X"02",X"B2",X"90",X"39",X"C3",X"92",X"69",X"59",X"90",X"90",
		X"88",X"82",X"90",X"19",X"2B",X"08",X"29",X"88",X"B0",X"0D",X"99",X"A2",X"F9",X"10",X"28",X"A1",
		X"A8",X"68",X"01",X"8F",X"79",X"92",X"2A",X"18",X"82",X"92",X"A9",X"2D",X"00",X"80",X"0A",X"79",
		X"88",X"18",X"02",X"88",X"29",X"9B",X"09",X"B9",X"84",X"98",X"A5",X"FA",X"19",X"00",X"00",X"A1",
		X"70",X"80",X"11",X"B1",X"90",X"0B",X"2E",X"08",X"19",X"B2",X"6C",X"48",X"08",X"17",X"89",X"1B",
		X"5A",X"19",X"19",X"92",X"09",X"8A",X"79",X"91",X"A2",X"A0",X"CF",X"3D",X"70",X"B9",X"38",X"B1",
		X"08",X"91",X"19",X"00",X"00",X"85",X"C1",X"12",X"B2",X"A1",X"90",X"68",X"E1",X"13",X"89",X"11",
		X"A2",X"9B",X"11",X"8A",X"1A",X"B2",X"F0",X"0A",X"88",X"B8",X"02",X"70",X"B0",X"89",X"AC",X"30",
		X"80",X"8B",X"58",X"23",X"D8",X"85",X"0B",X"1B",X"AA",X"78",X"00",X"02",X"02",X"A1",X"4A",X"40",
		X"D3",X"21",X"F4",X"B2",X"A8",X"19",X"1D",X"33",X"F8",X"7B",X"81",X"08",X"A2",X"0B",X"28",X"D3",
		X"91",X"A0",X"81",X"58",X"C1",X"00",X"90",X"18",X"49",X"B2",X"11",X"A1",X"53",X"88",X"2C",X"04",
		X"CA",X"38",X"C6",X"98",X"0B",X"0A",X"19",X"0D",X"1B",X"24",X"0C",X"01",X"C0",X"8A",X"28",X"A9",
		X"10",X"30",X"C4",X"49",X"59",X"82",X"82",X"A0",X"9F",X"29",X"20",X"28",X"A8",X"A7",X"8A",X"58",
		X"80",X"98",X"B3",X"37",X"A2",X"D8",X"A1",X"08",X"A0",X"81",X"09",X"19",X"8A",X"20",X"C1",X"24",
		X"E3",X"10",X"9A",X"9B",X"30",X"CB",X"21",X"9A",X"48",X"03",X"01",X"20",X"31",X"91",X"18",X"00",
		X"88",X"1A",X"19",X"81",X"88",X"08",X"0A",X"0C",X"28",X"9A",X"10",X"CA",X"08",X"88",X"B3",X"03",
		X"08",X"08",X"29",X"88",X"08",X"05",X"F3",X"98",X"88",X"18",X"2A",X"23",X"B1",X"D8",X"15",X"C8",
		X"49",X"7F",X"5C",X"03",X"A8",X"00",X"80",X"88",X"18",X"89",X"28",X"09",X"98",X"59",X"00",X"B3",
		X"90",X"19",X"A0",X"38",X"D3",X"B2",X"E5",X"A9",X"3B",X"19",X"4A",X"20",X"88",X"80",X"A2",X"82",
		X"89",X"81",X"0D",X"29",X"88",X"83",X"A0",X"91",X"09",X"6C",X"28",X"C1",X"59",X"B3",X"A1",X"88",
		X"81",X"08",X"20",X"80",X"30",X"A8",X"00",X"91",X"9A",X"38",X"91",X"91",X"C2",X"08",X"01",X"B1",
		X"0A",X"28",X"99",X"3A",X"28",X"1B",X"28",X"08",X"9A",X"48",X"0A",X"09",X"38",X"03",X"F1",X"09",
		X"83",X"88",X"19",X"A0",X"90",X"91",X"92",X"A0",X"01",X"80",X"39",X"08",X"08",X"87",X"FF",X"97",
		X"9F",X"6A",X"06",X"99",X"1A",X"92",X"A0",X"2C",X"3A",X"00",X"81",X"88",X"08",X"7B",X"38",X"91",
		X"88",X"01",X"B0",X"81",X"E3",X"A4",X"B1",X"98",X"0F",X"48",X"00",X"0B",X"20",X"D1",X"10",X"09",
		X"91",X"90",X"A7",X"A1",X"2A",X"94",X"0C",X"3A",X"A7",X"A0",X"1A",X"2A",X"19",X"09",X"01",X"93",
		X"A8",X"98",X"20",X"00",X"79",X"90",X"1B",X"A8",X"7A",X"D5",X"89",X"19",X"92",X"91",X"0B",X"28",
		X"B5",X"82",X"2F",X"10",X"A2",X"88",X"81",X"0B",X"82",X"A1",X"19",X"31",X"4F",X"3B",X"3A",X"19",
		X"A5",X"91",X"19",X"9A",X"83",X"98",X"92",X"A2",X"B2",X"8C",X"0A",X"4F",X"4A",X"1C",X"2A",X"80",
		X"79",X"88",X"1B",X"30",X"8A",X"38",X"1D",X"10",X"A3",X"00",X"6C",X"82",X"01",X"8A",X"32",X"82",
		X"8A",X"80",X"A0",X"8A",X"59",X"99",X"97",X"E2",X"8A",X"29",X"93",X"8A",X"19",X"A2",X"B4",X"B6",
		X"E2",X"09",X"02",X"A2",X"89",X"7D",X"01",X"81",X"98",X"0A",X"20",X"4C",X"69",X"91",X"89",X"88",
		X"28",X"2A",X"4A",X"90",X"19",X"89",X"08",X"29",X"8B",X"3A",X"28",X"9A",X"08",X"08",X"08",X"19",
		X"08",X"01",X"89",X"40",X"C3",X"B1",X"28",X"92",X"80",X"39",X"1C",X"18",X"83",X"A0",X"0A",X"28",
		X"0A",X"19",X"11",X"98",X"88",X"08",X"91",X"F7",X"E3",X"98",X"18",X"91",X"88",X"10",X"A1",X"80",
		X"90",X"81",X"88",X"18",X"83",X"80",X"80",X"81",X"99",X"10",X"80",X"80",X"80",X"81",X"00",X"80",
		X"10",X"A2",X"B0",X"81",X"A1",X"88",X"19",X"A2",X"8A",X"81",X"A0",X"01",X"1B",X"08",X"82",X"A0",
		X"39",X"19",X"10",X"B0",X"02",X"89",X"A2",X"80",X"A1",X"02",X"81",X"91",X"83",X"88",X"02",X"E1",
		X"09",X"09",X"08",X"08",X"18",X"91",X"90",X"8B",X"10",X"93",X"A9",X"01",X"A0",X"80",X"3F",X"77",
		X"F5",X"1F",X"11",X"B2",X"A9",X"95",X"92",X"0A",X"49",X"B3",X"9A",X"78",X"90",X"0A",X"2D",X"48",
		X"A8",X"12",X"C3",X"98",X"2A",X"97",X"A9",X"18",X"2C",X"07",X"A8",X"82",X"B1",X"00",X"A3",X"A1",
		X"98",X"2A",X"20",X"00",X"99",X"4D",X"10",X"02",X"BC",X"30",X"3A",X"F7",X"A8",X"29",X"08",X"08",
		X"98",X"23",X"F3",X"B3",X"A0",X"88",X"08",X"91",X"81",X"7F",X"49",X"B4",X"89",X"19",X"08",X"81",
		X"A4",X"98",X"0A",X"38",X"87",X"AA",X"4B",X"3D",X"3C",X"38",X"0A",X"2A",X"2B",X"7D",X"29",X"2A",
		X"19",X"18",X"08",X"00",X"88",X"08",X"08",X"00",X"09",X"08",X"1B",X"09",X"6D",X"3C",X"29",X"19",
		X"00",X"01",X"8C",X"5B",X"3A",X"00",X"80",X"29",X"80",X"89",X"0B",X"38",X"38",X"23",X"18",X"0B",
		X"19",X"3B",X"01",X"0A",X"F7",X"C1",X"09",X"2A",X"18",X"90",X"81",X"B4",X"0A",X"82",X"D0",X"79",
		X"A8",X"4C",X"39",X"08",X"09",X"01",X"90",X"1A",X"2A",X"38",X"2A",X"91",X"01",X"98",X"15",X"F7",
		X"C1",X"1D",X"6D",X"39",X"08",X"80",X"08",X"88",X"18",X"1D",X"38",X"09",X"08",X"92",X"0A",X"29",
		X"2A",X"08",X"2B",X"94",X"09",X"2B",X"1D",X"48",X"80",X"2A",X"2D",X"82",X"84",X"F2",X"89",X"4A",
		X"08",X"04",X"F4",X"B2",X"98",X"82",X"88",X"A8",X"38",X"88",X"8B",X"7A",X"0B",X"4A",X"28",X"89",
		X"4B",X"29",X"28",X"08",X"80",X"08",X"8A",X"99",X"7C",X"39",X"88",X"02",X"80",X"A2",X"8B",X"41",
		X"C5",X"B2",X"89",X"7D",X"91",X"3A",X"3D",X"11",X"98",X"81",X"0A",X"21",X"C0",X"3B",X"1B",X"21",
		X"91",X"01",X"F3",X"D4",X"A1",X"91",X"94",X"D2",X"90",X"82",X"A8",X"01",X"A0",X"4A",X"11",X"98",
		X"91",X"0A",X"28",X"03",X"1F",X"C5",X"3C",X"09",X"19",X"19",X"80",X"83",X"F1",X"11",X"B0",X"08",
		X"01",X"98",X"2B",X"1A",X"29",X"3C",X"21",X"2A",X"19",X"0A",X"4B",X"81",X"18",X"88",X"19",X"08",
		X"08",X"2A",X"08",X"A2",X"00",X"88",X"A6",X"B1",X"08",X"03",X"D1",X"A3",X"A1",X"B1",X"2B",X"00",
		X"2A",X"01",X"A3",X"80",X"8B",X"13",X"89",X"08",X"08",X"08",X"91",X"A2",X"08",X"A0",X"82",X"91",
		X"08",X"91",X"98",X"28",X"08",X"01",X"B1",X"08",X"0A",X"28",X"0A",X"28",X"91",X"0A",X"28",X"08",
		X"08",X"08",X"0A",X"28",X"0A",X"01",X"08",X"2A",X"0A",X"2A",X"01",X"08",X"08",X"0A",X"2B",X"38",
		X"99",X"4B",X"2A",X"08",X"28",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"0A",X"2A",X"2A",X"2A",X"08",X"2A",X"0A",X"23",X"89",X"B8",X"10",X"3C",
		X"13",X"B1",X"08",X"08",X"08",X"08",X"99",X"18",X"01",X"08",X"00",X"00",X"90",X"80",X"88",X"08",
		X"08",X"0A",X"09",X"00",X"80",X"08",X"28",X"08",X"08",X"08",X"08",X"19",X"08",X"08",X"0A",X"01",
		X"91",X"0A",X"08",X"01",X"08",X"08",X"08",X"08",X"08",X"91",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"98",X"08",X"01",X"98",X"08",X"01",X"08",X"08",X"08",X"08",X"00",X"88",X"08",X"08",
		X"0A",X"2A",X"2A",X"01",X"08",X"91",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"91",
		X"0A",X"08",X"28",X"A2",X"A2",X"08",X"0A",X"2A",X"28",X"08",X"08",X"08",X"08",X"08",X"98",X"08",
		X"28",X"08",X"08",X"91",X"08",X"08",X"08",X"08",X"08",X"0A",X"01",X"98",X"08",X"01",X"08",X"08",
		X"19",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"08",X"01",X"80",X"08",X"08",X"08",X"0A",X"09",
		X"3A",X"08",X"08",X"01",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"98",X"09",X"18",X"08",X"08",X"01",X"98",X"2A",X"28",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"98",X"28",X"91",
		X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"28",X"98",X"08",X"80",X"01",X"08",X"08",X"91",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"28",X"08",X"08",X"0A",X"08",X"28",
		X"08",X"08",X"08",X"08",X"08",X"08",X"91",X"08",X"08",X"0A",X"08",X"08",X"28",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"91",X"98",X"28",X"08",X"08",X"08",X"08",X"0A",X"2A",X"08",X"09",X"09",X"18",X"11",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"98",X"01",X"91",X"08",X"08",X"18",X"88",X"0A",X"2A",X"80",X"08",X"28",X"08",X"98",X"09",
		X"18",X"28",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"08",X"08",X"2A",
		X"28",X"08",X"08",X"00",X"88",X"08",X"08",X"08",X"08",X"08",X"98",X"08",X"28",X"08",X"0A",X"01",
		X"88",X"80",X"AF",X"FF",X"F1",X"23",X"50",X"18",X"D8",X"80",X"14",X"61",X"08",X"A9",X"AA",X"9A",
		X"9A",X"9B",X"FF",X"98",X"80",X"13",X"36",X"20",X"81",X"18",X"9B",X"FB",X"98",X"01",X"21",X"22",
		X"22",X"33",X"39",X"DA",X"88",X"00",X"11",X"12",X"53",X"35",X"20",X"DE",X"BA",X"A9",X"08",X"00",
		X"23",X"44",X"20",X"8C",X"BC",X"DA",X"90",X"00",X"21",X"23",X"53",X"19",X"DF",X"B0",X"01",X"13",
		X"24",X"42",X"89",X"AC",X"B8",X"99",X"8A",X"9B",X"B9",X"46",X"54",X"10",X"99",X"9A",X"BF",X"A9",
		X"80",X"00",X"12",X"11",X"12",X"43",X"43",X"42",X"23",X"60",X"09",X"CA",X"DA",X"BA",X"A9",X"80",
		X"02",X"12",X"22",X"22",X"42",X"12",X"26",X"10",X"00",X"B9",X"90",X"8D",X"CA",X"BB",X"A9",X"9B",
		X"23",X"8A",X"DC",X"AA",X"84",X"30",X"84",X"45",X"20",X"A9",X"AA",X"DB",X"9A",X"80",X"14",X"41",
		X"34",X"21",X"0B",X"DB",X"D8",X"88",X"01",X"14",X"53",X"42",X"89",X"BE",X"AC",X"9A",X"81",X"23",
		X"42",X"33",X"20",X"1C",X"DB",X"98",X"91",X"18",X"25",X"42",X"20",X"8C",X"BB",X"BE",X"9A",X"82",
		X"35",X"23",X"42",X"09",X"AC",X"DA",X"98",X"81",X"10",X"23",X"42",X"1A",X"CB",X"AB",X"9A",X"80",
		X"07",X"13",X"23",X"29",X"89",X"EB",X"AB",X"A0",X"83",X"43",X"62",X"19",X"AC",X"BE",X"00",X"09",
		X"10",X"33",X"31",X"18",X"99",X"00",X"89",X"83",X"FA",X"21",X"AD",X"D9",X"8D",X"01",X"32",X"46",
		X"11",X"12",X"28",X"82",X"E9",X"BB",X"BC",X"A9",X"81",X"24",X"20",X"B9",X"B9",X"FA",X"12",X"15",
		X"24",X"31",X"08",X"CB",X"AC",X"A8",X"90",X"51",X"22",X"32",X"32",X"90",X"AD",X"A1",X"BA",X"09",
		X"15",X"21",X"9D",X"D9",X"BA",X"CA",X"21",X"15",X"53",X"38",X"89",X"8D",X"BA",X"AA",X"93",X"31",
		X"12",X"63",X"20",X"AA",X"8D",X"0D",X"A4",X"23",X"EA",X"94",X"BB",X"08",X"28",X"97",X"31",X"23",
		X"11",X"11",X"F0",X"A8",X"CA",X"88",X"A9",X"72",X"1C",X"2A",X"08",X"1C",X"8D",X"02",X"39",X"11",
		X"25",X"B0",X"08",X"3B",X"F8",X"A0",X"8B",X"35",X"20",X"98",X"08",X"48",X"2B",X"B1",X"33",X"3F",
		X"A9",X"90",X"83",X"BC",X"0B",X"88",X"08",X"00",X"74",X"20",X"A9",X"1C",X"C8",X"88",X"12",X"13",
		X"0A",X"01",X"39",X"0A",X"0C",X"98",X"28",X"20",X"26",X"40",X"CB",X"D8",X"11",X"80",X"E8",X"01",
		X"11",X"02",X"10",X"B0",X"80",X"80",X"84",X"28",X"8A",X"08",X"AD",X"9B",X"82",X"61",X"AA",X"84",
		X"80",X"82",X"C1",X"02",X"A1",X"01",X"B9",X"14",X"88",X"D1",X"18",X"8A",X"08",X"42",X"12",X"F8",
		X"81",X"30",X"BB",X"91",X"28",X"80",X"CA",X"02",X"4A",X"89",X"21",X"39",X"0A",X"A1",X"22",X"A9",
		X"0A",X"82",X"99",X"09",X"08",X"01",X"0A",X"01",X"10",X"2C",X"98",X"18",X"88",X"10",X"01",X"10",
		X"8A",X"19",X"81",X"9A",X"08",X"08",X"21",X"08",X"28",X"09",X"10",X"8A",X"19",X"0A",X"08",X"08",
		X"08",X"08",X"28",X"98",X"08",X"08",X"01",X"08",X"18",X"88",X"0A",X"98",X"08",X"08",X"08",X"00",
		X"18",X"01",X"19",X"00",X"09",X"09",X"18",X"99",X"10",X"18",X"89",X"2A",X"28",X"80",X"08",X"08",
		X"18",X"18",X"89",X"08",X"89",X"0A",X"08",X"10",X"90",X"81",X"81",X"10",X"80",X"80",X"80",X"80",
		X"A0",X"10",X"80",X"8A",X"88",X"80",X"81",X"02",X"00",X"80",X"90",X"80",X"80",X"80",X"80",X"80",
		X"89",X"19",X"90",X"00",X"88",X"88",X"80",X"80",X"8A",X"88",X"80",X"B0",X"81",X"10",X"80",X"03",
		X"81",X"20",X"80",X"33",X"32",X"12",X"02",X"00",X"01",X"80",X"80",X"89",X"88",X"98",X"99",X"A9",
		X"88",X"A8",X"52",X"FB",X"00",X"76",X"32",X"73",X"61",X"AE",X"98",X"9A",X"A9",X"A8",X"F0",X"2C",
		X"20",X"F8",X"5B",X"82",X"90",X"11",X"50",X"98",X"03",X"90",X"17",X"0B",X"01",X"80",X"00",X"21",
		X"91",X"BD",X"03",X"0B",X"C0",X"90",X"61",X"E9",X"00",X"2A",X"95",X"C8",X"3D",X"82",X"A0",X"2B",
		X"80",X"04",X"0C",X"0B",X"91",X"93",X"38",X"F2",X"80",X"88",X"31",X"F9",X"21",X"02",X"D8",X"37",
		X"C8",X"80",X"08",X"23",X"9B",X"B0",X"92",X"27",X"0C",X"81",X"3D",X"39",X"99",X"83",X"00",X"B2",
		X"25",X"84",X"DA",X"98",X"13",X"3B",X"A0",X"73",X"F0",X"89",X"13",X"B9",X"6A",X"A2",X"91",X"2B",
		X"13",X"A0",X"B1",X"7A",X"C8",X"06",X"3D",X"98",X"18",X"92",X"02",X"8B",X"90",X"47",X"C9",X"11",
		X"09",X"B6",X"3F",X"80",X"10",X"A0",X"81",X"09",X"59",X"08",X"B2",X"06",X"8A",X"B1",X"2A",X"0B",
		X"68",X"95",X"1F",X"81",X"29",X"98",X"91",X"42",X"F9",X"02",X"80",X"28",X"C8",X"12",X"94",X"B8",
		X"B8",X"60",X"A1",X"9A",X"25",X"81",X"A2",X"8D",X"A0",X"04",X"2B",X"01",X"CB",X"06",X"99",X"13",
		X"B3",X"86",X"BB",X"93",X"00",X"E2",X"80",X"28",X"B8",X"27",X"28",X"8C",X"A0",X"A9",X"6A",X"A1",
		X"43",X"8C",X"B0",X"12",X"12",X"8C",X"94",X"11",X"AF",X"19",X"82",X"3B",X"92",X"11",X"9B",X"D4",
		X"99",X"10",X"27",X"2D",X"98",X"92",X"4B",X"9C",X"06",X"89",X"13",X"AB",X"12",X"A9",X"21",X"C2",
		X"89",X"4B",X"B3",X"B8",X"67",X"99",X"B1",X"22",X"6B",X"A9",X"93",X"30",X"F9",X"00",X"30",X"B0",
		X"89",X"23",X"1E",X"08",X"A2",X"50",X"98",X"85",X"90",X"D8",X"81",X"30",X"C9",X"98",X"10",X"54",
		X"9E",X"80",X"20",X"28",X"C0",X"82",X"09",X"D0",X"40",X"9B",X"10",X"93",X"08",X"2A",X"B4",X"B0",
		X"79",X"94",X"B0",X"2C",X"92",X"41",X"BF",X"13",X"A8",X"A1",X"82",X"36",X"9A",X"D9",X"00",X"10",
		X"B2",X"47",X"99",X"98",X"39",X"C9",X"03",X"20",X"22",X"BE",X"92",X"BA",X"54",X"0C",X"90",X"00",
		X"A1",X"12",X"48",X"6D",X"B0",X"21",X"81",X"98",X"98",X"20",X"8A",X"20",X"7A",X"2D",X"89",X"81",
		X"39",X"18",X"36",X"C8",X"9B",X"15",X"28",X"D0",X"1A",X"82",X"5A",X"0B",X"8D",X"85",X"20",X"CA",
		X"10",X"28",X"93",X"99",X"D0",X"78",X"88",X"01",X"10",X"C9",X"02",X"48",X"CB",X"90",X"14",X"88",
		X"28",X"09",X"9A",X"7B",X"B4",X"38",X"C9",X"23",X"99",X"91",X"32",X"29",X"D0",X"9F",X"11",X"91",
		X"90",X"3F",X"B3",X"10",X"06",X"81",X"0E",X"80",X"00",X"1C",X"82",X"1A",X"B3",X"7A",X"89",X"A1",
		X"39",X"38",X"A8",X"10",X"86",X"0B",X"D1",X"53",X"BF",X"81",X"08",X"10",X"89",X"19",X"20",X"11",
		X"1C",X"F8",X"20",X"A0",X"23",X"B9",X"70",X"88",X"A8",X"1A",X"A2",X"A1",X"3E",X"93",X"68",X"C2",
		X"11",X"A1",X"BC",X"8A",X"60",X"BB",X"36",X"88",X"18",X"8A",X"29",X"24",X"AC",X"69",X"A1",X"80",
		X"10",X"CA",X"19",X"13",X"B1",X"69",X"96",X"19",X"AA",X"A0",X"06",X"8B",X"02",X"19",X"38",X"1E",
		X"CB",X"14",X"24",X"19",X"F8",X"03",X"8B",X"93",X"11",X"CC",X"16",X"89",X"20",X"AB",X"40",X"99",
		X"19",X"A8",X"A0",X"40",X"B2",X"73",X"B0",X"C9",X"3B",X"11",X"28",X"08",X"1B",X"89",X"61",X"8F",
		X"12",X"C0",X"92",X"08",X"43",X"EB",X"82",X"A0",X"21",X"C5",X"4A",X"D0",X"28",X"00",X"28",X"A8",
		X"8C",X"30",X"E2",X"19",X"A0",X"00",X"89",X"51",X"20",X"E0",X"02",X"99",X"AB",X"85",X"22",X"F9",
		X"02",X"29",X"1B",X"A5",X"03",X"90",X"8A",X"2B",X"FB",X"48",X"22",X"98",X"8C",X"12",X"01",X"AD",
		X"C1",X"31",X"29",X"A1",X"00",X"F3",X"78",X"09",X"D8",X"19",X"13",X"9B",X"91",X"49",X"A0",X"80",
		X"60",X"AB",X"01",X"3A",X"87",X"AA",X"33",X"AE",X"91",X"21",X"68",X"09",X"C0",X"08",X"B4",X"AC",
		X"02",X"59",X"2A",X"80",X"12",X"8E",X"98",X"85",X"0B",X"19",X"42",X"98",X"AD",X"23",X"A1",X"0B",
		X"B3",X"02",X"63",X"AE",X"90",X"A0",X"29",X"92",X"39",X"E9",X"37",X"89",X"88",X"98",X"19",X"19",
		X"2A",X"70",X"90",X"22",X"3D",X"00",X"DB",X"A3",X"3F",X"91",X"10",X"53",X"AA",X"A2",X"19",X"DA",
		X"13",X"23",X"8E",X"BA",X"25",X"11",X"00",X"0C",X"C0",X"02",X"1D",X"00",X"A3",X"11",X"84",X"81",
		X"AD",X"89",X"3A",X"AE",X"91",X"21",X"32",X"F8",X"62",X"9A",X"18",X"A8",X"AB",X"24",X"BA",X"52",
		X"02",X"18",X"A8",X"72",X"F9",X"80",X"89",X"82",X"09",X"09",X"50",X"89",X"A3",X"48",X"92",X"B9",
		X"2C",X"95",X"12",X"7A",X"C0",X"00",X"10",X"8C",X"C8",X"90",X"33",X"90",X"12",X"82",X"08",X"F3",
		X"01",X"1C",X"F8",X"30",X"32",X"BA",X"09",X"D8",X"84",X"3B",X"D9",X"81",X"51",X"E8",X"20",X"08",
		X"40",X"C9",X"12",X"89",X"05",X"1B",X"A0",X"A8",X"01",X"8E",X"93",X"A9",X"26",X"10",X"89",X"9E",
		X"01",X"40",X"00",X"B1",X"29",X"90",X"08",X"4C",X"EB",X"31",X"9B",X"A2",X"73",X"98",X"32",X"BB",
		X"B8",X"24",X"6A",X"9C",X"81",X"01",X"B3",X"C8",X"2B",X"42",X"EA",X"51",X"90",X"00",X"22",X"BF",
		X"81",X"18",X"88",X"16",X"1A",X"DB",X"88",X"44",X"08",X"99",X"89",X"B0",X"25",X"2A",X"88",X"01",
		X"29",X"D2",X"3B",X"A9",X"A1",X"71",X"D9",X"02",X"20",X"01",X"F9",X"80",X"31",X"8A",X"17",X"2C",
		X"A8",X"90",X"01",X"9D",X"93",X"20",X"21",X"90",X"2A",X"40",X"BE",X"A0",X"43",X"51",X"B8",X"28",
		X"DA",X"9A",X"B9",X"33",X"70",X"B9",X"31",X"1B",X"F0",X"11",X"28",X"29",X"B0",X"A3",X"05",X"68",
		X"A8",X"A0",X"0D",X"8A",X"F0",X"41",X"02",X"09",X"9A",X"A9",X"22",X"58",X"9E",X"02",X"31",X"9A",
		X"C2",X"59",X"C9",X"3B",X"84",X"A8",X"81",X"18",X"21",X"97",X"98",X"10",X"9F",X"90",X"90",X"23",
		X"0A",X"9F",X"16",X"1A",X"10",X"8C",X"08",X"23",X"AE",X"89",X"40",X"80",X"91",X"0B",X"98",X"37",
		X"0C",X"91",X"81",X"10",X"09",X"30",X"01",X"8B",X"B0",X"8B",X"3D",X"F9",X"29",X"1D",X"24",X"23",
		X"C0",X"8D",X"94",X"4A",X"D1",X"00",X"91",X"18",X"8B",X"91",X"24",X"39",X"CA",X"01",X"97",X"90",
		X"1B",X"8B",X"D3",X"49",X"92",X"82",X"1E",X"00",X"86",X"0B",X"22",X"0B",X"9D",X"A8",X"C0",X"24",
		X"82",X"58",X"89",X"90",X"2B",X"18",X"B2",X"A2",X"3B",X"BB",X"F0",X"60",X"11",X"AA",X"EA",X"93",
		X"70",X"80",X"A0",X"20",X"1B",X"92",X"2A",X"0E",X"21",X"32",X"CC",X"14",X"88",X"A4",X"BC",X"BD",
		X"11",X"01",X"28",X"27",X"0B",X"81",X"68",X"B8",X"98",X"8A",X"85",X"9E",X"01",X"88",X"53",X"1A",
		X"A3",X"AD",X"00",X"00",X"59",X"A8",X"38",X"DB",X"83",X"21",X"28",X"07",X"09",X"8A",X"9B",X"D3",
		X"2B",X"2A",X"C3",X"41",X"39",X"F9",X"18",X"13",X"99",X"A1",X"3C",X"51",X"CB",X"0A",X"82",X"09",
		X"83",X"50",X"07",X"A8",X"08",X"29",X"AC",X"05",X"22",X"91",X"1D",X"A9",X"B8",X"03",X"BA",X"87",
		X"1A",X"11",X"B0",X"99",X"09",X"BF",X"07",X"02",X"11",X"AA",X"88",X"8D",X"24",X"30",X"FB",X"92",
		X"31",X"21",X"CF",X"91",X"12",X"28",X"AA",X"43",X"83",X"9C",X"AC",X"81",X"10",X"B2",X"91",X"EA",
		X"02",X"BB",X"53",X"43",X"2B",X"9B",X"B1",X"AD",X"14",X"CA",X"15",X"13",X"49",X"A8",X"E9",X"81",
		X"04",X"08",X"19",X"A2",X"14",X"02",X"FB",X"08",X"89",X"91",X"8D",X"08",X"41",X"D1",X"32",X"02",
		X"40",X"9C",X"A9",X"21",X"BD",X"B8",X"96",X"39",X"13",X"81",X"9F",X"C8",X"32",X"01",X"A9",X"9A",
		X"23",X"98",X"D2",X"70",X"A9",X"22",X"AA",X"25",X"AB",X"8A",X"22",X"F3",X"0A",X"81",X"1A",X"BF",
		X"17",X"08",X"09",X"01",X"10",X"89",X"A9",X"8F",X"A0",X"43",X"88",X"04",X"BB",X"CA",X"24",X"82",
		X"8B",X"98",X"08",X"D0",X"51",X"38",X"B1",X"C1",X"39",X"A1",X"13",X"73",X"0C",X"FB",X"82",X"01",
		X"08",X"35",X"A1",X"0A",X"06",X"0A",X"09",X"F0",X"00",X"10",X"8A",X"90",X"0B",X"92",X"0B",X"12",
		X"34",X"73",X"9A",X"B9",X"83",X"3F",X"F9",X"14",X"13",X"9A",X"A8",X"83",X"10",X"9F",X"02",X"10",
		X"09",X"B0",X"32",X"2F",X"CA",X"02",X"99",X"13",X"38",X"18",X"19",X"E9",X"44",X"8D",X"98",X"22",
		X"58",X"19",X"90",X"A0",X"88",X"CA",X"2B",X"9B",X"87",X"42",X"AA",X"81",X"6A",X"B8",X"2A",X"17",
		X"2B",X"B9",X"81",X"09",X"20",X"3B",X"B3",X"08",X"B4",X"81",X"AB",X"35",X"9A",X"FC",X"25",X"10",
		X"05",X"88",X"AA",X"9A",X"98",X"11",X"B5",X"4A",X"9B",X"83",X"12",X"D9",X"33",X"10",X"59",X"11",
		X"88",X"FB",X"02",X"83",X"2C",X"C9",X"89",X"90",X"21",X"09",X"43",X"87",X"AB",X"0C",X"C9",X"07",
		X"28",X"12",X"8C",X"99",X"14",X"10",X"0A",X"D8",X"08",X"21",X"08",X"5D",X"B8",X"38",X"0B",X"90",
		X"58",X"04",X"0C",X"A0",X"48",X"29",X"A9",X"99",X"44",X"00",X"C9",X"80",X"31",X"40",X"0F",X"90",
		X"A8",X"27",X"3C",X"80",X"09",X"88",X"9D",X"9A",X"37",X"49",X"9B",X"89",X"30",X"01",X"0A",X"49",
		X"82",X"BF",X"02",X"18",X"93",X"30",X"A1",X"BA",X"9C",X"84",X"18",X"39",X"FF",X"00",X"04",X"09",
		X"80",X"01",X"0A",X"A9",X"08",X"80",X"80",X"34",X"35",X"AC",X"2D",X"A8",X"80",X"86",X"42",X"90",
		X"29",X"BA",X"A9",X"BA",X"CB",X"B7",X"39",X"10",X"A2",X"3A",X"2A",X"D4",X"35",X"0C",X"92",X"09",
		X"99",X"AE",X"84",X"1B",X"08",X"13",X"8B",X"E0",X"34",X"8C",X"81",X"24",X"98",X"29",X"9D",X"8A",
		X"40",X"2B",X"12",X"32",X"FB",X"B1",X"02",X"33",X"4A",X"FA",X"08",X"00",X"41",X"AB",X"83",X"37",
		X"3B",X"98",X"D9",X"B8",X"30",X"A8",X"07",X"39",X"80",X"8D",X"A2",X"52",X"8B",X"03",X"1B",X"93",
		X"AA",X"9E",X"16",X"B9",X"39",X"22",X"9B",X"0B",X"34",X"EA",X"80",X"03",X"A9",X"B3",X"4B",X"72",
		X"29",X"98",X"DA",X"11",X"8C",X"93",X"22",X"03",X"20",X"28",X"99",X"BA",X"10",X"2C",X"9A",X"01",
		X"2C",X"A8",X"08",X"C4",X"28",X"03",X"1B",X"C9",X"A9",X"46",X"0A",X"04",X"88",X"B8",X"71",X"08",
		X"31",X"CB",X"9E",X"88",X"90",X"29",X"01",X"92",X"25",X"09",X"83",X"1B",X"C2",X"BC",X"89",X"23",
		X"41",X"93",X"20",X"8A",X"FB",X"13",X"23",X"BB",X"25",X"B4",X"1B",X"F0",X"80",X"80",X"99",X"D9",
		X"53",X"89",X"91",X"31",X"12",X"91",X"AA",X"FB",X"88",X"11",X"44",X"02",X"8B",X"BB",X"B5",X"CA",
		X"02",X"17",X"20",X"9C",X"88",X"8A",X"10",X"35",X"01",X"44",X"9E",X"A8",X"08",X"00",X"90",X"A1",
		X"10",X"80",X"30",X"C0",X"10",X"23",X"A2",X"C0",X"3B",X"CB",X"BC",X"96",X"30",X"30",X"90",X"14",
		X"0D",X"01",X"BD",X"84",X"22",X"99",X"BD",X"1A",X"AA",X"14",X"80",X"04",X"33",X"51",X"BB",X"CA",
		X"84",X"20",X"A2",X"8D",X"1B",X"A2",X"52",X"2C",X"F8",X"28",X"00",X"90",X"89",X"C0",X"02",X"3A",
		X"24",X"40",X"89",X"A1",X"A8",X"B8",X"30",X"C0",X"42",X"1D",X"AA",X"51",X"1B",X"0E",X"01",X"92",
		X"8A",X"50",X"19",X"91",X"31",X"99",X"1B",X"03",X"8D",X"AB",X"84",X"11",X"03",X"0C",X"10",X"DA",
		X"59",X"B1",X"40",X"83",X"8B",X"BB",X"D0",X"83",X"01",X"60",X"B0",X"A8",X"81",X"62",X"8A",X"91",
		X"3B",X"12",X"01",X"2A",X"9B",X"BC",X"02",X"08",X"19",X"A6",X"00",X"93",X"2A",X"A2",X"CB",X"0C",
		X"12",X"05",X"10",X"8B",X"FA",X"22",X"20",X"80",X"33",X"9D",X"B0",X"06",X"28",X"C9",X"88",X"23",
		X"BB",X"88",X"F0",X"10",X"33",X"89",X"80",X"B8",X"32",X"21",X"AF",X"B8",X"23",X"10",X"9A",X"00",
		X"88",X"50",X"8B",X"98",X"10",X"28",X"B8",X"21",X"A2",X"18",X"8C",X"19",X"A3",X"00",X"30",X"48",
		X"89",X"BC",X"A3",X"80",X"30",X"82",X"12",X"AB",X"A3",X"38",X"8B",X"B8",X"80",X"84",X"19",X"80",
		X"A9",X"81",X"2A",X"29",X"89",X"C0",X"C1",X"23",X"2A",X"04",X"88",X"22",X"2B",X"BB",X"B9",X"43",
		X"30",X"A2",X"0A",X"9C",X"08",X"12",X"AD",X"03",X"1A",X"52",X"AB",X"28",X"28",X"08",X"2A",X"28",
		X"9A",X"A9",X"08",X"08",X"4B",X"B8",X"03",X"B3",X"30",X"C0",X"82",X"82",X"80",X"81",X"2B",X"C0",
		X"B3",X"32",X"89",X"30",X"83",X"A8",X"C9",X"98",X"CA",X"24",X"33",X"0B",X"B8",X"C0",X"30",X"32",
		X"A0",X"80",X"18",X"20",X"80",X"AC",X"38",X"CB",X"A2",X"34",X"12",X"A9",X"00",X"C2",X"48",X"0C",
		X"AB",X"08",X"09",X"19",X"12",X"25",X"18",X"92",X"A9",X"AA",X"9A",X"2A",X"20",X"84",X"81",X"80",
		X"2A",X"81",X"AA",X"88",X"16",X"8A",X"0A",X"90",X"19",X"80",X"34",X"AB",X"28",X"9A",X"08",X"41",
		X"2E",X"90",X"81",X"50",X"8A",X"80",X"89",X"A0",X"8A",X"9A",X"95",X"40",X"81",X"01",X"18",X"83",
		X"8A",X"E8",X"88",X"A2",X"18",X"18",X"88",X"1A",X"28",X"05",X"19",X"9A",X"08",X"08",X"E8",X"28",
		X"A8",X"30",X"30",X"80",X"81",X"92",X"1B",X"B8",X"80",X"82",X"10",X"89",X"14",X"0A",X"C2",X"82",
		X"89",X"8B",X"C1",X"38",X"32",X"10",X"19",X"B8",X"CB",X"84",X"03",X"19",X"B1",X"19",X"A0",X"80",
		X"80",X"80",X"80",X"80",X"12",X"81",X"29",X"98",X"80",X"B1",X"A1",X"21",X"11",X"B8",X"80",X"80",
		X"01",X"11",X"09",X"C0",X"B8",X"08",X"82",X"1A",X"90",X"82",X"19",X"A2",X"10",X"C2",X"19",X"A0",
		X"01",X"A1",X"00",X"80",X"93",X"8B",X"80",X"B3",X"80",X"03",X"81",X"80",X"91",X"88",X"80",X"A2",
		X"03",X"89",X"AB",X"81",X"21",X"88",X"80",X"8A",X"94",X"8B",X"03",X"A2",X"B8",X"13",X"88",X"80",
		X"80",X"8A",X"9A",X"20",X"30",X"80",X"80",X"80",X"80",X"80",X"8B",X"80",X"80",X"81",X"81",X"19",
		X"10",X"80",X"82",X"82",X"89",X"AA",X"80",X"83",X"01",X"18",X"BB",X"82",X"10",X"A0",X"89",X"80",
		X"80",X"C1",X"33",X"89",X"82",X"A8",X"90",X"81",X"20",X"89",X"82",X"A2",X"80",X"80",X"00",X"00",
		X"82",X"B0",X"88",X"80",X"80",X"8A",X"90",X"84",X"08",X"81",X"0C",X"91",X"80",X"90",X"03",X"A8",
		X"80",X"20",X"B3",X"A2",X"00",X"88",X"80",X"81",X"8A",X"AA",X"2A",X"20",X"81",X"21",X"83",X"A8",
		X"80",X"90",X"80",X"80",X"80",X"A9",X"80",X"82",X"11",X"9A",X"90",X"30",X"80",X"00",X"88",X"80",
		X"80",X"80",X"8B",X"C0",X"30",X"C9",X"14",X"82",X"11",X"90",X"31",X"B9",X"CB",X"03",X"03",X"18",
		X"91",X"02",X"A9",X"80",X"00",X"9A",X"94",X"80",X"A9",X"80",X"81",X"20",X"A2",X"81",X"20",X"A0",
		X"1A",X"99",X"10",X"8A",X"88",X"80",X"19",X"80",X"81",X"02",X"8B",X"80",X"80",X"82",X"23",X"80",
		X"80",X"BA",X"91",X"89",X"81",X"33",X"A9",X"80",X"80",X"B3",X"88",X"92",X"A8",X"C8",X"03",X"A2",
		X"39",X"A4",X"31",X"09",X"CA",X"88",X"10",X"19",X"98",X"80",X"12",X"80",X"89",X"80",X"82",X"80",
		X"80",X"80",X"08",X"80",X"00",X"90",X"80",X"C0",X"03",X"89",X"11",X"09",X"B3",X"80",X"81",X"00",
		X"AA",X"9A",X"83",X"A8",X"20",X"B3",X"03",X"30",X"B8",X"80",X"80",X"A8",X"83",X"80",X"89",X"90",
		X"20",X"80",X"C1",X"31",X"98",X"80",X"80",X"8A",X"91",X"91",X"20",X"89",X"90",X"20",X"80",X"80",
		X"12",X"8B",X"B8",X"8A",X"80",X"83",X"12",X"A0",X"82",X"81",X"9B",X"28",X"A1",X"33",X"80",X"B0",
		X"80",X"90",X"80",X"80",X"A2",X"80",X"80",X"80",X"80",X"3A",X"9A",X"92",X"88",X"91",X"20",X"80",
		X"8B",X"80",X"82",X"10",X"8A",X"91",X"88",X"19",X"80",X"82",X"10",X"89",X"98",X"81",X"22",X"19",
		X"01",X"CA",X"88",X"08",X"00",X"38",X"28",X"80",X"0A",X"08",X"08",X"91",X"21",X"0A",X"98",X"A8",
		X"80",X"18",X"89",X"08",X"08",X"03",X"08",X"0B",X"38",X"21",X"9A",X"A9",X"12",X"08",X"08",X"9A",
		X"A2",X"48",X"10",X"9C",X"08",X"08",X"00",X"30",X"88",X"08",X"00",X"88",X"18",X"88",X"08",X"99",
		X"19",X"11",X"00",X"38",X"B8",X"A2",X"00",X"8B",X"09",X"19",X"48",X"08",X"A9",X"08",X"00",X"3A",
		X"09",X"38",X"0A",X"28",X"A8",X"18",X"21",X"2A",X"09",X"00",X"2B",X"09",X"08",X"B0",X"09",X"08",
		X"29",X"00",X"09",X"3A",X"09",X"80",X"11",X"08",X"98",X"88",X"38",X"19",X"10",X"9B",X"02",X"00",
		X"88",X"08",X"99",X"09",X"18",X"08",X"81",X"28",X"08",X"0A",X"88",X"19",X"31",X"89",X"A2",X"00",
		X"88",X"A0",X"28",X"A0",X"28",X"08",X"08",X"00",X"19",X"88",X"08",X"08",X"91",X"B8",X"08",X"08",
		X"19",X"08",X"19",X"0B",X"38",X"03",X"03",X"0A",X"90",X"09",X"A9",X"18",X"38",X"11",X"A8",X"08",
		X"00",X"00",X"98",X"08",X"0A",X"28",X"08",X"B8",X"03",X"18",X"88",X"00",X"88",X"9A",X"08",X"08",
		X"08",X"01",X"28",X"0C",X"08",X"28",X"28",X"08",X"0C",X"08",X"08",X"08",X"21",X"08",X"12",X"99",
		X"88",X"0A",X"01",X"08",X"08",X"08",X"0C",X"03",X"00",X"80",X"19",X"09",X"98",X"01",X"0A",X"89",
		X"28",X"88",X"11",X"08",X"08",X"98",X"01",X"A9",X"29",X"88",X"08",X"18",X"00",X"2A",X"28",X"18",
		X"10",X"8A",X"08",X"08",X"08",X"91",X"08",X"08",X"08",X"08",X"0A",X"2A",X"98",X"08",X"10",X"28",
		X"0C",X"30",X"80",X"80",X"A0",X"10",X"81",X"90",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",
		X"09",X"08",X"B1",X"69",X"93",X"E9",X"60",X"B2",X"8F",X"23",X"A9",X"29",X"F0",X"58",X"91",X"89",
		X"9B",X"71",X"A0",X"1B",X"B7",X"0A",X"19",X"A7",X"89",X"90",X"49",X"B2",X"3A",X"D2",X"3B",X"0A",
		X"B7",X"1B",X"1A",X"33",X"DA",X"41",X"C9",X"50",X"AA",X"41",X"BA",X"50",X"B9",X"41",X"B9",X"86",
		X"8A",X"95",X"0A",X"99",X"43",X"C8",X"90",X"5A",X"B3",X"4B",X"A1",X"5B",X"95",X"9B",X"48",X"A4",
		X"A9",X"48",X"C2",X"3C",X"89",X"32",X"B8",X"A8",X"70",X"A1",X"B9",X"78",X"98",X"94",X"0A",X"0A",
		X"07",X"99",X"08",X"A1",X"6A",X"81",X"8A",X"96",X"0B",X"18",X"A5",X"0B",X"09",X"16",X"A9",X"09",
		X"48",X"A9",X"25",X"A9",X"93",X"2C",X"89",X"42",X"D9",X"23",X"BB",X"17",X"99",X"89",X"69",X"90",
		X"93",X"2D",X"09",X"05",X"A9",X"84",X"8A",X"93",X"2C",X"89",X"50",X"B8",X"84",X"1C",X"09",X"15",
		X"A9",X"2B",X"95",X"2D",X"08",X"94",X"0B",X"81",X"4B",X"98",X"58",X"A8",X"85",X"8A",X"94",X"1C",
		X"81",X"4B",X"98",X"15",X"A9",X"1A",X"87",X"8A",X"18",X"A1",X"6B",X"81",X"A8",X"41",X"C0",X"19",
		X"A1",X"69",X"91",X"9A",X"26",X"B8",X"1A",X"24",X"C8",X"80",X"4A",X"A0",X"59",X"99",X"14",X"AA",
		X"05",X"99",X"89",X"58",X"A8",X"85",X"0B",X"00",X"B2",X"7B",X"00",X"A3",X"2D",X"09",X"05",X"A9",
		X"09",X"25",X"B8",X"89",X"50",X"B9",X"16",X"A8",X"19",X"A1",X"7A",X"91",X"98",X"32",X"D0",X"0A",
		X"05",X"9A",X"08",X"49",X"90",X"A3",X"6C",X"08",X"84",X"9A",X"1A",X"16",X"A8",X"0A",X"23",X"C8",
		X"91",X"6A",X"90",X"95",X"8B",X"04",X"9A",X"83",X"1D",X"85",X"9A",X"13",X"C8",X"3B",X"02",X"B2",
		X"1D",X"40",X"D1",X"3C",X"84",X"9A",X"22",X"D8",X"38",X"B0",X"59",X"A0",X"93",X"3C",X"82",X"B9",
		X"44",X"D0",X"1A",X"94",X"2C",X"82",X"9B",X"26",X"A9",X"19",X"95",X"0B",X"19",X"97",X"8A",X"09",
		X"23",X"C8",X"29",X"A9",X"17",X"8A",X"18",X"99",X"34",X"C8",X"90",X"69",X"91",X"8B",X"07",X"99",
		X"09",X"31",X"C0",X"98",X"58",X"A1",X"99",X"60",X"B1",X"8A",X"33",X"E8",X"81",X"4B",X"89",X"41",
		X"C8",X"30",X"BA",X"36",X"B9",X"85",X"8A",X"93",X"2D",X"83",X"0D",X"13",X"C9",X"48",X"B2",X"3D",
		X"82",X"1B",X"88",X"58",X"A8",X"84",X"1C",X"88",X"32",X"C9",X"84",X"1C",X"93",X"2C",X"A3",X"5C",
		X"88",X"30",X"B9",X"86",X"0A",X"0A",X"84",X"3E",X"01",X"A9",X"42",X"D0",X"0A",X"15",X"A9",X"18",
		X"99",X"50",X"A0",X"8A",X"42",X"C8",X"83",X"2D",X"09",X"15",X"B9",X"05",X"9A",X"82",X"2B",X"A0",
		X"79",X"99",X"15",X"A9",X"09",X"23",X"D9",X"14",X"A8",X"99",X"60",X"B1",X"8A",X"43",X"E0",X"0A",
		X"14",X"AA",X"03",X"0B",X"98",X"78",X"A8",X"22",X"D0",X"4A",X"A1",X"4B",X"94",X"8B",X"06",X"9A",
		X"2A",X"93",X"4C",X"81",X"89",X"91",X"7A",X"81",X"8A",X"86",X"8A",X"1A",X"14",X"A9",X"0A",X"35",
		X"C8",X"80",X"49",X"90",X"A0",X"79",X"90",X"A3",X"2C",X"09",X"96",X"0B",X"09",X"23",X"C9",X"05",
		X"9A",X"85",X"8A",X"88",X"59",X"A8",X"40",X"B9",X"33",X"D9",X"40",X"C1",X"2C",X"12",X"C0",X"3B",
		X"96",X"9A",X"04",X"9A",X"04",X"AA",X"32",X"C9",X"04",X"8A",X"0A",X"43",X"D8",X"81",X"4B",X"81",
		X"8B",X"87",X"0B",X"10",X"B2",X"6B",X"81",X"A9",X"43",X"E0",X"1A",X"85",X"99",X"88",X"48",X"A9",
		X"32",X"C0",X"98",X"68",X"A1",X"A8",X"68",X"B8",X"13",X"9B",X"86",X"8A",X"91",X"6A",X"92",X"A9",
		X"34",X"D0",X"89",X"40",X"B8",X"04",X"8A",X"98",X"68",X"A8",X"05",X"9A",X"81",X"4A",X"A8",X"41",
		X"B8",X"A2",X"7A",X"90",X"A5",X"0B",X"09",X"32",X"C8",X"93",X"4C",X"00",X"B0",X"79",X"91",X"9A",
		X"51",X"C0",X"0A",X"41",X"B8",X"0A",X"50",X"A9",X"05",X"99",X"90",X"6A",X"90",X"4B",X"94",X"8B",
		X"32",X"D9",X"58",X"A8",X"21",X"B9",X"14",X"A9",X"92",X"5A",X"99",X"16",X"AA",X"14",X"AB",X"34",
		X"C9",X"04",X"8A",X"91",X"5A",X"99",X"32",X"C9",X"24",X"C9",X"14",X"B9",X"84",X"1B",X"0A",X"07",
		X"9A",X"29",X"A5",X"1C",X"09",X"13",X"A9",X"91",X"7A",X"98",X"48",X"A9",X"15",X"A9",X"88",X"50",
		X"B1",X"A8",X"79",X"91",X"8A",X"07",X"9A",X"28",X"A8",X"41",X"C0",X"0A",X"15",X"A9",X"1A",X"24",
		X"B8",X"98",X"79",X"90",X"93",X"1C",X"80",X"4A",X"A2",X"4B",X"A0",X"69",X"A8",X"40",X"B9",X"24",
		X"C9",X"40",X"B0",X"4A",X"B3",X"3D",X"93",X"2C",X"89",X"15",X"A8",X"89",X"50",X"B1",X"A8",X"78",
		X"A1",X"99",X"40",X"B9",X"15",X"99",X"89",X"41",X"B9",X"96",X"0A",X"98",X"50",X"B9",X"23",X"BB",
		X"43",X"D9",X"40",X"B9",X"16",X"A9",X"81",X"3B",X"80",X"B4",X"5C",X"89",X"24",X"B8",X"1C",X"16",
		X"A9",X"10",X"B0",X"40",X"B1",X"0A",X"A5",X"3D",X"01",X"A9",X"51",X"C0",X"1B",X"07",X"A8",X"09",
		X"13",X"B9",X"84",X"0A",X"A3",X"4C",X"A3",X"4C",X"92",X"2D",X"04",X"AA",X"31",X"C9",X"40",X"B8",
		X"22",X"C8",X"59",X"B4",X"0C",X"21",X"C2",X"1C",X"03",X"9A",X"80",X"59",X"99",X"24",X"C8",X"83",
		X"0B",X"A3",X"6A",X"91",X"B0",X"79",X"98",X"93",X"3D",X"82",X"8B",X"85",X"1C",X"01",X"B2",X"4B",
		X"98",X"06",X"9A",X"85",X"99",X"88",X"58",X"A0",X"8A",X"51",X"B8",X"90",X"69",X"91",X"9A",X"51",
		X"C8",X"03",X"9B",X"06",X"9A",X"82",X"3B",X"88",X"B6",X"2C",X"88",X"48",X"A0",X"A1",X"7A",X"98",
		X"04",X"99",X"0A",X"34",X"C0",X"0B",X"26",X"B8",X"1B",X"07",X"99",X"88",X"30",X"A8",X"A4",X"2C",
		X"92",X"4B",X"A1",X"5B",X"A2",X"5A",X"99",X"05",X"99",X"94",X"0B",X"96",X"9A",X"04",X"9A",X"84",
		X"0A",X"A2",X"4B",X"98",X"69",X"A0",X"59",X"A1",X"A1",X"5A",X"92",X"8A",X"A1",X"51",X"B1",X"0A",
		X"10",X"98",X"BC",X"57",X"B8",X"18",X"89",X"85",X"1C",X"08",X"95",X"0B",X"18",X"A2",X"5B",X"98",
		X"24",X"C8",X"83",X"1C",X"90",X"69",X"98",X"94",X"0B",X"94",X"1B",X"A6",X"0B",X"91",X"49",X"98",
		X"A4",X"3D",X"08",X"85",X"9A",X"82",X"2C",X"88",X"58",X"A9",X"15",X"A8",X"8A",X"50",X"A9",X"85",
		X"8A",X"80",X"5A",X"99",X"50",X"A9",X"05",X"A9",X"84",X"8B",X"84",X"0B",X"91",X"5A",X"80",X"B4",
		X"3D",X"08",X"94",X"0C",X"84",X"8A",X"93",X"2B",X"8A",X"51",X"BA",X"51",X"C0",X"93",X"2C",X"89",
		X"25",X"B8",X"89",X"68",X"A9",X"24",X"B8",X"98",X"78",X"A0",X"91",X"4A",X"99",X"86",X"8A",X"19",
		X"95",X"0B",X"1A",X"97",X"8A",X"19",X"85",X"99",X"09",X"86",X"99",X"19",X"94",X"0B",X"80",X"48",
		X"B1",X"B3",X"7A",X"98",X"85",X"99",X"92",X"3C",X"94",X"0C",X"85",X"99",X"80",X"3A",X"A8",X"50",
		X"B9",X"34",X"C8",X"91",X"5A",X"91",X"A0",X"7A",X"89",X"13",X"AB",X"25",X"B8",X"90",X"79",X"90",
		X"91",X"3B",X"A8",X"78",X"A8",X"14",X"B9",X"83",X"2D",X"91",X"4A",X"A0",X"69",X"98",X"85",X"A8",
		X"91",X"4A",X"98",X"85",X"8A",X"89",X"26",X"B8",X"0A",X"50",X"B8",X"14",X"B9",X"82",X"4B",X"88",
		X"A4",X"4C",X"89",X"32",X"C9",X"16",X"AA",X"83",X"2C",X"91",X"4A",X"99",X"15",X"A9",X"91",X"7A",
		X"91",X"A3",X"2C",X"89",X"25",X"A9",X"1B",X"87",X"8A",X"19",X"96",X"8A",X"93",X"1B",X"09",X"86",
		X"8A",X"09",X"15",X"AA",X"85",X"8A",X"95",X"8A",X"80",X"49",X"98",X"93",X"3D",X"98",X"68",X"A0",
		X"90",X"7A",X"80",X"98",X"48",X"A0",X"92",X"3C",X"08",X"B3",X"7A",X"92",X"9B",X"07",X"99",X"88",
		X"48",X"A0",X"92",X"3B",X"8B",X"27",X"A9",X"83",X"2D",X"94",X"0C",X"21",X"D1",X"3C",X"84",X"9A",
		X"13",X"C9",X"13",X"A9",X"93",X"3C",X"A1",X"79",X"A1",X"A2",X"4C",X"88",X"23",X"B9",X"99",X"70",
		X"B2",X"8C",X"25",X"B8",X"1B",X"25",X"B9",X"1A",X"25",X"B8",X"1B",X"87",X"8A",X"1A",X"15",X"B8",
		X"80",X"4A",X"98",X"24",X"C8",X"83",X"0B",X"A6",X"0B",X"86",X"9A",X"04",X"A9",X"93",X"2B",X"00",
		X"D2",X"5B",X"80",X"A3",X"4D",X"08",X"94",X"1B",X"00",X"B8",X"78",X"A1",X"98",X"58",X"A1",X"A8",
		X"68",X"B1",X"0B",X"26",X"A9",X"1A",X"05",X"99",X"19",X"A2",X"6B",X"82",X"9A",X"94",X"4C",X"82",
		X"9A",X"16",X"A9",X"19",X"95",X"0B",X"88",X"48",X"B1",X"5A",X"A8",X"41",X"B9",X"05",X"AA",X"59",
		X"A3",X"0C",X"22",X"D8",X"49",X"A0",X"4A",X"A2",X"4B",X"89",X"15",X"A9",X"88",X"68",X"A0",X"90",
		X"59",X"91",X"B8",X"60",X"B1",X"0B",X"07",X"9A",X"19",X"13",X"BA",X"15",X"B9",X"58",X"B0",X"5A",
		X"98",X"22",X"B9",X"85",X"8B",X"06",X"AA",X"31",X"D0",X"4A",X"98",X"49",X"98",X"05",X"99",X"0A",
		X"24",X"C8",X"82",X"2C",X"90",X"59",X"99",X"32",X"CA",X"50",X"B9",X"50",X"B8",X"49",X"B3",X"3D",
		X"94",X"0B",X"09",X"16",X"A9",X"18",X"A0",X"69",X"91",X"99",X"40",X"B1",X"A8",X"79",X"90",X"94",
		X"0B",X"18",X"B5",X"2C",X"90",X"30",X"B0",X"A3",X"6C",X"88",X"48",X"B8",X"58",X"A9",X"23",X"BA",
		X"06",X"9A",X"95",X"1B",X"09",X"95",X"1C",X"01",X"9A",X"87",X"89",X"00",X"89",X"92",X"6B",X"82",
		X"B9",X"61",X"C0",X"1A",X"94",X"1B",X"08",X"94",X"1C",X"92",X"3B",X"B5",X"1C",X"85",X"A9",X"13",
		X"C9",X"22",X"BA",X"42",X"C8",X"83",X"2D",X"92",X"4B",X"98",X"87",X"99",X"09",X"24",X"C0",X"1A",
		X"A3",X"5B",X"92",X"AA",X"44",X"C8",X"19",X"93",X"3D",X"01",X"C0",X"6A",X"91",X"2B",X"94",X"0B",
		X"92",X"4A",X"99",X"07",X"99",X"09",X"31",X"C0",X"93",X"2C",X"98",X"68",X"A9",X"06",X"99",X"0A",
		X"32",X"C9",X"15",X"AA",X"04",X"8B",X"93",X"3C",X"98",X"50",X"B9",X"68",X"A9",X"14",X"A8",X"1A",
		X"A3",X"7B",X"82",X"9B",X"27",X"A9",X"1A",X"06",X"A9",X"19",X"04",X"A9",X"80",X"48",X"A8",X"94",
		X"3D",X"00",X"B4",X"2C",X"80",X"A5",X"0A",X"88",X"95",X"0A",X"01",X"AA",X"17",X"9A",X"29",X"A3",
		X"5C",X"80",X"93",X"2D",X"08",X"93",X"3D",X"00",X"B3",X"4C",X"09",X"86",X"99",X"88",X"48",X"A9",
		X"23",X"BB",X"27",X"AA",X"85",X"0B",X"1A",X"06",X"9A",X"19",X"85",X"8A",X"08",X"A5",X"1B",X"98",
		X"68",X"A8",X"04",X"9A",X"88",X"58",X"A8",X"85",X"8A",X"92",X"3B",X"B1",X"7A",X"A1",X"5A",X"A3",
		X"1D",X"13",X"C9",X"14",X"AA",X"14",X"AA",X"23",X"CA",X"06",X"99",X"1A",X"15",X"B9",X"03",X"8C",
		X"05",X"9A",X"83",X"1B",X"98",X"78",X"A9",X"40",X"B8",X"59",X"A8",X"14",X"A8",X"8A",X"51",X"C8",
		X"49",X"A0",X"4A",X"A2",X"3D",X"84",X"9A",X"85",X"9A",X"04",X"9B",X"32",X"C9",X"40",X"B9",X"25",
		X"A9",X"1B",X"17",X"A8",X"08",X"98",X"41",X"C1",X"1A",X"98",X"68",X"A1",X"8B",X"27",X"B8",X"1A",
		X"23",X"C9",X"13",X"AB",X"34",X"CA",X"16",X"A8",X"90",X"5A",X"98",X"59",X"99",X"31",X"B9",X"24",
		X"C8",X"92",X"5B",X"88",X"94",X"2C",X"08",X"A5",X"0B",X"09",X"07",X"9A",X"2A",X"86",X"8A",X"09",
		X"84",X"0B",X"09",X"87",X"8A",X"10",X"A9",X"17",X"A8",X"19",X"93",X"1C",X"92",X"3C",X"94",X"0B",
		X"93",X"3D",X"89",X"34",X"C9",X"04",X"8B",X"84",X"0B",X"88",X"68",X"B0",X"5A",X"A1",X"4A",X"A2",
		X"3C",X"98",X"40",X"B1",X"8B",X"62",X"D0",X"1B",X"15",X"A9",X"81",X"3B",X"A0",X"69",X"A0",X"59",
		X"A8",X"22",X"C8",X"82",X"4B",X"89",X"95",X"3E",X"01",X"99",X"93",X"5C",X"01",X"A9",X"69",X"91",
		X"8A",X"15",X"A9",X"18",X"99",X"42",X"C0",X"89",X"68",X"A8",X"83",X"2D",X"09",X"14",X"A9",X"88",
		X"59",X"98",X"94",X"2D",X"01",X"B1",X"6B",X"81",X"A0",X"6A",X"80",X"8A",X"25",X"B8",X"80",X"49",
		X"B0",X"59",X"A1",X"4C",X"83",X"8C",X"04",X"9A",X"04",X"AA",X"32",X"D9",X"14",X"99",X"0A",X"26",
		X"B8",X"2A",X"A2",X"7B",X"88",X"03",X"9B",X"06",X"9A",X"04",X"9A",X"82",X"3C",X"89",X"25",X"BA",
		X"15",X"AA",X"14",X"AB",X"25",X"BA",X"33",X"E8",X"49",X"A1",X"3C",X"91",X"4A",X"89",X"86",X"99",
		X"19",X"93",X"3D",X"00",X"9A",X"27",X"A8",X"1A",X"94",X"1C",X"10",X"B1",X"6A",X"98",X"04",X"99",
		X"89",X"41",X"B8",X"93",X"4C",X"89",X"25",X"B9",X"2C",X"24",X"B9",X"88",X"68",X"A1",X"9A",X"52",
		X"C0",X"1B",X"97",X"8A",X"18",X"A1",X"5A",X"91",X"A1",X"5A",X"90",X"94",X"0B",X"88",X"50",X"B9",
		X"16",X"AA",X"14",X"B9",X"31",X"D0",X"4A",X"A2",X"3D",X"93",X"1C",X"84",X"8A",X"92",X"4B",X"82",
		X"9C",X"07",X"8A",X"10",X"B0",X"59",X"90",X"98",X"58",X"A0",X"92",X"4C",X"00",X"B3",X"4C",X"88",
		X"04",X"9A",X"80",X"59",X"91",X"A9",X"78",X"A1",X"A8",X"69",X"90",X"91",X"4A",X"91",X"B0",X"79",
		X"91",X"A0",X"5A",X"A1",X"4A",X"98",X"05",X"A9",X"82",X"3C",X"88",X"95",X"1C",X"18",X"A1",X"6B",
		X"82",X"B0",X"6A",X"90",X"3A",X"98",X"87",X"99",X"09",X"31",X"BA",X"26",X"AA",X"83",X"2C",X"90",
		X"69",X"A8",X"48",X"B8",X"68",X"B0",X"30",X"B8",X"94",X"1B",X"0A",X"07",X"99",X"1B",X"25",X"BA",
		X"15",X"AA",X"14",X"A9",X"90",X"79",X"91",X"A0",X"59",X"A8",X"30",X"B9",X"06",X"8A",X"88",X"58",
		X"A0",X"A0",X"79",X"91",X"8B",X"26",X"A9",X"19",X"A2",X"5A",X"92",X"99",X"93",X"5C",X"01",X"A9",
		X"68",X"B8",X"31",X"B9",X"06",X"9A",X"14",X"B9",X"86",X"9A",X"04",X"9A",X"84",X"0B",X"91",X"59",
		X"99",X"04",X"9B",X"32",X"E8",X"48",X"A9",X"14",X"9A",X"92",X"5B",X"89",X"16",X"A9",X"2B",X"95",
		X"2C",X"81",X"A2",X"3C",X"89",X"15",X"A9",X"88",X"68",X"A9",X"14",X"A9",X"93",X"3C",X"99",X"51",
		X"BA",X"17",X"A9",X"04",X"A9",X"84",X"8A",X"91",X"4A",X"99",X"26",X"B8",X"89",X"68",X"A8",X"84",
		X"0B",X"88",X"58",X"A1",X"A8",X"79",X"91",X"A0",X"5A",X"98",X"04",X"8A",X"00",X"B1",X"7A",X"81",
		X"8A",X"93",X"5B",X"89",X"23",X"C9",X"85",X"1C",X"00",X"A1",X"6A",X"99",X"32",X"D8",X"49",X"A3",
		X"1D",X"83",X"0B",X"93",X"3E",X"84",X"AA",X"40",X"B0",X"4A",X"A0",X"59",X"98",X"85",X"99",X"92",
		X"4B",X"89",X"15",X"A9",X"91",X"5A",X"99",X"33",X"CA",X"07",X"9A",X"83",X"1B",X"98",X"68",X"A9",
		X"24",X"B8",X"8A",X"61",X"C0",X"89",X"33",X"D0",X"1B",X"85",X"8A",X"1A",X"06",X"A9",X"81",X"5A",
		X"98",X"84",X"1C",X"08",X"94",X"1C",X"18",X"A2",X"4B",X"88",X"A4",X"4D",X"01",X"A9",X"50",X"B1",
		X"0B",X"15",X"A9",X"1A",X"16",X"A9",X"09",X"33",X"E0",X"91",X"4A",X"A0",X"49",X"B2",X"4B",X"A5",
		X"0C",X"03",X"B9",X"58",X"B1",X"4B",X"88",X"95",X"0B",X"80",X"59",X"A8",X"58",X"B0",X"49",X"B0",
		X"69",X"90",X"92",X"3D",X"09",X"85",X"8A",X"18",X"99",X"41",X"B0",X"1D",X"07",X"99",X"1A",X"04",
		X"9A",X"10",X"B1",X"7A",X"91",X"90",X"4A",X"98",X"13",X"B0",X"A8",X"70",X"B8",X"85",X"8A",X"91",
		X"5A",X"99",X"24",X"B8",X"0B",X"37",X"B8",X"0A",X"41",X"B8",X"1B",X"87",X"8A",X"20",X"AA",X"07",
		X"99",X"28",X"B0",X"7A",X"80",X"92",X"2C",X"09",X"05",X"99",X"09",X"96",X"0B",X"19",X"85",X"9A",
		X"81",X"5A",X"91",X"A1",X"5B",X"88",X"84",X"8A",X"90",X"7A",X"89",X"14",X"A9",X"80",X"5A",X"98",
		X"48",X"A9",X"32",X"CA",X"25",X"AB",X"16",X"AA",X"14",X"AA",X"23",X"D9",X"32",X"D8",X"83",X"1C",
		X"83",X"1B",X"99",X"60",X"B9",X"50",X"B9",X"41",X"B9",X"85",X"0B",X"94",X"1B",X"89",X"51",X"C8",
		X"84",X"0B",X"1A",X"97",X"89",X"09",X"95",X"0B",X"19",X"95",X"1C",X"08",X"95",X"0B",X"08",X"93",
		X"3D",X"00",X"9A",X"17",X"99",X"18",X"A8",X"79",X"91",X"A1",X"4B",X"88",X"85",X"8A",X"09",X"05",
		X"99",X"92",X"3C",X"98",X"58",X"B8",X"69",X"A0",X"30",X"B0",X"A0",X"79",X"A8",X"48",X"A8",X"59",
		X"A8",X"31",X"B9",X"87",X"8A",X"94",X"0B",X"80",X"6A",X"98",X"13",X"AB",X"25",X"BA",X"25",X"B9",
		X"81",X"6A",X"98",X"04",X"9B",X"05",X"99",X"91",X"5B",X"89",X"16",X"A9",X"81",X"3A",X"99",X"07",
		X"99",X"89",X"41",X"C1",X"1B",X"A3",X"6B",X"81",X"A9",X"60",X"B8",X"03",X"8A",X"A2",X"7A",X"88",
		X"95",X"8B",X"85",X"8A",X"81",X"3A",X"A9",X"35",X"B8",X"99",X"78",X"A1",X"8B",X"44",X"C8",X"19",
		X"92",X"4C",X"00",X"A1",X"5A",X"A8",X"40",X"A9",X"15",X"A9",X"92",X"3B",X"B2",X"6A",X"B1",X"6A",
		X"98",X"48",X"A9",X"40",X"A9",X"05",X"99",X"8A",X"43",X"D0",X"1B",X"07",X"A9",X"19",X"84",X"0B",
		X"09",X"05",X"99",X"89",X"41",X"B8",X"93",X"4C",X"A3",X"4D",X"83",X"0B",X"89",X"41",X"B0",X"B2",
		X"7A",X"91",X"A4",X"1C",X"88",X"40",X"B9",X"07",X"99",X"1A",X"85",X"8A",X"88",X"48",X"A9",X"15",
		X"A8",X"8A",X"51",X"B8",X"93",X"3D",X"90",X"69",X"A8",X"22",X"BA",X"41",X"C9",X"50",X"B8",X"85",
		X"8A",X"09",X"15",X"A9",X"89",X"50",X"A0",X"A0",X"79",X"98",X"83",X"0B",X"92",X"4B",X"A8",X"60",
		X"A8",X"A3",X"5C",X"09",X"85",X"8A",X"01",X"B9",X"61",X"B0",X"8A",X"34",X"C0",X"8A",X"42",X"C0",
		X"8A",X"43",X"D0",X"89",X"32",X"D0",X"0A",X"16",X"A8",X"1A",X"94",X"1C",X"08",X"85",X"9A",X"08",
		X"59",X"A8",X"31",X"C8",X"5A",X"94",X"8C",X"13",X"BA",X"32",X"C9",X"05",X"99",X"93",X"2C",X"A5",
		X"0B",X"94",X"1C",X"83",X"1C",X"93",X"1B",X"A4",X"4C",X"90",X"49",X"A8",X"23",X"C9",X"05",X"9A",
		X"85",X"8A",X"90",X"58",X"A8",X"94",X"1B",X"0A",X"87",X"8A",X"10",X"AA",X"37",X"B8",X"80",X"49",
		X"A8",X"85",X"0B",X"18",X"B2",X"7A",X"92",X"9A",X"35",X"C8",X"09",X"31",X"C8",X"84",X"8A",X"1A",
		X"07",X"99",X"91",X"4B",X"08",X"A3",X"5C",X"82",X"B8",X"68",X"A1",X"8A",X"24",X"C0",X"1B",X"86",
		X"8A",X"19",X"95",X"8A",X"92",X"3B",X"99",X"51",X"BA",X"35",X"B9",X"91",X"7A",X"88",X"84",X"8B",
		X"82",X"3C",X"89",X"07",X"99",X"1A",X"86",X"9A",X"08",X"22",X"C0",X"09",X"A4",X"4C",X"01",X"A9",
		X"50",X"B1",X"99",X"68",X"A8",X"84",X"8B",X"85",X"8A",X"84",X"8A",X"0A",X"17",X"A9",X"2A",X"84",
		X"0C",X"19",X"04",X"A9",X"84",X"8B",X"86",X"8A",X"88",X"59",X"98",X"04",X"A9",X"93",X"2B",X"A8",
		X"78",X"B0",X"5A",X"A2",X"3C",X"94",X"8B",X"23",X"E8",X"49",X"A0",X"21",X"B0",X"90",X"69",X"98",
		X"94",X"1B",X"90",X"69",X"A0",X"93",X"4C",X"81",X"A9",X"60",X"B8",X"30",X"C8",X"40",X"C8",X"48",
		X"B2",X"3C",X"A2",X"4B",X"98",X"58",X"B0",X"59",X"A8",X"23",X"C9",X"85",X"8A",X"09",X"25",X"B9",
		X"95",X"0A",X"08",X"B4",X"3C",X"81",X"B0",X"79",X"91",X"8B",X"26",X"B8",X"2A",X"A4",X"3D",X"82",
		X"B0",X"59",X"A0",X"82",X"2B",X"01",X"D8",X"60",X"B1",X"0B",X"16",X"B8",X"09",X"48",X"A8",X"31",
		X"B8",X"A3",X"5B",X"A9",X"71",X"B0",X"98",X"69",X"A8",X"23",X"B9",X"A4",X"3C",X"A0",X"69",X"99",
		X"15",X"AA",X"04",X"9B",X"24",X"BA",X"32",X"D9",X"15",X"A9",X"81",X"4A",X"B1",X"6A",X"89",X"05",
		X"99",X"89",X"33",X"D8",X"1B",X"17",X"A8",X"1A",X"83",X"3E",X"01",X"B0",X"6A",X"88",X"83",X"0B",
		X"89",X"34",X"C0",X"8A",X"35",X"C0",X"1B",X"86",X"8A",X"10",X"B8",X"79",X"90",X"82",X"8B",X"15",
		X"B9",X"40",X"C8",X"48",X"A0",X"92",X"4B",X"88",X"95",X"0B",X"91",X"5A",X"89",X"05",X"AA",X"41",
		X"C9",X"14",X"A8",X"98",X"58",X"A0",X"A3",X"5C",X"08",X"94",X"0B",X"92",X"3B",X"A9",X"52",X"B0",
		X"1E",X"06",X"9A",X"81",X"3A",X"91",X"B3",X"5B",X"A8",X"68",X"A0",X"94",X"0B",X"94",X"1C",X"95",
		X"0B",X"84",X"9B",X"48",X"B3",X"1D",X"21",X"C1",X"3C",X"95",X"99",X"82",X"1B",X"88",X"58",X"A8",
		X"94",X"2C",X"09",X"86",X"8A",X"19",X"96",X"99",X"90",X"59",X"90",X"98",X"69",X"91",X"99",X"40",
		X"B1",X"A0",X"7A",X"81",X"A8",X"69",X"90",X"89",X"23",X"C8",X"0A",X"41",X"B0",X"1A",X"B2",X"79",
		X"91",X"09",X"A9",X"71",X"B0",X"8A",X"60",X"B0",X"92",X"4B",X"98",X"41",X"C8",X"94",X"2C",X"88",
		X"30",X"D8",X"58",X"A0",X"93",X"1C",X"89",X"42",X"C0",X"98",X"68",X"A0",X"89",X"40",X"B0",X"98",
		X"79",X"90",X"94",X"0B",X"09",X"25",X"B9",X"92",X"5A",X"98",X"96",X"8A",X"1A",X"07",X"A9",X"00",
		X"3A",X"B2",X"5B",X"A2",X"4B",X"A2",X"4B",X"A0",X"69",X"99",X"23",X"C9",X"32",X"D9",X"40",X"B9",
		X"25",X"B8",X"89",X"50",X"A0",X"0B",X"87",X"8A",X"28",X"A9",X"51",X"C1",X"0B",X"16",X"A9",X"1A",
		X"05",X"A8",X"09",X"31",X"B8",X"A3",X"5B",X"A8",X"78",X"A1",X"A0",X"6A",X"98",X"13",X"9A",X"0B",
		X"45",X"C0",X"90",X"5A",X"98",X"13",X"BA",X"16",X"A9",X"92",X"4B",X"A2",X"5B",X"99",X"42",X"C0",
		X"8A",X"43",X"D0",X"0A",X"86",X"8A",X"10",X"A9",X"34",X"C8",X"1B",X"34",X"C9",X"14",X"A9",X"94",
		X"0A",X"0A",X"17",X"A8",X"0A",X"15",X"A9",X"80",X"4A",X"A1",X"5A",X"A0",X"5A",X"98",X"48",X"A8",
		X"85",X"8A",X"91",X"4A",X"99",X"17",X"A8",X"0A",X"15",X"B9",X"05",X"99",X"09",X"85",X"8A",X"0A",
		X"25",X"B8",X"1B",X"07",X"8B",X"29",X"93",X"2D",X"91",X"4A",X"98",X"23",X"C9",X"87",X"99",X"80",
		X"4A",X"98",X"31",X"BA",X"07",X"9A",X"84",X"0B",X"85",X"9B",X"14",X"9A",X"92",X"4A",X"91",X"C1",
		X"7A",X"92",X"9A",X"41",X"C0",X"0A",X"41",X"B0",X"1A",X"A1",X"79",X"91",X"0A",X"90",X"79",X"91",
		X"0B",X"06",X"9A",X"08",X"30",X"C8",X"58",X"B1",X"3C",X"84",X"A9",X"49",X"B1",X"5A",X"98",X"21",
		X"A9",X"86",X"8B",X"05",X"AA",X"23",X"D8",X"49",X"A8",X"31",X"B9",X"84",X"3D",X"81",X"B2",X"6A",
		X"91",X"B0",X"79",X"91",X"99",X"32",X"D8",X"83",X"1B",X"90",X"59",X"A8",X"58",X"A9",X"24",X"C0",
		X"90",X"5A",X"98",X"31",X"C9",X"24",X"BA",X"07",X"99",X"90",X"59",X"98",X"93",X"3D",X"81",X"A1",
		X"5A",X"99",X"05",X"8A",X"10",X"C0",X"7A",X"92",X"8A",X"83",X"3D",X"01",X"99",X"93",X"4B",X"82",
		X"C9",X"78",X"A1",X"8A",X"42",X"D0",X"09",X"22",X"C0",X"98",X"58",X"A1",X"99",X"68",X"A0",X"92",
		X"3D",X"88",X"31",X"C8",X"83",X"2C",X"8A",X"42",X"CA",X"34",X"BA",X"06",X"9A",X"88",X"50",X"B8",
		X"04",X"9B",X"06",X"9A",X"84",X"0B",X"80",X"4A",X"A2",X"4B",X"A0",X"79",X"A0",X"4A",X"A4",X"8B",
		X"23",X"C9",X"05",X"A9",X"04",X"A9",X"81",X"5A",X"91",X"9A",X"36",X"B8",X"2A",X"A1",X"7A",X"81",
		X"B0",X"69",X"98",X"84",X"8A",X"00",X"B3",X"5B",X"81",X"B8",X"79",X"98",X"04",X"9A",X"08",X"48",
		X"C2",X"2D",X"84",X"99",X"81",X"3B",X"99",X"35",X"C9",X"14",X"AA",X"32",X"D9",X"32",X"D8",X"85",
		X"8A",X"92",X"2B",X"89",X"42",X"C9",X"86",X"8A",X"88",X"58",X"A0",X"A2",X"5B",X"98",X"24",X"B8",
		X"98",X"78",X"A1",X"8B",X"26",X"B8",X"1A",X"87",X"99",X"08",X"94",X"0B",X"10",X"B1",X"7A",X"81",
		X"9A",X"25",X"B8",X"88",X"48",X"A9",X"24",X"B9",X"86",X"9A",X"04",X"9A",X"85",X"99",X"88",X"59",
		X"98",X"94",X"1B",X"0A",X"24",X"B8",X"A1",X"79",X"A2",X"9A",X"35",X"C9",X"04",X"9A",X"85",X"8B",
		X"05",X"AA",X"31",X"B9",X"05",X"99",X"98",X"51",X"C0",X"2A",X"A1",X"7A",X"92",X"9A",X"42",X"C8",
		X"80",X"49",X"A8",X"59",X"A0",X"5A",X"A1",X"4A",X"A0",X"48",X"B8",X"40",X"A8",X"A4",X"2C",X"91",
		X"5A",X"A0",X"31",X"C9",X"24",X"BA",X"06",X"9B",X"15",X"AA",X"04",X"8B",X"85",X"8A",X"93",X"2C",
		X"09",X"87",X"99",X"09",X"05",X"A9",X"80",X"49",X"90",X"A2",X"6B",X"82",X"B9",X"43",X"D8",X"09",
		X"32",X"D8",X"03",X"8C",X"05",X"9B",X"14",X"B9",X"31",X"C9",X"32",X"BA",X"87",X"8A",X"2A",X"95",
		X"1C",X"01",X"B0",X"7A",X"81",X"A8",X"58",X"A0",X"90",X"59",X"A2",X"8B",X"17",X"A9",X"2A",X"85",
		X"A9",X"03",X"9A",X"82",X"3C",X"89",X"34",X"D8",X"49",X"A8",X"58",X"A9",X"22",X"AB",X"07",X"8A",
		X"92",X"4B",X"88",X"94",X"2C",X"00",X"9B",X"17",X"8A",X"10",X"9A",X"83",X"7B",X"82",X"B8",X"79",
		X"98",X"11",X"A9",X"05",X"99",X"91",X"5A",X"A0",X"5A",X"90",X"4A",X"A3",X"1D",X"85",X"9A",X"13",
		X"BA",X"15",X"A9",X"82",X"3C",X"A2",X"5A",X"99",X"16",X"A9",X"09",X"41",X"C0",X"0A",X"06",X"99",
		X"09",X"85",X"99",X"0A",X"34",X"C8",X"0A",X"51",X"C0",X"1B",X"06",X"99",X"09",X"04",X"9A",X"09",
		X"58",X"A8",X"14",X"BA",X"24",X"B9",X"84",X"0B",X"A5",X"1B",X"89",X"35",X"C9",X"14",X"AA",X"14",
		X"AB",X"07",X"99",X"09",X"30",X"B9",X"34",X"CA",X"24",X"AA",X"83",X"2C",X"99",X"53",X"D0",X"0B",
		X"26",X"B8",X"1B",X"24",X"A9",X"1B",X"85",X"2D",X"01",X"A9",X"51",X"C0",X"1A",X"95",X"0B",X"19",
		X"04",X"9A",X"80",X"59",X"A8",X"69",X"A8",X"32",X"C8",X"2A",X"A2",X"7A",X"81",X"9A",X"85",X"1B",
		X"01",X"C8",X"68",X"A1",X"A0",X"5A",X"90",X"84",X"9A",X"30",X"D2",X"2D",X"03",X"AA",X"32",X"D8",
		X"03",X"8B",X"95",X"1B",X"A3",X"5C",X"88",X"31",X"C9",X"05",X"99",X"89",X"50",X"A9",X"84",X"2D",
		X"08",X"94",X"0B",X"09",X"15",X"A9",X"0A",X"51",X"B0",X"0C",X"17",X"A9",X"08",X"21",X"B9",X"05",
		X"9A",X"05",X"AA",X"40",X"C0",X"4A",X"98",X"13",X"A9",X"90",X"79",X"91",X"9A",X"51",X"C1",X"99",
		X"50",X"B1",X"0A",X"95",X"1C",X"09",X"31",X"B9",X"07",X"99",X"0A",X"33",X"D0",X"98",X"58",X"A0",
		X"90",X"5A",X"A0",X"59",X"A8",X"58",X"A1",X"99",X"41",X"C0",X"0A",X"24",X"B8",X"98",X"79",X"98",
		X"13",X"B9",X"92",X"6A",X"98",X"85",X"8A",X"0A",X"16",X"A8",X"0B",X"17",X"A9",X"28",X"B1",X"6A",
		X"90",X"02",X"9B",X"33",X"D9",X"32",X"D8",X"49",X"B4",X"8B",X"32",X"E1",X"2C",X"03",X"B8",X"5A",
		X"A1",X"4A",X"88",X"94",X"0A",X"89",X"42",X"C0",X"1C",X"85",X"0B",X"19",X"96",X"8A",X"80",X"4A",
		X"98",X"32",X"D0",X"98",X"68",X"A0",X"0A",X"84",X"2C",X"01",X"B9",X"43",X"D0",X"19",X"A8",X"78",
		X"A0",X"92",X"3C",X"89",X"40",X"A9",X"86",X"8A",X"19",X"94",X"3E",X"00",X"A1",X"4A",X"90",X"92",
		X"3D",X"92",X"3B",X"B3",X"5C",X"91",X"4B",X"89",X"33",X"C9",X"93",X"5B",X"88",X"A7",X"0B",X"84",
		X"8B",X"81",X"5A",X"90",X"A3",X"4C",X"01",X"C0",X"69",X"A2",X"A8",X"59",X"98",X"83",X"1C",X"08",
		X"94",X"1B",X"A1",X"6A",X"98",X"24",X"C0",X"8A",X"35",X"C8",X"09",X"40",X"B8",X"85",X"8A",X"0A",
		X"34",X"C0",X"98",X"58",X"A0",X"A3",X"3C",X"A3",X"3D",X"A3",X"3C",X"A1",X"59",X"B0",X"58",X"B8",
		X"58",X"A9",X"23",X"C9",X"32",X"D9",X"24",X"BA",X"15",X"AA",X"05",X"9A",X"83",X"2C",X"09",X"96",
		X"0B",X"18",X"A3",X"4C",X"81",X"A9",X"51",X"C0",X"90",X"69",X"91",X"A8",X"40",X"B0",X"0B",X"43",
		X"CA",X"05",X"8B",X"85",X"8A",X"81",X"4B",X"89",X"06",X"99",X"89",X"41",X"B0",X"8B",X"45",X"C8",
		X"09",X"24",X"C8",X"19",X"94",X"1B",X"00",X"B0",X"79",X"98",X"84",X"0B",X"88",X"40",X"B9",X"16",
		X"A9",X"85",X"9A",X"85",X"99",X"92",X"3B",X"99",X"33",X"E8",X"59",X"B4",X"8B",X"23",X"D8",X"30",
		X"C8",X"22",X"B8",X"93",X"4C",X"0A",X"07",X"9A",X"83",X"1B",X"A2",X"5A",X"A0",X"69",X"A8",X"14",
		X"B9",X"05",X"AA",X"14",X"AA",X"85",X"0B",X"18",X"A5",X"0B",X"90",X"69",X"98",X"85",X"99",X"93",
		X"1B",X"0B",X"27",X"A8",X"0A",X"17",X"A9",X"09",X"31",X"B8",X"A4",X"3C",X"82",X"C8",X"51",X"C0",
		X"1B",X"15",X"B8",X"89",X"42",X"C8",X"81",X"3A",X"98",X"A4",X"6B",X"93",X"BA",X"70",X"B8",X"22",
		X"C9",X"23",X"B8",X"98",X"79",X"90",X"92",X"4C",X"89",X"15",X"A9",X"09",X"32",X"C0",X"A8",X"78",
		X"A8",X"04",X"AA",X"14",X"A9",X"92",X"5A",X"91",X"9B",X"27",X"9A",X"29",X"A3",X"5C",X"80",X"92",
		X"3D",X"09",X"05",X"9A",X"82",X"3C",X"00",X"B3",X"5C",X"90",X"30",X"B1",X"A9",X"70",X"B8",X"84",
		X"1B",X"09",X"A7",X"0B",X"1A",X"24",X"B9",X"1B",X"52",X"C9",X"04",X"99",X"92",X"4C",X"89",X"17",
		X"A8",X"08",X"A3",X"3C",X"81",X"B0",X"69",X"99",X"05",X"99",X"91",X"5A",X"90",X"92",X"5C",X"00",
		X"A0",X"59",X"90",X"8A",X"34",X"C0",X"8A",X"42",X"D0",X"09",X"30",X"B0",X"A2",X"6A",X"99",X"16",
		X"A9",X"29",X"B2",X"7A",X"92",X"9A",X"33",X"D8",X"1B",X"16",X"99",X"09",X"05",X"A9",X"84",X"8A",
		X"90",X"69",X"99",X"14",X"A9",X"80",X"49",X"B2",X"4C",X"92",X"3D",X"92",X"3B",X"A0",X"69",X"A8",
		X"59",X"99",X"31",X"BA",X"35",X"BA",X"15",X"AA",X"15",X"BA",X"50",X"B9",X"40",X"B8",X"23",X"C8",
		X"91",X"7A",X"80",X"A3",X"2C",X"89",X"33",X"D9",X"04",X"8A",X"92",X"4B",X"99",X"35",X"C8",X"93",
		X"4C",X"81",X"A9",X"60",X"B0",X"90",X"69",X"90",X"A1",X"6A",X"98",X"22",X"C8",X"04",X"AA",X"23",
		X"C8",X"92",X"4B",X"B5",X"1D",X"04",X"A9",X"03",X"9A",X"80",X"59",X"B0",X"69",X"A8",X"31",X"BA",
		X"34",X"BB",X"17",X"9A",X"83",X"1C",X"95",X"0B",X"92",X"4A",X"99",X"06",X"A8",X"0A",X"26",X"B8",
		X"1A",X"86",X"9A",X"19",X"13",X"BA",X"85",X"1B",X"09",X"A7",X"1C",X"10",X"B0",X"69",X"90",X"0A",
		X"04",X"8A",X"18",X"B1",X"79",X"91",X"0B",X"85",X"1C",X"08",X"94",X"1C",X"80",X"39",X"A9",X"68",
		X"A8",X"48",X"A9",X"06",X"99",X"1A",X"84",X"0B",X"08",X"A6",X"0A",X"09",X"95",X"1C",X"09",X"05",
		X"99",X"90",X"59",X"90",X"A1",X"5A",X"80",X"B1",X"7A",X"88",X"84",X"8A",X"09",X"86",X"99",X"88",
		X"48",X"A9",X"24",X"B9",X"95",X"0B",X"93",X"4C",X"88",X"86",X"99",X"88",X"31",X"C8",X"85",X"8A",
		X"90",X"69",X"A8",X"22",X"BA",X"68",X"B1",X"4C",X"84",X"9A",X"82",X"2B",X"91",X"5A",X"90",X"A6",
		X"0B",X"11",X"C8",X"68",X"A1",X"8A",X"15",X"A9",X"19",X"95",X"0B",X"09",X"24",X"B9",X"84",X"0C",
		X"83",X"2D",X"09",X"05",X"99",X"0A",X"87",X"8A",X"10",X"A9",X"68",X"A1",X"99",X"33",X"D0",X"0A",
		X"85",X"0B",X"88",X"40",X"A9",X"86",X"8A",X"93",X"2D",X"94",X"1C",X"83",X"0B",X"92",X"4B",X"99",
		X"34",X"D9",X"40",X"B8",X"14",X"AB",X"25",X"AA",X"83",X"4C",X"81",X"A9",X"60",X"B1",X"0B",X"87",
		X"8A",X"09",X"15",X"B8",X"09",X"48",X"A8",X"31",X"D8",X"59",X"A1",X"3C",X"90",X"59",X"91",X"A8",
		X"69",X"98",X"03",X"9A",X"91",X"6A",X"89",X"86",X"99",X"09",X"31",X"C0",X"92",X"4B",X"99",X"34",
		X"C8",X"90",X"79",X"A8",X"30",X"B9",X"50",X"C1",X"3B",X"B6",X"0B",X"80",X"48",X"A0",X"99",X"60",
		X"B8",X"03",X"8C",X"15",X"AA",X"14",X"BA",X"24",X"A9",X"89",X"42",X"C0",X"A0",X"79",X"91",X"99",
		X"50",X"C1",X"0B",X"15",X"9A",X"28",X"99",X"83",X"5C",X"01",X"A9",X"25",X"C0",X"90",X"59",X"A8",
		X"04",X"99",X"92",X"3B",X"A9",X"70",X"B9",X"33",X"CA",X"15",X"9A",X"1B",X"26",X"A9",X"0A",X"34",
		X"C0",X"98",X"58",X"B2",X"0C",X"16",X"A9",X"80",X"38",X"A8",X"91",X"7A",X"88",X"94",X"0B",X"88",
		X"68",X"A9",X"14",X"A9",X"82",X"2B",X"B3",X"7B",X"90",X"5A",X"A2",X"3D",X"84",X"9A",X"85",X"99",
		X"82",X"1B",X"91",X"6A",X"98",X"13",X"AA",X"93",X"6B",X"99",X"60",X"B8",X"85",X"8A",X"80",X"49",
		X"B0",X"6A",X"98",X"48",X"A1",X"A8",X"68",X"A8",X"03",X"9A",X"91",X"7A",X"88",X"94",X"2D",X"80",
		X"3A",X"A0",X"69",X"99",X"13",X"A8",X"A8",X"78",X"A1",X"A0",X"7A",X"90",X"03",X"A9",X"92",X"4B",
		X"88",X"A7",X"0A",X"98",X"34",X"C8",X"18",X"9A",X"04",X"2B",X"02",X"A9",X"9C",X"55",X"C0",X"19",
		X"A0",X"7A",X"81",X"A8",X"40",X"B1",X"99",X"42",X"C0",X"0B",X"16",X"9A",X"1A",X"15",X"A9",X"88",
		X"69",X"98",X"04",X"9A",X"88",X"58",X"98",X"90",X"7A",X"80",X"A2",X"3C",X"92",X"3D",X"93",X"1C",
		X"85",X"9A",X"21",X"C0",X"4A",X"A0",X"48",X"A0",X"91",X"6A",X"91",X"A2",X"4C",X"80",X"A3",X"4C",
		X"91",X"3A",X"B1",X"7A",X"89",X"22",X"BA",X"26",X"A9",X"0A",X"25",X"B9",X"04",X"9A",X"93",X"4C",
		X"92",X"3D",X"91",X"5A",X"98",X"84",X"0B",X"80",X"59",X"A9",X"26",X"A9",X"0A",X"34",X"C9",X"03",
		X"8C",X"23",X"E8",X"49",X"A0",X"49",X"A8",X"23",X"B8",X"0B",X"87",X"0B",X"20",X"AB",X"45",X"C0",
		X"88",X"38",X"B8",X"24",X"B9",X"89",X"53",X"D0",X"19",X"A9",X"61",X"B8",X"29",X"B0",X"78",X"A1",
		X"99",X"50",X"B0",X"89",X"50",X"B1",X"A8",X"79",X"98",X"21",X"B9",X"68",X"B0",X"49",X"B1",X"5A",
		X"A1",X"4B",X"93",X"0C",X"05",X"B9",X"48",X"A8",X"05",X"A8",X"90",X"59",X"90",X"8A",X"51",X"B0",
		X"0B",X"07",X"99",X"1A",X"14",X"B8",X"0A",X"35",X"C8",X"88",X"40",X"B1",X"A8",X"78",X"A8",X"03",
		X"9B",X"87",X"8A",X"81",X"2A",X"88",X"A3",X"7B",X"88",X"85",X"9A",X"85",X"99",X"82",X"1C",X"84",
		X"9B",X"41",X"C8",X"31",X"C9",X"23",X"C9",X"14",X"AA",X"86",X"8A",X"09",X"40",X"B0",X"92",X"4B",
		X"A8",X"68",X"A9",X"06",X"99",X"88",X"59",X"98",X"85",X"99",X"0A",X"15",X"A9",X"88",X"41",X"C1",
		X"8A",X"41",X"C9",X"14",X"9A",X"09",X"41",X"BA",X"15",X"9B",X"07",X"99",X"0A",X"15",X"A9",X"83",
		X"0B",X"90",X"79",X"91",X"A8",X"68",X"A0",X"1B",X"87",X"99",X"18",X"89",X"82",X"4B",X"82",X"A9",
		X"92",X"7A",X"80",X"A3",X"4D",X"08",X"94",X"0B",X"88",X"40",X"B9",X"34",X"C8",X"93",X"2C",X"89",
		X"51",X"C0",X"90",X"6A",X"98",X"49",X"99",X"15",X"A9",X"2A",X"96",X"0C",X"19",X"13",X"B9",X"1B",
		X"17",X"99",X"1A",X"86",X"99",X"88",X"30",X"B8",X"86",X"8A",X"90",X"58",X"A8",X"92",X"6B",X"81",
		X"B1",X"7A",X"91",X"09",X"A2",X"5A",X"90",X"93",X"2D",X"94",X"1C",X"82",X"1B",X"A4",X"3D",X"92",
		X"2C",X"84",X"8C",X"21",X"C1",X"3D",X"03",X"AA",X"23",X"C9",X"23",X"C9",X"40",X"C8",X"31",X"C8",
		X"13",X"AA",X"92",X"7A",X"98",X"48",X"A9",X"15",X"AA",X"04",X"8B",X"95",X"0A",X"08",X"B4",X"5C",
		X"81",X"09",X"98",X"25",X"B8",X"18",X"B0",X"79",X"98",X"85",X"99",X"18",X"A0",X"68",X"B2",X"0C",
		X"06",X"9A",X"19",X"85",X"99",X"88",X"31",X"B8",X"A5",X"2C",X"08",X"A4",X"2C",X"80",X"94",X"0B",
		X"89",X"42",X"B9",X"96",X"0B",X"95",X"1C",X"09",X"14",X"A9",X"89",X"50",X"B9",X"41",X"C8",X"30",
		X"BA",X"51",X"B8",X"90",X"79",X"91",X"8B",X"35",X"C0",X"1B",X"05",X"9A",X"82",X"2C",X"93",X"3C",
		X"98",X"40",X"C0",X"5A",X"98",X"49",X"99",X"23",X"B8",X"A0",X"79",X"91",X"B2",X"6B",X"80",X"A5",
		X"0B",X"08",X"85",X"8B",X"82",X"3C",X"A2",X"5A",X"B2",X"4B",X"A5",X"0C",X"83",X"0A",X"98",X"68",
		X"A1",X"A1",X"5A",X"91",X"B0",X"79",X"91",X"8A",X"83",X"4C",X"01",X"99",X"93",X"4C",X"09",X"86",
		X"99",X"88",X"48",X"A9",X"05",X"9A",X"05",X"AA",X"05",X"9A",X"84",X"8A",X"94",X"1B",X"90",X"69",
		X"A8",X"48",X"A8",X"85",X"8A",X"88",X"40",X"C8",X"31",X"B0",X"B1",X"7A",X"88",X"94",X"2C",X"80",
		X"A5",X"0B",X"92",X"4A",X"99",X"07",X"99",X"91",X"4A",X"98",X"05",X"9A",X"09",X"16",X"A9",X"80",
		X"49",X"B0",X"69",X"B1",X"4B",X"94",X"0C",X"04",X"AA",X"23",X"C8",X"82",X"2C",X"80",X"49",X"B0",
		X"69",X"A8",X"31",X"B9",X"06",X"9B",X"14",X"9A",X"90",X"68",X"A1",X"9A",X"36",X"C8",X"29",X"98",
		X"40",X"B0",X"0A",X"50",X"B8",X"84",X"1B",X"08",X"B6",X"2D",X"09",X"30",X"B9",X"25",X"AA",X"86",
		X"99",X"94",X"0B",X"84",X"8B",X"84",X"1C",X"09",X"23",X"C8",X"90",X"79",X"91",X"A8",X"69",X"98",
		X"11",X"B9",X"50",X"B8",X"23",X"C8",X"2C",X"87",X"99",X"19",X"93",X"2C",X"01",X"99",X"92",X"7A",
		X"81",X"89",X"A0",X"68",X"A1",X"9A",X"52",X"D0",X"1B",X"15",X"A9",X"18",X"99",X"42",X"C0",X"89",
		X"25",X"C0",X"1B",X"06",X"A8",X"1A",X"85",X"99",X"09",X"05",X"9A",X"81",X"3A",X"9A",X"43",X"CA",
		X"15",X"AA",X"15",X"AA",X"05",X"A9",X"84",X"8A",X"88",X"58",X"A0",X"A3",X"4C",X"88",X"85",X"8A",
		X"1A",X"86",X"99",X"89",X"50",X"B1",X"0B",X"17",X"A9",X"09",X"32",X"C0",X"90",X"5A",X"A1",X"5B",
		X"90",X"59",X"A8",X"30",X"B9",X"50",X"C0",X"4A",X"94",X"9B",X"23",X"C9",X"23",X"C8",X"92",X"5B",
		X"82",X"B9",X"53",X"D8",X"1A",X"86",X"99",X"18",X"A8",X"33",X"D0",X"0A",X"34",X"D9",X"22",X"C0",
		X"4A",X"A1",X"4B",X"A2",X"4B",X"82",X"C0",X"69",X"A1",X"89",X"24",X"C0",X"0A",X"86",X"8A",X"09",
		X"14",X"B8",X"93",X"3D",X"92",X"3C",X"92",X"3D",X"93",X"2C",X"91",X"4A",X"A8",X"58",X"B8",X"41",
		X"B9",X"85",X"0B",X"88",X"50",X"B8",X"93",X"5C",X"88",X"84",X"0B",X"10",X"C0",X"79",X"91",X"99",
		X"24",X"C0",X"89",X"32",X"D9",X"23",X"BA",X"86",X"8A",X"94",X"1B",X"91",X"5A",X"A8",X"41",X"B9",
		X"85",X"8B",X"86",X"99",X"91",X"59",X"A1",X"99",X"68",X"A1",X"8A",X"85",X"0B",X"11",X"C0",X"6A",
		X"81",X"A9",X"50",X"B0",X"80",X"5A",X"98",X"85",X"8A",X"09",X"40",X"B8",X"05",X"9A",X"84",X"0C",
		X"82",X"2B",X"8A",X"17",X"A8",X"1A",X"93",X"5C",X"80",X"94",X"0C",X"83",X"1B",X"89",X"41",X"BA",
		X"07",X"8B",X"85",X"8A",X"81",X"3B",X"B3",X"5B",X"A3",X"2E",X"04",X"B9",X"48",X"B2",X"3D",X"94",
		X"0B",X"80",X"59",X"90",X"99",X"51",X"B8",X"91",X"59",X"90",X"B2",X"7A",X"91",X"A2",X"3C",X"81",
		X"B1",X"7A",X"98",X"21",X"A0",X"A0",X"79",X"98",X"84",X"8A",X"1A",X"97",X"8A",X"1A",X"14",X"A9",
		X"91",X"6A",X"88",X"95",X"8A",X"09",X"31",X"C0",X"98",X"79",X"98",X"83",X"1B",X"0B",X"36",X"B9",
		X"95",X"0B",X"80",X"59",X"A8",X"23",X"CA",X"50",X"C1",X"3D",X"03",X"BA",X"32",X"C9",X"24",X"B8",
		X"2C",X"06",X"9A",X"19",X"85",X"8A",X"18",X"A0",X"69",X"91",X"9A",X"42",X"D0",X"1A",X"85",X"8B",
		X"19",X"23",X"CA",X"33",X"D9",X"23",X"C9",X"05",X"99",X"89",X"34",X"C8",X"92",X"3B",X"9A",X"27",
		X"A9",X"81",X"5B",X"98",X"58",X"A8",X"85",X"8A",X"92",X"4C",X"01",X"B9",X"60",X"B1",X"1C",X"05",
		X"9A",X"19",X"85",X"8A",X"91",X"4A",X"98",X"58",X"A1",X"9A",X"43",X"D0",X"08",X"99",X"26",X"A9",
		X"19",X"94",X"2D",X"88",X"30",X"B9",X"68",X"B0",X"5A",X"98",X"31",X"B9",X"86",X"8A",X"91",X"5A",
		X"A2",X"3C",X"98",X"33",X"C8",X"1B",X"97",X"1C",X"01",X"9A",X"16",X"A9",X"1A",X"32",X"C8",X"82",
		X"3B",X"B8",X"70",X"B9",X"50",X"C0",X"4A",X"A1",X"4A",X"98",X"31",X"C9",X"14",X"AA",X"06",X"AA",
		X"32",X"D8",X"30",X"C8",X"48",X"A8",X"05",X"9A",X"83",X"1D",X"03",X"B8",X"4C",X"13",X"C9",X"40",
		X"B9",X"40",X"A9",X"15",X"A9",X"88",X"69",X"A8",X"40",X"B8",X"84",X"0A",X"0A",X"07",X"99",X"0A",
		X"16",X"A9",X"19",X"93",X"4C",X"81",X"A0",X"5A",X"90",X"93",X"3E",X"01",X"99",X"93",X"6B",X"81",
		X"8B",X"17",X"9A",X"19",X"04",X"9A",X"09",X"33",X"D0",X"1C",X"07",X"9A",X"28",X"A1",X"4B",X"88",
		X"84",X"8B",X"05",X"9A",X"82",X"3C",X"A2",X"5B",X"98",X"40",X"A9",X"05",X"9A",X"95",X"0C",X"13",
		X"B9",X"88",X"78",X"A1",X"99",X"40",X"B9",X"15",X"9B",X"24",X"D8",X"4A",X"93",X"8B",X"14",X"B9",
		X"84",X"1C",X"10",X"B1",X"7A",X"80",X"0A",X"84",X"1C",X"10",X"A9",X"34",X"C0",X"89",X"41",X"C0",
		X"0A",X"41",X"C0",X"90",X"59",X"90",X"A2",X"4B",X"98",X"24",X"C9",X"40",X"D0",X"4A",X"80",X"A2",
		X"4B",X"82",X"BA",X"44",X"C8",X"29",X"A3",X"4D",X"08",X"94",X"0B",X"82",X"2B",X"A1",X"7A",X"98",
		X"23",X"C8",X"93",X"4C",X"89",X"06",X"99",X"89",X"58",X"A8",X"84",X"1C",X"00",X"A3",X"2D",X"00",
		X"A0",X"79",X"91",X"89",X"89",X"51",X"C1",X"0B",X"24",X"B9",X"83",X"1D",X"85",X"8B",X"04",X"9A",
		X"85",X"8A",X"88",X"59",X"98",X"03",X"9A",X"92",X"5B",X"8A",X"43",X"D9",X"15",X"B9",X"14",X"AB",
		X"15",X"A9",X"93",X"3C",X"98",X"58",X"A9",X"05",X"99",X"92",X"3C",X"A5",X"1C",X"83",X"0C",X"80",
		X"5A",X"89",X"14",X"A8",X"8A",X"27",X"B8",X"1A",X"06",X"A9",X"08",X"21",X"BA",X"34",X"B8",X"A0",
		X"78",X"A2",X"9B",X"36",X"B9",X"2A",X"95",X"1C",X"01",X"99",X"92",X"7A",X"81",X"8A",X"84",X"1C",
		X"18",X"A3",X"3D",X"90",X"49",X"A8",X"58",X"A9",X"40",X"AA",X"33",X"CA",X"42",X"D9",X"14",X"9A",
		X"09",X"41",X"C8",X"84",X"8A",X"96",X"8B",X"04",X"9A",X"82",X"3B",X"9A",X"44",X"C8",X"94",X"0A",
		X"A0",X"79",X"91",X"99",X"40",X"B8",X"84",X"0A",X"98",X"79",X"99",X"23",X"B9",X"94",X"1C",X"95",
		X"0B",X"09",X"07",X"A8",X"1A",X"85",X"8B",X"08",X"48",X"A8",X"85",X"8A",X"89",X"68",X"A8",X"04",
		X"9B",X"15",X"AA",X"04",X"8A",X"90",X"69",X"91",X"A8",X"69",X"A1",X"89",X"23",X"C0",X"0B",X"86",
		X"1C",X"18",X"A2",X"5C",X"08",X"84",X"9A",X"1A",X"33",X"CA",X"15",X"A9",X"93",X"3C",X"8A",X"42",
		X"C9",X"05",X"8A",X"89",X"33",X"C8",X"0B",X"07",X"8A",X"28",X"C2",X"5C",X"08",X"93",X"2C",X"88",
		X"30",X"C8",X"58",X"A9",X"24",X"B8",X"90",X"69",X"A0",X"93",X"2C",X"00",X"B2",X"7B",X"08",X"A5",
		X"1C",X"18",X"A4",X"0B",X"19",X"85",X"99",X"89",X"41",X"B0",X"8B",X"71",X"B0",X"8A",X"51",X"C0",
		X"91",X"4A",X"A0",X"49",X"99",X"24",X"B9",X"94",X"2C",X"90",X"6A",X"98",X"14",X"A9",X"92",X"5B",
		X"88",X"96",X"8B",X"82",X"3C",X"A3",X"3C",X"A3",X"3C",X"B4",X"3E",X"03",X"B9",X"31",X"C9",X"04",
		X"1C",X"09",X"24",X"C8",X"2B",X"06",X"A9",X"08",X"30",X"B1",X"9A",X"70",X"B1",X"A1",X"5B",X"90",
		X"48",X"A1",X"B8",X"70",X"B1",X"0B",X"06",X"99",X"92",X"3C",X"90",X"59",X"A8",X"31",X"BA",X"07",
		X"99",X"1B",X"26",X"B8",X"09",X"48",X"B8",X"32",X"CA",X"34",X"C9",X"23",X"CA",X"33",X"D9",X"32",
		X"D9",X"32",X"C0",X"A2",X"5B",X"89",X"24",X"BA",X"86",X"0B",X"09",X"33",X"D8",X"93",X"3D",X"89",
		X"33",X"D8",X"93",X"3D",X"88",X"05",X"9A",X"0A",X"43",X"D0",X"1A",X"A3",X"6B",X"81",X"A9",X"68",
		X"A0",X"91",X"4A",X"98",X"14",X"A9",X"93",X"4D",X"00",X"A3",X"3E",X"09",X"85",X"8A",X"18",X"A1",
		X"6A",X"92",X"B0",X"69",X"A0",X"83",X"0C",X"81",X"4A",X"A0",X"59",X"A8",X"48",X"A9",X"06",X"8B",
		X"82",X"3C",X"A4",X"1C",X"84",X"8A",X"88",X"31",X"C0",X"A2",X"7A",X"98",X"22",X"B8",X"A8",X"70",
		X"B2",X"A9",X"60",X"B0",X"90",X"5A",X"90",X"94",X"1B",X"08",X"B4",X"5C",X"01",X"9A",X"24",X"C8",
		X"1A",X"33",X"D9",X"03",X"8B",X"85",X"0B",X"91",X"7A",X"92",X"8B",X"17",X"A9",X"2A",X"94",X"1B",
		X"09",X"96",X"0B",X"1A",X"15",X"A9",X"09",X"33",X"E0",X"89",X"58",X"A8",X"84",X"8A",X"88",X"58",
		X"A1",X"8B",X"43",X"D8",X"88",X"58",X"A8",X"84",X"8A",X"91",X"5A",X"A0",X"59",X"A8",X"23",X"C9",
		X"85",X"0B",X"93",X"3C",X"A3",X"3E",X"95",X"9A",X"04",X"9A",X"82",X"3B",X"81",X"D2",X"5B",X"88",
		X"95",X"0B",X"09",X"15",X"A9",X"93",X"2B",X"A8",X"78",X"A1",X"A8",X"79",X"A0",X"49",X"A0",X"49",
		X"B2",X"3C",X"A3",X"3E",X"84",X"A9",X"30",X"C1",X"3B",X"99",X"35",X"B8",X"98",X"78",X"A0",X"91",
		X"4A",X"90",X"A5",X"1C",X"88",X"40",X"B0",X"91",X"6A",X"91",X"A9",X"51",X"B0",X"1C",X"86",X"8A",
		X"10",X"B8",X"60",X"B1",X"8A",X"25",X"B8",X"1A",X"94",X"2C",X"88",X"22",X"C9",X"50",X"B9",X"58",
		X"A8",X"30",X"D0",X"49",X"B2",X"3B",X"B2",X"6A",X"90",X"93",X"2C",X"88",X"94",X"4C",X"81",X"B1",
		X"7A",X"90",X"83",X"8B",X"82",X"4B",X"B1",X"79",X"A8",X"31",X"B0",X"0C",X"17",X"A9",X"1A",X"15",
		X"A9",X"81",X"3B",X"99",X"51",X"BA",X"42",X"CA",X"26",X"A9",X"1A",X"86",X"8A",X"09",X"22",X"B8",
		X"A2",X"7A",X"98",X"85",X"0B",X"10",X"AA",X"27",X"A8",X"18",X"9A",X"17",X"A8",X"09",X"13",X"BA",
		X"07",X"99",X"92",X"3B",X"B2",X"5A",X"A8",X"68",X"A8",X"85",X"8A",X"88",X"22",X"D9",X"50",X"B8",
		X"13",X"B9",X"96",X"0B",X"94",X"0C",X"13",X"C8",X"49",X"B2",X"4C",X"88",X"30",X"A9",X"05",X"99",
		X"98",X"79",X"90",X"93",X"2D",X"09",X"14",X"B9",X"23",X"C8",X"A1",X"7A",X"88",X"84",X"8A",X"1A",
		X"87",X"99",X"08",X"93",X"1C",X"09",X"24",X"B8",X"98",X"79",X"99",X"32",X"C9",X"14",X"A9",X"90",
		X"69",X"90",X"A3",X"3D",X"09",X"85",X"1C",X"01",X"A9",X"41",X"C0",X"1A",X"94",X"2C",X"01",X"C0",
		X"58",X"B2",X"A8",X"58",X"B1",X"91",X"5B",X"88",X"84",X"0B",X"89",X"60",X"B1",X"99",X"78",X"A1",
		X"99",X"33",X"E0",X"89",X"32",X"C8",X"84",X"8A",X"91",X"6A",X"90",X"94",X"0B",X"09",X"06",X"9A",
		X"83",X"1B",X"8A",X"43",X"D9",X"86",X"8A",X"09",X"23",X"C8",X"93",X"3D",X"89",X"41",X"BA",X"16",
		X"A9",X"80",X"59",X"A8",X"05",X"9A",X"95",X"0B",X"94",X"1B",X"90",X"59",X"98",X"93",X"4C",X"01",
		X"B9",X"36",X"C0",X"1A",X"95",X"0B",X"88",X"40",X"B8",X"05",X"99",X"90",X"6A",X"80",X"A3",X"3E",
		X"80",X"39",X"B1",X"5A",X"A0",X"59",X"98",X"93",X"3E",X"00",X"A2",X"5B",X"92",X"A9",X"50",X"B0",
		X"90",X"79",X"91",X"99",X"40",X"C1",X"98",X"58",X"A8",X"82",X"3C",X"A1",X"6A",X"89",X"04",X"9A",
		X"84",X"0B",X"93",X"3D",X"92",X"3C",X"A3",X"3D",X"91",X"4A",X"B4",X"2D",X"83",X"0B",X"94",X"0B",
		X"96",X"0B",X"91",X"5A",X"98",X"05",X"99",X"89",X"40",X"A8",X"92",X"6B",X"81",X"B0",X"79",X"A1",
		X"91",X"3B",X"B3",X"5B",X"A0",X"69",X"A0",X"49",X"A8",X"31",X"C9",X"15",X"A8",X"90",X"6A",X"89",
		X"14",X"A9",X"0A",X"25",X"B8",X"1C",X"16",X"A8",X"1A",X"92",X"5C",X"01",X"B0",X"69",X"A1",X"90",
		X"49",X"A1",X"A0",X"69",X"91",X"8A",X"06",X"A9",X"08",X"40",X"B0",X"8A",X"60",X"B8",X"30",X"C8",
		X"58",X"B0",X"49",X"B0",X"58",X"A9",X"14",X"A9",X"82",X"2B",X"8B",X"37",X"A9",X"1B",X"43",X"D9",
		X"13",X"AC",X"33",X"D9",X"15",X"A9",X"09",X"32",X"D8",X"84",X"8A",X"09",X"33",X"DA",X"16",X"A8",
		X"90",X"5A",X"98",X"04",X"99",X"0A",X"07",X"99",X"1A",X"85",X"0C",X"10",X"A0",X"59",X"A1",X"0A",
		X"92",X"59",X"91",X"89",X"8A",X"07",X"8A",X"29",X"B3",X"7B",X"81",X"B3",X"3D",X"91",X"4A",X"A0",
		X"59",X"99",X"32",X"C9",X"15",X"B8",X"88",X"58",X"A9",X"05",X"99",X"0A",X"17",X"A8",X"0A",X"15",
		X"B8",X"1B",X"16",X"A9",X"09",X"40",X"A9",X"05",X"9A",X"83",X"1C",X"95",X"8B",X"14",X"BA",X"41",
		X"D1",X"2A",X"A2",X"4C",X"88",X"30",X"A9",X"15",X"AB",X"33",X"D9",X"32",X"D8",X"83",X"1B",X"0A",
		X"87",X"8A",X"1A",X"25",X"B9",X"2B",X"87",X"99",X"09",X"30",X"C8",X"58",X"B8",X"58",X"A0",X"93",
		X"1B",X"A2",X"6A",X"99",X"24",X"B8",X"A1",X"7A",X"98",X"15",X"B8",X"09",X"32",X"D0",X"98",X"58",
		X"A1",X"9A",X"60",X"B1",X"A0",X"79",X"91",X"8A",X"85",X"8A",X"18",X"A3",X"3D",X"89",X"40",X"A9",
		X"06",X"9A",X"04",X"9B",X"14",X"AA",X"14",X"AA",X"85",X"0B",X"0A",X"35",X"C8",X"80",X"5A",X"91",
		X"A1",X"6B",X"01",X"B0",X"6A",X"80",X"A2",X"4B",X"90",X"95",X"8A",X"88",X"32",X"C0",X"9A",X"70",
		X"B1",X"0B",X"17",X"A9",X"2A",X"85",X"9A",X"18",X"93",X"3D",X"08",X"A4",X"2C",X"09",X"86",X"9A",
		X"03",X"8B",X"85",X"8B",X"86",X"99",X"83",X"8B",X"09",X"34",X"C8",X"91",X"59",X"A9",X"25",X"B8",
		X"91",X"6A",X"98",X"86",X"99",X"00",X"B1",X"59",X"A1",X"A0",X"79",X"91",X"99",X"24",X"C8",X"2B",
		X"86",X"99",X"88",X"30",X"A8",X"94",X"1B",X"98",X"79",X"A1",X"4A",X"B2",X"4B",X"A3",X"2C",X"91",
		X"5B",X"95",X"8C",X"22",X"C8",X"38",X"B8",X"58",X"A8",X"86",X"99",X"80",X"3A",X"A3",X"3D",X"A2",
		X"4A",X"A8",X"50",X"B9",X"16",X"A9",X"88",X"58",X"A1",X"A8",X"68",X"A0",X"93",X"1C",X"0A",X"17",
		X"A8",X"09",X"04",X"A9",X"93",X"2B",X"8B",X"45",X"C0",X"89",X"25",X"C8",X"18",X"A0",X"69",X"91",
		X"A0",X"49",X"98",X"92",X"5B",X"80",X"A3",X"4D",X"00",X"A1",X"5A",X"90",X"93",X"2C",X"89",X"32",
		X"C9",X"87",X"8A",X"94",X"0A",X"89",X"33",X"C8",X"99",X"78",X"A8",X"30",X"D0",X"49",X"B0",X"59",
		X"A8",X"40",X"A8",X"93",X"3D",X"09",X"86",X"99",X"18",X"B2",X"5A",X"90",X"A4",X"1B",X"98",X"68",
		X"A9",X"33",X"D9",X"05",X"99",X"0A",X"24",X"B8",X"1C",X"25",X"B8",X"89",X"50",X"B8",X"22",X"C9",
		X"32",X"D9",X"58",X"A9",X"24",X"B9",X"83",X"2C",X"89",X"16",X"A8",X"1B",X"87",X"99",X"19",X"85",
		X"9A",X"81",X"3B",X"A2",X"5B",X"A2",X"5B",X"98",X"31",X"C9",X"17",X"A9",X"00",X"3A",X"B2",X"5B",
		X"98",X"58",X"A8",X"85",X"8B",X"82",X"3B",X"99",X"87",X"8A",X"28",X"9B",X"07",X"0B",X"11",X"9A",
		X"94",X"4C",X"81",X"A0",X"69",X"A0",X"94",X"0A",X"0A",X"16",X"A9",X"80",X"5A",X"98",X"85",X"8A",
		X"09",X"24",X"BA",X"85",X"1C",X"09",X"05",X"9A",X"83",X"0B",X"A3",X"5B",X"A0",X"79",X"98",X"04",
		X"AA",X"04",X"8B",X"09",X"41",X"B9",X"07",X"A8",X"89",X"50",X"B1",X"98",X"5A",X"98",X"40",X"B9",
		X"06",X"99",X"0A",X"25",X"B8",X"0A",X"35",X"C8",X"09",X"31",X"B9",X"93",X"5B",X"8A",X"34",X"C8",
		X"A4",X"3D",X"08",X"95",X"8A",X"88",X"48",X"A1",X"B0",X"78",X"A1",X"9A",X"52",X"C8",X"09",X"22",
		X"C0",X"98",X"68",X"A1",X"A1",X"4B",X"91",X"4B",X"A4",X"2D",X"82",X"1B",X"89",X"51",X"B8",X"95",
		X"0B",X"93",X"3D",X"90",X"48",X"AA",X"25",X"B8",X"92",X"5B",X"89",X"87",X"9A",X"02",X"1C",X"85",
		X"9A",X"83",X"1C",X"09",X"32",X"D8",X"83",X"1C",X"84",X"8B",X"86",X"8A",X"91",X"5A",X"90",X"92",
		X"3C",X"80",X"B4",X"4C",X"01",X"B9",X"60",X"B1",X"8A",X"42",X"D8",X"02",X"0A",X"89",X"42",X"C0",
		X"A2",X"5B",X"81",X"B8",X"78",X"A1",X"A0",X"59",X"A0",X"82",X"2C",X"09",X"87",X"99",X"1A",X"86",
		X"8A",X"01",X"B0",X"69",X"A1",X"90",X"4A",X"98",X"31",X"BA",X"17",X"AA",X"23",X"C9",X"23",X"C8",
		X"91",X"5A",X"A1",X"5B",X"98",X"41",X"C0",X"93",X"1B",X"90",X"79",X"90",X"A2",X"5C",X"82",X"9A",
		X"25",X"B8",X"1A",X"95",X"1C",X"08",X"84",X"8A",X"1A",X"86",X"8B",X"08",X"59",X"99",X"14",X"AA",
		X"15",X"AA",X"05",X"A9",X"83",X"1C",X"88",X"58",X"A9",X"32",X"C9",X"86",X"8A",X"1A",X"87",X"99",
		X"09",X"22",X"C0",X"1B",X"06",X"99",X"19",X"A4",X"1C",X"08",X"38",X"B9",X"35",X"BA",X"06",X"8A",
		X"89",X"50",X"AA",X"15",X"A9",X"88",X"68",X"A8",X"83",X"1C",X"88",X"58",X"A9",X"32",X"C8",X"A5",
		X"1B",X"90",X"40",X"B8",X"A4",X"3C",X"89",X"17",X"A8",X"90",X"59",X"A1",X"A2",X"4C",X"88",X"85",
		X"8A",X"09",X"23",X"D0",X"98",X"79",X"90",X"90",X"4A",X"89",X"13",X"9A",X"A1",X"79",X"90",X"A3",
		X"5C",X"82",X"B8",X"79",X"90",X"90",X"38",X"B2",X"9B",X"61",X"B9",X"14",X"AB",X"17",X"A9",X"03",
		X"9A",X"93",X"3C",X"0A",X"87",X"8A",X"10",X"C1",X"6A",X"91",X"99",X"41",X"B0",X"8A",X"51",X"B8",
		X"94",X"1B",X"90",X"69",X"A1",X"A2",X"5B",X"89",X"85",X"0B",X"09",X"40",X"B0",X"B2",X"7A",X"90",
		X"95",X"0B",X"92",X"4B",X"A0",X"69",X"A8",X"58",X"A8",X"83",X"1C",X"88",X"58",X"A8",X"94",X"1B",
		X"89",X"50",X"B9",X"42",X"D9",X"23",X"B9",X"92",X"6B",X"88",X"06",X"A9",X"1A",X"06",X"9A",X"1A",
		X"23",X"C9",X"32",X"D9",X"40",X"C1",X"3B",X"A5",X"8B",X"05",X"A8",X"88",X"49",X"98",X"84",X"0B",
		X"0A",X"35",X"B8",X"1C",X"06",X"99",X"89",X"40",X"A9",X"15",X"B9",X"84",X"1C",X"92",X"3B",X"A0",
		X"79",X"A8",X"31",X"C8",X"04",X"9A",X"93",X"4B",X"A8",X"68",X"A9",X"58",X"B0",X"48",X"B9",X"50",
		X"A9",X"85",X"89",X"0A",X"86",X"0B",X"01",X"98",X"A0",X"52",X"D0",X"19",X"A1",X"59",X"A1",X"A1",
		X"6A",X"91",X"A2",X"5C",X"81",X"A3",X"2D",X"88",X"48",X"A8",X"05",X"A8",X"89",X"41",X"C0",X"1B",
		X"87",X"8A",X"19",X"95",X"8A",X"09",X"22",X"BA",X"26",X"B9",X"23",X"D9",X"23",X"C8",X"82",X"2C",
		X"A5",X"1B",X"A4",X"1C",X"85",X"9A",X"13",X"D8",X"49",X"A1",X"3B",X"A1",X"5A",X"A0",X"59",X"98",
		X"84",X"8A",X"88",X"58",X"A9",X"24",X"BA",X"06",X"99",X"91",X"4A",X"91",X"B1",X"7A",X"92",X"89",
		X"A3",X"5C",X"81",X"A0",X"6A",X"80",X"98",X"58",X"A8",X"83",X"1C",X"09",X"33",X"E0",X"89",X"33",
		X"D0",X"0A",X"87",X"99",X"18",X"A8",X"68",X"A1",X"0B",X"87",X"99",X"08",X"11",X"B8",X"58",X"B0",
		X"49",X"B2",X"4C",X"93",X"0C",X"13",X"C0",X"3C",X"03",X"C0",X"4B",X"93",X"1C",X"84",X"9A",X"05",
		X"A9",X"85",X"99",X"80",X"3A",X"98",X"85",X"1C",X"00",X"A4",X"2E",X"08",X"03",X"A9",X"0A",X"42",
		X"C8",X"80",X"6A",X"89",X"04",X"9A",X"83",X"2D",X"92",X"4B",X"99",X"34",X"B8",X"A8",X"78",X"A1",
		X"8B",X"43",X"E0",X"80",X"3A",X"98",X"86",X"8A",X"1A",X"87",X"99",X"1A",X"86",X"99",X"00",X"A1",
		X"4A",X"91",X"8A",X"87",X"8A",X"1A",X"23",X"BB",X"27",X"B8",X"83",X"0B",X"91",X"6A",X"A0",X"59",
		X"90",X"A2",X"5B",X"88",X"94",X"1C",X"08",X"96",X"8A",X"09",X"05",X"A8",X"90",X"6A",X"92",X"A9",
		X"50",X"B0",X"80",X"49",X"A8",X"05",X"9A",X"80",X"6A",X"89",X"85",X"0B",X"01",X"B0",X"79",X"90",
		X"91",X"3B",X"89",X"06",X"A8",X"90",X"69",X"A1",X"A0",X"69",X"A2",X"A8",X"59",X"90",X"A4",X"1B",
		X"89",X"33",X"D9",X"58",X"B1",X"4B",X"A2",X"4C",X"80",X"4A",X"90",X"95",X"0B",X"88",X"40",X"B9",
		X"25",X"B9",X"87",X"99",X"88",X"31",X"C0",X"0A",X"25",X"C0",X"90",X"49",X"A8",X"31",X"C8",X"86",
		X"99",X"91",X"4A",X"90",X"95",X"8A",X"10",X"C8",X"78",X"A1",X"0A",X"93",X"4C",X"81",X"8A",X"16",
		X"A9",X"09",X"31",X"B0",X"99",X"62",X"D0",X"1B",X"06",X"9A",X"19",X"13",X"C0",X"91",X"4B",X"90",
		X"6A",X"89",X"23",X"D8",X"83",X"0B",X"90",X"68",X"A8",X"95",X"1C",X"09",X"23",X"D0",X"91",X"4B",
		X"88",X"95",X"0B",X"1A",X"87",X"8A",X"1A",X"86",X"8A",X"01",X"9A",X"07",X"99",X"09",X"04",X"99",
		X"88",X"31",X"C0",X"A4",X"2C",X"09",X"86",X"8A",X"00",X"A8",X"68",X"A0",X"91",X"4A",X"99",X"16",
		X"B8",X"09",X"58",X"B0",X"04",X"9B",X"06",X"9B",X"23",X"C9",X"31",X"D8",X"38",X"B1",X"5B",X"93",
		X"2E",X"03",X"B9",X"40",X"C1",X"3B",X"A1",X"6A",X"88",X"84",X"99",X"88",X"40",X"B9",X"24",X"B8",
		X"99",X"60",X"B8",X"93",X"6C",X"88",X"13",X"BA",X"25",X"B9",X"85",X"8A",X"88",X"59",X"A8",X"58",
		X"B8",X"32",X"D8",X"49",X"B2",X"4B",X"A5",X"8B",X"14",X"C8",X"49",X"A0",X"49",X"A8",X"23",X"C8",
		X"09",X"58",X"A0",X"98",X"68",X"A8",X"04",X"A9",X"28",X"C1",X"6A",X"92",X"A9",X"41",X"C0",X"0A",
		X"41",X"B0",X"90",X"6A",X"80",X"A4",X"0B",X"09",X"58",X"A9",X"24",X"B8",X"0B",X"44",X"D0",X"0A",
		X"32",X"D0",X"91",X"4B",X"98",X"58",X"A8",X"48",X"B0",X"5A",X"98",X"14",X"B9",X"84",X"0B",X"89",
		X"60",X"B8",X"32",X"D8",X"83",X"1C",X"09",X"86",X"0B",X"01",X"B8",X"79",X"91",X"99",X"34",X"D0",
		X"19",X"A1",X"6A",X"92",X"A9",X"41",X"B8",X"88",X"68",X"A0",X"91",X"5B",X"08",X"A3",X"4D",X"09",
		X"13",X"BA",X"41",X"D0",X"4A",X"93",X"AA",X"58",X"B1",X"4B",X"A1",X"6A",X"89",X"31",X"C8",X"48",
		X"B0",X"5A",X"A2",X"3C",X"94",X"8B",X"01",X"4B",X"82",X"B9",X"70",X"B1",X"A0",X"69",X"A2",X"99",
		X"32",X"D8",X"2A",X"A5",X"2C",X"82",X"A9",X"41",X"C0",X"92",X"3C",X"91",X"5B",X"89",X"40",X"B8",
		X"03",X"0D",X"84",X"0B",X"0A",X"27",X"A9",X"1A",X"48",X"A8",X"84",X"0C",X"09",X"58",X"A1",X"0B",
		X"26",X"B8",X"1B",X"17",X"A9",X"2B",X"06",X"9A",X"19",X"13",X"B8",X"92",X"4B",X"B4",X"2D",X"83",
		X"1C",X"80",X"38",X"C0",X"14",X"BB",X"17",X"A8",X"92",X"3C",X"81",X"B3",X"4C",X"80",X"A3",X"3D",
		X"01",X"A9",X"52",X"D8",X"2A",X"94",X"2D",X"00",X"92",X"1C",X"04",X"A9",X"83",X"1D",X"08",X"31",
		X"C0",X"1B",X"06",X"8B",X"20",X"A8",X"90",X"79",X"92",X"9A",X"94",X"3E",X"18",X"94",X"9A",X"03",
		X"8B",X"84",X"1D",X"80",X"38",X"B2",X"B0",X"7A",X"93",X"B0",X"58",X"B0",X"94",X"0A",X"98",X"34",
		X"C0",X"A2",X"5C",X"80",X"85",X"A9",X"83",X"1B",X"0B",X"17",X"9A",X"19",X"31",X"E8",X"48",X"B0",
		X"49",X"A0",X"4A",X"A0",X"59",X"A8",X"05",X"A9",X"01",X"3B",X"B6",X"8B",X"23",X"E8",X"30",X"C0",
		X"03",X"A9",X"91",X"6A",X"81",X"8B",X"35",X"D1",X"89",X"22",X"D0",X"1A",X"14",X"AA",X"83",X"2C",
		X"10",X"B2",X"7B",X"80",X"95",X"9A",X"04",X"9A",X"81",X"3B",X"08",X"A6",X"0C",X"10",X"B4",X"2E",
		X"10",X"A2",X"3C",X"92",X"A0",X"59",X"A1",X"93",X"1D",X"19",X"05",X"AA",X"2A",X"25",X"BA",X"3B",
		X"26",X"B9",X"1A",X"50",X"B1",X"A5",X"8B",X"01",X"3B",X"B2",X"5B",X"B1",X"69",X"A8",X"22",X"BA",
		X"42",X"F1",X"2B",X"93",X"1C",X"96",X"8B",X"03",X"9A",X"03",X"2B",X"81",X"9A",X"41",X"E1",X"19",
		X"91",X"4A",X"B3",X"1E",X"23",X"D0",X"00",X"3B",X"A1",X"95",X"0C",X"19",X"21",X"B9",X"15",X"BB",
		X"15",X"0D",X"19",X"21",X"C8",X"31",X"C8",X"31",X"D1",X"94",X"8C",X"10",X"03",X"AB",X"10",X"84",
		X"BA",X"2A",X"32",X"E1",X"09",X"3A",X"C1",X"59",X"B3",X"2B",X"A0",X"23",X"B8",X"0A",X"69",X"B2",
		X"1B",X"23",X"BB",X"3A",X"32",X"BA",X"23",X"BA",X"05",X"9B",X"23",X"BB",X"33",X"BA",X"20",X"3E",
		X"10",X"8A",X"23",X"BA",X"39",X"A2",X"4E",X"10",X"80",X"2B",X"91",X"0A",X"23",X"E1",X"19",X"91",
		X"3E",X"11",X"A1",X"3D",X"18",X"03",X"BA",X"10",X"10",X"A0",X"08",X"84",X"AC",X"21",X"90",X"10",
		X"D2",X"00",X"09",X"00",X"1A",X"08",X"4B",X"A3",X"9B",X"33",X"BB",X"30",X"1A",X"08",X"10",X"B1",
		X"03",X"B8",X"03",X"BA",X"20",X"1A",X"92",X"1A",X"00",X"1D",X"20",X"83",X"BA",X"21",X"90",X"3B",
		X"80",X"81",X"0B",X"10",X"84",X"B8",X"80",X"3B",X"80",X"00",X"90",X"82",X"89",X"80",X"84",X"B8",
		X"19",X"03",X"BB",X"38",X"03",X"BB",X"31",X"89",X"08",X"29",X"A1",X"03",X"B8",X"03",X"BA",X"32",
		X"B8",X"00",X"1C",X"10",X"12",X"D1",X"80",X"3B",X"A2",X"18",X"90",X"81",X"2D",X"10",X"80",X"10",
		X"E2",X"08",X"81",X"0C",X"20",X"88",X"29",X"B2",X"99",X"00",X"09",X"81",X"00",X"80",X"80",X"80",
		X"80",X"88",X"91",X"92",X"80",X"80",X"88",X"92",X"80",X"80",X"88",X"09",X"80",X"82",X"89",X"80",
		X"82",X"89",X"80",X"82",X"89",X"10",X"80",X"91",X"80",X"80",X"91",X"08",X"A2",X"00",X"99",X"80",
		X"10",X"08",X"80",X"08",X"80",X"80",X"80",X"89",X"88",X"81",X"01",X"80",X"A0",X"90",X"00",X"80",
		X"01",X"B1",X"80",X"A0",X"12",X"89",X"81",X"00",X"80",X"80",X"80",X"A9",X"01",X"01",X"81",X"90",
		X"81",X"08",X"90",X"88",X"81",X"10",X"91",X"98",X"80",X"00",X"88",X"A2",X"89",X"80",X"08",X"80",
		X"10",X"80",X"B0",X"00",X"81",X"90",X"A0",X"82",X"10",X"81",X"98",X"92",X"19",X"80",X"80",X"A8",
		X"11",X"99",X"81",X"19",X"98",X"03",X"A8",X"83",X"88",X"98",X"02",X"89",X"11",X"90",X"81",X"88",
		X"00",X"88",X"80",X"81",X"98",X"01",X"08",X"B2",X"18",X"98",X"00",X"80",X"80",X"08",X"A0",X"08",
		X"88",X"02",X"0A",X"91",X"19",X"89",X"01",X"88",X"83",X"08",X"A0",X"20",X"B9",X"02",X"09",X"90",
		X"00",X"A0",X"82",X"00",X"92",X"81",X"81",X"89",X"81",X"81",X"A0",X"A2",X"01",X"A0",X"82",X"89",
		X"83",X"99",X"91",X"01",X"A0",X"91",X"98",X"82",X"00",X"B9",X"12",X"80",X"80",X"A8",X"90",X"80",
		X"80",X"80",X"01",X"90",X"20",X"A1",X"00",X"80",X"91",X"88",X"00",X"80",X"91",X"81",X"09",X"98",
		X"18",X"08",X"00",X"80",X"98",X"12",X"88",X"91",X"88",X"80",X"80",X"80",X"89",X"11",X"90",X"80",
		X"89",X"11",X"90",X"80",X"A0",X"91",X"08",X"88",X"81",X"80",X"90",X"02",X"08",X"89",X"01",X"A0",
		X"00",X"18",X"9A",X"21",X"0C",X"08",X"20",X"88",X"28",X"08",X"98",X"01",X"19",X"08",X"18",X"88",
		X"19",X"08",X"08",X"10",X"89",X"80",X"19",X"08",X"18",X"89",X"18",X"08",X"08",X"08",X"08",X"98",
		X"20",X"88",X"08",X"99",X"11",X"0A",X"88",X"11",X"08",X"98",X"28",X"08",X"08",X"0A",X"08",X"28",
		X"99",X"80",X"20",X"A8",X"02",X"18",X"88",X"08",X"0A",X"81",X"18",X"0B",X"11",X"19",X"90",X"18",
		X"0A",X"01",X"08",X"9A",X"21",X"08",X"98",X"2A",X"08",X"20",X"18",X"98",X"08",X"98",X"01",X"08",
		X"08",X"08",X"08",X"98",X"10",X"0A",X"29",X"88",X"01",X"08",X"08",X"00",X"88",X"80",X"28",X"88",
		X"80",X"1A",X"08",X"08",X"08",X"21",X"8B",X"91",X"08",X"89",X"08",X"29",X"80",X"18",X"8A",X"01",
		X"18",X"08",X"0A",X"08",X"09",X"19",X"88",X"08",X"10",X"88",X"09",X"18",X"18",X"08",X"08",X"09",
		X"08",X"18",X"08",X"80",X"10",X"91",X"09",X"88",X"28",X"08",X"09",X"00",X"18",X"09",X"08",X"00",
		X"00",X"09",X"18",X"09",X"88",X"18",X"19",X"88",X"08",X"0A",X"80",X"20",X"09",X"19",X"08",X"00",
		X"09",X"0A",X"08",X"10",X"98",X"08",X"08",X"01",X"0A",X"08",X"08",X"08",X"01",X"08",X"08",X"0A",
		X"89",X"19",X"18",X"18",X"08",X"28",X"18",X"09",X"08",X"08",X"09",X"88",X"28",X"08",X"08",X"08",
		X"18",X"08",X"81",X"09",X"09",X"08",X"00",X"8A",X"92",X"20",X"9A",X"88",X"10",X"89",X"11",X"19",
		X"98",X"20",X"88",X"98",X"28",X"0A",X"80",X"28",X"89",X"01",X"0A",X"88",X"08",X"10",X"89",X"10",
		X"1A",X"80",X"28",X"08",X"98",X"01",X"89",X"00",X"18",X"90",X"18",X"09",X"88",X"20",X"8A",X"01",
		X"19",X"88",X"11",X"1A",X"98",X"10",X"8A",X"01",X"08",X"0A",X"28",X"08",X"08",X"08",X"98",X"00",
		X"19",X"18",X"08",X"0A",X"08",X"80",X"28",X"0A",X"2A",X"28",X"08",X"08",X"18",X"88",X"00",X"09",
		X"10",X"88",X"00",X"08",X"09",X"09",X"08",X"08",X"08",X"0A",X"01",X"0A",X"08",X"2A",X"88",X"80",
		X"11",X"08",X"80",X"9A",X"BB",X"09",X"01",X"64",X"18",X"99",X"9A",X"88",X"08",X"08",X"A8",X"43",
		X"20",X"BA",X"CE",X"13",X"71",X"08",X"8A",X"A0",X"81",X"00",X"9A",X"08",X"89",X"AB",X"67",X"01",
		X"89",X"8C",X"98",X"01",X"10",X"9F",X"BA",X"27",X"13",X"0A",X"9B",X"B0",X"85",X"19",X"9F",X"A0",
		X"34",X"41",X"8A",X"BC",X"80",X"41",X"9B",X"CA",X"33",X"72",X"18",X"BC",X"90",X"19",X"A8",X"86",
		X"01",X"40",X"1B",X"B8",X"9B",X"F9",X"23",X"22",X"31",X"8A",X"B9",X"BF",X"F0",X"31",X"22",X"98",
		X"89",X"09",X"FD",X"84",X"11",X"2A",X"89",X"83",X"BF",X"B1",X"70",X"18",X"B8",X"94",X"2C",X"C8",
		X"52",X"00",X"DA",X"03",X"4B",X"C8",X"33",X"29",X"EA",X"04",X"2D",X"A2",X"13",X"1C",X"B8",X"25",
		X"AB",X"95",X"21",X"AD",X"81",X"48",X"D9",X"32",X"18",X"D9",X"05",X"0C",X"92",X"21",X"8D",X"91",
		X"48",X"B9",X"33",X"09",X"E8",X"14",X"AB",X"85",X"28",X"AC",X"03",X"2C",X"A8",X"62",X"AA",X"A2",
		X"30",X"E8",X"05",X"0A",X"A8",X"40",X"B9",X"05",X"2B",X"9A",X"26",X"BB",X"28",X"70",X"B8",X"03",
		X"8E",X"01",X"12",X"D8",X"82",X"4E",X"82",X"85",X"AB",X"11",X"3D",X"A2",X"13",X"9E",X"18",X"38",
		X"F1",X"20",X"2D",X"80",X"31",X"F0",X"28",X"5B",X"B2",X"12",X"E8",X"20",X"3A",X"E2",X"02",X"AD",
		X"21",X"01",X"D1",X"82",X"8D",X"11",X"96",X"B9",X"02",X"1E",X"82",X"85",X"AB",X"28",X"3C",X"A3",
		X"01",X"1F",X"18",X"29",X"C2",X"19",X"6B",X"88",X"20",X"D0",X"29",X"6A",X"A1",X"82",X"BA",X"38",
		X"50",X"E1",X"82",X"9B",X"11",X"87",X"A9",X"82",X"0C",X"01",X"86",X"9A",X"00",X"1A",X"91",X"04",
		X"0D",X"19",X"28",X"C1",X"18",X"6B",X"0A",X"30",X"C0",X"19",X"79",X"98",X"01",X"A9",X"28",X"78",
		X"B0",X"82",X"9A",X"18",X"51",X"C1",X"A1",X"89",X"80",X"27",X"A8",X"A1",X"1A",X"91",X"87",X"0A",
		X"88",X"1A",X"90",X"07",X"1C",X"1A",X"18",X"90",X"84",X"3C",X"1B",X"00",X"A8",X"00",X"71",X"A8",
		X"90",X"B1",X"0A",X"72",X"B2",X"B8",X"90",X"90",X"37",X"80",X"AA",X"0B",X"29",X"97",X"3A",X"1B",
		X"AA",X"10",X"86",X"5A",X"1A",X"A9",X"92",X"8A",X"72",X"92",X"C9",X"A1",X"80",X"17",X"08",X"0B",
		X"A9",X"10",X"83",X"69",X"3A",X"E8",X"81",X"88",X"51",X"93",X"CB",X"90",X"28",X"97",X"19",X"2C",
		X"99",X"00",X"80",X"78",X"82",X"C9",X"81",X"80",X"97",X"88",X"1A",X"9A",X"2A",X"29",X"70",X"81",
		X"BA",X"A2",X"81",X"97",X"00",X"0B",X"AB",X"30",X"29",X"78",X"01",X"BB",X"B4",X"01",X"E6",X"91",
		X"09",X"A9",X"29",X"1E",X"78",X"00",X"A9",X"82",X"91",X"B7",X"80",X"89",X"99",X"28",X"2A",X"3A",
		X"23",X"D0",X"B2",X"C3",X"BA",X"71",X"2A",X"8D",X"18",X"0A",X"97",X"02",X"A9",X"B0",X"18",X"1E",
		X"79",X"29",X"8B",X"01",X"82",X"A3",X"A5",X"99",X"89",X"19",X"3F",X"95",X"02",X"9A",X"B2",X"80",
		X"9C",X"61",X"39",X"DA",X"11",X"81",X"D3",X"03",X"8B",X"BA",X"20",X"5A",X"03",X"08",X"89",X"F1",
		X"83",X"AA",X"B7",X"30",X"AA",X"A1",X"0A",X"9F",X"70",X"2A",X"AA",X"21",X"89",X"A7",X"94",X"99",
		X"B0",X"10",X"3A",X"91",X"03",X"99",X"D2",X"81",X"BA",X"E4",X"44",X"AC",X"80",X"08",X"8A",X"07",
		X"29",X"B8",X"A2",X"10",X"92",X"B7",X"A3",X"C0",X"93",X"80",X"BA",X"A5",X"60",X"99",X"B2",X"18",
		X"C0",X"A7",X"85",X"AA",X"92",X"00",X"8A",X"85",X"2A",X"9A",X"A1",X"42",X"9B",X"B6",X"96",X"A8",
		X"92",X"90",X"A8",X"B7",X"04",X"B9",X"A4",X"90",X"99",X"32",X"6A",X"AB",X"10",X"20",X"89",X"10",
		X"4A",X"9C",X"28",X"5B",X"0E",X"05",X"95",X"B0",X"A2",X"91",X"B0",X"B7",X"04",X"AA",X"A3",X"91",
		X"99",X"58",X"28",X"AE",X"10",X"10",X"A1",X"04",X"89",X"BB",X"12",X"2A",X"96",X"01",X"1E",X"A0",
		X"21",X"1C",X"C4",X"97",X"A1",X"B1",X"81",X"A8",X"A7",X"97",X"A8",X"91",X"92",X"99",X"28",X"38",
		X"AC",X"00",X"11",X"C4",X"A5",X"90",X"B8",X"81",X"19",X"11",X"59",X"0D",X"98",X"20",X"8A",X"68",
		X"20",X"BD",X"01",X"01",X"B2",X"B7",X"01",X"E1",X"A3",X"90",X"B6",X"93",X"9A",X"A0",X"10",X"0C",
		X"49",X"79",X"8A",X"09",X"28",X"90",X"23",X"08",X"DA",X"83",X"88",X"B7",X"83",X"0C",X"B0",X"18",
		X"2D",X"4A",X"79",X"0B",X"08",X"10",X"98",X"32",X"18",X"E9",X"92",X"00",X"C6",X"93",X"89",X"C8",
		X"10",X"1B",X"3A",X"78",X"0C",X"09",X"28",X"8A",X"41",X"20",X"CB",X"92",X"01",X"D4",X"97",X"90",
		X"B8",X"82",X"88",X"93",X"32",X"0F",X"9A",X"20",X"1C",X"5A",X"69",X"0B",X"09",X"28",X"88",X"23",
		X"01",X"F9",X"92",X"00",X"C5",X"A5",X"90",X"B0",X"81",X"0A",X"84",X"20",X"0E",X"8A",X"38",X"1D",
		X"48",X"39",X"8C",X"91",X"01",X"98",X"26",X"80",X"D8",X"92",X"81",X"C5",X"93",X"90",X"D0",X"81",
		X"88",X"93",X"31",X"0F",X"99",X"28",X"1B",X"49",X"79",X"1D",X"08",X"18",X"0A",X"48",X"39",X"9C",
		X"81",X"01",X"B2",X"07",X"80",X"D0",X"92",X"80",X"C4",X"84",X"98",X"C0",X"81",X"09",X"94",X"12",
		X"8C",X"A9",X"20",X"1E",X"38",X"69",X"0C",X"09",X"28",X"0C",X"48",X"38",X"9C",X"81",X"00",X"A9",
		X"61",X"01",X"D9",X"82",X"91",X"C3",X"06",X"90",X"C8",X"82",X"91",X"D4",X"83",X"98",X"C8",X"10",
		X"0A",X"94",X"31",X"8D",X"9A",X"38",X"1D",X"11",X"79",X"1C",X"09",X"29",X"1C",X"38",X"69",X"0C",
		X"08",X"18",X"0C",X"59",X"39",X"8B",X"08",X"10",X"9C",X"68",X"39",X"9B",X"00",X"00",X"AA",X"72",
		X"08",X"AB",X"93",X"92",X"E0",X"42",X"82",X"E9",X"82",X"91",X"C0",X"35",X"91",X"BA",X"A4",X"91",
		X"C2",X"17",X"90",X"B8",X"93",X"A1",X"D3",X"87",X"90",X"B1",X"A2",X"91",X"C4",X"96",X"90",X"B0",
		X"92",X"80",X"C4",X"95",X"90",X"B0",X"81",X"88",X"B5",X"96",X"89",X"A0",X"92",X"88",X"B7",X"94",
		X"98",X"B1",X"92",X"88",X"B6",X"83",X"8A",X"B8",X"01",X"0B",X"97",X"11",X"0C",X"A9",X"28",X"2C",
		X"03",X"79",X"1C",X"89",X"29",X"2C",X"11",X"69",X"1C",X"89",X"29",X"1B",X"48",X"79",X"0B",X"0A",
		X"39",X"1C",X"5A",X"59",X"0B",X"09",X"28",X"0B",X"69",X"39",X"8C",X"00",X"00",X"8B",X"68",X"38",
		X"AB",X"80",X"00",X"A8",X"72",X"00",X"D9",X"92",X"92",X"C2",X"25",X"90",X"D8",X"92",X"80",X"B5",
		X"97",X"90",X"B0",X"92",X"91",X"C5",X"95",X"A1",X"C1",X"91",X"91",X"A5",X"93",X"A0",X"C0",X"82",
		X"98",X"A6",X"01",X"89",X"B9",X"10",X"09",X"06",X"39",X"8B",X"BA",X"48",X"0C",X"30",X"78",X"0B",
		X"8B",X"28",X"0D",X"79",X"49",X"0C",X"08",X"18",X"0B",X"59",X"49",X"0C",X"08",X"19",X"1B",X"60",
		X"19",X"8C",X"08",X"18",X"88",X"42",X"09",X"9C",X"88",X"29",X"98",X"72",X"1A",X"9C",X"80",X"1A",
		X"93",X"37",X"09",X"C9",X"80",X"18",X"B6",X"85",X"88",X"C0",X"90",X"00",X"C6",X"82",X"88",X"C0",
		X"80",X"80",X"A6",X"83",X"99",X"C0",X"81",X"88",X"B7",X"83",X"89",X"C0",X"80",X"09",X"A7",X"83",
		X"98",X"C8",X"00",X"08",X"A5",X"03",X"0B",X"B9",X"08",X"1A",X"E6",X"03",X"0B",X"AB",X"28",X"1B",
		X"94",X"33",X"5D",X"8B",X"18",X"19",X"A9",X"70",X"49",X"9A",X"92",X"90",X"A9",X"34",X"06",X"A9",
		X"98",X"2A",X"0C",X"94",X"18",X"58",X"98",X"81",X"A9",X"B9",X"05",X"08",X"68",X"1A",X"2A",X"9A",
		X"CA",X"96",X"08",X"31",X"28",X"2B",X"AD",X"B9",X"91",X"49",X"26",X"22",X"09",X"C9",X"A9",X"A9",
		X"B8",X"32",X"64",X"11",X"88",X"0B",X"BD",X"C8",X"90",X"02",X"42",X"52",X"10",X"99",X"CB",X"A9",
		X"AB",X"10",X"61",X"38",X"11",X"22",X"10",X"C9",X"BC",X"D9",X"89",X"02",X"15",X"11",X"28",X"01",
		X"CB",X"98",X"92",X"A0",X"C1",X"20",X"CA",X"90",X"17",X"13",X"99",X"08",X"0B",X"A0",X"83",X"09",
		X"49",X"19",X"9A",X"9B",X"02",X"40",X"01",X"20",X"9C",X"B0",X"12",X"00",X"80",X"94",X"80",X"B8",
		X"81",X"0B",X"19",X"10",X"08",X"81",X"92",X"80",X"A9",X"10",X"8B",X"B0",X"20",X"31",X"02",X"89",
		X"89",X"A9",X"C0",X"30",X"80",X"01",X"11",X"00",X"98",X"A9",X"80",X"08",X"81",X"11",X"81",X"11",
		X"98",X"A8",X"98",X"90",X"82",X"11",X"00",X"81",X"A8",X"80",X"80",X"99",X"80",X"83",X"81",X"99",
		X"10",X"A1",X"91",X"91",X"88",X"90",X"91",X"21",X"80",X"90",X"99",X"90",X"12",X"80",X"80",X"19",
		X"89",X"08",X"10",X"80",X"91",X"01",X"98",X"A9",X"19",X"03",X"84",X"A8",X"98",X"00",X"81",X"98",
		X"98",X"20",X"19",X"80",X"80",X"80",X"81",X"88",X"00",X"09",X"98",X"20",X"00",X"09",X"89",X"B0",
		X"80",X"80",X"03",X"08",X"A9",X"8A",X"20",X"81",X"90",X"02",X"08",X"00",X"A8",X"91",X"87",X"99",
		X"39",X"90",X"92",X"B0",X"B4",X"85",X"8B",X"31",X"A0",X"3F",X"90",X"1A",X"32",X"A8",X"88",X"08",
		X"2A",X"0B",X"88",X"2A",X"0B",X"3B",X"40",X"14",X"38",X"AC",X"0A",X"FD",X"93",X"2A",X"72",X"12",
		X"0D",X"8A",X"9C",X"A3",X"0B",X"73",X"14",X"9C",X"98",X"BB",X"41",X"C6",X"29",X"2B",X"8A",X"BB",
		X"71",X"A7",X"09",X"9A",X"19",X"A2",X"58",X"58",X"B9",X"C2",X"9A",X"54",X"92",X"8B",X"BB",X"29",
		X"A7",X"69",X"1A",X"A8",X"91",X"90",X"71",X"08",X"E0",X"80",X"0B",X"71",X"A1",X"B8",X"1A",X"2A",
		X"27",X"90",X"8C",X"18",X"08",X"A7",X"1A",X"1C",X"10",X"90",X"92",X"7A",X"09",X"A2",X"91",X"9A",
		X"71",X"A0",X"B2",X"0A",X"09",X"46",X"B1",X"AA",X"39",X"09",X"B7",X"4C",X"0A",X"20",X"A0",X"00",
		X"7A",X"09",X"92",X"98",X"1B",X"72",X"D0",X"81",X"8A",X"10",X"97",X"98",X"89",X"29",X"91",X"94",
		X"3F",X"19",X"00",X"A2",X"0A",X"78",X"A0",X"92",X"99",X"28",X"97",X"A0",X"98",X"2B",X"10",X"A7",
		X"0B",X"2A",X"18",X"A3",X"9A",X"78",X"98",X"82",X"A8",X"2A",X"17",X"A1",X"B9",X"3B",X"39",X"A7",
		X"1B",X"2C",X"18",X"92",X"9B",X"71",X"99",X"A3",X"A0",X"4A",X"B7",X"92",X"9B",X"08",X"49",X"99",
		X"58",X"19",X"B0",X"83",X"B8",X"A7",X"21",X"CC",X"28",X"29",X"92",X"3C",X"5A",X"B8",X"85",X"89",
		X"39",X"A5",X"99",X"99",X"30",X"91",X"2A",X"79",X"B8",X"02",X"A0",X"C6",X"81",X"1C",X"88",X"10",
		X"8B",X"21",X"84",X"0B",X"81",X"19",X"AC",X"91",X"04",X"20",X"28",X"A0",X"9D",X"9C",X"09",X"15",
		X"18",X"48",X"11",X"9A",X"FA",X"89",X"84",X"13",X"22",X"29",X"B9",X"FB",X"A9",X"10",X"34",X"52",
		X"18",X"9B",X"99",X"DB",X"C8",X"24",X"33",X"12",X"18",X"AB",X"D9",X"CD",X"98",X"24",X"22",X"31",
		X"29",X"CA",X"A9",X"BE",X"A9",X"14",X"33",X"42",X"09",X"BA",X"80",X"CC",X"B8",X"91",X"34",X"63",
		X"20",X"BB",X"BB",X"BC",X"CB",X"08",X"32",X"73",X"43",X"31",X"11",X"AA",X"FB",X"AC",X"AA",X"B0",
		X"14",X"41",X"21",X"12",X"08",X"90",X"11",X"CC",X"EA",X"08",X"22",X"53",X"10",X"9A",X"1A",X"DA",
		X"B9",X"10",X"A8",X"07",X"21",X"28",X"10",X"A0",X"AA",X"0E",X"80",X"81",X"90",X"03",X"64",X"00",
		X"90",X"9D",X"BA",X"CA",X"AA",X"98",X"22",X"54",X"53",X"23",X"00",X"89",X"D9",X"DA",X"AA",X"AA",
		X"03",X"54",X"13",X"31",X"0A",X"CC",X"A9",X"90",X"99",X"88",X"25",X"35",X"21",X"89",X"8A",X"AB",
		X"E0",X"B9",X"09",X"C3",X"87",X"21",X"32",X"28",X"CB",X"9B",X"0B",X"89",X"AA",X"AC",X"00",X"54",
		X"33",X"12",X"09",X"B9",X"B8",X"AB",X"FA",X"08",X"00",X"36",X"31",X"09",X"88",X"0A",X"AB",X"08",
		X"BC",X"B3",X"13",X"53",X"44",X"00",X"AB",X"AA",X"AC",X"A8",X"8B",X"88",X"44",X"33",X"52",X"08",
		X"AA",X"BA",X"AB",X"BE",X"8A",X"02",X"04",X"52",X"11",X"90",X"89",X"BA",X"81",X"99",X"AD",X"82",
		X"20",X"36",X"21",X"9C",X"A9",X"98",X"D9",X"88",X"B8",X"84",X"33",X"61",X"31",X"08",X"AA",X"90",
		X"99",X"DA",X"AA",X"08",X"04",X"44",X"01",X"11",X"8B",X"CB",X"99",X"BA",X"9B",X"83",X"04",X"62",
		X"30",X"08",X"AA",X"8A",X"9B",X"AB",X"B9",X"B0",X"33",X"44",X"33",X"18",X"9A",X"99",X"B8",X"B8",
		X"D9",X"80",X"06",X"23",X"31",X"9A",X"9B",X"AA",X"98",X"CB",X"A9",X"00",X"45",X"24",X"22",X"09",
		X"AB",X"AB",X"9C",X"BA",X"9B",X"84",X"24",X"35",X"11",X"00",X"9B",X"99",X"BA",X"AB",X"89",X"01",
		X"35",X"41",X"10",X"98",X"C9",X"8A",X"AA",X"E8",X"B0",X"33",X"64",X"18",X"1A",X"C1",X"58",X"DA",
		X"9D",X"A1",X"50",X"52",X"20",X"BD",X"B9",X"D3",X"83",X"32",X"39",X"8F",X"CA",X"86",X"84",X"00",
		X"9C",X"8B",X"0C",X"72",X"01",X"9A",X"D8",X"80",X"87",X"11",X"9C",X"89",X"08",X"04",X"29",X"3C",
		X"B9",X"04",X"B9",X"72",X"99",X"A0",X"88",X"0A",X"17",X"01",X"AC",X"08",X"3A",X"B6",X"29",X"0B",
		X"90",X"83",X"DA",X"72",X"98",X"B0",X"10",X"8C",X"97",X"29",X"9B",X"20",X"0A",X"A0",X"72",X"AB",
		X"A6",X"89",X"88",X"07",X"8A",X"98",X"59",X"98",X"00",X"7A",X"98",X"04",X"AA",X"29",X"16",X"B9",
		X"00",X"4C",X"82",X"90",X"5C",X"00",X"82",X"C0",X"3B",X"86",X"A8",X"08",X"2B",X"02",X"BA",X"70",
		X"A0",X"82",X"8A",X"1A",X"B7",X"3E",X"00",X"01",X"A8",X"09",X"17",X"AA",X"28",X"29",X"B2",X"8A",
		X"70",X"D1",X"00",X"1B",X"01",X"A1",X"7A",X"A2",X"82",X"AA",X"28",X"B7",X"0C",X"10",X"01",X"B8",
		X"2A",X"17",X"B9",X"28",X"2A",X"B3",X"8B",X"71",X"D1",X"08",X"2B",X"82",X"99",X"79",X"A2",X"91",
		X"0C",X"10",X"93",X"3F",X"81",X"02",X"B9",X"28",X"B7",X"0C",X"10",X"00",X"B0",X"19",X"07",X"AA",
		X"39",X"2A",X"A2",X"0D",X"70",X"C1",X"00",X"0B",X"11",X"A1",X"6B",X"92",X"92",X"AA",X"39",X"A7",
		X"0C",X"28",X"00",X"B1",X"1A",X"17",X"AA",X"28",X"1A",X"A4",X"9A",X"52",X"C8",X"08",X"5B",X"A2",
		X"0A",X"78",X"B1",X"19",X"2C",X"01",X"98",X"79",X"B3",X"81",X"9A",X"29",X"B7",X"2E",X"01",X"80",
		X"90",X"09",X"87",X"9B",X"30",X"90",X"91",X"A9",X"70",X"C1",X"18",X"89",X"18",X"88",X"79",X"A2",
		X"88",X"0A",X"18",X"98",X"78",X"B2",X"00",X"1E",X"00",X"80",X"7A",X"A3",X"90",X"89",X"18",X"91",
		X"7A",X"91",X"81",X"9A",X"18",X"A7",X"2E",X"10",X"92",X"A8",X"09",X"17",X"B9",X"38",X"88",X"90",
		X"89",X"70",X"D2",X"09",X"19",X"88",X"81",X"7A",X"92",X"A2",X"8B",X"11",X"A8",X"79",X"A3",X"91",
		X"0D",X"00",X"80",X"7A",X"92",X"91",X"8B",X"28",X"93",X"5D",X"01",X"A3",X"9B",X"2A",X"A7",X"2E",
		X"11",X"91",X"A8",X"09",X"17",X"A9",X"39",X"80",X"A0",X"8A",X"71",X"D2",X"88",X"09",X"08",X"93",
		X"6C",X"01",X"A1",X"0A",X"08",X"A7",X"0B",X"28",X"81",X"A8",X"08",X"97",X"8B",X"39",X"11",X"D0",
		X"0A",X"44",X"D0",X"19",X"2A",X"90",X"89",X"70",X"C2",X"88",X"1A",X"08",X"90",X"79",X"92",X"A2",
		X"8B",X"08",X"A7",X"2E",X"10",X"81",X"A8",X"0A",X"37",X"B8",X"2A",X"28",X"B0",X"89",X"71",X"D1",
		X"08",X"19",X"90",X"91",X"7A",X"92",X"90",X"1B",X"08",X"A7",X"1C",X"10",X"92",X"9A",X"00",X"A7",
		X"0C",X"20",X"91",X"A8",X"09",X"27",X"B8",X"2A",X"39",X"A8",X"89",X"71",X"D2",X"88",X"19",X"90",
		X"90",X"79",X"91",X"92",X"8B",X"80",X"A7",X"2D",X"10",X"92",X"99",X"89",X"87",X"0B",X"29",X"10",
		X"B0",X"99",X"73",X"E0",X"19",X"18",X"A0",X"89",X"78",X"A1",X"08",X"1A",X"88",X"91",X"79",X"91",
		X"92",X"0C",X"80",X"96",X"1D",X"10",X"92",X"99",X"88",X"87",X"8B",X"39",X"01",X"B8",X"89",X"47",
		X"B8",X"19",X"28",X"B8",X"09",X"71",X"D1",X"08",X"1A",X"88",X"80",X"79",X"91",X"92",X"0B",X"90",
		X"95",X"6C",X"81",X"92",X"8A",X"80",X"97",X"0B",X"01",X"92",X"A9",X"09",X"87",X"0B",X"29",X"28",
		X"B9",X"09",X"47",X"B8",X"2A",X"28",X"B8",X"0A",X"73",X"E0",X"19",X"29",X"A0",X"88",X"78",X"B2",
		X"08",X"1B",X"88",X"91",X"78",X"B2",X"82",X"8D",X"08",X"81",X"7A",X"92",X"92",X"8C",X"00",X"A4",
		X"5C",X"01",X"A2",X"8B",X"08",X"87",X"0C",X"11",X"91",X"99",X"89",X"07",X"0C",X"28",X"82",X"B8",
		X"0A",X"27",X"9A",X"28",X"00",X"B8",X"0A",X"37",X"A9",X"2A",X"49",X"B0",X"89",X"72",X"D0",X"19",
		X"29",X"A8",X"88",X"71",X"D1",X"08",X"19",X"90",X"90",X"79",X"A2",X"80",X"0A",X"88",X"92",X"7A",
		X"92",X"92",X"8C",X"08",X"94",X"5C",X"82",X"92",X"9B",X"08",X"97",X"1D",X"10",X"81",X"99",X"09",
		X"87",X"0B",X"10",X"81",X"B8",X"09",X"07",X"0C",X"28",X"00",X"B8",X"1A",X"17",X"99",X"19",X"38",
		X"D0",X"88",X"27",X"A9",X"2A",X"28",X"B8",X"88",X"72",X"D0",X"19",X"29",X"A0",X"98",X"70",X"B1",
		X"08",X"1A",X"90",X"A0",X"70",X"B2",X"81",X"0D",X"08",X"92",X"7A",X"92",X"92",X"8C",X"08",X"94",
		X"5C",X"01",X"A2",X"8B",X"08",X"97",X"1C",X"10",X"92",X"A9",X"09",X"87",X"0B",X"28",X"01",X"C8",
		X"88",X"07",X"99",X"2A",X"38",X"C8",X"09",X"37",X"B8",X"2A",X"39",X"C0",X"89",X"71",X"C1",X"09",
		X"2A",X"90",X"98",X"70",X"B2",X"80",X"1C",X"80",X"90",X"78",X"B2",X"81",X"0C",X"08",X"93",X"7A",
		X"91",X"92",X"8B",X"80",X"A7",X"2C",X"01",X"92",X"9B",X"09",X"97",X"2D",X"10",X"81",X"A8",X"89",
		X"07",X"0C",X"10",X"00",X"A8",X"0A",X"27",X"A8",X"08",X"28",X"B8",X"89",X"72",X"D0",X"19",X"29",
		X"A0",X"98",X"71",X"C1",X"09",X"2A",X"90",X"90",X"70",X"C1",X"00",X"0A",X"90",X"91",X"79",X"91",
		X"93",X"8C",X"88",X"03",X"5C",X"81",X"92",X"8B",X"88",X"A7",X"3E",X"10",X"92",X"99",X"89",X"07",
		X"0B",X"00",X"01",X"B8",X"8A",X"27",X"99",X"19",X"48",X"C0",X"88",X"35",X"C8",X"19",X"28",X"B0",
		X"99",X"72",X"D1",X"09",X"3A",X"A0",X"98",X"71",X"C0",X"00",X"1A",X"90",X"90",X"78",X"A1",X"81",
		X"0B",X"90",X"94",X"7B",X"81",X"92",X"8B",X"88",X"97",X"2C",X"00",X"82",X"9A",X"89",X"87",X"2D",
		X"01",X"81",X"A9",X"09",X"87",X"0B",X"10",X"01",X"C8",X"09",X"17",X"99",X"08",X"20",X"C8",X"09",
		X"17",X"A8",X"1A",X"30",X"D0",X"88",X"25",X"B8",X"1A",X"48",X"B8",X"89",X"54",X"C0",X"09",X"39",
		X"B0",X"98",X"71",X"C0",X"18",X"19",X"A0",X"A8",X"72",X"D1",X"08",X"1A",X"90",X"98",X"71",X"C1",
		X"80",X"2C",X"80",X"91",X"69",X"90",X"81",X"1C",X"80",X"91",X"79",X"90",X"93",X"0C",X"88",X"83",
		X"6B",X"80",X"93",X"0D",X"08",X"95",X"2D",X"01",X"92",X"8B",X"09",X"87",X"1C",X"01",X"92",X"9A",
		X"0A",X"87",X"1C",X"10",X"82",X"B9",X"09",X"87",X"0B",X"18",X"12",X"C9",X"1A",X"07",X"89",X"09",
		X"22",X"D8",X"89",X"27",X"99",X"09",X"21",X"C8",X"09",X"35",X"B8",X"0A",X"40",X"C0",X"98",X"52",
		X"C0",X"09",X"39",X"B0",X"A9",X"73",X"D0",X"08",X"3A",X"A0",X"A8",X"71",X"B0",X"81",X"3D",X"91",
		X"A0",X"78",X"90",X"91",X"2C",X"88",X"94",X"4B",X"80",X"93",X"0C",X"89",X"97",X"2C",X"00",X"93",
		X"9A",X"89",X"97",X"2C",X"08",X"03",X"AA",X"0A",X"07",X"0A",X"09",X"22",X"C9",X"8A",X"46",X"A8",
		X"0A",X"30",X"B8",X"9B",X"73",X"C0",X"88",X"49",X"A0",X"A8",X"70",X"A0",X"80",X"3B",X"A0",X"A1",
		X"70",X"A1",X"B3",X"2C",X"98",X"B7",X"3B",X"80",X"A4",X"8B",X"0A",X"97",X"2B",X"09",X"04",X"AA",
		X"0B",X"27",X"89",X"1B",X"23",X"C8",X"AA",X"72",X"A8",X"0A",X"48",X"A8",X"A9",X"71",X"A1",X"A0",
		X"4A",X"98",X"B2",X"78",X"88",X"A2",X"2B",X"8A",X"C7",X"2A",X"88",X"93",X"0B",X"8A",X"A7",X"3B",
		X"1B",X"86",X"99",X"8A",X"07",X"88",X"0B",X"22",X"A9",X"9C",X"62",X"A0",X"99",X"38",X"A0",X"BA",
		X"73",X"A1",X"C0",X"3A",X"89",X"D3",X"69",X"80",X"B2",X"1A",X"0B",X"C7",X"19",X"09",X"93",X"89",
		X"8C",X"07",X"80",X"0B",X"02",X"90",X"AD",X"35",X"98",X"0B",X"20",X"90",X"BC",X"71",X"80",X"A9",
		X"20",X"98",X"C8",X"70",X"80",X"A8",X"28",X"8A",X"C2",X"79",X"00",X"A0",X"08",X"0A",X"C4",X"49",
		X"08",X"B2",X"09",X"0C",X"B7",X"10",X"0A",X"91",X"88",X"8C",X"97",X"18",X"09",X"91",X"88",X"8D",
		X"96",X"18",X"09",X"91",X"88",X"8C",X"95",X"20",X"88",X"A0",X"80",X"8E",X"92",X"50",X"00",X"B8",
		X"00",X"0D",X"B0",X"62",X"00",X"99",X"88",X"09",X"E9",X"06",X"10",X"09",X"98",X"00",X"BD",X"81",
		X"61",X"00",X"A8",X"80",X"8B",X"D8",X"05",X"30",X"08",X"A8",X"88",X"AE",X"A0",X"27",X"10",X"09",
		X"88",X"89",X"BD",X"91",X"27",X"18",X"08",X"08",X"9A",X"CB",X"00",X"13",X"71",X"01",X"89",X"9C",
		X"9A",X"A0",X"80",X"37",X"32",X"19",X"AA",X"BA",X"CA",X"B8",X"25",X"15",X"40",X"00",X"99",X"AC",
		X"AB",X"A8",X"15",X"21",X"33",X"14",X"0B",X"AD",X"99",X"DA",X"81",X"33",X"00",X"00",X"53",X"21",
		X"AC",X"AB",X"CD",X"A0",X"23",X"12",X"81",X"11",X"00",X"22",X"C0",X"9D",X"9A",X"A8",X"BB",X"98",
		X"71",X"22",X"24",X"48",X"98",X"8B",X"0E",X"99",X"A1",X"40",X"09",X"B0",X"3B",X"88",X"97",X"32",
		X"18",X"90",X"B9",X"0F",X"8A",X"20",X"08",X"83",X"83",X"19",X"BB",X"80",X"80",X"80",X"82",X"34",
		X"08",X"A8",X"C8",X"AB",X"A8",X"94",X"33",X"42",X"20",X"9C",X"BB",X"D9",X"90",X"01",X"54",X"22",
		X"18",X"9A",X"CA",X"BC",X"99",X"21",X"43",X"22",X"00",X"89",X"9A",X"C8",X"80",X"81",X"12",X"11",
		X"08",X"A9",X"9A",X"80",X"81",X"00",X"88",X"88",X"03",X"10",X"98",X"89",X"98",X"8B",X"84",X"13",
		X"10",X"00",X"A0",X"A9",X"A0",X"82",X"11",X"08",X"98",X"00",X"A2",X"80",X"81",X"20",X"A9",X"B8",
		X"81",X"10",X"A1",X"82",X"00",X"88",X"80",X"88",X"99",X"80",X"82",X"10",X"80",X"80",X"80",X"08",
		X"80",X"A0",X"82",X"A0",X"10",X"02",X"98",X"B8",X"80",X"90",X"11",X"00",X"01",X"A0",X"80",X"A9",
		X"80",X"80",X"80",X"11",X"00",X"80",X"89",X"80",X"80",X"80",X"80",X"80",X"80",X"88",X"01",X"90",
		X"B8",X"00",X"83",X"80",X"80",X"80",X"80",X"08",X"A0",X"80",X"90",X"00",X"10",X"B8",X"82",X"1A",
		X"88",X"10",X"3B",X"E4",X"1A",X"1A",X"20",X"B5",X"2B",X"C7",X"98",X"2C",X"92",X"C0",X"49",X"B0",
		X"57",X"1C",X"90",X"10",X"C9",X"09",X"04",X"03",X"5A",X"91",X"C0",X"0E",X"98",X"08",X"75",X"AA",
		X"02",X"2C",X"98",X"AA",X"37",X"4A",X"D0",X"40",X"AA",X"08",X"A2",X"71",X"E8",X"21",X"0C",X"00",
		X"A0",X"70",X"D1",X"01",X"8B",X"11",X"C5",X"2D",X"82",X"91",X"98",X"1C",X"44",X"D0",X"2B",X"18",
		X"08",X"B6",X"3E",X"01",X"91",X"98",X"0B",X"72",X"D8",X"39",X"98",X"28",X"C7",X"0D",X"21",X"A9",
		X"03",X"B9",X"79",X"B5",X"8A",X"82",X"1D",X"14",X"B8",X"29",X"98",X"21",X"E4",X"1D",X"03",X"A9",
		X"02",X"A9",X"78",X"C3",X"1B",X"93",X"0E",X"41",X"D1",X"2A",X"B2",X"5B",X"05",X"C9",X"5A",X"A0",
		X"30",X"E5",X"8D",X"30",X"A9",X"22",X"BB",X"70",X"C3",X"09",X"B3",X"2F",X"42",X"D9",X"48",X"B8",
		X"4A",X"34",X"DB",X"50",X"D0",X"5C",X"33",X"E9",X"59",X"D1",X"4B",X"33",X"F8",X"49",X"B8",X"58",
		X"C5",X"9C",X"31",X"AB",X"34",X"C8",X"5A",X"92",X"8B",X"97",X"A9",X"69",X"D2",X"3A",X"C3",X"09",
		X"7B",X"D3",X"4C",X"B4",X"08",X"6D",X"C5",X"2C",X"A3",X"83",X"4E",X"B5",X"0A",X"A2",X"04",X"3F",
		X"A4",X"0A",X"A3",X"1C",X"6A",X"B2",X"29",X"C0",X"6A",X"A6",X"AA",X"30",X"AC",X"30",X"C7",X"0D",
		X"02",X"8B",X"03",X"E5",X"2D",X"A3",X"0C",X"03",X"C5",X"2D",X"A1",X"3B",X"94",X"B3",X"4C",X"99",
		X"30",X"D3",X"88",X"6B",X"0B",X"03",X"B2",X"0C",X"79",X"88",X"A4",X"A9",X"3B",X"78",X"B1",X"92",
		X"9A",X"0A",X"73",X"C8",X"A3",X"0A",X"29",X"A5",X"80",X"0C",X"29",X"08",X"81",X"2B",X"20",X"09",
		X"C0",X"21",X"8D",X"90",X"78",X"88",X"01",X"1B",X"B8",X"11",X"90",X"83",X"42",X"A9",X"9A",X"CA",
		X"88",X"24",X"07",X"18",X"A9",X"88",X"9A",X"A9",X"26",X"12",X"01",X"18",X"AC",X"CA",X"9B",X"04",
		X"43",X"31",X"01",X"2F",X"B8",X"AA",X"89",X"03",X"81",X"88",X"82",X"A1",X"90",X"81",X"90",X"80",
		X"81",X"90",X"80",X"80",X"80",X"80",X"80",X"81",X"90",X"80",X"80",X"80",X"80",X"81",X"88",X"81",
		X"90",X"80",X"82",X"9A",X"12",X"A0",X"8B",X"32",X"89",X"A2",X"80",X"80",X"01",X"A0",X"80",X"39",
		X"A0",X"0C",X"03",X"80",X"84",X"0C",X"8E",X"93",X"31",X"13",X"BD",X"61",X"A9",X"0B",X"E0",X"AE",
		X"84",X"51",X"88",X"00",X"08",X"C8",X"88",X"21",X"BF",X"E9",X"36",X"19",X"80",X"00",X"03",X"8F",
		X"F9",X"26",X"89",X"91",X"00",X"90",X"00",X"91",X"19",X"BF",X"96",X"39",X"B0",X"28",X"C9",X"44",
		X"9B",X"09",X"D0",X"71",X"A9",X"10",X"98",X"23",X"BF",X"93",X"20",X"AA",X"15",X"2B",X"F9",X"35",
		X"9B",X"82",X"28",X"98",X"F0",X"58",X"B0",X"20",X"88",X"1C",X"B6",X"2B",X"92",X"19",X"83",X"F9",
		X"41",X"C0",X"28",X"80",X"0C",X"04",X"9A",X"28",X"01",X"98",X"1E",X"05",X"AA",X"21",X"08",X"00",
		X"F0",X"6A",X"A1",X"10",X"80",X"BC",X"61",X"B8",X"10",X"29",X"A9",X"04",X"0D",X"02",X"00",X"B8",
		X"7B",X"95",X"99",X"10",X"1A",X"10",X"F2",X"3D",X"81",X"10",X"90",X"D1",X"5A",X"A2",X"81",X"88",
		X"0E",X"25",X"C9",X"38",X"09",X"A5",X"8B",X"21",X"A1",X"B5",X"1B",X"2F",X"15",X"D9",X"21",X"09",
		X"2F",X"05",X"9C",X"11",X"00",X"8B",X"20",X"00",X"C2",X"1B",X"59",X"81",X"F3",X"3F",X"01",X"81",
		X"83",X"F9",X"5A",X"A3",X"00",X"91",X"AB",X"70",X"A8",X"84",X"0A",X"8C",X"43",X"D9",X"22",X"AA",
		X"34",X"F0",X"39",X"99",X"40",X"A6",X"D9",X"5A",X"92",X"02",X"E3",X"8D",X"48",X"91",X"B5",X"88",
		X"89",X"85",X"9A",X"83",X"2D",X"84",X"B0",X"2A",X"1B",X"07",X"91",X"BB",X"78",X"B0",X"23",X"F3",
		X"9C",X"5A",X"01",X"E4",X"2C",X"81",X"08",X"90",X"19",X"A7",X"88",X"8D",X"50",X"D0",X"06",X"C8",
		X"4D",X"12",X"A3",X"D1",X"29",X"80",X"B3",X"2D",X"1A",X"41",X"C3",X"9E",X"31",X"A9",X"06",X"A8",
		X"2B",X"83",X"A1",X"B8",X"79",X"18",X"C0",X"38",X"AA",X"51",X"A8",X"2E",X"12",X"99",X"95",X"89",
		X"28",X"F2",X"19",X"98",X"58",X"90",X"8A",X"21",X"9B",X"24",X"98",X"3F",X"83",X"90",X"B1",X"38",
		X"11",X"F8",X"28",X"8D",X"50",X"A1",X"1D",X"01",X"00",X"C3",X"08",X"00",X"C8",X"12",X"8B",X"31",
		X"82",X"9F",X"81",X"3B",X"B5",X"19",X"39",X"F0",X"10",X"98",X"38",X"83",X"AF",X"81",X"10",X"91",
		X"80",X"59",X"E0",X"08",X"10",X"19",X"01",X"0A",X"C9",X"04",X"10",X"A2",X"10",X"1F",X"B8",X"24",
		X"0A",X"11",X"B4",X"1F",X"98",X"13",X"81",X"9B",X"42",X"AB",X"AB",X"36",X"3A",X"B0",X"50",X"AA",
		X"9B",X"27",X"8A",X"02",X"11",X"0D",X"A0",X"19",X"80",X"30",X"20",X"1A",X"B1",X"DD",X"82",X"31",
		X"82",X"03",X"1E",X"C8",X"91",X"89",X"32",X"60",X"9C",X"83",X"09",X"BA",X"A4",X"68",X"B8",X"32",
		X"8A",X"92",X"01",X"8F",X"C1",X"38",X"88",X"02",X"40",X"C8",X"03",X"8D",X"C0",X"03",X"0A",X"10",
		X"61",X"AA",X"81",X"19",X"CB",X"96",X"18",X"91",X"03",X"0D",X"19",X"31",X"BC",X"08",X"19",X"A8",
		X"17",X"3A",X"A1",X"01",X"99",X"AB",X"40",X"9D",X"13",X"39",X"B8",X"04",X"2B",X"D9",X"41",X"B8",
		X"B3",X"58",X"B9",X"92",X"2A",X"0C",X"27",X"89",X"98",X"03",X"9A",X"B0",X"52",X"9B",X"01",X"08",
		X"98",X"95",X"0B",X"8A",X"21",X"90",X"89",X"30",X"89",X"81",X"88",X"80",X"A4",X"98",X"80",X"81",
		X"90",X"80",X"00",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"90",X"80",X"80",X"80",
		X"80",X"81",X"91",X"91",X"90",X"80",X"80",X"80",X"81",X"90",X"80",X"80",X"80",X"80",X"00",X"90",
		X"80",X"81",X"90",X"81",X"88",X"80",X"08",X"08",X"80",X"81",X"90",X"81",X"91",X"91",X"91",X"91",
		X"90",X"81",X"80",X"91",X"91",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"81",X"90",X"80",X"80",X"81",X"81",X"98",X"89",X"82",X"81",X"02",X"8A",
		X"99",X"82",X"80",X"80",X"03",X"08",X"C0",X"B1",X"10",X"A0",X"1B",X"78",X"4C",X"0B",X"19",X"4A",
		X"00",X"38",X"A5",X"98",X"AD",X"10",X"4D",X"11",X"4A",X"4F",X"09",X"01",X"91",X"22",X"1B",X"8C",
		X"A9",X"B4",X"E6",X"32",X"BB",X"9D",X"03",X"83",X"F1",X"51",X"AC",X"99",X"24",X"28",X"F8",X"41",
		X"9A",X"C0",X"32",X"2D",X"B2",X"50",X"AB",X"B4",X"32",X"AF",X"84",X"29",X"CA",X"14",X"19",X"BB",
		X"53",X"2E",X"B1",X"23",X"9B",X"B2",X"51",X"1F",X"91",X"21",X"BB",X"31",X"11",X"AF",X"11",X"10",
		X"C0",X"19",X"02",X"3D",X"C0",X"34",X"AB",X"80",X"40",X"00",X"F8",X"31",X"8F",X"01",X"00",X"92",
		X"8C",X"02",X"2A",X"B1",X"21",X"9A",X"50",X"F0",X"12",X"9C",X"03",X"0A",X"96",X"8C",X"83",X"19",
		X"B0",X"40",X"B9",X"50",X"AC",X"24",X"9A",X"94",X"1D",X"83",X"3C",X"C1",X"48",X"A9",X"22",X"AA",
		X"15",X"99",X"D3",X"4B",X"98",X"40",X"D1",X"11",X"A9",X"94",X"1B",X"80",X"29",X"C4",X"18",X"C8",
		X"14",X"A9",X"00",X"2B",X"93",X"48",X"F0",X"03",X"A9",X"19",X"2B",X"05",X"88",X"B1",X"95",X"A0",
		X"0B",X"38",X"1B",X"07",X"B4",X"F1",X"3B",X"0A",X"22",X"D2",X"82",X"A0",X"D2",X"3A",X"A8",X"40",
		X"AA",X"17",X"A8",X"80",X"83",X"B0",X"0A",X"5C",X"20",X"03",X"CF",X"14",X"9A",X"82",X"2C",X"83",
		X"2B",X"D2",X"3C",X"08",X"20",X"C1",X"82",X"8A",X"59",X"0F",X"14",X"A9",X"01",X"2E",X"03",X"8A",
		X"94",X"98",X"0A",X"48",X"B1",X"13",X"E8",X"38",X"1F",X"04",X"A8",X"81",X"1A",X"80",X"39",X"B4",
		X"D2",X"2D",X"10",X"80",X"92",X"88",X"18",X"BB",X"70",X"90",X"B2",X"49",X"B0",X"7A",X"94",X"B8",
		X"4B",X"10",X"A1",X"82",X"89",X"48",X"DA",X"60",X"99",X"82",X"1B",X"03",X"0C",X"82",X"C3",X"8A",
		X"4B",X"84",X"88",X"93",X"88",X"1F",X"15",X"D0",X"93",X"0B",X"28",X"11",X"8F",X"85",X"99",X"80",
		X"28",X"A2",X"19",X"09",X"F4",X"1B",X"09",X"21",X"D2",X"29",X"9A",X"5B",X"03",X"B1",X"98",X"38",
		X"1B",X"97",X"09",X"F2",X"4B",X"98",X"22",X"B8",X"93",X"5B",X"1F",X"06",X"A9",X"00",X"2A",X"81",
		X"19",X"1A",X"E4",X"1A",X"09",X"03",X"C1",X"18",X"89",X"3F",X"12",X"A8",X"80",X"28",X"88",X"A3",
		X"31",X"FE",X"41",X"A8",X"80",X"39",X"A9",X"60",X"98",X"F2",X"3B",X"89",X"22",X"A9",X"02",X"3B",
		X"9F",X"15",X"A8",X"88",X"38",X"8A",X"04",X"9A",X"12",X"F1",X"29",X"9A",X"41",X"C2",X"81",X"10",
		X"FB",X"52",X"9B",X"94",X"2B",X"88",X"31",X"BA",X"3D",X"32",X"D8",X"28",X"0A",X"21",X"91",X"B0",
		X"7F",X"04",X"A8",X"08",X"2A",X"94",X"88",X"08",X"8F",X"23",X"AA",X"83",X"2C",X"80",X"13",X"BB",
		X"33",X"BF",X"20",X"19",X"B3",X"0A",X"58",X"90",X"15",X"FA",X"79",X"88",X"01",X"98",X"19",X"11",
		X"A8",X"03",X"F8",X"38",X"88",X"92",X"98",X"49",X"80",X"03",X"FB",X"78",X"98",X"02",X"8A",X"1A",
		X"24",X"C8",X"11",X"2F",X"95",X"89",X"90",X"29",X"82",X"90",X"00",X"2F",X"A6",X"89",X"88",X"20",
		X"A0",X"00",X"1A",X"01",X"A5",X"E0",X"4A",X"80",X"93",X"9A",X"48",X"90",X"12",X"CF",X"23",X"9A",
		X"A4",X"2C",X"18",X"92",X"1A",X"89",X"43",X"F9",X"59",X"89",X"84",X"99",X"29",X"80",X"12",X"CF",
		X"23",X"9A",X"93",X"2B",X"08",X"A4",X"09",X"89",X"34",X"FA",X"50",X"99",X"93",X"2C",X"01",X"88",
		X"12",X"9F",X"96",X"0B",X"81",X"10",X"A1",X"99",X"40",X"A9",X"03",X"4F",X"A5",X"09",X"99",X"31",
		X"A8",X"08",X"30",X"98",X"F8",X"58",X"90",X"91",X"19",X"08",X"A3",X"2A",X"99",X"15",X"8F",X"85",
		X"89",X"B1",X"58",X"A8",X"12",X"8A",X"01",X"D9",X"58",X"88",X"91",X"2B",X"04",X"99",X"03",X"0D",
		X"94",X"B9",X"58",X"90",X"B2",X"4A",X"80",X"11",X"A1",X"0B",X"7E",X"B6",X"1A",X"89",X"23",X"BA",
		X"12",X"19",X"80",X"B0",X"31",X"DC",X"25",X"9A",X"81",X"3A",X"93",X"80",X"8B",X"51",X"A4",X"FD",
		X"50",X"98",X"91",X"28",X"8A",X"83",X"10",X"9D",X"02",X"83",X"DC",X"32",X"90",X"A9",X"58",X"92",
		X"09",X"A1",X"20",X"85",X"FE",X"32",X"98",X"A9",X"60",X"B0",X"10",X"19",X"88",X"81",X"09",X"3F",
		X"A5",X"0A",X"2A",X"93",X"09",X"01",X"89",X"94",X"19",X"A0",X"BF",X"35",X"B8",X"1A",X"32",X"E0",
		X"39",X"92",X"89",X"08",X"88",X"23",X"FD",X"50",X"A1",X"A0",X"39",X"93",X"99",X"18",X"11",X"C9",
		X"44",X"FC",X"32",X"90",X"A8",X"30",X"A2",X"89",X"38",X"92",X"C9",X"18",X"07",X"CC",X"22",X"02",
		X"DB",X"34",X"88",X"A0",X"10",X"80",X"A0",X"2A",X"2C",X"F9",X"78",X"08",X"B1",X"48",X"80",X"98",
		X"28",X"A1",X"8A",X"01",X"33",X"FF",X"22",X"88",X"B8",X"40",X"80",X"89",X"19",X"11",X"98",X"A0",
		X"2F",X"F3",X"18",X"1B",X"02",X"11",X"1B",X"C0",X"14",X"8A",X"C9",X"13",X"11",X"DF",X"14",X"88",
		X"8A",X"13",X"90",X"1A",X"91",X"00",X"89",X"0C",X"21",X"FE",X"40",X"81",X"A8",X"22",X"28",X"B9",
		X"9D",X"14",X"2B",X"B8",X"18",X"29",X"84",X"F9",X"68",X"81",X"A9",X"21",X"18",X"A9",X"11",X"A8",
		X"2D",X"D2",X"2A",X"E1",X"22",X"39",X"F8",X"32",X"1B",X"B2",X"1B",X"81",X"A8",X"85",X"4F",X"D3",
		X"28",X"1A",X"B3",X"18",X"10",X"B0",X"88",X"11",X"0C",X"D8",X"31",X"1F",X"B5",X"28",X"0B",X"01",
		X"80",X"48",X"A8",X"91",X"0A",X"02",X"0F",X"00",X"1E",X"B4",X"48",X"0A",X"91",X"28",X"38",X"A0",
		X"BB",X"23",X"0A",X"9C",X"08",X"48",X"F9",X"78",X"00",X"A8",X"3A",X"93",X"10",X"9B",X"B4",X"31",
		X"DB",X"92",X"08",X"27",X"CC",X"24",X"81",X"99",X"9A",X"54",X"8B",X"80",X"18",X"A9",X"93",X"08",
		X"B8",X"0E",X"13",X"11",X"29",X"88",X"D5",X"49",X"88",X"90",X"AB",X"28",X"E8",X"28",X"08",X"07",
		X"1D",X"92",X"02",X"08",X"C8",X"25",X"8B",X"88",X"02",X"AA",X"9B",X"51",X"08",X"BC",X"37",X"89",
		X"09",X"13",X"8B",X"84",X"22",X"C8",X"C0",X"18",X"88",X"80",X"FD",X"22",X"11",X"09",X"80",X"24",
		X"9A",X"B8",X"03",X"98",X"9A",X"09",X"18",X"98",X"21",X"21",X"20",X"EA",X"81",X"21",X"2B",X"8C",
		X"31",X"3A",X"89",X"00",X"09",X"0A",X"28",X"08",X"B8",X"25",X"09",X"AA",X"94",X"10",X"98",X"82",
		X"10",X"A9",X"12",X"8A",X"C8",X"01",X"19",X"98",X"08",X"12",X"89",X"82",X"10",X"A2",X"11",X"00",
		X"A9",X"A0",X"B0",X"90",X"03",X"19",X"A2",X"A3",X"09",X"80",X"13",X"0C",X"CA",X"20",X"30",X"80",
		X"80",X"01",X"10",X"80",X"A8",X"90",X"80",X"80",X"89",X"88",X"2A",X"81",X"10",X"01",X"80",X"82",
		X"80",X"89",X"88",X"90",X"89",X"90",X"20",X"80",X"80",X"80",X"80",X"81",X"80",X"9A",X"02",X"00",
		X"90",X"81",X"09",X"82",X"19",X"A0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"01",X"91",X"80",X"98",X"82",X"1A",X"90",X"80",X"80",X"80",X"80",X"80",X"81",X"90",X"80",X"80",
		X"80",X"00",X"91",X"80",X"90",X"81",X"08",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"89",X"10",X"00",X"90",X"00",X"91",X"91",X"88",X"81",X"90",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"80",X"81",X"80",X"92",X"98",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"91",X"88",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"80",X"00",X"88",
		X"00",X"88",X"08",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"90",X"80",
		X"81",X"80",X"91",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"81",X"80",X"00",X"88",X"80",X"80",X"90",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"90",X"00",X"90",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"90",X"81",X"90",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",
		X"81",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"18",X"09",X"0C",X"19",X"4A",X"D3",X"41",X"88",X"A2",
		X"F0",X"C0",X"17",X"84",X"54",X"9F",X"CA",X"84",X"31",X"08",X"9A",X"A0",X"09",X"64",X"AD",X"D1",
		X"70",X"A8",X"02",X"3F",X"B2",X"22",X"9C",X"02",X"08",X"01",X"9F",X"01",X"39",X"E0",X"48",X"90",
		X"1A",X"B1",X"50",X"BA",X"42",X"A8",X"31",X"FB",X"61",X"C9",X"22",X"A9",X"48",X"0E",X"85",X"0C",
		X"94",X"1B",X"01",X"00",X"F1",X"39",X"B8",X"69",X"91",X"2A",X"0F",X"58",X"9A",X"05",X"A8",X"39",
		X"9A",X"14",X"C2",X"B3",X"8A",X"50",X"A9",X"94",X"81",X"E1",X"18",X"82",X"B6",X"E2",X"3C",X"82",
		X"A1",X"02",X"90",X"E2",X"19",X"A0",X"11",X"C5",X"91",X"D3",X"0C",X"11",X"98",X"04",X"A9",X"19",
		X"3F",X"4B",X"01",X"92",X"90",X"90",X"2E",X"23",X"D8",X"13",X"AB",X"4B",X"29",X"05",X"D0",X"11",
		X"8A",X"18",X"09",X"1B",X"59",X"A6",X"88",X"F5",X"99",X"08",X"2A",X"11",X"2F",X"12",X"C1",X"A4",
		X"B1",X"18",X"9A",X"6B",X"3C",X"3A",X"85",X"A2",X"E5",X"A1",X"B0",X"5C",X"28",X"1C",X"30",X"C5",
		X"D1",X"01",X"88",X"3F",X"29",X"4D",X"11",X"81",X"94",X"F4",X"91",X"A8",X"3B",X"28",X"5F",X"21",
		X"A2",X"D3",X"90",X"01",X"C2",X"0B",X"6C",X"28",X"82",X"8B",X"11",X"8B",X"B7",X"88",X"31",X"F1",
		X"2C",X"08",X"3B",X"03",X"8C",X"86",X"9B",X"86",X"9A",X"50",X"D0",X"5D",X"88",X"6C",X"12",X"0F",
		X"24",X"C9",X"05",X"B2",X"81",X"F2",X"4C",X"91",X"4B",X"18",X"4D",X"05",X"C8",X"85",X"B1",X"2A",
		X"D2",X"02",X"E1",X"3A",X"28",X"D0",X"11",X"8B",X"85",X"00",X"99",X"A1",X"31",X"F9",X"58",X"18",
		X"B9",X"21",X"2E",X"82",X"02",X"8B",X"C1",X"24",X"BC",X"21",X"48",X"BC",X"01",X"49",X"B0",X"14",
		X"00",X"D9",X"82",X"29",X"98",X"24",X"0B",X"CA",X"14",X"81",X"A0",X"30",X"8A",X"BA",X"10",X"21",
		X"01",X"83",X"2B",X"9C",X"E0",X"01",X"08",X"23",X"01",X"2E",X"B9",X"00",X"B1",X"18",X"45",X"81",
		X"00",X"BD",X"89",X"A9",X"38",X"33",X"63",X"A1",X"9E",X"99",X"8B",X"04",X"29",X"14",X"19",X"30",
		X"EA",X"00",X"B0",X"1B",X"A6",X"38",X"05",X"08",X"88",X"DB",X"82",X"B8",X"31",X"04",X"3A",X"91",
		X"3A",X"D1",X"B9",X"33",X"CC",X"13",X"21",X"49",X"D0",X"4C",X"BD",X"99",X"A0",X"BB",X"17",X"88",
		X"83",X"02",X"40",X"93",X"42",X"18",X"13",X"54",X"09",X"01",X"39",X"C9",X"B8",X"39",X"EA",X"80",
		X"8B",X"BD",X"92",X"0C",X"99",X"08",X"80",X"C9",X"11",X"90",X"C1",X"91",X"09",X"03",X"80",X"80",
		X"08",X"80",X"80",X"00",X"91",X"20",X"80",X"80",X"12",X"80",X"81",X"08",X"08",X"92",X"10",X"89",
		X"11",X"91",X"91",X"81",X"08",X"91",X"88",X"08",X"90",X"81",X"89",X"09",X"80",X"88",X"80",X"80",
		X"90",X"80",X"80",X"80",X"01",X"80",X"90",X"00",X"80",X"81",X"00",X"89",X"19",X"88",X"80",X"80",
		X"80",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"08",X"18",X"1A",X"88",X"10",X"80",
		X"80",X"80",X"98",X"08",X"82",X"A1",X"80",X"90",X"81",X"90",X"80",X"80",X"80",X"A2",X"A2",X"80",
		X"80",X"89",X"19",X"91",X"82",X"8B",X"30",X"80",X"A0",X"1A",X"08",X"20",X"81",X"B8",X"80",X"81",
		X"11",X"83",X"00",X"D0",X"B8",X"A2",X"A6",X"13",X"82",X"D0",X"A9",X"8A",X"A8",X"83",X"53",X"24",
		X"AF",X"89",X"89",X"2B",X"98",X"72",X"13",X"B8",X"BB",X"A3",X"9B",X"C3",X"16",X"78",X"1A",X"8D",
		X"19",X"80",X"89",X"06",X"38",X"3A",X"CA",X"8A",X"93",X"AB",X"47",X"29",X"6A",X"9A",X"80",X"A1",
		X"99",X"33",X"70",X"3C",X"9D",X"18",X"A1",X"92",X"86",X"21",X"9B",X"0F",X"08",X"1B",X"11",X"24",
		X"97",X"A8",X"B0",X"8A",X"29",X"28",X"71",X"08",X"B1",X"E0",X"92",X"A2",X"02",X"6A",X"4B",X"8B",
		X"81",X"C2",X"94",X"95",X"01",X"9B",X"1E",X"1A",X"18",X"00",X"25",X"A5",X"A9",X"A9",X"1A",X"19",
		X"20",X"37",X"82",X"C0",X"C9",X"18",X"0A",X"38",X"33",X"24",X"D8",X"D8",X"00",X"89",X"00",X"36",
		X"02",X"9A",X"D8",X"08",X"0A",X"19",X"34",X"37",X"8B",X"9A",X"1A",X"19",X"0E",X"30",X"51",X"2B",
		X"0E",X"81",X"90",X"B0",X"00",X"52",X"48",X"B8",X"C0",X"90",X"8B",X"0B",X"75",X"83",X"A9",X"AB",
		X"2B",X"0A",X"29",X"17",X"34",X"8D",X"0B",X"89",X"8A",X"12",X"64",X"82",X"1F",X"0C",X"88",X"93",
		X"13",X"73",X"E0",X"B8",X"90",X"3A",X"29",X"55",X"2D",X"9C",X"01",X"12",X"A8",X"B7",X"21",X"E9",
		X"A2",X"23",X"9C",X"90",X"61",X"3F",X"99",X"22",X"09",X"D0",X"14",X"01",X"F9",X"02",X"3A",X"AB",
		X"14",X"31",X"AF",X"91",X"32",X"CA",X"82",X"38",X"1B",X"9B",X"24",X"3C",X"B0",X"14",X"90",X"0A",
		X"6F",X"10",X"01",X"C1",X"81",X"0A",X"28",X"4F",X"00",X"10",X"B1",X"82",X"99",X"38",X"5F",X"82",
		X"82",X"C8",X"10",X"09",X"20",X"A0",X"E4",X"09",X"8A",X"58",X"8A",X"13",X"92",X"F8",X"39",X"1E",
		X"12",X"98",X"83",X"A3",X"F8",X"5A",X"89",X"04",X"A9",X"02",X"2E",X"83",X"A1",X"A0",X"4B",X"00",
		X"18",X"A5",X"93",X"F8",X"4A",X"1B",X"14",X"C0",X"02",X"8B",X"3C",X"21",X"B1",X"91",X"2C",X"18",
		X"38",X"D5",X"C1",X"2C",X"2A",X"02",X"A1",X"93",X"89",X"4F",X"11",X"A0",X"A4",X"89",X"81",X"3C",
		X"86",X"D1",X"19",X"0A",X"20",X"90",X"84",X"A0",X"8E",X"6A",X"81",X"92",X"99",X"20",X"0A",X"97",
		X"D1",X"19",X"1B",X"21",X"98",X"84",X"98",X"3F",X"28",X"A1",X"A4",X"89",X"01",X"1B",X"87",X"E1",
		X"2A",X"09",X"03",X"A8",X"03",X"8B",X"5F",X"12",X"B0",X"81",X"1A",X"82",X"19",X"B7",X"B9",X"6A",
		X"08",X"93",X"98",X"01",X"1B",X"6F",X"04",X"B0",X"08",X"19",X"00",X"01",X"A1",X"0F",X"38",X"91",
		X"B2",X"19",X"08",X"4A",X"2B",X"F6",X"99",X"19",X"10",X"91",X"81",X"8A",X"7E",X"03",X"A0",X"90",
		X"29",X"09",X"21",X"A4",X"F0",X"3B",X"19",X"81",X"00",X"A2",X"2A",X"3F",X"A7",X"99",X"19",X"10",
		X"88",X"03",X"90",X"EA",X"79",X"81",X"A1",X"19",X"08",X"10",X"96",X"F0",X"3A",X"09",X"82",X"80",
		X"91",X"29",X"3F",X"A6",X"98",X"09",X"02",X"99",X"12",X"99",X"6F",X"11",X"91",X"99",X"20",X"89",
		X"11",X"94",X"F9",X"59",X"80",X"91",X"19",X"80",X"29",X"96",X"E0",X"29",X"08",X"92",X"80",X"90",
		X"28",X"1B",X"F5",X"99",X"2A",X"83",X"89",X"02",X"89",X"5E",X"96",X"99",X"19",X"01",X"89",X"11",
		X"90",X"4F",X"83",X"90",X"99",X"21",X"8A",X"13",X"90",X"1F",X"00",X"95",X"BA",X"40",X"89",X"10",
		X"02",X"BF",X"49",X"93",X"B8",X"38",X"89",X"38",X"83",X"AF",X"39",X"A6",X"B9",X"30",X"89",X"20",
		X"82",X"9F",X"28",X"B7",X"A9",X"20",X"88",X"01",X"00",X"2F",X"81",X"94",X"BB",X"41",X"99",X"12",
		X"80",X"3F",X"B7",X"98",X"09",X"01",X"09",X"83",X"90",X"2D",X"C6",X"98",X"2B",X"82",X"08",X"91",
		X"28",X"20",X"F9",X"29",X"5B",X"B4",X"19",X"80",X"10",X"88",X"0F",X"28",X"95",X"BA",X"58",X"88",
		X"01",X"08",X"2F",X"95",X"98",X"09",X"01",X"88",X"01",X"80",X"01",X"F9",X"38",X"2B",X"B4",X"18",
		X"98",X"30",X"80",X"4F",X"A4",X"92",X"BB",X"50",X"89",X"03",X"88",X"18",X"F0",X"19",X"4B",X"C4",
		X"08",X"88",X"38",X"88",X"2F",X"82",X"92",X"AB",X"41",X"8A",X"12",X"08",X"86",X"FA",X"79",X"92",
		X"A0",X"18",X"80",X"00",X"01",X"9C",X"B7",X"89",X"3B",X"A5",X"88",X"80",X"10",X"89",X"4F",X"83",
		X"98",X"1B",X"21",X"98",X"83",X"80",X"09",X"2F",X"01",X"A5",X"AD",X"40",X"90",X"92",X"00",X"81",
		X"F9",X"69",X"92",X"A8",X"39",X"80",X"81",X"00",X"A4",X"DB",X"78",X"92",X"A9",X"39",X"08",X"82",
		X"01",X"A4",X"FA",X"69",X"81",X"A0",X"29",X"88",X"11",X"82",X"B4",X"F9",X"48",X"80",X"A0",X"3A",
		X"88",X"12",X"82",X"B5",X"FA",X"58",X"80",X"A1",X"2A",X"08",X"01",X"02",X"B3",X"FC",X"68",X"91",
		X"A0",X"29",X"08",X"82",X"01",X"A0",X"CD",X"78",X"91",X"99",X"38",X"90",X"92",X"11",X"8B",X"3F",
		X"01",X"82",X"AF",X"31",X"A0",X"91",X"20",X"1A",X"4F",X"B5",X"09",X"09",X"83",X"98",X"08",X"11",
		X"3B",X"91",X"F0",X"19",X"4A",X"E3",X"19",X"09",X"03",X"00",X"93",X"FE",X"40",X"A1",X"99",X"38",
		X"80",X"91",X"22",X"AA",X"5F",X"93",X"08",X"0C",X"13",X"A0",X"0A",X"22",X"18",X"B3",X"F9",X"39",
		X"3B",X"F2",X"3A",X"89",X"04",X"00",X"98",X"0F",X"01",X"83",X"AF",X"22",X"A0",X"89",X"40",X"08",
		X"98",X"F1",X"18",X"2A",X"D3",X"2A",X"09",X"85",X"08",X"89",X"2F",X"82",X"81",X"8E",X"13",X"98",
		X"0A",X"31",X"00",X"92",X"FB",X"40",X"08",X"E1",X"39",X"88",X"82",X"10",X"0B",X"3F",X"C5",X"09",
		X"09",X"94",X"89",X"19",X"83",X"18",X"98",X"8F",X"12",X"A2",X"9F",X"22",X"98",X"89",X"50",X"80",
		X"B3",X"CD",X"40",X"91",X"8C",X"31",X"A1",X"99",X"42",X"8A",X"95",X"DB",X"50",X"91",X"A9",X"31",
		X"A0",X"90",X"41",X"0A",X"A5",X"CD",X"31",X"91",X"9B",X"41",X"A1",X"A8",X"51",X"0A",X"A4",X"BF",
		X"30",X"91",X"8C",X"22",X"90",X"99",X"42",X"89",X"A1",X"6F",X"92",X"00",X"0C",X"03",X"09",X"89",
		X"13",X"01",X"BB",X"7A",X"F2",X"19",X"18",X"C2",X"28",X"8A",X"94",X"10",X"0B",X"94",X"BF",X"30",
		X"92",X"9C",X"23",X"80",X"BB",X"52",X"08",X"AA",X"32",X"FA",X"20",X"20",X"F8",X"32",X"9A",X"A2",
		X"32",X"0C",X"A1",X"7C",X"B2",X"20",X"0B",X"B6",X"18",X"8B",X"03",X"21",X"AC",X"83",X"1F",X"91",
		X"03",X"0F",X"82",X"28",X"8B",X"94",X"20",X"9A",X"85",X"BF",X"21",X"92",X"9D",X"23",X"98",X"9A",
		X"33",X"18",X"BE",X"12",X"1C",X"B1",X"23",X"0E",X"A3",X"40",X"99",X"B8",X"52",X"89",X"92",X"9F",
		X"94",X"91",X"1F",X"03",X"09",X"99",X"14",X"00",X"BB",X"12",X"29",X"F8",X"12",X"19",X"D8",X"33",
		X"0A",X"BA",X"25",X"10",X"B8",X"5D",X"E2",X"28",X"88",X"B3",X"38",X"AA",X"A5",X"31",X"8D",X"B3",
		X"10",X"3F",X"B2",X"30",X"8B",X"C3",X"50",X"8A",X"99",X"23",X"19",X"A9",X"5A",X"F8",X"49",X"10",
		X"D0",X"48",X"88",X"B1",X"41",X"0A",X"D0",X"20",X"00",X"F8",X"38",X"00",X"C8",X"32",X"09",X"A8",
		X"80",X"30",X"98",X"87",X"BF",X"03",X"81",X"8E",X"03",X"08",X"8C",X"05",X"00",X"AB",X"12",X"08",
		X"1E",X"A4",X"00",X"0B",X"A4",X"20",X"8A",X"81",X"80",X"98",X"21",X"80",X"1F",X"F2",X"28",X"0C",
		X"A5",X"18",X"99",X"03",X"29",X"BA",X"02",X"08",X"39",X"FA",X"40",X"00",X"F8",X"31",X"19",X"A0",
		X"08",X"19",X"01",X"99",X"24",X"FF",X"30",X"82",X"D8",X"31",X"89",X"A8",X"51",X"8A",X"B8",X"40",
		X"90",X"2D",X"C3",X"10",X"2B",X"D1",X"31",X"0A",X"91",X"1A",X"01",X"12",X"BD",X"3E",X"F1",X"38",
		X"08",X"C1",X"48",X"08",X"C0",X"32",X"1C",X"C0",X"21",X"99",X"04",X"CB",X"22",X"11",X"BF",X"13",
		X"01",X"AA",X"02",X"09",X"80",X"1A",X"82",X"AF",X"F3",X"10",X"0C",X"94",X"29",X"09",X"B3",X"42",
		X"AD",X"91",X"10",X"9A",X"17",X"BD",X"21",X"02",X"AD",X"13",X"00",X"9B",X"12",X"00",X"89",X"1A",
		X"81",X"2B",X"FF",X"31",X"08",X"E0",X"31",X"08",X"88",X"2B",X"A3",X"09",X"8B",X"C3",X"0A",X"27",
		X"4B",X"F8",X"30",X"19",X"F0",X"31",X"89",X"B1",X"31",X"8A",X"99",X"10",X"9C",X"AA",X"27",X"08",
		X"99",X"26",X"0B",X"12",X"90",X"9B",X"03",X"8B",X"D9",X"54",X"18",X"FB",X"41",X"08",X"C9",X"33",
		X"09",X"C8",X"30",X"08",X"88",X"1B",X"85",X"9F",X"C4",X"01",X"8B",X"95",X"19",X"08",X"91",X"11",
		X"1A",X"B9",X"28",X"1C",X"B3",X"73",X"FB",X"21",X"12",X"CB",X"23",X"82",X"9C",X"02",X"81",X"88",
		X"19",X"09",X"A1",X"3F",X"F2",X"10",X"0C",X"A5",X"28",X"80",X"99",X"00",X"22",X"8D",X"A0",X"10",
		X"AA",X"37",X"4F",X"A2",X"11",X"0B",X"B2",X"31",X"1A",X"B9",X"31",X"28",X"98",X"10",X"1B",X"F8",
		X"4E",X"A4",X"08",X"2A",X"B3",X"38",X"03",X"8D",X"98",X"12",X"58",X"C9",X"81",X"89",X"88",X"73",
		X"FB",X"22",X"11",X"BB",X"83",X"42",X"9D",X"91",X"12",X"8A",X"10",X"98",X"B9",X"81",X"78",X"F9",
		X"22",X"10",X"D9",X"21",X"32",X"9D",X"A8",X"32",X"08",X"A9",X"00",X"9A",X"C0",X"63",X"3F",X"E1",
		X"20",X"19",X"C0",X"03",X"28",X"CA",X"03",X"39",X"99",X"92",X"0B",X"BA",X"24",X"34",X"FF",X"12",
		X"01",X"AA",X"82",X"32",X"8C",X"B0",X"41",X"8A",X"90",X"00",X"9B",X"A8",X"33",X"52",X"EF",X"12",
		X"01",X"9C",X"82",X"32",X"9E",X"91",X"31",X"9B",X"80",X"10",X"9D",X"80",X"42",X"0B",X"F8",X"23",
		X"19",X"C9",X"05",X"20",X"BB",X"83",X"40",X"CA",X"82",X"00",X"BB",X"A2",X"71",X"09",X"E9",X"32",
		X"18",X"BB",X"26",X"11",X"CA",X"84",X"30",X"BF",X"82",X"19",X"99",X"81",X"23",X"9D",X"98",X"43",
		X"8D",X"80",X"34",X"0D",X"A1",X"33",X"8C",X"D0",X"21",X"89",X"C8",X"02",X"30",X"C8",X"82",X"18",
		X"88",X"93",X"52",X"EA",X"84",X"38",X"BC",X"A2",X"20",X"8E",X"82",X"02",X"80",X"9A",X"83",X"28",
		X"B9",X"36",X"1D",X"A0",X"43",X"AB",X"88",X"10",X"98",X"B8",X"00",X"30",X"8C",X"00",X"30",X"8A",
		X"94",X"51",X"DA",X"03",X"49",X"BA",X"01",X"19",X"B8",X"08",X"19",X"40",X"09",X"98",X"88",X"38",
		X"08",X"48",X"BC",X"34",X"28",X"C9",X"82",X"98",X"89",X"89",X"12",X"80",X"18",X"9A",X"83",X"80",
		X"80",X"30",X"CB",X"86",X"28",X"9B",X"08",X"4B",X"A0",X"A1",X"81",X"10",X"81",X"08",X"B9",X"03",
		X"08",X"81",X"2B",X"A8",X"06",X"89",X"88",X"82",X"98",X"80",X"80",X"A9",X"32",X"1A",X"90",X"C1",
		X"02",X"80",X"84",X"BB",X"91",X"33",X"0A",X"88",X"91",X"88",X"80",X"80",X"C1",X"24",X"8B",X"A8",
		X"92",X"10",X"80",X"82",X"89",X"A8",X"24",X"89",X"98",X"84",X"89",X"A0",X"80",X"80",X"00",X"99",
		X"A0",X"10",X"88",X"83",X"00",X"88",X"80",X"12",X"89",X"88",X"91",X"2A",X"90",X"82",X"89",X"80",
		X"80",X"8A",X"90",X"82",X"10",X"80",X"81",X"88",X"12",X"A2",X"B3",X"89",X"91",X"88",X"90",X"81",
		X"80",X"9A",X"22",X"AB",X"B0",X"31",X"1A",X"02",X"80",X"81",X"02",X"A8",X"81",X"88",X"90",X"81",
		X"90",X"80",X"81",X"90",X"80",X"08",X"B8",X"84",X"80",X"80",X"80",X"81",X"00",X"80",X"82",X"A8",
		X"80",X"09",X"80",X"80",X"80",X"80",X"80",X"C0",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",
		X"19",X"00",X"80",X"08",X"28",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",
		X"08",X"01",X"98",X"09",X"1A",X"22",X"B4",X"B1",X"19",X"1D",X"AC",X"F0",X"1C",X"80",X"A9",X"90",
		X"10",X"52",X"03",X"49",X"60",X"12",X"A6",X"0A",X"20",X"93",X"1C",X"20",X"B5",X"80",X"0F",X"1A",
		X"80",X"C3",X"9C",X"3B",X"00",X"00",X"69",X"11",X"B1",X"0A",X"89",X"A9",X"BB",X"CA",X"E9",X"18",
		X"2B",X"6E",X"11",X"A5",X"A9",X"3A",X"90",X"84",X"33",X"17",X"01",X"02",X"9A",X"DB",X"AB",X"EA",
		X"A8",X"83",X"74",X"41",X"30",X"81",X"D9",X"AF",X"8B",X"A1",X"85",X"31",X"51",X"11",X"9C",X"CD",
		X"A9",X"83",X"35",X"32",X"20",X"DD",X"BA",X"80",X"24",X"33",X"12",X"1F",X"AC",X"A8",X"02",X"43",
		X"35",X"0B",X"FA",X"98",X"11",X"33",X"32",X"0F",X"CA",X"80",X"12",X"41",X"30",X"DB",X"BA",X"11",
		X"34",X"35",X"0C",X"AD",X"90",X"12",X"21",X"50",X"BB",X"C9",X"00",X"33",X"17",X"0B",X"AB",X"A0",
		X"14",X"12",X"50",X"C9",X"C8",X"81",X"21",X"34",X"8B",X"BE",X"88",X"12",X"14",X"38",X"BC",X"C9",
		X"81",X"32",X"44",X"9A",X"BC",X"99",X"22",X"25",X"39",X"9B",X"D8",X"A1",X"13",X"31",X"0A",X"8A",
		X"B9",X"92",X"30",X"00",X"83",X"B3",X"A8",X"80",X"88",X"88",X"12",X"92",X"9B",X"9A",X"B2",X"96",
		X"89",X"19",X"82",X"D0",X"AA",X"58",X"81",X"98",X"9A",X"0E",X"12",X"83",X"10",X"2B",X"0B",X"C2",
		X"80",X"51",X"28",X"9A",X"BA",X"08",X"21",X"43",X"88",X"9B",X"98",X"80",X"80",X"12",X"82",X"90",
		X"98",X"09",X"98",X"89",X"10",X"12",X"12",X"88",X"A8",X"B8",X"80",X"80",X"80",X"08",X"80",X"82",
		X"11",X"00",X"98",X"B8",X"A9",X"81",X"81",X"10",X"8A",X"81",X"82",X"01",X"10",X"80",X"B8",X"80",
		X"80",X"80",X"89",X"98",X"80",X"81",X"20",X"80",X"89",X"90",X"81",X"10",X"80",X"80",X"A8",X"81",
		X"10",X"80",X"80",X"80",X"A2",X"80",X"81",X"88",X"80",X"89",X"82",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"91",X"90",X"80",X"80",
		X"08",X"19",X"3B",X"08",X"80",X"80",X"80",X"08",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"91",X"90",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"67",X"E3",X"00",X"08",X"00",X"20",X"00",X"00",X"00",X"60",X"FF",X"FF",X"00",X"20",X"00",
		X"20",X"00",X"60",X"FF",X"FF",X"00",X"20",X"00",X"40",X"00",X"60",X"FF",X"FF",X"00",X"20",X"00",
		X"60",X"00",X"60",X"FF",X"FF",X"00",X"20",X"00",X"80",X"00",X"60",X"FF",X"FF",X"00",X"20",X"00",
		X"A0",X"00",X"60",X"FF",X"FF",X"00",X"20",X"00",X"C0",X"00",X"60",X"FF",X"FF",X"00",X"00",X"00",
		X"1E",X"49",X"00",X"30",X"C0",X"00",X"20",X"00",X"20",X"00",X"60",X"3D",X"E0",X"00",X"E0",X"FF",
		X"FF",X"07",X"00",X"E0",X"00",X"00",X"00",X"00",X"94",X"03",X"05",X"00",X"00",X"3E",X"81",X"32",
		X"00",X"F6",X"3A",X"00",X"F6",X"FE",X"00",X"CA",X"74",X"E0",X"FE",X"01",X"CA",X"74",X"E0",X"FE",
		X"09",X"C2",X"62",X"E0",X"00",X"3E",X"81",X"32",X"00",X"F8",X"3A",X"00",X"F8",X"FE",X"00",X"CA",
		X"8C",X"E0",X"FE",X"01",X"CA",X"8C",X"E0",X"FE",X"09",X"C2",X"7A",X"E0",X"00",X"3E",X"81",X"32",
		X"00",X"FE",X"3A",X"00",X"FE",X"FE",X"00",X"CA",X"A4",X"E0",X"FE",X"01",X"CA",X"A4",X"E0",X"FE",
		X"09",X"C2",X"92",X"E0",X"00",X"3E",X"82",X"32",X"00",X"FA",X"3A",X"00",X"FA",X"FE",X"00",X"CA",
		X"BC",X"E0",X"FE",X"01",X"CA",X"BC",X"E0",X"FE",X"09",X"C2",X"AA",X"E0",X"00",X"18",X"FE",X"3E",
		X"FE",X"32",X"01",X"F8",X"3E",X"01",X"32",X"02",X"F8",X"3E",X"80",X"32",X"00",X"F8",X"3A",X"00",
		X"F8",X"FE",X"00",X"CA",X"E0",X"E0",X"FE",X"01",X"CA",X"E0",X"E0",X"FE",X"09",X"C2",X"CE",X"E0",
		X"00",X"3A",X"04",X"F8",X"C9",X"3E",X"FE",X"32",X"01",X"F8",X"3E",X"F0",X"32",X"02",X"F8",X"3E",
		X"80",X"32",X"00",X"F8",X"3A",X"00",X"F8",X"FE",X"00",X"CA",X"06",X"E1",X"FE",X"01",X"CA",X"06",
		X"E1",X"FE",X"09",X"C2",X"F4",X"E0",X"00",X"21",X"03",X"F8",X"7E",X"A7",X"4F",X"06",X"00",X"11",
		X"01",X"F6",X"23",X"12",X"13",X"28",X"02",X"ED",X"B0",X"36",X"0D",X"EB",X"36",X"20",X"C9",X"18",
		X"1D",X"4E",X"3E",X"84",X"32",X"00",X"FE",X"3A",X"00",X"FE",X"FE",X"00",X"CA",X"39",X"E1",X"FE",
		X"01",X"CA",X"39",X"E1",X"FE",X"09",X"C2",X"27",X"E1",X"00",X"FE",X"09",X"28",X"E4",X"3A",X"01",
		X"FE",X"0F",X"30",X"DE",X"79",X"32",X"01",X"FE",X"3E",X"86",X"32",X"00",X"FE",X"3A",X"00",X"FE",
		X"FE",X"00",X"CA",X"5F",X"E1",X"FE",X"01",X"CA",X"5F",X"E1",X"FE",X"09",X"C2",X"4D",X"E1",X"00",
		X"23",X"10",X"BE",X"C9",X"DB",X"04",X"E6",X"80",X"32",X"7F",X"FF",X"C9",X"21",X"8B",X"FF",X"7E",
		X"A7",X"C8",X"23",X"CD",X"E3",X"E1",X"18",X"F7",X"7C",X"CD",X"7D",X"E1",X"7D",X"F5",X"0F",X"0F",
		X"0F",X"0F",X"CD",X"86",X"E1",X"F1",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"07",X"C6",X"30",
		X"18",X"51",X"06",X"01",X"3E",X"20",X"CD",X"E3",X"E1",X"10",X"F9",X"C9",X"3A",X"7F",X"FF",X"A7",
		X"C8",X"3E",X"84",X"32",X"00",X"FE",X"3A",X"00",X"FE",X"FE",X"00",X"CA",X"B8",X"E1",X"FE",X"01",
		X"CA",X"B8",X"E1",X"FE",X"09",X"C2",X"A6",X"E1",X"00",X"FE",X"09",X"28",X"E4",X"3A",X"01",X"FE",
		X"0F",X"30",X"DE",X"3E",X"0C",X"32",X"01",X"FE",X"3E",X"86",X"32",X"00",X"FE",X"3A",X"00",X"FE",
		X"FE",X"00",X"CA",X"DF",X"E1",X"FE",X"01",X"CA",X"DF",X"E1",X"FE",X"09",X"C2",X"CD",X"E1",X"00",
		X"C9",X"3E",X"0D",X"CD",X"49",X"E2",X"FE",X"0D",X"C0",X"D9",X"79",X"A7",X"20",X"0A",X"36",X"20",
		X"0C",X"DD",X"34",X"00",X"23",X"36",X"0D",X"3C",X"0F",X"30",X"09",X"36",X"20",X"0C",X"DD",X"34",
		X"00",X"23",X"36",X"0D",X"79",X"32",X"01",X"F6",X"3E",X"82",X"32",X"00",X"F6",X"3A",X"00",X"F6",
		X"FE",X"00",X"CA",X"1F",X"E2",X"FE",X"01",X"CA",X"1F",X"E2",X"FE",X"09",X"C2",X"0D",X"E2",X"00",
		X"DD",X"36",X"00",X"00",X"21",X"7C",X"FF",X"34",X"7E",X"FE",X"12",X"38",X"02",X"36",X"12",X"3A",
		X"7F",X"FF",X"A7",X"D9",X"C8",X"D9",X"23",X"34",X"7E",X"FE",X"3D",X"38",X"02",X"36",X"3D",X"21",
		X"02",X"F6",X"41",X"04",X"CD",X"21",X"E1",X"D9",X"C9",X"D9",X"DD",X"21",X"01",X"F6",X"21",X"02",
		X"F6",X"DD",X"4E",X"00",X"06",X"00",X"09",X"77",X"DD",X"34",X"00",X"D9",X"C9",X"11",X"01",X"01",
		X"CD",X"B3",X"E2",X"06",X"5A",X"21",X"7B",X"E2",X"C5",X"CD",X"8E",X"E2",X"C1",X"10",X"F6",X"C9",
		X"11",X"03",X"01",X"CD",X"B3",X"E2",X"06",X"50",X"C3",X"65",X"E2",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"CD",X"B3",X"E2",X"01",X"10",
		X"00",X"79",X"32",X"01",X"F6",X"11",X"02",X"F6",X"ED",X"B0",X"3E",X"84",X"32",X"00",X"F6",X"3A",
		X"00",X"F6",X"FE",X"00",X"CA",X"B1",X"E2",X"FE",X"01",X"CA",X"B1",X"E2",X"FE",X"09",X"C2",X"9F",
		X"E2",X"00",X"C9",X"7B",X"32",X"01",X"F6",X"7A",X"32",X"02",X"F6",X"3E",X"83",X"32",X"00",X"F6",
		X"3A",X"00",X"F6",X"FE",X"00",X"CA",X"D2",X"E2",X"FE",X"01",X"CA",X"D2",X"E2",X"FE",X"09",X"C2",
		X"C0",X"E2",X"00",X"C9",X"3E",X"7F",X"32",X"02",X"F6",X"3E",X"01",X"32",X"01",X"F6",X"3E",X"84",
		X"32",X"00",X"F6",X"3A",X"00",X"F6",X"FE",X"00",X"CA",X"F5",X"E2",X"FE",X"01",X"CA",X"F5",X"E2",
		X"FE",X"09",X"C2",X"E3",X"E2",X"00",X"C9",X"06",X"00",X"00",X"10",X"FD",X"0D",X"20",X"F8",X"C9",
		X"D6",X"30",X"D8",X"FE",X"0A",X"3F",X"D0",X"FE",X"11",X"D8",X"FE",X"17",X"3F",X"D8",X"D6",X"07",
		X"C9",X"EB",X"36",X"00",X"23",X"36",X"00",X"2B",X"1A",X"CD",X"00",X"E3",X"38",X"09",X"ED",X"6F",
		X"23",X"ED",X"6F",X"2B",X"13",X"18",X"F1",X"23",X"23",X"EB",X"7E",X"FE",X"0D",X"C8",X"FE",X"30",
		X"C9",X"78",X"A7",X"C8",X"D5",X"C5",X"11",X"02",X"FA",X"7E",X"12",X"23",X"13",X"10",X"FA",X"C1",
		X"48",X"CB",X"39",X"30",X"04",X"0C",X"3E",X"20",X"12",X"79",X"32",X"01",X"FA",X"3E",X"89",X"32",
		X"00",X"FA",X"3A",X"00",X"FA",X"FE",X"00",X"CA",X"64",X"E3",X"FE",X"01",X"CA",X"64",X"E3",X"FE",
		X"09",X"C2",X"52",X"E3",X"00",X"D1",X"C9",X"31",X"00",X"F6",X"3E",X"80",X"32",X"00",X"F6",X"3A",
		X"00",X"F6",X"FE",X"00",X"CA",X"81",X"E3",X"FE",X"01",X"CA",X"81",X"E3",X"FE",X"09",X"C2",X"6F",
		X"E3",X"00",X"3E",X"80",X"32",X"00",X"FE",X"3A",X"00",X"FE",X"FE",X"00",X"CA",X"99",X"E3",X"FE",
		X"01",X"CA",X"99",X"E3",X"FE",X"09",X"C2",X"87",X"E3",X"00",X"AF",X"32",X"03",X"FE",X"3E",X"40",
		X"32",X"01",X"FE",X"3E",X"4E",X"32",X"02",X"FE",X"3E",X"82",X"32",X"00",X"FE",X"3A",X"00",X"FE",
		X"FE",X"00",X"CA",X"BF",X"E3",X"FE",X"01",X"CA",X"BF",X"E3",X"FE",X"09",X"C2",X"AD",X"E3",X"00",
		X"3E",X"15",X"32",X"01",X"FE",X"3E",X"83",X"32",X"00",X"FE",X"3A",X"00",X"FE",X"FE",X"00",X"CA",
		X"DC",X"E3",X"FE",X"01",X"CA",X"DC",X"E3",X"FE",X"09",X"C2",X"CA",X"E3",X"00",X"21",X"1F",X"E1",
		X"06",X"02",X"CD",X"21",X"E1",X"AF",X"32",X"7C",X"FF",X"32",X"7D",X"FF",X"CD",X"7C",X"E8",X"CD",
		X"F8",X"E3",X"AF",X"32",X"7F",X"FF",X"18",X"F7",X"21",X"80",X"E5",X"AF",X"32",X"03",X"E0",X"32",
		X"7F",X"FF",X"32",X"01",X"F6",X"CD",X"6F",X"E1",X"CD",X"E5",X"E0",X"3A",X"04",X"F8",X"FE",X"0D",
		X"28",X"E6",X"21",X"BD",X"E4",X"CD",X"19",X"E5",X"A7",X"28",X"11",X"FE",X"7F",X"CA",X"9F",X"E4",
		X"21",X"5C",X"E5",X"AF",X"32",X"01",X"F6",X"CD",X"6F",X"E1",X"18",X"CC",X"EB",X"21",X"79",X"E4",
		X"E5",X"21",X"47",X"E4",X"79",X"FE",X"09",X"D2",X"76",X"E4",X"3D",X"07",X"85",X"6F",X"3E",X"00",
		X"8C",X"67",X"7E",X"23",X"66",X"6F",X"E9",X"6A",X"E4",X"6A",X"E4",X"76",X"E4",X"76",X"E4",X"57",
		X"E4",X"57",X"E4",X"57",X"E4",X"57",X"E4",X"EB",X"7E",X"FE",X"54",X"28",X"03",X"FE",X"49",X"C0",
		X"7E",X"32",X"41",X"E0",X"23",X"7E",X"FE",X"2C",X"23",X"C9",X"EB",X"7E",X"FE",X"34",X"CA",X"60",
		X"E4",X"FE",X"32",X"C0",X"18",X"EA",X"AF",X"EB",X"C9",X"20",X"17",X"79",X"32",X"04",X"E0",X"E5",
		X"06",X"00",X"11",X"05",X"E0",X"CD",X"11",X"E3",X"28",X"1B",X"30",X"0C",X"04",X"F1",X"23",X"E5",
		X"18",X"F3",X"21",X"6D",X"E5",X"C3",X"23",X"E4",X"E1",X"21",X"4B",X"E5",X"C3",X"23",X"E4",X"79",
		X"32",X"04",X"E0",X"18",X"06",X"04",X"F1",X"78",X"32",X"03",X"E0",X"E5",X"3A",X"04",X"E0",X"07",
		X"5F",X"16",X"00",X"21",X"FB",X"E4",X"19",X"EB",X"CD",X"14",X"E6",X"D1",X"E9",X"52",X"00",X"42",
		X"50",X"57",X"00",X"42",X"50",X"52",X"00",X"32",X"4B",X"57",X"00",X"32",X"4B",X"52",X"00",X"34",
		X"4B",X"57",X"00",X"34",X"4B",X"52",X"00",X"38",X"4B",X"57",X"00",X"38",X"4B",X"52",X"00",X"44",
		X"55",X"4D",X"50",X"00",X"50",X"44",X"55",X"4D",X"50",X"00",X"54",X"52",X"41",X"53",X"00",X"50",
		X"55",X"54",X"00",X"45",X"44",X"49",X"54",X"00",X"3F",X"00",X"FF",X"5D",X"E0",X"FD",X"EB",X"8E",
		X"EB",X"FD",X"EB",X"8E",X"EB",X"FD",X"EB",X"8E",X"EB",X"FD",X"EB",X"8E",X"EB",X"3F",X"F3",X"28",
		X"F3",X"D7",X"F2",X"D0",X"F1",X"23",X"EE",X"D9",X"ED",X"0E",X"00",X"11",X"04",X"F8",X"7E",X"FE",
		X"FF",X"28",X"18",X"A7",X"28",X"15",X"47",X"1A",X"B8",X"20",X"04",X"13",X"23",X"18",X"EF",X"23",
		X"7E",X"FE",X"FF",X"C8",X"A7",X"20",X"F8",X"23",X"0C",X"18",X"E0",X"1A",X"FE",X"2C",X"28",X"07",
		X"FE",X"0D",X"20",X"EC",X"3E",X"7F",X"C9",X"AF",X"13",X"EB",X"C9",X"2A",X"20",X"4E",X"55",X"4D",
		X"45",X"52",X"49",X"43",X"20",X"65",X"72",X"72",X"6F",X"72",X"0D",X"00",X"2A",X"20",X"43",X"4F",
		X"4D",X"4D",X"41",X"4E",X"44",X"20",X"65",X"72",X"72",X"6F",X"72",X"0D",X"00",X"2A",X"20",X"50",
		X"41",X"52",X"41",X"4D",X"45",X"54",X"45",X"52",X"20",X"65",X"72",X"72",X"6F",X"72",X"0D",X"00",
		X"0D",X"2A",X"20",X"49",X"4E",X"50",X"55",X"54",X"20",X"43",X"4F",X"4D",X"4D",X"41",X"4E",X"44",
		X"0D",X"00",X"0D",X"2A",X"4E",X"6F",X"2D",X"65",X"72",X"61",X"73",X"65",X"20",X"72",X"6F",X"6D",
		X"20",X"3D",X"20",X"00",X"0D",X"2A",X"45",X"72",X"61",X"73",X"65",X"20",X"72",X"6F",X"6D",X"0D",
		X"00",X"20",X"52",X"4F",X"4D",X"20",X"20",X"44",X"41",X"54",X"41",X"20",X"20",X"43",X"4D",X"50",
		X"20",X"20",X"44",X"41",X"54",X"41",X"20",X"20",X"20",X"20",X"52",X"4F",X"4D",X"20",X"4E",X"4F",
		X"2E",X"3D",X"00",X"52",X"4F",X"4D",X"20",X"4E",X"4F",X"2E",X"3D",X"00",X"20",X"20",X"20",X"45",
		X"72",X"72",X"6F",X"72",X"73",X"3D",X"00",X"20",X"43",X"68",X"65",X"63",X"6B",X"2D",X"73",X"75",
		X"6D",X"3D",X"00",X"20",X"20",X"20",X"42",X"6C",X"61",X"6E",X"6B",X"0D",X"00",X"7C",X"BA",X"C0",
		X"7D",X"BB",X"C9",X"A7",X"ED",X"52",X"23",X"C9",X"23",X"7C",X"B5",X"2B",X"C9",X"7D",X"02",X"03",
		X"7C",X"02",X"03",X"C9",X"1A",X"6F",X"13",X"1A",X"67",X"C9",X"CD",X"39",X"E6",X"21",X"00",X"00",
		X"22",X"4D",X"E0",X"7D",X"32",X"3F",X"E0",X"2A",X"05",X"E0",X"22",X"49",X"E0",X"22",X"4F",X"E0",
		X"3A",X"03",X"E0",X"A7",X"C0",X"F1",X"3E",X"01",X"C9",X"21",X"40",X"E0",X"3A",X"04",X"E0",X"FE",
		X"07",X"36",X"00",X"38",X"02",X"36",X"10",X"3D",X"CB",X"3F",X"28",X"05",X"07",X"C6",X"02",X"18",
		X"0B",X"5F",X"3A",X"41",X"E0",X"FE",X"34",X"20",X"01",X"1C",X"7B",X"07",X"21",X"6B",X"E6",X"5F",
		X"16",X"00",X"19",X"7E",X"23",X"66",X"6F",X"22",X"45",X"E0",X"C9",X"20",X"00",X"00",X"02",X"00",
		X"08",X"00",X"10",X"00",X"20",X"CD",X"7B",X"E6",X"C3",X"00",X"E7",X"CD",X"1A",X"E6",X"FE",X"01",
		X"20",X"23",X"2A",X"49",X"E0",X"11",X"00",X"E0",X"CD",X"FD",X"E5",X"38",X"07",X"21",X"FF",X"FF",
		X"22",X"49",X"E0",X"23",X"EB",X"2A",X"45",X"E0",X"22",X"47",X"E0",X"2B",X"19",X"22",X"4B",X"E0",
		X"3E",X"01",X"D8",X"AF",X"C9",X"FE",X"02",X"20",X"21",X"EB",X"2A",X"07",X"E0",X"22",X"4B",X"E0",
		X"CD",X"03",X"E6",X"38",X"EB",X"22",X"47",X"E0",X"EB",X"2A",X"45",X"E0",X"1B",X"CD",X"FD",X"E5",
		X"3E",X"00",X"30",X"01",X"3C",X"32",X"3F",X"E0",X"AF",X"C9",X"EB",X"2A",X"07",X"E0",X"22",X"4B",
		X"E0",X"CD",X"03",X"E6",X"38",X"CA",X"22",X"47",X"E0",X"2A",X"09",X"E0",X"22",X"4D",X"E0",X"EB",
		X"2A",X"45",X"E0",X"2B",X"CD",X"FD",X"E5",X"3E",X"01",X"38",X"DA",X"2A",X"47",X"E0",X"19",X"EB",
		X"2A",X"45",X"E0",X"CD",X"FD",X"E5",X"3E",X"00",X"30",X"CB",X"3C",X"18",X"C8",X"CD",X"D0",X"E7",
		X"A7",X"C0",X"21",X"05",X"E0",X"06",X"3A",X"36",X"00",X"23",X"10",X"FB",X"3A",X"3F",X"E0",X"A7",
		X"28",X"2A",X"3A",X"04",X"E0",X"FE",X"05",X"3E",X"00",X"30",X"5B",X"ED",X"5B",X"45",X"E0",X"2A",
		X"47",X"E0",X"2B",X"CD",X"FD",X"E5",X"D2",X"37",X"E8",X"44",X"4D",X"2A",X"4D",X"E0",X"09",X"DA",
		X"A0",X"E6",X"CD",X"FD",X"E5",X"3E",X"01",X"D0",X"AF",X"32",X"3F",X"E0",X"3A",X"04",X"E0",X"FE",
		X"05",X"21",X"56",X"E0",X"3E",X"01",X"38",X"02",X"3E",X"07",X"77",X"01",X"05",X"E0",X"2A",X"47",
		X"E0",X"CD",X"0D",X"E6",X"2A",X"4D",X"E0",X"CD",X"0D",X"E6",X"EB",X"2A",X"45",X"E0",X"19",X"22",
		X"4D",X"E0",X"2A",X"49",X"E0",X"CD",X"0D",X"E6",X"2A",X"4F",X"E0",X"CD",X"0D",X"E6",X"21",X"56",
		X"E0",X"35",X"20",X"DA",X"AF",X"C9",X"01",X"05",X"E0",X"ED",X"5B",X"45",X"E0",X"2A",X"4D",X"E0",
		X"00",X"00",X"00",X"01",X"80",X"00",X"01",X"70",X"81",X"70",X"0C",X"00",X"8D",X"70",X"05",X"40",
		X"92",X"B0",X"01",X"C8",X"94",X"78",X"09",X"90",X"9E",X"08",X"1F",X"FF",X"BE",X"08",X"0D",X"FF",
		X"CC",X"08",X"01",X"2F",X"9E",X"08",X"09",X"FF",X"CD",X"38",X"07",X"FF",X"D5",X"38",X"07",X"FF",
		X"DD",X"38",X"01",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"E8",X"10",X"E8",X"72",X"E8",X"28",X"E8",X"8F",
		X"E8",X"CF",X"E9",X"33",X"E9",X"C5",X"EC",X"8B",X"EC",X"8B",X"F1",X"06",X"F2",X"CC",X"E8",X"27",
		X"E8",X"27",X"E8",X"27",X"E8",X"27",X"E8",X"27",X"E8",X"27",X"E8",X"27",X"E8",X"27",X"E8",X"27",
		X"76",X"BC",X"51",X"00",X"52",X"36",X"53",X"00",X"51",X"00",X"52",X"38",X"53",X"00",X"58",X"0F",
		X"59",X"0F",X"10",X"25",X"C0",X"77",X"03",X"FF",X"76",X"A7",X"51",X"00",X"53",X"00",X"50",X"00",
		X"52",X"00",X"56",X"00",X"59",X"08",X"18",X"08",X"10",X"59",X"0B",X"18",X"0B",X"10",X"59",X"0C",
		X"18",X"0C",X"10",X"59",X"0E",X"18",X"0E",X"10",X"59",X"0F",X"18",X"0F",X"10",X"59",X"0D",X"18",
		X"0D",X"08",X"59",X"0B",X"18",X"0D",X"08",X"59",X"09",X"18",X"09",X"08",X"59",X"07",X"18",X"07",
		X"08",X"59",X"05",X"18",X"05",X"08",X"59",X"03",X"18",X"03",X"08",X"58",X"00",X"59",X"00",X"77",
		X"18",X"FF",X"76",X"BD",X"53",X"00",X"52",X"43",X"59",X"10",X"5B",X"00",X"5C",X"10",X"1D",X"09",
		X"20",X"52",X"53",X"59",X"10",X"1D",X"09",X"E0",X"52",X"00",X"59",X"00",X"77",X"02",X"FF",X"76",
		X"A7",X"50",X"00",X"51",X"00",X"52",X"00",X"53",X"00",X"56",X"0B",X"59",X"00",X"18",X"00",X"08",
		X"59",X"02",X"18",X"02",X"08",X"59",X"04",X"18",X"04",X"08",X"59",X"06",X"18",X"06",X"08",X"59",
		X"08",X"18",X"08",X"08",X"59",X"0A",X"18",X"0A",X"08",X"59",X"0C",X"18",X"0C",X"08",X"59",X"0E",
		X"18",X"0E",X"08",X"59",X"0F",X"18",X"0F",X"08",X"58",X"00",X"59",X"00",X"77",X"18",X"FF",X"76",
		X"BC",X"51",X"00",X"52",X"2B",X"53",X"00",X"59",X"08",X"18",X"08",X"08",X"59",X"0A",X"18",X"0A",
		X"08",X"59",X"0C",X"18",X"0C",X"08",X"59",X"0E",X"18",X"0E",X"08",X"59",X"0D",X"18",X"0D",X"08",
		X"59",X"0C",X"18",X"0C",X"08",X"59",X"0B",X"18",X"0B",X"08",X"59",X"0A",X"18",X"0A",X"08",X"59",
		X"09",X"18",X"09",X"08",X"59",X"08",X"18",X"08",X"08",X"59",X"07",X"18",X"07",X"08",X"59",X"06",
		X"18",X"06",X"08",X"59",X"05",X"18",X"05",X"08",X"59",X"04",X"18",X"04",X"08",X"59",X"03",X"18",
		X"03",X"08",X"59",X"02",X"18",X"02",X"08",X"59",X"01",X"18",X"01",X"08",X"58",X"00",X"59",X"00",
		X"77",X"03",X"FF",X"66",X"BC",X"41",X"00",X"43",X"00",X"42",X"9F",X"6C",X"14",X"6D",X"14",X"6E",
		X"14",X"68",X"0F",X"69",X"0F",X"00",X"BD",X"0C",X"00",X"00",X"18",X"68",X"0F",X"69",X"0F",X"00",
		X"BD",X"18",X"68",X"0F",X"69",X"0F",X"00",X"BD",X"18",X"68",X"0F",X"69",X"0F",X"00",X"BD",X"18",
		X"42",X"7E",X"68",X"0F",X"69",X"0F",X"00",X"9F",X"18",X"42",X"9F",X"68",X"0F",X"69",X"0F",X"00",
		X"BD",X"18",X"42",X"7E",X"68",X"0F",X"69",X"0F",X"00",X"9F",X"18",X"42",X"77",X"68",X"0F",X"69",
		X"0F",X"00",X"8E",X"0C",X"00",X"00",X"18",X"42",X"77",X"68",X"0F",X"69",X"0F",X"00",X"8E",X"18",
		X"68",X"0F",X"69",X"0F",X"00",X"8E",X"18",X"68",X"0F",X"69",X"0F",X"00",X"8E",X"18",X"42",X"5E",
		X"68",X"0F",X"69",X"0F",X"00",X"77",X"18",X"42",X"77",X"68",X"0F",X"69",X"0F",X"00",X"8E",X"18",
		X"42",X"5E",X"68",X"0F",X"69",X"0F",X"00",X"77",X"18",X"42",X"4F",X"68",X"0F",X"69",X"0F",X"00",
		X"5E",X"60",X"67",X"03",X"FF",X"66",X"BC",X"41",X"00",X"43",X"01",X"6C",X"14",X"6D",X"14",X"6E",
		X"14",X"42",X"65",X"68",X"0F",X"69",X"0F",X"00",X"B3",X"40",X"68",X"0F",X"69",X"0F",X"00",X"B3",
		X"20",X"68",X"0F",X"69",X"0F",X"00",X"77",X"40",X"68",X"0F",X"69",X"0F",X"00",X"77",X"20",X"42",
		X"DD",X"68",X"0F",X"69",X"0F",X"00",X"8E",X"40",X"68",X"0F",X"69",X"0F",X"00",X"8E",X"20",X"49",
		X"0F",X"68",X"0F",X"00",X"9F",X"20",X"68",X"0F",X"00",X"8E",X"20",X"49",X"00",X"68",X"0F",X"69",
		X"0F",X"00",X"9F",X"20",X"42",X"65",X"48",X"0F",X"49",X"0F",X"00",X"B3",X"60",X"00",X"B3",X"60",
		X"48",X"00",X"49",X"00",X"67",X"03",X"FF",X"66",X"8F",X"43",X"0E",X"45",X"0A",X"4B",X"02",X"4C",
		X"01",X"4D",X"09",X"49",X"10",X"4A",X"10",X"00",X"00",X"30",X"00",X"00",X"30",X"FE",X"EA",X"27",
		X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",
		X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",
		X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",
		X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"4A",X"10",X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",
		X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",
		X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",
		X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",
		X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",
		X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",
		X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",
		X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",
		X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"06",
		X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"1C",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"4A",X"10",X"06",X"01",X"1C",X"06",X"01",X"1C",X"FE",X"EC",X"8B",X"66",X"9F",X"4B",X"03",X"4C",
		X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",
		X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",
		X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",
		X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",
		X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",
		X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",
		X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",
		X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",X"4B",
		X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",
		X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",
		X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",
		X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",
		X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",
		X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",
		X"06",X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",
		X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",
		X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",
		X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",
		X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",
		X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",
		X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",
		X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",
		X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",
		X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",
		X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",
		X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",
		X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",
		X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",
		X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"06",X"01",X"1C",X"4B",X"03",
		X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",
		X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",X"4A",X"10",X"06",X"01",X"0E",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"0F",
		X"4A",X"10",X"06",X"01",X"0E",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"4A",X"10",X"06",X"01",X"0E",
		X"06",X"01",X"1C",X"FE",X"EC",X"8B",X"66",X"B8",X"41",X"00",X"43",X"00",X"45",X"01",X"6D",X"14",
		X"6C",X"14",X"6E",X"14",X"FE",X"F2",X"39",X"48",X"00",X"49",X"00",X"6A",X"00",X"04",X"00",X"24",
		X"40",X"9F",X"42",X"7E",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"45",X"02",X"04",X"7D",X"24",X"6A",
		X"00",X"04",X"00",X"24",X"40",X"8E",X"42",X"77",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"7D",
		X"24",X"6A",X"00",X"04",X"00",X"24",X"48",X"00",X"49",X"00",X"40",X"7E",X"42",X"6A",X"68",X"0F",
		X"69",X"0F",X"6A",X"0F",X"04",X"7D",X"24",X"40",X"6A",X"42",X"59",X"48",X"0F",X"49",X"0F",X"6A",
		X"00",X"04",X"00",X"24",X"6A",X"0F",X"04",X"7D",X"24",X"40",X"77",X"42",X"5E",X"48",X"0F",X"49",
		X"0F",X"6A",X"00",X"04",X"00",X"24",X"45",X"01",X"6A",X"0F",X"04",X"DD",X"24",X"6A",X"00",X"04",
		X"00",X"24",X"6A",X"0F",X"04",X"DD",X"24",X"6A",X"00",X"04",X"00",X"24",X"6A",X"0F",X"04",X"DD",
		X"24",X"48",X"00",X"49",X"00",X"6A",X"00",X"04",X"00",X"24",X"6A",X"0F",X"04",X"DD",X"24",X"FE",
		X"F2",X"39",X"48",X"00",X"49",X"00",X"6A",X"00",X"04",X"00",X"24",X"40",X"59",X"42",X"47",X"68",
		X"0F",X"69",X"0F",X"6A",X"0F",X"45",X"02",X"04",X"7D",X"24",X"40",X"5E",X"42",X"4F",X"68",X"0F",
		X"69",X"0F",X"6A",X"00",X"04",X"00",X"24",X"40",X"6A",X"42",X"59",X"68",X"0F",X"69",X"0F",X"6A",
		X"0F",X"04",X"7D",X"24",X"40",X"77",X"42",X"5E",X"68",X"0F",X"69",X"0F",X"6A",X"00",X"04",X"00",
		X"24",X"40",X"6A",X"42",X"59",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"7D",X"24",X"6A",X"00",
		X"04",X"00",X"24",X"40",X"7E",X"42",X"6A",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"7D",X"24",
		X"6A",X"00",X"04",X"00",X"24",X"40",X"8E",X"42",X"77",X"48",X"0F",X"49",X"0F",X"45",X"01",X"6A",
		X"0F",X"04",X"DD",X"24",X"6A",X"00",X"04",X"00",X"24",X"6A",X"0F",X"04",X"DD",X"24",X"6A",X"00",
		X"04",X"00",X"24",X"6A",X"0F",X"04",X"DD",X"24",X"6A",X"00",X"04",X"00",X"24",X"48",X"00",X"49",
		X"00",X"6A",X"00",X"04",X"00",X"24",X"67",X"07",X"FF",X"40",X"BD",X"42",X"9F",X"68",X"0F",X"69",
		X"0F",X"6A",X"00",X"04",X"00",X"24",X"40",X"8E",X"42",X"77",X"48",X"0F",X"49",X"0F",X"6A",X"0F",
		X"04",X"DD",X"24",X"6A",X"00",X"04",X"00",X"24",X"6A",X"0F",X"04",X"DD",X"24",X"48",X"00",X"49",
		X"00",X"40",X"BD",X"42",X"9F",X"68",X"0F",X"69",X"0F",X"6A",X"00",X"04",X"00",X"24",X"40",X"77",
		X"42",X"5E",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"DD",X"24",X"6A",X"00",X"04",X"00",X"24",
		X"6A",X"0F",X"04",X"DD",X"24",X"48",X"00",X"49",X"00",X"68",X"0F",X"69",X"0F",X"04",X"DD",X"24",
		X"40",X"6A",X"42",X"59",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"65",X"24",X"6A",X"00",X"04",
		X"00",X"24",X"40",X"77",X"42",X"5E",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"65",X"24",X"6A",
		X"00",X"04",X"00",X"24",X"40",X"B3",X"42",X"8E",X"48",X"0F",X"49",X"0F",X"6A",X"0F",X"04",X"65",
		X"24",X"6A",X"00",X"04",X"00",X"24",X"6A",X"0F",X"04",X"65",X"24",X"FD",X"66",X"BC",X"41",X"00",
		X"43",X"00",X"6C",X"14",X"6D",X"14",X"6E",X"14",X"42",X"9F",X"68",X"0F",X"69",X"0F",X"00",X"BD",
		X"1C",X"68",X"00",X"69",X"00",X"00",X"00",X"1C",X"42",X"BD",X"68",X"0F",X"69",X"0F",X"00",X"EE",
		X"1C",X"42",X"9F",X"68",X"0F",X"69",X"0F",X"00",X"BD",X"1C",X"42",X"7E",X"68",X"0F",X"69",X"0F",
		X"00",X"9F",X"1C",X"68",X"00",X"69",X"00",X"00",X"00",X"1C",X"42",X"9F",X"68",X"0F",X"69",X"0F",
		X"00",X"BD",X"1C",X"42",X"7E",X"68",X"0F",X"69",X"0F",X"00",X"9F",X"1C",X"42",X"6A",X"68",X"0F",
		X"69",X"0F",X"00",X"7E",X"C0",X"67",X"03",X"FF",X"CD",X"E1",X"E1",X"3E",X"01",X"32",X"7F",X"FF",
		X"CD",X"42",X"F3",X"C3",X"9C",X"E1",X"7E",X"E6",X"7F",X"FE",X"20",X"D0",X"3E",X"20",X"C9",X"CD",
		X"E1",X"E1",X"21",X"30",X"30",X"22",X"80",X"FF",X"CD",X"D6",X"F3",X"2A",X"E5",X"FF",X"3A",X"03",
		X"E0",X"A7",X"28",X"09",X"2A",X"05",X"E0",X"22",X"E5",X"FF",X"22",X"E7",X"FF",X"EB",X"21",X"FF",
		X"00",X"19",X"EB",X"3A",X"03",X"E0",X"FE",X"02",X"38",X"04",X"ED",X"5B",X"07",X"E0",X"ED",X"53",
		X"07",X"E0",X"11",X"8B",X"FF",X"E5",X"E5",X"3A",X"03",X"E0",X"FE",X"03",X"38",X"0C",X"2A",X"09",
		X"E0",X"E5",X"01",X"10",X"00",X"09",X"22",X"09",X"E0",X"E1",X"CD",X"05",X"F4",X"CD",X"34",X"F4",
		X"E1",X"06",X"10",X"4E",X"CD",X"1D",X"F4",X"23",X"10",X"F9",X"06",X"04",X"CD",X"C4",X"F3",X"E1",
		X"06",X"10",X"CD",X"36",X"F3",X"12",X"23",X"13",X"10",X"F8",X"E5",X"CD",X"CB",X"F3",X"CD",X"6C",
		X"E1",X"D1",X"2A",X"07",X"E0",X"A7",X"ED",X"52",X"EB",X"30",X"B7",X"22",X"E5",X"FF",X"C9",X"11",
		X"8B",X"FF",X"06",X"5A",X"3E",X"20",X"12",X"13",X"10",X"FC",X"C9",X"3A",X"7E",X"FF",X"3D",X"32",
		X"7E",X"FF",X"C0",X"CD",X"9C",X"E1",X"3E",X"3C",X"32",X"7E",X"FF",X"21",X"6E",X"FF",X"3A",X"80",
		X"FF",X"FE",X"39",X"28",X"14",X"3C",X"32",X"80",X"FF",X"77",X"3A",X"81",X"FF",X"2B",X"32",X"81",
		X"FF",X"77",X"21",X"5C",X"FF",X"CD",X"6F",X"E1",X"C9",X"3E",X"30",X"77",X"32",X"80",X"FF",X"3A",
		X"81",X"FF",X"3C",X"18",X"E8",X"D9",X"01",X"4B",X"00",X"11",X"8C",X"FF",X"21",X"8B",X"FF",X"3E",
		X"20",X"77",X"ED",X"B0",X"3E",X"0D",X"77",X"23",X"3E",X"00",X"77",X"D9",X"C9",X"13",X"79",X"1F",
		X"1F",X"1F",X"1F",X"CD",X"27",X"F4",X"79",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"07",X"C6",
		X"30",X"12",X"13",X"C9",X"13",X"CD",X"3D",X"F4",X"3E",X"2D",X"12",X"13",X"C9",X"4C",X"CD",X"1E",
		X"F4",X"4D",X"C3",X"1E",X"F4",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"F7",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"DF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"E6",X"E1",X"E6",X"E1",X"85",X"E1",
		X"E6",X"E1",X"0D",X"EB",X"4F",X"ED",X"00",X"01",X"E6",X"E1",X"76",X"E1",X"0B",X"E4",X"F2",X"E3",
		X"00",X"00",X"2A",X"20",X"49",X"4E",X"50",X"55",X"54",X"20",X"43",X"4F",X"4D",X"4D",X"41",X"4E",
		X"44",X"20",X"0D",X"73",X"3D",X"31",X"32",X"41",X"37",X"20",X"43",X"68",X"65",X"63",X"6B",X"2D",
		X"73",X"75",X"6D",X"3D",X"45",X"30",X"30",X"30",X"0D",X"20",X"39",X"31",X"20",X"36",X"39",X"20",
		X"30",X"38",X"20",X"46",X"39",X"20",X"31",X"31",X"20",X"20",X"20",X"20",X"7C",X"20",X"22",X"20",
		X"20",X"49",X"20",X"7C",X"20",X"30",X"20",X"20",X"69",X"20",X"79",X"20",X"20",X"20",X"0D",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"40",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"40",X"FF",X"00",
		X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"00",X"FF",X"80",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"0E",X"FE",X"F0",X"07",X"38",X"4B",X"57",X"2C",X"49",X"2C",X"30",X"0D",X"30",X"0D",X"30",X"2C",
		X"33",X"0D",X"46",X"2C",X"33",X"41",X"30",X"30",X"0D",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FD",X"00",X"FD",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"EE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"7F",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FB",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"EB",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"09",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"40",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"40",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"0F",X"8E",X"00",X"FF",X"BD",X"FC",X"18",X"86",X"BF",X"C6",X"07",X"BD",X"FC",X"5A",X"86",X"13",
		X"C6",X"0F",X"BD",X"FC",X"5A",X"BD",X"FC",X"2D",X"7F",X"20",X"00",X"0F",X"BD",X"FB",X"C8",X"96",
		X"BD",X"2B",X"07",X"BD",X"FE",X"63",X"86",X"FF",X"97",X"BD",X"0E",X"CE",X"00",X"00",X"DF",X"D2",
		X"96",X"80",X"26",X"0B",X"DE",X"84",X"D6",X"8C",X"BD",X"FD",X"5E",X"DF",X"84",X"97",X"80",X"7C",
		X"00",X"D3",X"96",X"81",X"26",X"0B",X"DE",X"86",X"D6",X"8D",X"BD",X"FD",X"5E",X"DF",X"86",X"97",
		X"81",X"7C",X"00",X"D3",X"96",X"82",X"26",X"0B",X"DE",X"88",X"D6",X"8E",X"BD",X"FD",X"5E",X"DF",
		X"88",X"97",X"82",X"7C",X"00",X"D3",X"96",X"83",X"26",X"0B",X"DE",X"8A",X"D6",X"8F",X"BD",X"FD",
		X"5E",X"DF",X"8A",X"97",X"83",X"96",X"A8",X"27",X"08",X"7F",X"00",X"A8",X"C6",X"08",X"BD",X"FC",
		X"BC",X"96",X"A9",X"27",X"08",X"7F",X"00",X"A9",X"C6",X"09",X"BD",X"FC",X"BC",X"96",X"AA",X"27",
		X"08",X"7F",X"00",X"AA",X"C6",X"0A",X"BD",X"FC",X"BC",X"96",X"AB",X"27",X"08",X"7F",X"00",X"AB",
		X"C6",X"18",X"BD",X"FC",X"D5",X"96",X"AC",X"27",X"08",X"7F",X"00",X"AC",X"C6",X"19",X"BD",X"FC",
		X"D5",X"96",X"AD",X"27",X"08",X"7F",X"00",X"AD",X"C6",X"1A",X"BD",X"FC",X"D5",X"96",X"BF",X"16",
		X"9A",X"D8",X"0F",X"97",X"D8",X"54",X"24",X"09",X"D6",X"CC",X"C1",X"03",X"26",X"03",X"5C",X"D7",
		X"BD",X"C6",X"0F",X"BD",X"FC",X"60",X"7E",X"FA",X"9B",X"96",X"C2",X"B7",X"08",X"01",X"96",X"C3",
		X"B7",X"08",X"02",X"7C",X"00",X"BE",X"96",X"C0",X"4C",X"97",X"C0",X"44",X"24",X"32",X"DE",X"C4",
		X"09",X"27",X"1E",X"DF",X"C4",X"DE",X"C8",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C2",X"DE",
		X"C6",X"09",X"27",X"15",X"DF",X"C6",X"DE",X"CA",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C3",
		X"3B",X"86",X"01",X"9A",X"BF",X"97",X"BF",X"20",X"E6",X"86",X"02",X"9A",X"BF",X"97",X"BF",X"3B",
		X"96",X"C8",X"81",X"20",X"25",X"09",X"DE",X"C8",X"A6",X"00",X"97",X"C2",X"08",X"DF",X"C8",X"96",
		X"CA",X"81",X"20",X"25",X"09",X"DE",X"CA",X"A6",X"00",X"97",X"C3",X"08",X"DF",X"CA",X"96",X"C0",
		X"84",X"0E",X"26",X"CC",X"7C",X"00",X"C1",X"3B",X"96",X"C1",X"27",X"3E",X"7A",X"00",X"C1",X"96",
		X"80",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"80",X"96",X"81",X"27",X"06",X"4C",X"27",X"03",
		X"7A",X"00",X"81",X"96",X"82",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"82",X"96",X"83",X"27",
		X"06",X"4C",X"27",X"03",X"7A",X"00",X"83",X"CE",X"00",X"06",X"A6",X"AD",X"27",X"09",X"4A",X"26",
		X"04",X"6C",X"A7",X"A6",X"B3",X"A7",X"AD",X"09",X"26",X"F0",X"39",X"B7",X"20",X"00",X"C6",X"0E",
		X"BD",X"FC",X"A2",X"84",X"3F",X"97",X"BD",X"3B",X"CE",X"FF",X"FF",X"DF",X"00",X"C6",X"4F",X"08",
		X"86",X"00",X"A7",X"80",X"08",X"5A",X"26",X"FA",X"86",X"13",X"97",X"D8",X"39",X"BD",X"FC",X"45",
		X"86",X"BF",X"97",X"BC",X"C6",X"FF",X"D7",X"82",X"D7",X"83",X"D7",X"B1",X"D7",X"B2",X"D7",X"B3",
		X"C6",X"17",X"7E",X"FC",X"60",X"86",X"BF",X"97",X"BB",X"C6",X"FF",X"D7",X"80",X"D7",X"81",X"D7",
		X"AE",X"D7",X"AF",X"D7",X"B0",X"C6",X"07",X"7E",X"FC",X"60",X"7C",X"00",X"BE",X"20",X"04",X"0F",
		X"7F",X"00",X"BE",X"37",X"36",X"C1",X"10",X"2A",X"19",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",
		X"08",X"D7",X"03",X"5C",X"32",X"97",X"02",X"96",X"BE",X"27",X"FC",X"D7",X"03",X"5A",X"D7",X"03",
		X"33",X"39",X"86",X"15",X"97",X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"10",X"20",X"E3",X"37",X"20",
		X"E4",X"37",X"86",X"15",X"97",X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"14",X"20",X"0D",X"C1",X"10",
		X"2A",X"EF",X"37",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"0C",X"4F",X"97",X"03",X"97",X"00",
		X"D7",X"03",X"96",X"02",X"5F",X"D7",X"03",X"5A",X"D7",X"00",X"33",X"39",X"0F",X"BD",X"FC",X"A2",
		X"C6",X"09",X"7F",X"00",X"BE",X"84",X"1F",X"81",X"10",X"2A",X"08",X"4A",X"81",X"07",X"2B",X"03",
		X"BD",X"FC",X"8E",X"0E",X"39",X"0F",X"BD",X"FC",X"91",X"C6",X"11",X"20",X"E5",X"17",X"84",X"0F",
		X"81",X"08",X"2A",X"08",X"A6",X"94",X"AB",X"98",X"A7",X"94",X"20",X"67",X"CB",X"38",X"DE",X"CE",
		X"A6",X"05",X"36",X"DE",X"D2",X"AB",X"94",X"A7",X"94",X"32",X"2B",X"0C",X"24",X"02",X"6C",X"98",
		X"BD",X"FC",X"5F",X"5C",X"A6",X"94",X"20",X"4B",X"25",X"F6",X"6A",X"98",X"20",X"F2",X"6F",X"8C",
		X"DE",X"CE",X"C1",X"A0",X"2B",X"02",X"08",X"08",X"08",X"08",X"08",X"C1",X"C0",X"2B",X"08",X"17",
		X"84",X"0F",X"81",X"08",X"2B",X"01",X"08",X"86",X"01",X"39",X"DF",X"CE",X"DE",X"D2",X"6A",X"90",
		X"27",X"DC",X"C1",X"A0",X"2A",X"10",X"C4",X"1F",X"A6",X"94",X"36",X"DE",X"CE",X"A6",X"03",X"BD",
		X"FC",X"5F",X"0E",X"32",X"08",X"39",X"C1",X"C0",X"2A",X"93",X"A6",X"90",X"44",X"A6",X"94",X"25",
		X"02",X"A6",X"98",X"C4",X"1F",X"BD",X"FC",X"5F",X"0E",X"DE",X"CE",X"A6",X"04",X"39",X"26",X"CA",
		X"DF",X"CE",X"E6",X"00",X"2A",X"03",X"7E",X"FE",X"15",X"C4",X"3F",X"C1",X"20",X"2A",X"11",X"A6",
		X"01",X"BD",X"FC",X"5F",X"0E",X"E6",X"00",X"08",X"08",X"58",X"2B",X"E4",X"A6",X"00",X"08",X"39",
		X"C4",X"1F",X"17",X"84",X"0F",X"26",X"31",X"A6",X"01",X"97",X"CF",X"A6",X"02",X"97",X"CE",X"BD",
		X"FE",X"56",X"DC",X"CE",X"04",X"DD",X"CE",X"E6",X"00",X"C4",X"1F",X"5C",X"5C",X"BD",X"FE",X"56",
		X"7C",X"00",X"CF",X"26",X"03",X"7C",X"00",X"CE",X"BD",X"FE",X"56",X"CB",X"07",X"86",X"09",X"BD",
		X"FC",X"60",X"0E",X"E6",X"00",X"08",X"20",X"BF",X"80",X"08",X"2B",X"29",X"DD",X"D0",X"84",X"03",
		X"C1",X"30",X"2B",X"02",X"8B",X"03",X"16",X"A6",X"01",X"CE",X"00",X"00",X"3A",X"D6",X"D0",X"C1",
		X"04",X"2A",X"0B",X"A6",X"B4",X"A7",X"AE",X"DE",X"CE",X"D6",X"D1",X"7E",X"FD",X"6F",X"A7",X"B4",
		X"DE",X"CE",X"7E",X"FD",X"75",X"4C",X"27",X"17",X"5C",X"C1",X"10",X"2A",X"09",X"96",X"BB",X"A4",
		X"01",X"97",X"BB",X"7E",X"FD",X"71",X"96",X"BC",X"A4",X"01",X"97",X"BC",X"7E",X"FD",X"71",X"C1",
		X"10",X"2A",X"09",X"96",X"BB",X"AA",X"01",X"97",X"BB",X"7E",X"FD",X"71",X"96",X"BC",X"AA",X"01",
		X"97",X"BC",X"7E",X"FD",X"71",X"C1",X"F0",X"2A",X"17",X"A6",X"01",X"EE",X"02",X"3C",X"DE",X"D2",
		X"E7",X"8C",X"4C",X"A7",X"90",X"32",X"A7",X"94",X"32",X"A7",X"98",X"DE",X"CE",X"86",X"01",X"39",
		X"5C",X"27",X"12",X"DE",X"D2",X"5C",X"26",X"10",X"DC",X"CE",X"A7",X"9C",X"E7",X"A0",X"DE",X"CE",
		X"EE",X"01",X"86",X"01",X"39",X"86",X"FF",X"39",X"A6",X"9C",X"E6",X"A0",X"DD",X"CE",X"DE",X"CE",
		X"08",X"08",X"08",X"86",X"01",X"39",X"96",X"CF",X"BD",X"FC",X"5F",X"5C",X"96",X"CE",X"BD",X"FC",
		X"60",X"5C",X"39",X"26",X"09",X"BD",X"FC",X"18",X"7F",X"00",X"D9",X"7E",X"FC",X"2D",X"81",X"10",
		X"2B",X"03",X"7E",X"FE",X"EB",X"81",X"03",X"2A",X"35",X"97",X"CC",X"96",X"D8",X"8A",X"01",X"16",
		X"C4",X"FE",X"D7",X"D8",X"C6",X"0F",X"BD",X"FC",X"60",X"86",X"05",X"7F",X"00",X"BE",X"D6",X"BE",
		X"27",X"FC",X"4A",X"26",X"F6",X"D6",X"CC",X"58",X"58",X"CE",X"E7",X"80",X"3A",X"3C",X"EE",X"00",
		X"DF",X"C8",X"38",X"EE",X"02",X"DF",X"C4",X"96",X"BF",X"84",X"02",X"97",X"BF",X"39",X"81",X"06",
		X"27",X"C7",X"81",X"09",X"27",X"C3",X"97",X"CD",X"96",X"D8",X"8A",X"02",X"16",X"C4",X"FD",X"D7",
		X"D8",X"C6",X"0F",X"BD",X"FC",X"60",X"86",X"05",X"7F",X"00",X"BE",X"D6",X"BE",X"27",X"FC",X"4A",
		X"26",X"F6",X"D6",X"CD",X"58",X"58",X"CE",X"E7",X"80",X"3A",X"3C",X"EE",X"00",X"DF",X"CA",X"38",
		X"EE",X"02",X"DF",X"C6",X"96",X"BF",X"84",X"01",X"97",X"BF",X"39",X"16",X"58",X"CE",X"E7",X"C8",
		X"3A",X"EE",X"00",X"81",X"15",X"2A",X"33",X"97",X"A6",X"DF",X"88",X"7F",X"00",X"82",X"7F",X"00",
		X"8E",X"C6",X"BC",X"DA",X"BC",X"D7",X"BC",X"39",X"DF",X"8A",X"97",X"A7",X"7F",X"00",X"83",X"7F",
		X"00",X"8F",X"86",X"98",X"9A",X"BC",X"97",X"BC",X"39",X"DF",X"86",X"97",X"A5",X"7F",X"00",X"81",
		X"7F",X"00",X"8D",X"86",X"80",X"9A",X"BB",X"97",X"BB",X"39",X"81",X"18",X"27",X"1F",X"81",X"20",
		X"27",X"26",X"3C",X"36",X"BD",X"FC",X"18",X"BD",X"FC",X"2D",X"32",X"38",X"97",X"A4",X"DF",X"84",
		X"7F",X"00",X"8C",X"7F",X"00",X"80",X"86",X"98",X"9A",X"BB",X"97",X"BB",X"39",X"D6",X"BA",X"54",
		X"25",X"FA",X"C6",X"01",X"D7",X"BA",X"20",X"C1",X"7F",X"00",X"BA",X"7E",X"FC",X"45",X"4D",X"50",
		X"20",X"4C",X"49",X"53",X"54",X"20",X"50",X"41",X"47",X"45",X"20",X"3D",X"20",X"FF",X"00",X"0D",
		X"0D",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"0B",X"00",X"FE",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FA",X"80",X"FA",X"80",X"FA",X"80",X"FA",X"80",X"FC",X"0B",X"FA",X"80",X"FB",X"59",X"FA",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
