library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  20479) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"C3",X"69",X"00",X"FF",X"FF",X"FF",X"C3",X"00",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"0E",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"1A",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"2D",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"E6",X"0A",X"AF",X"21",X"00",X"A8",X"06",X"08",X"77",
		X"23",X"10",X"FC",X"3E",X"9B",X"32",X"03",X"98",X"3A",X"01",X"98",X"CB",X"57",X"CA",X"01",X"04",
		X"21",X"00",X"88",X"11",X"00",X"8C",X"FD",X"21",X"8D",X"00",X"C3",X"3B",X"01",X"FD",X"21",X"94",
		X"00",X"C3",X"18",X"02",X"21",X"9A",X"00",X"C3",X"4B",X"02",X"52",X"41",X"4D",X"20",X"31",X"47",
		X"48",X"4A",X"4B",X"00",X"21",X"00",X"80",X"11",X"00",X"88",X"FD",X"21",X"B1",X"00",X"C3",X"3B",
		X"01",X"21",X"B7",X"00",X"C3",X"4B",X"02",X"32",X"43",X"20",X"52",X"4F",X"4D",X"20",X"20",X"20",
		X"00",X"21",X"00",X"00",X"DD",X"21",X"CB",X"00",X"C3",X"14",X"01",X"21",X"D1",X"00",X"C3",X"4B",
		X"02",X"32",X"45",X"00",X"21",X"00",X"10",X"DD",X"21",X"DE",X"00",X"C3",X"14",X"01",X"21",X"E4",
		X"00",X"C3",X"4B",X"02",X"32",X"46",X"00",X"21",X"00",X"20",X"DD",X"21",X"F1",X"00",X"C3",X"14",
		X"01",X"21",X"F7",X"00",X"C3",X"4B",X"02",X"32",X"48",X"00",X"21",X"00",X"30",X"DD",X"21",X"04",
		X"01",X"C3",X"14",X"01",X"21",X"0A",X"01",X"C3",X"4B",X"02",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"C3",X"1A",X"14",X"01",X"00",X"10",X"AF",X"16",X"FF",X"86",X"5F",X"7A",X"A6",X"57",X"7B",
		X"23",X"0D",X"C2",X"1A",X"01",X"08",X"3A",X"00",X"70",X"08",X"10",X"EE",X"FE",X"FF",X"C2",X"33",
		X"01",X"DD",X"E9",X"7A",X"FE",X"FF",X"C2",X"6C",X"02",X"DD",X"E9",X"DD",X"21",X"42",X"01",X"C3",
		X"82",X"01",X"44",X"4D",X"36",X"00",X"23",X"7D",X"BB",X"C2",X"44",X"01",X"08",X"3A",X"00",X"B0",
		X"08",X"7C",X"BA",X"C2",X"44",X"01",X"69",X"60",X"01",X"55",X"00",X"DD",X"21",X"62",X"01",X"C3",
		X"93",X"01",X"01",X"AA",X"55",X"DD",X"21",X"6C",X"01",X"C3",X"D5",X"01",X"01",X"FF",X"AA",X"DD",
		X"21",X"76",X"01",X"C3",X"93",X"01",X"01",X"00",X"FF",X"DD",X"21",X"80",X"01",X"C3",X"D5",X"01",
		X"FD",X"E9",X"06",X"00",X"70",X"7E",X"B8",X"C2",X"72",X"02",X"08",X"3A",X"00",X"B0",X"08",X"10",
		X"F3",X"DD",X"E9",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",
		X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"D9",X"7E",X"A8",X"C2",X"72",X"02",X"71",X"7E",X"A9",
		X"C2",X"72",X"02",X"23",X"7D",X"BB",X"C2",X"A8",X"01",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",
		X"C2",X"A8",X"01",X"D9",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",
		X"7A",X"D9",X"57",X"DD",X"E9",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",
		X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"D9",X"EB",X"2B",X"7E",X"A8",X"C2",X"72",
		X"02",X"71",X"7E",X"A9",X"C2",X"72",X"02",X"08",X"3A",X"00",X"B0",X"08",X"7D",X"BB",X"C2",X"EB",
		X"01",X"7C",X"BA",X"C2",X"EB",X"01",X"D9",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",
		X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"DD",X"E9",X"21",X"00",X"88",X"11",X"00",X"8C",X"06",X"10",
		X"DD",X"21",X"27",X"02",X"C3",X"38",X"02",X"21",X"00",X"90",X"11",X"00",X"94",X"06",X"00",X"DD",
		X"21",X"36",X"02",X"C3",X"38",X"02",X"FD",X"E9",X"70",X"23",X"7D",X"BB",X"C2",X"38",X"02",X"08",
		X"3A",X"00",X"B0",X"08",X"7C",X"BA",X"C2",X"38",X"02",X"DD",X"E9",X"EB",X"21",X"6E",X"8B",X"1A",
		X"B7",X"CA",X"69",X"02",X"D6",X"30",X"F2",X"5B",X"02",X"3E",X"10",X"77",X"08",X"3A",X"00",X"B0",
		X"08",X"01",X"E0",X"FF",X"09",X"13",X"C3",X"4F",X"02",X"EB",X"23",X"E9",X"3A",X"00",X"B0",X"C3",
		X"6C",X"02",X"3A",X"00",X"B0",X"C3",X"72",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2F",X"31",X"80",X"80",X"F5",X"3A",X"00",X"B0",X"F1",X"CD",X"83",X"05",X"F5",X"3A",X"00",X"B0",
		X"F1",X"D7",X"00",X"E7",X"04",X"04",X"01",X"E7",X"04",X"08",X"02",X"E7",X"04",X"0C",X"03",X"E7",
		X"04",X"10",X"04",X"3E",X"9B",X"32",X"03",X"98",X"3E",X"88",X"32",X"03",X"A0",X"F5",X"3A",X"00",
		X"B0",X"F1",X"3E",X"10",X"32",X"02",X"98",X"CF",X"60",X"20",X"50",X"4F",X"52",X"54",X"20",X"41",
		X"20",X"31",X"00",X"21",X"30",X"40",X"CD",X"DF",X"04",X"3A",X"00",X"98",X"CD",X"C2",X"04",X"3E",
		X"00",X"32",X"02",X"98",X"CF",X"60",X"40",X"50",X"4F",X"52",X"54",X"20",X"41",X"20",X"32",X"00",
		X"21",X"50",X"40",X"CD",X"DF",X"04",X"3A",X"00",X"98",X"CD",X"C2",X"04",X"CF",X"68",X"60",X"50",
		X"4F",X"52",X"54",X"20",X"42",X"00",X"21",X"70",X"40",X"CD",X"DF",X"04",X"3A",X"01",X"98",X"CD",
		X"C2",X"04",X"CF",X"68",X"80",X"50",X"4F",X"52",X"54",X"20",X"43",X"00",X"21",X"90",X"40",X"CD",
		X"DF",X"04",X"3A",X"02",X"98",X"CD",X"C2",X"04",X"CF",X"40",X"A8",X"37",X"20",X"36",X"20",X"35",
		X"20",X"34",X"20",X"33",X"20",X"32",X"20",X"31",X"20",X"30",X"00",X"CF",X"50",X"B0",X"42",X"49",
		X"54",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"53",X"00",X"2E",X"00",X"2D",X"20",X"FD",X"C3",
		X"2D",X"04",X"06",X"08",X"07",X"F5",X"E6",X"01",X"F6",X"30",X"CD",X"6B",X"05",X"AF",X"CD",X"6B",
		X"05",X"F5",X"3A",X"00",X"B0",X"F1",X"F1",X"10",X"EB",X"C9",X"F5",X"AF",X"C3",X"E3",X"04",X"F5",
		X"3A",X"E5",X"80",X"94",X"3D",X"67",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"1D",
		X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"D5",X"11",X"00",X"88",X"19",X"D1",X"F1",X"C9",
		X"E3",X"F5",X"C5",X"D5",X"56",X"23",X"5E",X"23",X"EB",X"CD",X"DA",X"04",X"1A",X"13",X"B7",X"CA",
		X"18",X"05",X"CD",X"6B",X"05",X"C3",X"0C",X"05",X"EB",X"D1",X"C1",X"F1",X"E3",X"C9",X"0E",X"03",
		X"C3",X"2A",X"05",X"0E",X"00",X"C3",X"2A",X"05",X"0E",X"01",X"F5",X"C5",X"D5",X"E5",X"CD",X"DA",
		X"04",X"78",X"3D",X"20",X"02",X"CB",X"81",X"1A",X"CB",X"40",X"20",X"05",X"07",X"07",X"07",X"07",
		X"1B",X"13",X"E6",X"0F",X"C2",X"56",X"05",X"CB",X"41",X"CA",X"58",X"05",X"3E",X"20",X"CB",X"49",
		X"C2",X"64",X"05",X"C3",X"61",X"05",X"CB",X"81",X"C6",X"30",X"FE",X"3A",X"DA",X"61",X"05",X"C6",
		X"07",X"CD",X"6B",X"05",X"10",X"CB",X"E1",X"D1",X"C1",X"F1",X"C9",X"C5",X"D6",X"30",X"F2",X"73",
		X"05",X"3E",X"10",X"77",X"01",X"E0",X"FF",X"09",X"7C",X"FE",X"88",X"30",X"04",X"01",X"00",X"04",
		X"09",X"C1",X"C9",X"F5",X"C5",X"E5",X"21",X"00",X"88",X"0E",X"04",X"3E",X"10",X"CD",X"A8",X"05",
		X"21",X"00",X"90",X"0E",X"01",X"CD",X"A7",X"05",X"3E",X"00",X"32",X"03",X"A8",X"32",X"05",X"A8",
		X"32",X"04",X"A8",X"E1",X"C1",X"F1",X"C9",X"AF",X"06",X"00",X"77",X"23",X"10",X"FC",X"0D",X"20",
		X"F9",X"C9",X"F5",X"C5",X"D5",X"E5",X"50",X"E5",X"CD",X"DA",X"04",X"3E",X"20",X"CD",X"6B",X"05",
		X"10",X"F9",X"E1",X"7D",X"C6",X"08",X"6F",X"42",X"0D",X"20",X"EC",X"E1",X"D1",X"C1",X"F1",X"C9",
		X"E3",X"F5",X"C5",X"D5",X"56",X"23",X"5E",X"23",X"EB",X"CD",X"DF",X"04",X"1A",X"13",X"B7",X"CA",
		X"E8",X"05",X"CD",X"6B",X"05",X"C3",X"DC",X"05",X"EB",X"D1",X"C1",X"F1",X"E3",X"C9",X"F5",X"C5",
		X"D5",X"E5",X"CD",X"DF",X"04",X"0E",X"01",X"C3",X"31",X"05",X"21",X"00",X"00",X"22",X"58",X"81",
		X"22",X"5E",X"81",X"21",X"E2",X"80",X"06",X"24",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"E1",X"7E",
		X"23",X"E5",X"11",X"00",X"00",X"06",X"20",X"C3",X"37",X"06",X"E1",X"7E",X"23",X"E5",X"47",X"0F",
		X"0F",X"E6",X"3E",X"4F",X"78",X"06",X"00",X"21",X"01",X"90",X"09",X"77",X"C9",X"E1",X"46",X"23",
		X"5E",X"16",X"00",X"23",X"7E",X"23",X"E5",X"21",X"01",X"90",X"19",X"19",X"77",X"23",X"23",X"10",
		X"FB",X"C9",X"21",X"01",X"90",X"19",X"19",X"77",X"23",X"23",X"10",X"FB",X"C9",X"DF",X"FF",X"CF",
		X"10",X"F8",X"3B",X"31",X"39",X"38",X"31",X"20",X"53",X"54",X"45",X"52",X"4E",X"20",X"45",X"4C",
		X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"00",X"C9",X"AF",
		X"32",X"1E",X"86",X"3A",X"12",X"81",X"B7",X"28",X"1C",X"DF",X"F1",X"CF",X"18",X"F0",X"43",X"52",
		X"45",X"44",X"49",X"54",X"53",X"20",X"5B",X"20",X"00",X"21",X"F0",X"68",X"11",X"12",X"81",X"06",
		X"02",X"CD",X"1E",X"05",X"C9",X"DF",X"F3",X"CF",X"18",X"F0",X"49",X"4E",X"53",X"45",X"52",X"54",
		X"20",X"43",X"4F",X"49",X"4E",X"00",X"C9",X"AF",X"32",X"1D",X"86",X"DF",X"0B",X"CF",X"20",X"00",
		X"31",X"53",X"54",X"00",X"21",X"08",X"10",X"11",X"4F",X"81",X"06",X"06",X"CD",X"28",X"05",X"CF",
		X"58",X"00",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"00",X"21",X"08",X"68",
		X"11",X"13",X"81",X"06",X"06",X"CD",X"28",X"05",X"3A",X"22",X"86",X"FE",X"02",X"C0",X"CF",X"D0",
		X"00",X"32",X"4E",X"44",X"00",X"21",X"08",X"C0",X"11",X"52",X"81",X"06",X"06",X"CD",X"28",X"05",
		X"C9",X"DF",X"F5",X"CF",X"18",X"F0",X"4C",X"49",X"56",X"45",X"53",X"20",X"4C",X"45",X"46",X"54",
		X"20",X"5B",X"20",X"00",X"21",X"F0",X"80",X"11",X"28",X"86",X"06",X"02",X"CD",X"1E",X"05",X"C9",
		X"DF",X"7E",X"CF",X"40",X"78",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"00",X"21",X"78",X"78",
		X"11",X"27",X"86",X"06",X"01",X"CD",X"28",X"05",X"CF",X"80",X"78",X"20",X"55",X"50",X"00",X"C9",
		X"3A",X"12",X"81",X"B7",X"C8",X"21",X"B8",X"00",X"01",X"05",X"20",X"CD",X"B2",X"05",X"E7",X"05",
		X"17",X"05",X"3A",X"12",X"81",X"FE",X"01",X"20",X"40",X"CF",X"18",X"B8",X"50",X"55",X"53",X"48",
		X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"CF",X"68",X"C8",X"5B",X"20",X"4F",X"52",X"20",X"5B",
		X"00",X"CF",X"30",X"D8",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"41",X"4E",X"4F",X"54",X"48",
		X"45",X"52",X"20",X"43",X"4F",X"49",X"4E",X"00",X"C9",X"CF",X"48",X"B8",X"50",X"55",X"53",X"48",
		X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"CF",X"68",X"C8",X"5B",X"20",X"4F",
		X"52",X"20",X"5B",X"00",X"CF",X"28",X"D8",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",
		X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"06",X"05",X"C5",
		X"E7",X"05",X"17",X"01",X"3E",X"05",X"CD",X"CF",X"14",X"E7",X"05",X"17",X"02",X"3E",X"05",X"CD",
		X"CF",X"14",X"E7",X"05",X"17",X"03",X"3E",X"05",X"CD",X"CF",X"14",X"E7",X"05",X"17",X"04",X"3E",
		X"05",X"CD",X"CF",X"14",X"E7",X"05",X"17",X"05",X"3E",X"05",X"CD",X"CF",X"14",X"E7",X"05",X"17",
		X"06",X"3E",X"05",X"CD",X"CF",X"14",X"E7",X"05",X"17",X"07",X"3E",X"05",X"CD",X"CF",X"14",X"E7",
		X"05",X"17",X"00",X"3E",X"05",X"CD",X"CF",X"14",X"C1",X"10",X"B4",X"C9",X"F5",X"3A",X"1F",X"86",
		X"B7",X"28",X"09",X"3A",X"01",X"98",X"E6",X"02",X"28",X"11",X"F1",X"C9",X"3A",X"9A",X"86",X"B7",
		X"28",X"09",X"3A",X"01",X"98",X"E6",X"02",X"28",X"02",X"F1",X"C9",X"F1",X"F3",X"32",X"00",X"A0",
		X"AF",X"32",X"01",X"A0",X"E3",X"E3",X"3E",X"08",X"32",X"01",X"A0",X"FB",X"C9",X"D9",X"ED",X"5B",
		X"18",X"86",X"19",X"29",X"19",X"29",X"19",X"29",X"19",X"29",X"29",X"19",X"29",X"29",X"19",X"29",
		X"29",X"19",X"29",X"19",X"29",X"29",X"19",X"29",X"19",X"29",X"19",X"11",X"2F",X"6A",X"19",X"22",
		X"18",X"86",X"7C",X"D9",X"C9",X"FD",X"E1",X"DD",X"21",X"46",X"82",X"DD",X"CB",X"00",X"C6",X"DD",
		X"CB",X"00",X"CE",X"CD",X"1F",X"09",X"31",X"90",X"80",X"FD",X"E9",X"FD",X"E1",X"DD",X"21",X"18",
		X"82",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"1F",X"09",X"31",X"B8",X"80",X"DD",
		X"21",X"55",X"81",X"DD",X"CB",X"00",X"C6",X"CD",X"08",X"09",X"CD",X"33",X"09",X"FD",X"E9",X"D9",
		X"21",X"47",X"0A",X"CD",X"ED",X"08",X"D9",X"D0",X"CD",X"08",X"09",X"CD",X"33",X"09",X"37",X"C9",
		X"D9",X"21",X"57",X"0A",X"CD",X"ED",X"08",X"D9",X"D0",X"CD",X"08",X"09",X"CD",X"33",X"09",X"37",
		X"DD",X"CB",X"00",X"E6",X"C9",X"E1",X"D9",X"21",X"67",X"0A",X"CD",X"ED",X"08",X"D9",X"D2",X"DC",
		X"08",X"DD",X"22",X"DA",X"80",X"CD",X"1F",X"09",X"CD",X"C8",X"09",X"37",X"E9",X"E1",X"D9",X"21",
		X"3F",X"0A",X"C3",X"CA",X"08",X"E1",X"D9",X"21",X"35",X"0A",X"C3",X"CA",X"08",X"E5",X"D1",X"7E",
		X"23",X"66",X"6F",X"B4",X"C8",X"7E",X"B7",X"28",X"06",X"13",X"13",X"D5",X"E1",X"18",X"F0",X"E5",
		X"DD",X"E1",X"DD",X"CB",X"00",X"C6",X"37",X"C9",X"D9",X"DD",X"E5",X"E1",X"DD",X"2A",X"DA",X"80",
		X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"CB",X"00",X"DE",X"E5",X"DD",X"E1",X"D9",X"C9",X"D9",
		X"DD",X"CB",X"00",X"CE",X"DD",X"E5",X"E1",X"22",X"DA",X"80",X"AF",X"06",X"0F",X"23",X"77",X"10",
		X"FC",X"D9",X"C9",X"D9",X"DD",X"E5",X"E1",X"22",X"D8",X"80",X"AF",X"06",X"0C",X"23",X"77",X"10",
		X"FC",X"D9",X"C9",X"21",X"00",X"00",X"39",X"31",X"68",X"80",X"FD",X"E5",X"FD",X"2A",X"DA",X"80",
		X"FD",X"22",X"DE",X"80",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"C9",X"21",X"00",X"00",X"39",X"31",
		X"68",X"80",X"DD",X"2A",X"DA",X"80",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"2A",X"DE",X"80",X"7C",
		X"B5",X"28",X"0C",X"DD",X"2A",X"DE",X"80",X"21",X"00",X"00",X"22",X"DE",X"80",X"18",X"04",X"DD",
		X"2A",X"DA",X"80",X"CD",X"98",X"09",X"DD",X"CB",X"00",X"46",X"28",X"F7",X"DD",X"22",X"DA",X"80",
		X"DD",X"66",X"0F",X"DD",X"6E",X"0E",X"F9",X"C9",X"D9",X"01",X"2E",X"00",X"DD",X"09",X"DD",X"E5",
		X"E1",X"01",X"0C",X"86",X"B7",X"ED",X"42",X"38",X"04",X"DD",X"21",X"18",X"82",X"D9",X"C9",X"DD",
		X"2A",X"DA",X"80",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"CD",X"5B",X"09",X"DD",X"2A",X"DA",
		X"80",X"DD",X"CB",X"00",X"6E",X"20",X"F3",X"C9",X"D9",X"D1",X"01",X"2E",X"00",X"DD",X"E5",X"E1",
		X"09",X"F9",X"D5",X"D9",X"C9",X"CD",X"E5",X"09",X"D9",X"2A",X"DA",X"80",X"06",X"10",X"AF",X"77",
		X"23",X"10",X"FC",X"D9",X"C9",X"DD",X"2A",X"DA",X"80",X"DD",X"CB",X"00",X"5E",X"C8",X"DD",X"CB",
		X"00",X"9E",X"D9",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"06",X"0D",X"AF",X"77",X"23",X"10",X"FC",
		X"DD",X"77",X"01",X"DD",X"77",X"01",X"D9",X"C9",X"CD",X"69",X"0C",X"DD",X"21",X"18",X"82",X"AF",
		X"DD",X"77",X"00",X"DD",X"21",X"74",X"82",X"DD",X"77",X"00",X"CD",X"98",X"09",X"30",X"02",X"18",
		X"F6",X"DD",X"21",X"55",X"81",X"11",X"0D",X"00",X"06",X"0F",X"DD",X"77",X"00",X"DD",X"19",X"10",
		X"F9",X"CD",X"6F",X"0C",X"C9",X"CA",X"84",X"F8",X"84",X"26",X"85",X"54",X"85",X"00",X"00",X"82",
		X"85",X"B0",X"85",X"DE",X"85",X"00",X"00",X"62",X"81",X"6F",X"81",X"7C",X"81",X"89",X"81",X"96",
		X"81",X"A3",X"81",X"B0",X"81",X"00",X"00",X"BD",X"81",X"CA",X"81",X"D7",X"81",X"E4",X"81",X"F1",
		X"81",X"FE",X"81",X"0B",X"82",X"00",X"00",X"74",X"82",X"A2",X"82",X"D0",X"82",X"FE",X"82",X"2C",
		X"83",X"5A",X"83",X"88",X"83",X"B6",X"83",X"E4",X"83",X"12",X"84",X"40",X"84",X"6E",X"84",X"00",
		X"00",X"3E",X"11",X"CD",X"0C",X"08",X"CD",X"83",X"05",X"CD",X"BC",X"0A",X"CD",X"F1",X"06",X"3A",
		X"22",X"86",X"3D",X"06",X"03",X"28",X"07",X"06",X"05",X"3E",X"04",X"CD",X"0C",X"08",X"C5",X"CD",
		X"FA",X"05",X"CD",X"10",X"07",X"3E",X"0C",X"CD",X"AF",X"09",X"21",X"70",X"38",X"01",X"03",X"0E",
		X"CD",X"B2",X"05",X"3E",X"05",X"CD",X"AF",X"09",X"C1",X"10",X"E3",X"C9",X"3A",X"27",X"86",X"FE",
		X"02",X"20",X"15",X"3A",X"02",X"98",X"E6",X"08",X"20",X"0E",X"3E",X"00",X"32",X"02",X"98",X"3E",
		X"FF",X"32",X"07",X"A8",X"32",X"06",X"A8",X"C9",X"3E",X"10",X"32",X"02",X"98",X"3E",X"00",X"32",
		X"07",X"A8",X"32",X"06",X"A8",X"C9",X"F5",X"3A",X"00",X"B0",X"AF",X"32",X"01",X"A8",X"3C",X"32",
		X"01",X"A8",X"3A",X"06",X"81",X"CB",X"0F",X"32",X"06",X"81",X"DA",X"47",X"0C",X"3A",X"07",X"81",
		X"B7",X"C2",X"44",X"0C",X"CD",X"46",X"0C",X"3C",X"32",X"07",X"81",X"ED",X"73",X"DC",X"80",X"31",
		X"40",X"80",X"08",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"D9",X"C5",X"D5",X"E5",X"21",
		X"A2",X"86",X"34",X"3A",X"A2",X"86",X"FE",X"3D",X"20",X"09",X"36",X"00",X"2A",X"A3",X"86",X"23",
		X"22",X"A3",X"86",X"3A",X"9A",X"86",X"B7",X"C2",X"87",X"0B",X"21",X"55",X"81",X"11",X"40",X"90",
		X"06",X"08",X"C5",X"CB",X"46",X"CC",X"04",X"0E",X"01",X"06",X"00",X"09",X"3A",X"27",X"86",X"FE",
		X"02",X"20",X"1E",X"3A",X"02",X"98",X"E6",X"08",X"20",X"17",X"7E",X"3D",X"3D",X"12",X"23",X"13",
		X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"23",X"23",X"23",X"13",X"7E",X"3C",X"3C",X"12",X"18",
		X"11",X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"23",X"23",X"23",X"13",
		X"7E",X"12",X"23",X"13",X"C1",X"10",X"BB",X"21",X"BD",X"81",X"11",X"61",X"90",X"06",X"07",X"C5",
		X"CB",X"46",X"CC",X"04",X"0E",X"01",X"06",X"00",X"09",X"3A",X"27",X"86",X"FE",X"02",X"20",X"17",
		X"3A",X"02",X"98",X"E6",X"08",X"20",X"10",X"7E",X"C6",X"06",X"12",X"01",X"06",X"00",X"09",X"13",
		X"13",X"7E",X"C6",X"04",X"C3",X"C5",X"0B",X"7E",X"C6",X"08",X"12",X"01",X"06",X"00",X"09",X"13",
		X"13",X"7E",X"2F",X"C6",X"F1",X"12",X"23",X"13",X"13",X"C1",X"10",X"C3",X"3A",X"E5",X"80",X"21",
		X"04",X"90",X"06",X"1B",X"77",X"23",X"23",X"10",X"FB",X"2A",X"E2",X"80",X"ED",X"5B",X"E4",X"80",
		X"19",X"22",X"E4",X"80",X"CD",X"20",X"32",X"21",X"74",X"82",X"06",X"0D",X"C5",X"CB",X"7E",X"C4",
		X"75",X"0C",X"11",X"2E",X"00",X"19",X"C1",X"10",X"F3",X"CD",X"CB",X"0F",X"21",X"18",X"82",X"46",
		X"CB",X"90",X"CB",X"40",X"C4",X"9A",X"0C",X"CB",X"D0",X"CB",X"58",X"C4",X"40",X"0D",X"21",X"46",
		X"82",X"06",X"15",X"C5",X"46",X"CB",X"40",X"C4",X"9A",X"0C",X"CB",X"58",X"C4",X"40",X"0D",X"11",
		X"2E",X"00",X"19",X"C1",X"10",X"ED",X"CD",X"13",X"0E",X"CD",X"73",X"0E",X"E1",X"D1",X"C1",X"D9",
		X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"08",X"ED",X"7B",X"DC",X"80",X"AF",X"32",X"07",
		X"81",X"CD",X"46",X"0C",X"F1",X"C9",X"C9",X"ED",X"73",X"E0",X"80",X"31",X"D8",X"80",X"C5",X"D5",
		X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"CD",X"73",X"0E",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",
		X"E1",X"D1",X"C1",X"ED",X"7B",X"E0",X"80",X"F1",X"C9",X"3E",X"FF",X"32",X"06",X"81",X"C9",X"3E",
		X"00",X"32",X"06",X"81",X"C9",X"CB",X"4E",X"C8",X"CB",X"5E",X"C0",X"E5",X"01",X"05",X"00",X"09",
		X"5E",X"23",X"56",X"13",X"13",X"13",X"23",X"23",X"46",X"23",X"23",X"7E",X"C6",X"04",X"6F",X"78",
		X"C6",X"04",X"67",X"1A",X"CD",X"DF",X"04",X"77",X"E1",X"C9",X"E5",X"23",X"5E",X"23",X"56",X"D5",
		X"FD",X"E1",X"23",X"CB",X"68",X"28",X"05",X"35",X"20",X"02",X"CB",X"A8",X"23",X"CB",X"60",X"28",
		X"6D",X"35",X"20",X"6A",X"CB",X"F8",X"23",X"5E",X"23",X"56",X"13",X"13",X"13",X"13",X"13",X"1A",
		X"B7",X"C2",X"D5",X"0C",X"13",X"1A",X"B7",X"C2",X"CE",X"0C",X"CB",X"A0",X"CB",X"B8",X"EB",X"23",
		X"7E",X"23",X"66",X"6F",X"EB",X"72",X"2B",X"73",X"13",X"13",X"1A",X"CB",X"7F",X"28",X"3D",X"4F",
		X"C5",X"FD",X"7E",X"03",X"FD",X"AE",X"04",X"4F",X"FD",X"7E",X"04",X"B7",X"F2",X"F0",X"0C",X"2F",
		X"1F",X"CB",X"19",X"1F",X"CB",X"19",X"FD",X"7E",X"09",X"FD",X"AE",X"0A",X"47",X"FD",X"7E",X"0A",
		X"B7",X"F2",X"05",X"0D",X"2F",X"1F",X"CB",X"18",X"1F",X"CB",X"18",X"78",X"B1",X"C1",X"CB",X"3F",
		X"CB",X"3F",X"4F",X"1A",X"CB",X"BF",X"91",X"F2",X"1B",X"0D",X"AF",X"3C",X"2B",X"77",X"CB",X"50",
		X"28",X"1B",X"CB",X"48",X"CA",X"3D",X"0D",X"23",X"23",X"23",X"E5",X"5E",X"23",X"56",X"2A",X"E2",
		X"80",X"19",X"EB",X"E1",X"73",X"FD",X"73",X"05",X"23",X"72",X"FD",X"72",X"06",X"E1",X"70",X"C9",
		X"CB",X"48",X"C8",X"E5",X"DD",X"E1",X"CB",X"78",X"28",X"14",X"CB",X"BE",X"DD",X"66",X"06",X"DD",
		X"6E",X"05",X"23",X"23",X"23",X"7E",X"FD",X"77",X"07",X"23",X"7E",X"FD",X"77",X"08",X"CB",X"50",
		X"CA",X"00",X"0E",X"DD",X"7E",X"07",X"FD",X"77",X"05",X"DD",X"7E",X"08",X"FD",X"77",X"06",X"DD",
		X"7E",X"09",X"FD",X"77",X"0B",X"DD",X"7E",X"0A",X"FD",X"77",X"0C",X"FD",X"E5",X"E1",X"23",X"FD",
		X"CB",X"00",X"4E",X"28",X"07",X"35",X"20",X"04",X"FD",X"CB",X"00",X"8E",X"23",X"FD",X"CB",X"00",
		X"56",X"28",X"07",X"35",X"20",X"04",X"FD",X"CB",X"00",X"96",X"FD",X"CB",X"00",X"76",X"20",X"60",
		X"FD",X"CB",X"00",X"5E",X"20",X"5A",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"09",
		X"EB",X"2B",X"73",X"DD",X"73",X"07",X"23",X"72",X"DD",X"72",X"08",X"FD",X"CB",X"00",X"66",X"20",
		X"0F",X"7A",X"FE",X"09",X"38",X"06",X"FE",X"F1",X"30",X"02",X"18",X"04",X"FD",X"CB",X"00",X"F6",
		X"23",X"23",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"2B",X"73",X"DD",
		X"73",X"09",X"23",X"72",X"DD",X"72",X"0A",X"FD",X"CB",X"00",X"66",X"20",X"13",X"7E",X"FE",X"13",
		X"30",X"04",X"3E",X"13",X"18",X"06",X"FE",X"D4",X"38",X"06",X"3E",X"D3",X"77",X"DD",X"77",X"0A",
		X"DD",X"E5",X"E1",X"C9",X"AF",X"E5",X"DD",X"E1",X"DD",X"77",X"06",X"DD",X"77",X"0C",X"C9",X"00",
		X"00",X"00",X"00",X"DD",X"21",X"18",X"82",X"FD",X"21",X"74",X"82",X"3A",X"21",X"86",X"6F",X"DD",
		X"4E",X"0A",X"D9",X"3A",X"20",X"86",X"6F",X"DD",X"4E",X"08",X"06",X"0D",X"FD",X"7E",X"00",X"E6",
		X"41",X"EE",X"41",X"20",X"37",X"FD",X"56",X"06",X"FD",X"5E",X"05",X"1A",X"67",X"13",X"1A",X"D9",
		X"85",X"1F",X"67",X"FD",X"7E",X"0A",X"91",X"30",X"02",X"ED",X"44",X"BC",X"D9",X"30",X"1D",X"7C",
		X"85",X"1F",X"67",X"FD",X"7E",X"08",X"91",X"30",X"02",X"ED",X"44",X"BC",X"30",X"0E",X"DD",X"7E",
		X"0D",X"FD",X"56",X"0C",X"B2",X"DD",X"77",X"0D",X"FD",X"CB",X"0D",X"C6",X"11",X"2E",X"00",X"FD",
		X"19",X"10",X"B9",X"21",X"08",X"81",X"7E",X"23",X"46",X"A8",X"4F",X"3A",X"00",X"98",X"2F",X"77",
		X"2B",X"70",X"A1",X"E6",X"C0",X"23",X"23",X"CB",X"7F",X"28",X"01",X"34",X"23",X"CB",X"77",X"28",
		X"01",X"34",X"CD",X"C0",X"0E",X"CD",X"26",X"0F",X"C9",X"3A",X"12",X"81",X"C6",X"99",X"27",X"32",
		X"12",X"81",X"C9",X"47",X"B7",X"C8",X"3E",X"FF",X"32",X"1E",X"86",X"3A",X"12",X"81",X"FE",X"99",
		X"C8",X"80",X"27",X"30",X"02",X"3E",X"99",X"32",X"12",X"81",X"3E",X"05",X"CD",X"0C",X"08",X"C9",
		X"D9",X"11",X"0A",X"81",X"3A",X"0C",X"81",X"4F",X"21",X"6B",X"0F",X"CD",X"E5",X"0E",X"79",X"32",
		X"0C",X"81",X"11",X"0B",X"81",X"3A",X"0D",X"81",X"4F",X"21",X"9B",X"0F",X"CD",X"E5",X"0E",X"79",
		X"32",X"0D",X"81",X"D9",X"C9",X"3A",X"02",X"98",X"2F",X"E6",X"06",X"CB",X"3F",X"47",X"28",X"08",
		X"D5",X"11",X"0C",X"00",X"19",X"10",X"FD",X"D1",X"1A",X"B7",X"C8",X"09",X"AF",X"86",X"08",X"79",
		X"FE",X"0B",X"20",X"09",X"D5",X"11",X"0C",X"00",X"AF",X"ED",X"52",X"4F",X"D1",X"0C",X"23",X"08",
		X"EB",X"35",X"CD",X"1C",X"0F",X"EB",X"20",X"E5",X"CD",X"A3",X"0E",X"C9",X"F5",X"3A",X"0E",X"81",
		X"3C",X"32",X"0E",X"81",X"F1",X"C9",X"3A",X"11",X"81",X"B7",X"28",X"25",X"3A",X"10",X"81",X"B7",
		X"28",X"05",X"3D",X"32",X"10",X"81",X"C9",X"3A",X"0F",X"81",X"B7",X"28",X"0E",X"3E",X"00",X"32",
		X"02",X"A8",X"32",X"0F",X"81",X"3E",X"0C",X"32",X"10",X"81",X"C9",X"3E",X"00",X"32",X"11",X"81",
		X"C9",X"3A",X"0E",X"81",X"B7",X"C8",X"3D",X"32",X"0E",X"81",X"3E",X"FF",X"32",X"11",X"81",X"32",
		X"0F",X"81",X"32",X"02",X"A8",X"3E",X"04",X"32",X"10",X"81",X"C9",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"3A",X"1F",X"86",X"B7",X"C2",
		X"C3",X"46",X"DD",X"21",X"0C",X"86",X"21",X"00",X"98",X"CD",X"30",X"10",X"DD",X"23",X"23",X"CD",
		X"30",X"10",X"DD",X"23",X"23",X"CD",X"30",X"10",X"3A",X"27",X"86",X"FE",X"02",X"C0",X"3A",X"02",
		X"98",X"E6",X"08",X"C0",X"21",X"0F",X"86",X"DD",X"21",X"10",X"86",X"DD",X"CB",X"00",X"56",X"CB",
		X"8E",X"28",X"02",X"CB",X"CE",X"3A",X"0F",X"86",X"E6",X"C7",X"6F",X"3A",X"10",X"86",X"E6",X"38",
		X"B5",X"32",X"0F",X"86",X"21",X"11",X"86",X"DD",X"21",X"0F",X"86",X"DD",X"CB",X"00",X"46",X"CB",
		X"A6",X"28",X"02",X"CB",X"E6",X"21",X"11",X"86",X"CB",X"46",X"CB",X"B6",X"C8",X"CB",X"F6",X"C9",
		X"DD",X"7E",X"00",X"DD",X"46",X"03",X"57",X"7E",X"2F",X"4F",X"7A",X"A1",X"DD",X"77",X"06",X"DD",
		X"70",X"00",X"DD",X"71",X"03",X"C9",X"CD",X"C5",X"08",X"30",X"FB",X"DD",X"36",X"03",X"64",X"3A",
		X"2C",X"86",X"21",X"91",X"86",X"77",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"6E",X"20",X"29",
		X"DD",X"36",X"03",X"64",X"DD",X"CB",X"00",X"EE",X"21",X"91",X"86",X"35",X"20",X"1B",X"3A",X"23",
		X"86",X"21",X"2B",X"86",X"BE",X"30",X"0B",X"21",X"23",X"86",X"34",X"FD",X"21",X"DB",X"29",X"CD",
		X"43",X"09",X"21",X"91",X"86",X"3A",X"2C",X"86",X"77",X"CD",X"5B",X"09",X"18",X"CC",X"AF",X"32",
		X"23",X"86",X"21",X"B0",X"10",X"3A",X"2A",X"86",X"BE",X"28",X"0B",X"3E",X"FF",X"BE",X"C8",X"11",
		X"06",X"00",X"19",X"C3",X"95",X"10",X"23",X"01",X"05",X"00",X"11",X"2B",X"86",X"ED",X"B0",X"C9",
		X"01",X"02",X"15",X"30",X"D0",X"00",X"02",X"03",X"10",X"30",X"12",X"01",X"03",X"03",X"10",X"30",
		X"22",X"01",X"04",X"03",X"10",X"30",X"22",X"01",X"05",X"03",X"0F",X"40",X"32",X"01",X"06",X"03",
		X"0E",X"40",X"32",X"01",X"07",X"03",X"0D",X"40",X"42",X"01",X"08",X"04",X"0C",X"50",X"42",X"01",
		X"09",X"04",X"09",X"50",X"42",X"01",X"0A",X"04",X"09",X"50",X"42",X"01",X"0B",X"04",X"06",X"60",
		X"42",X"01",X"0C",X"04",X"06",X"60",X"42",X"01",X"0D",X"04",X"06",X"60",X"52",X"01",X"0E",X"05",
		X"06",X"70",X"52",X"01",X"0F",X"05",X"06",X"70",X"52",X"01",X"10",X"05",X"06",X"70",X"52",X"01",
		X"11",X"05",X"06",X"90",X"52",X"01",X"12",X"05",X"06",X"A0",X"52",X"01",X"13",X"05",X"06",X"B0",
		X"52",X"01",X"14",X"05",X"06",X"E0",X"62",X"01",X"15",X"05",X"06",X"F0",X"62",X"01",X"FF",X"00",
		X"00",X"01",X"00",X"00",X"10",X"08",X"09",X"27",X"05",X"10",X"08",X"09",X"25",X"05",X"00",X"01",
		X"34",X"11",X"00",X"00",X"01",X"00",X"00",X"08",X"10",X"09",X"24",X"05",X"08",X"10",X"09",X"26",
		X"05",X"00",X"01",X"47",X"11",X"00",X"00",X"01",X"00",X"00",X"08",X"10",X"09",X"64",X"05",X"08",
		X"10",X"09",X"66",X"05",X"00",X"01",X"5A",X"11",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"04",
		X"38",X"01",X"01",X"00",X"04",X"B8",X"02",X"01",X"00",X"04",X"F8",X"03",X"01",X"00",X"04",X"38",
		X"02",X"01",X"00",X"04",X"B8",X"03",X"01",X"00",X"04",X"F8",X"01",X"01",X"00",X"04",X"38",X"03",
		X"01",X"00",X"04",X"B8",X"01",X"01",X"00",X"04",X"F8",X"02",X"01",X"00",X"05",X"37",X"01",X"01",
		X"00",X"05",X"B7",X"02",X"01",X"00",X"05",X"F7",X"03",X"01",X"00",X"05",X"37",X"02",X"01",X"00",
		X"05",X"B7",X"01",X"01",X"00",X"05",X"F7",X"03",X"01",X"00",X"05",X"36",X"01",X"01",X"00",X"05",
		X"B6",X"02",X"01",X"00",X"05",X"F6",X"03",X"00",X"00",X"00",X"00",X"CD",X"C5",X"08",X"D2",X"7F",
		X"09",X"DD",X"E5",X"CD",X"9F",X"08",X"D2",X"55",X"13",X"FD",X"E1",X"CD",X"B1",X"13",X"CD",X"D7",
		X"13",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"FD",X"CB",X"00",X"D6",X"DD",X"E5",X"CD",
		X"5B",X"09",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"55",X"13",X"FD",X"CB",X"00",X"76",X"C2",
		X"55",X"13",X"FD",X"CB",X"00",X"4E",X"CC",X"1D",X"12",X"DD",X"7E",X"0A",X"FE",X"16",X"DA",X"DE",
		X"12",X"FE",X"D0",X"D2",X"DE",X"12",X"FD",X"E5",X"CD",X"5B",X"09",X"18",X"D5",X"FD",X"CB",X"00",
		X"DE",X"DD",X"7E",X"0A",X"E6",X"0E",X"FE",X"02",X"C2",X"AE",X"12",X"DD",X"7E",X"0A",X"CB",X"67",
		X"CA",X"AE",X"12",X"3A",X"E5",X"80",X"47",X"DD",X"7E",X"08",X"90",X"47",X"E6",X"0E",X"FE",X"0C",
		X"C2",X"AE",X"12",X"78",X"CB",X"67",X"CA",X"AE",X"12",X"FD",X"36",X"01",X"07",X"FD",X"CB",X"00",
		X"CE",X"DD",X"CB",X"00",X"A6",X"CD",X"B7",X"12",X"FE",X"02",X"20",X"27",X"FD",X"36",X"09",X"01",
		X"FD",X"36",X"0A",X"FF",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"42",X"11",X"DD",
		X"CB",X"0B",X"5E",X"28",X"04",X"FD",X"36",X"0A",X"FE",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",
		X"36",X"04",X"01",X"FE",X"03",X"20",X"27",X"FD",X"36",X"09",X"FF",X"FD",X"36",X"0A",X"00",X"FD",
		X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"55",X"11",X"DD",X"CB",X"0B",X"5E",X"28",X"04",
		X"FD",X"36",X"0A",X"01",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",
		X"00",X"9E",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"CB",X"0B",X"DE",X"3E",X"6C",X"FD",X"BE",X"06",
		X"28",X"07",X"3E",X"6B",X"FD",X"BE",X"06",X"20",X"0E",X"3A",X"61",X"81",X"FD",X"BE",X"0C",X"38",
		X"03",X"3E",X"03",X"C9",X"3E",X"02",X"C9",X"3E",X"00",X"DD",X"CB",X"0B",X"9E",X"C9",X"FD",X"36",
		X"09",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"CB",
		X"00",X"9E",X"01",X"01",X"03",X"CD",X"73",X"17",X"3E",X"0E",X"CD",X"0C",X"08",X"DD",X"CB",X"0C",
		X"96",X"DD",X"CB",X"00",X"A6",X"21",X"68",X"11",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",
		X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"66",X"28",X"39",X"DD",X"66",X"02",X"DD",
		X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"CB",X"00",X"76",X"20",X"2A",X"3E",X"FF",X"32",X"05",X"A8",
		X"3E",X"03",X"CD",X"AF",X"09",X"3E",X"00",X"32",X"05",X"A8",X"3E",X"04",X"CD",X"AF",X"09",X"3E",
		X"FF",X"32",X"03",X"A8",X"3E",X"02",X"CD",X"AF",X"09",X"3E",X"00",X"32",X"03",X"A8",X"3E",X"04",
		X"CD",X"AF",X"09",X"18",X"C1",X"3E",X"00",X"32",X"03",X"A8",X"32",X"05",X"A8",X"DD",X"66",X"02",
		X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",
		X"03",X"00",X"FD",X"36",X"04",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"08",X"00",X"FD",X"36",
		X"06",X"00",X"FD",X"36",X"0C",X"00",X"DD",X"CB",X"00",X"96",X"3E",X"FF",X"CD",X"AF",X"09",X"CD",
		X"D5",X"09",X"CD",X"3D",X"08",X"CB",X"47",X"28",X"0C",X"FD",X"21",X"4E",X"2E",X"CD",X"43",X"09",
		X"CD",X"5B",X"09",X"18",X"FB",X"FD",X"21",X"CB",X"11",X"CD",X"43",X"09",X"CD",X"5B",X"09",X"18",
		X"FB",X"FD",X"36",X"08",X"EB",X"CD",X"3D",X"08",X"E6",X"03",X"FD",X"36",X"0A",X"53",X"FE",X"00",
		X"28",X"0C",X"FD",X"36",X"0A",X"93",X"FE",X"01",X"28",X"04",X"FD",X"36",X"0A",X"73",X"DD",X"36",
		X"04",X"FF",X"DD",X"36",X"03",X"01",X"C9",X"21",X"2F",X"11",X"FD",X"75",X"05",X"FD",X"74",X"06",
		X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"E5",X"3E",X"10",X"77",X"2B",X"77",X"3E",
		X"FF",X"32",X"9B",X"86",X"E1",X"3E",X"13",X"CD",X"0C",X"08",X"C9",X"E5",X"3A",X"9B",X"86",X"B7",
		X"28",X"15",X"3E",X"10",X"77",X"2B",X"77",X"3E",X"00",X"32",X"9B",X"86",X"3E",X"13",X"CD",X"0C",
		X"08",X"01",X"01",X"03",X"CD",X"73",X"17",X"E1",X"C9",X"76",X"3E",X"00",X"32",X"01",X"A8",X"32",
		X"02",X"A8",X"32",X"03",X"A8",X"32",X"04",X"A8",X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"9B",
		X"32",X"03",X"98",X"3E",X"88",X"32",X"03",X"A0",X"31",X"68",X"80",X"21",X"68",X"80",X"0E",X"08",
		X"CD",X"A7",X"05",X"3E",X"FF",X"32",X"08",X"81",X"32",X"09",X"81",X"21",X"FA",X"14",X"11",X"13",
		X"81",X"01",X"3C",X"00",X"ED",X"B0",X"31",X"68",X"80",X"21",X"00",X"90",X"0E",X"01",X"CD",X"A7",
		X"05",X"CD",X"87",X"14",X"CD",X"7D",X"14",X"CD",X"36",X"15",X"3E",X"08",X"CD",X"A4",X"14",X"CD",
		X"B3",X"17",X"3E",X"04",X"CD",X"A4",X"14",X"CD",X"0F",X"1B",X"C3",X"61",X"14",X"3A",X"01",X"98",
		X"2F",X"E6",X"03",X"C0",X"3E",X"99",X"C9",X"E1",X"22",X"1A",X"86",X"32",X"1C",X"86",X"CD",X"08",
		X"0A",X"CD",X"65",X"08",X"AF",X"32",X"07",X"81",X"3E",X"FF",X"32",X"01",X"A8",X"2A",X"1A",X"86",
		X"3A",X"1C",X"86",X"E9",X"D5",X"E5",X"C5",X"F5",X"DD",X"2A",X"DA",X"80",X"DD",X"CB",X"00",X"EE",
		X"DD",X"36",X"03",X"1E",X"CD",X"3D",X"08",X"CD",X"57",X"2F",X"3A",X"1E",X"86",X"B7",X"C4",X"6F",
		X"06",X"DD",X"CB",X"00",X"6E",X"20",X"ED",X"F1",X"3D",X"20",X"DC",X"C1",X"E1",X"D1",X"C9",X"D5",
		X"E5",X"C5",X"F5",X"DD",X"2A",X"DA",X"80",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"03",X"01",X"CD",
		X"3D",X"08",X"CD",X"57",X"2F",X"3A",X"1E",X"86",X"B7",X"C4",X"6F",X"06",X"DD",X"CB",X"00",X"6E",
		X"20",X"ED",X"F1",X"3D",X"20",X"DC",X"C1",X"E1",X"D1",X"C9",X"02",X"04",X"40",X"47",X"4A",X"4C",
		X"01",X"99",X"10",X"4F",X"42",X"45",X"01",X"61",X"20",X"45",X"4C",X"50",X"01",X"17",X"80",X"4D",
		X"59",X"4B",X"00",X"98",X"60",X"41",X"50",X"48",X"00",X"85",X"70",X"4A",X"56",X"43",X"00",X"65",
		X"50",X"52",X"4F",X"42",X"00",X"03",X"30",X"4A",X"4D",X"48",X"00",X"02",X"20",X"44",X"41",X"4E",
		X"00",X"01",X"10",X"57",X"48",X"50",X"CD",X"83",X"05",X"CD",X"4D",X"06",X"CD",X"6F",X"06",X"CD",
		X"A7",X"06",X"DF",X"2A",X"E7",X"06",X"07",X"03",X"E7",X"08",X"0D",X"02",X"E7",X"05",X"15",X"05",
		X"CF",X"38",X"28",X"5B",X"20",X"54",X"4F",X"50",X"20",X"31",X"30",X"20",X"53",X"43",X"4F",X"52",
		X"45",X"53",X"20",X"5B",X"00",X"11",X"13",X"81",X"21",X"38",X"38",X"3E",X"01",X"08",X"D5",X"EB",
		X"7E",X"23",X"B6",X"23",X"B6",X"EB",X"D1",X"C8",X"E5",X"D5",X"08",X"32",X"00",X"80",X"08",X"06",
		X"02",X"11",X"00",X"80",X"CD",X"28",X"05",X"01",X"00",X"20",X"09",X"D1",X"06",X"06",X"CD",X"28",
		X"05",X"13",X"13",X"13",X"01",X"00",X"30",X"09",X"CD",X"DA",X"04",X"06",X"03",X"3E",X"20",X"CD",
		X"6B",X"05",X"10",X"F9",X"06",X"03",X"1A",X"13",X"CD",X"6B",X"05",X"10",X"F9",X"E1",X"01",X"10",
		X"00",X"09",X"08",X"C6",X"01",X"27",X"FE",X"11",X"DA",X"6D",X"15",X"3E",X"01",X"CD",X"A4",X"14",
		X"C3",X"30",X"07",X"3A",X"27",X"86",X"B7",X"C8",X"CD",X"2E",X"17",X"0E",X"0A",X"11",X"13",X"81",
		X"E5",X"D5",X"06",X"03",X"1A",X"BE",X"38",X"11",X"20",X"04",X"13",X"23",X"10",X"F6",X"D1",X"21",
		X"06",X"00",X"19",X"EB",X"E1",X"0D",X"20",X"E8",X"C9",X"D1",X"D5",X"CD",X"66",X"17",X"0D",X"28",
		X"16",X"06",X"00",X"21",X"00",X"00",X"09",X"29",X"09",X"29",X"E5",X"19",X"2B",X"54",X"5D",X"01",
		X"06",X"00",X"09",X"EB",X"C1",X"ED",X"B8",X"D1",X"E1",X"01",X"03",X"00",X"ED",X"B0",X"D5",X"CD",
		X"83",X"05",X"CD",X"BC",X"0A",X"CD",X"A7",X"06",X"DF",X"1A",X"CF",X"20",X"28",X"43",X"4F",X"4E",
		X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"00",X"21",X"28",X"D8",X"11",X"27",X"86",X"06",X"01",X"CD",X"28",X"05",X"E7",
		X"0F",X"07",X"04",X"CF",X"28",X"38",X"59",X"4F",X"55",X"20",X"20",X"48",X"41",X"56",X"45",X"20",
		X"20",X"4A",X"4F",X"49",X"4E",X"45",X"44",X"20",X"20",X"54",X"48",X"45",X"00",X"CF",X"30",X"48",
		X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"20",X"44",X"52",X"49",X"56",
		X"45",X"52",X"53",X"00",X"CF",X"50",X"58",X"48",X"41",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"46",
		X"41",X"4D",X"45",X"00",X"E7",X"03",X"0F",X"05",X"CF",X"28",X"78",X"45",X"4E",X"54",X"45",X"52",
		X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"20",X"5B",
		X"00",X"CF",X"70",X"88",X"5B",X"5B",X"5B",X"00",X"E7",X"03",X"16",X"07",X"CF",X"10",X"B0",X"55",
		X"53",X"45",X"20",X"53",X"54",X"49",X"43",X"4B",X"20",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",
		X"47",X"45",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"00",X"CF",X"10",X"C0",X"54",X"48",X"45",
		X"4E",X"20",X"50",X"52",X"45",X"53",X"53",X"20",X"53",X"41",X"57",X"20",X"54",X"4F",X"20",X"53",
		X"54",X"4F",X"52",X"45",X"20",X"49",X"54",X"00",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",
		X"FB",X"21",X"88",X"70",X"CD",X"DA",X"04",X"D1",X"06",X"03",X"0E",X"41",X"3E",X"FF",X"32",X"1A",
		X"86",X"CD",X"3B",X"17",X"20",X"FB",X"79",X"E5",X"CD",X"6B",X"05",X"C5",X"3E",X"09",X"CD",X"CF",
		X"14",X"C1",X"E1",X"3A",X"1A",X"86",X"3D",X"32",X"1A",X"86",X"C8",X"CD",X"3B",X"17",X"20",X"05",
		X"CD",X"41",X"17",X"18",X"DC",X"79",X"12",X"13",X"CD",X"6B",X"05",X"10",X"CF",X"C9",X"3A",X"27",
		X"86",X"FE",X"02",X"21",X"52",X"81",X"C8",X"21",X"4F",X"81",X"C9",X"3A",X"0F",X"86",X"E6",X"08",
		X"C9",X"F5",X"D5",X"3A",X"0F",X"86",X"57",X"79",X"CB",X"62",X"28",X"0A",X"C6",X"01",X"FE",X"5B",
		X"38",X"10",X"3E",X"40",X"18",X"0C",X"CB",X"6A",X"28",X"08",X"D6",X"01",X"FE",X"40",X"30",X"02",
		X"3E",X"5A",X"4F",X"D1",X"F1",X"C9",X"79",X"FE",X"0A",X"3E",X"0F",X"CA",X"0C",X"08",X"3E",X"0F",
		X"C3",X"0C",X"08",X"3A",X"1F",X"86",X"B7",X"C0",X"3E",X"FF",X"32",X"1D",X"86",X"1E",X"04",X"CD",
		X"2E",X"17",X"23",X"23",X"23",X"CB",X"38",X"08",X"04",X"2B",X"1D",X"10",X"FC",X"08",X"30",X"08",
		X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"79",X"86",X"27",X"77",X"D0",X"2B",X"1D",X"C8",
		X"0E",X"01",X"18",X"F4",X"21",X"28",X"86",X"7E",X"C6",X"01",X"27",X"77",X"3E",X"05",X"CD",X"0C",
		X"08",X"AF",X"C9",X"CD",X"83",X"05",X"3E",X"00",X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"FF",
		X"32",X"03",X"A8",X"CD",X"4D",X"06",X"CD",X"6F",X"06",X"DF",X"02",X"CF",X"40",X"00",X"53",X"54",
		X"45",X"52",X"4E",X"20",X"20",X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"00",X"DF",X"14",
		X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"E7",
		X"07",X"04",X"07",X"CF",X"10",X"20",X"41",X"56",X"4F",X"49",X"44",X"20",X"54",X"48",X"45",X"20",
		X"52",X"4F",X"42",X"42",X"45",X"52",X"53",X"20",X"41",X"4E",X"44",X"20",X"4F",X"54",X"48",X"45",
		X"52",X"00",X"CF",X"20",X"30",X"48",X"41",X"5A",X"41",X"52",X"44",X"53",X"20",X"20",X"50",X"49",
		X"43",X"4B",X"20",X"55",X"50",X"20",X"41",X"4C",X"4C",X"20",X"54",X"48",X"45",X"00",X"CF",X"18",
		X"40",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"53",X"20",X"59",X"4F",X"55",X"20",X"43",X"41",X"4E",
		X"20",X"41",X"4E",X"44",X"20",X"47",X"45",X"54",X"20",X"49",X"54",X"00",X"CF",X"28",X"50",X"54",
		X"4F",X"20",X"54",X"48",X"45",X"20",X"42",X"41",X"4E",X"4B",X"20",X"46",X"4F",X"52",X"20",X"42",
		X"4F",X"4E",X"55",X"53",X"00",X"CD",X"3F",X"19",X"CF",X"20",X"C0",X"5B",X"5B",X"5B",X"5B",X"20",
		X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"4D",X"45",X"44",X"20",X"42",X"59",X"20",X"5B",X"5B",
		X"5B",X"5B",X"00",X"CF",X"10",X"D0",X"43",X"48",X"52",X"49",X"53",X"20",X"4F",X"42",X"45",X"52",
		X"54",X"48",X"5B",X"5B",X"47",X"55",X"4E",X"41",X"52",X"53",X"20",X"4C",X"49",X"43",X"49",X"54",
		X"49",X"53",X"00",X"06",X"05",X"C5",X"DF",X"10",X"E7",X"0C",X"0B",X"07",X"3E",X"05",X"CD",X"CF",
		X"14",X"DF",X"11",X"E7",X"0C",X"0B",X"06",X"3E",X"05",X"CD",X"CF",X"14",X"DF",X"12",X"E7",X"0C",
		X"0B",X"05",X"3E",X"05",X"CD",X"CF",X"14",X"DF",X"13",X"E7",X"0C",X"0B",X"04",X"3E",X"05",X"CD",
		X"CF",X"14",X"DF",X"14",X"E7",X"0C",X"0B",X"03",X"3E",X"05",X"CD",X"CF",X"14",X"DF",X"15",X"E7",
		X"0C",X"0B",X"02",X"3E",X"05",X"CD",X"CF",X"14",X"DF",X"16",X"E7",X"0C",X"0B",X"01",X"3E",X"05",
		X"CD",X"CF",X"14",X"DF",X"17",X"E7",X"0C",X"0B",X"00",X"3E",X"05",X"CD",X"CF",X"14",X"C1",X"10",
		X"A4",X"CF",X"20",X"C0",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CF",X"10",X"D0",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"C3",X"30",X"07",X"11",
		X"8B",X"88",X"21",X"FB",X"19",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"AB",X"88",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"CB",X"88",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"EB",X"88",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"0B",X"89",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"2B",X"89",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"4B",X"89",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"6B",X"89",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"8B",X"89",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"AB",X"89",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"CB",X"89",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"EB",X"89",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"0B",X"8A",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"2B",X"8A",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"4B",X"8A",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"6B",X"8A",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"8B",X"8A",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"AB",X"8A",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"CB",X"8A",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"EB",X"8A",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"0B",X"8B",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"2B",X"8B",X"01",X"0C",X"00",
		X"ED",X"B0",X"11",X"4B",X"8B",X"01",X"0C",X"00",X"ED",X"B0",X"C9",X"10",X"10",X"10",X"10",X"10",
		X"F5",X"F4",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"F5",X"F6",X"F6",X"F4",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"F5",X"F6",X"F6",X"F6",X"F6",X"F4",X"10",X"10",X"10",X"10",
		X"10",X"F5",X"F6",X"F6",X"10",X"10",X"F6",X"F6",X"F4",X"10",X"10",X"10",X"F5",X"F6",X"F6",X"F6",
		X"10",X"23",X"F6",X"F6",X"F6",X"F4",X"10",X"84",X"85",X"85",X"F6",X"F6",X"1F",X"1B",X"F6",X"F6",
		X"85",X"85",X"C8",X"10",X"10",X"10",X"79",X"F6",X"24",X"1E",X"F6",X"7B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"79",X"F6",X"10",X"11",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",
		X"29",X"12",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"11",X"10",X"F6",X"7B",
		X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"27",X"15",X"F6",X"7B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"79",X"F6",X"10",X"18",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",
		X"23",X"24",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"19",X"10",X"F6",X"7B",
		X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"18",X"1F",X"F6",X"7B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"79",X"F6",X"24",X"24",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",
		X"10",X"10",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"1F",X"24",X"F6",X"7B",
		X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"17",X"15",X"F6",X"7B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"79",X"F6",X"10",X"17",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",
		X"10",X"10",X"F6",X"7B",X"10",X"10",X"10",X"10",X"10",X"10",X"79",X"F6",X"F6",X"F6",X"F6",X"7B",
		X"10",X"10",X"10",X"10",X"10",X"10",X"86",X"85",X"85",X"85",X"85",X"7A",X"10",X"10",X"10",X"CD",
		X"A8",X"46",X"AF",X"32",X"27",X"86",X"32",X"39",X"86",X"21",X"22",X"86",X"06",X"01",X"70",X"21",
		X"27",X"86",X"36",X"01",X"23",X"CD",X"4B",X"30",X"23",X"36",X"00",X"23",X"36",X"01",X"3E",X"00",
		X"32",X"92",X"86",X"21",X"9D",X"8A",X"22",X"95",X"86",X"3E",X"04",X"32",X"30",X"86",X"CD",X"AD",
		X"30",X"CD",X"08",X"0A",X"CD",X"FA",X"05",X"3E",X"00",X"32",X"1F",X"86",X"CD",X"0C",X"08",X"3E",
		X"FF",X"32",X"9A",X"86",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",
		X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",X"07",X"CF",X"20",X"30",X"59",
		X"4F",X"55",X"20",X"43",X"41",X"4E",X"20",X"4F",X"4E",X"4C",X"59",X"20",X"47",X"4F",X"20",X"54",
		X"48",X"52",X"55",X"20",X"41",X"4E",X"00",X"CF",X"30",X"40",X"49",X"4E",X"54",X"45",X"52",X"53",
		X"45",X"43",X"54",X"49",X"4F",X"4E",X"20",X"49",X"4E",X"20",X"54",X"48",X"45",X"00",X"CF",X"20",
		X"50",X"44",X"49",X"52",X"45",X"43",X"54",X"49",X"4F",X"4E",X"20",X"54",X"48",X"41",X"54",X"20",
		X"54",X"48",X"45",X"20",X"41",X"52",X"52",X"4F",X"57",X"00",X"CF",X"18",X"60",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"20",X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"46",X"45",X"57",X"20",X"53",
		X"45",X"43",X"4F",X"4E",X"44",X"53",X"00",X"CF",X"28",X"70",X"54",X"48",X"45",X"20",X"41",X"52",
		X"52",X"4F",X"57",X"53",X"20",X"57",X"49",X"4C",X"4C",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",
		X"00",X"CD",X"D3",X"26",X"CD",X"E3",X"46",X"3E",X"4C",X"32",X"D3",X"8A",X"32",X"D3",X"89",X"3E",
		X"4D",X"32",X"53",X"8A",X"32",X"53",X"89",X"3E",X"05",X"CD",X"A4",X"14",X"DF",X"9F",X"3E",X"06",
		X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"DF",X"9C",X"3E",X"4D",X"32",X"D3",X"8A",X"32",
		X"D3",X"89",X"3E",X"4C",X"32",X"53",X"8A",X"32",X"53",X"89",X"3E",X"03",X"CD",X"A4",X"14",X"DF",
		X"9F",X"3E",X"06",X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"DF",X"9C",X"3E",X"4C",X"32",
		X"D3",X"8A",X"32",X"D3",X"89",X"3E",X"4D",X"32",X"53",X"8A",X"32",X"53",X"89",X"3E",X"00",X"CD",
		X"0C",X"08",X"3E",X"02",X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",
		X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",X"04",X"CF",
		X"28",X"30",X"44",X"52",X"4F",X"50",X"20",X"41",X"20",X"53",X"41",X"57",X"48",X"4F",X"52",X"53",
		X"45",X"20",X"54",X"4F",X"20",X"47",X"4F",X"00",X"CF",X"30",X"40",X"54",X"48",X"52",X"55",X"20",
		X"41",X"4E",X"20",X"49",X"4E",X"54",X"45",X"52",X"53",X"45",X"43",X"54",X"49",X"4F",X"4E",X"00",
		X"CF",X"28",X"50",X"4F",X"52",X"20",X"54",X"4F",X"20",X"42",X"4C",X"4F",X"57",X"20",X"55",X"50",
		X"20",X"41",X"20",X"52",X"4F",X"42",X"42",X"45",X"52",X"00",X"CF",X"30",X"60",X"42",X"4C",X"4F",
		X"57",X"49",X"4E",X"47",X"20",X"55",X"50",X"20",X"41",X"20",X"52",X"4F",X"42",X"42",X"45",X"52",
		X"00",X"CF",X"30",X"70",X"53",X"43",X"4F",X"52",X"45",X"53",X"20",X"20",X"32",X"30",X"30",X"20",
		X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"CD",X"D3",X"26",X"CD",X"E3",X"46",X"3E",X"4C",
		X"32",X"D3",X"89",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",X"32",
		X"42",X"90",X"3E",X"93",X"32",X"43",X"90",X"32",X"47",X"90",X"DD",X"21",X"40",X"90",X"3E",X"0C",
		X"32",X"45",X"90",X"3E",X"03",X"32",X"46",X"90",X"06",X"25",X"0E",X"01",X"16",X"36",X"3E",X"07",
		X"CD",X"0C",X"08",X"1E",X"30",X"DD",X"70",X"00",X"DD",X"71",X"04",X"C5",X"DD",X"E5",X"3E",X"01",
		X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"3E",X"66",X"B8",X"20",X"0A",X"3E",X"02",X"CD",X"0C",
		X"08",X"3E",X"2F",X"32",X"53",X"8A",X"3E",X"66",X"B9",X"28",X"01",X"0C",X"3E",X"66",X"B9",X"20",
		X"1C",X"1D",X"7B",X"B7",X"C2",X"5C",X"1D",X"3E",X"00",X"DD",X"77",X"04",X"DD",X"72",X"05",X"14",
		X"3E",X"39",X"BA",X"20",X"08",X"3E",X"36",X"57",X"3E",X"10",X"32",X"53",X"8A",X"3E",X"86",X"B8",
		X"20",X"0A",X"3E",X"02",X"CD",X"0C",X"08",X"3E",X"2F",X"32",X"D3",X"89",X"3E",X"F1",X"B8",X"20",
		X"A4",X"3E",X"00",X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",
		X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",
		X"09",X"06",X"01",X"CF",X"30",X"30",X"55",X"53",X"45",X"20",X"54",X"48",X"45",X"20",X"53",X"45",
		X"43",X"4F",X"4E",X"44",X"20",X"47",X"45",X"41",X"52",X"00",X"CF",X"20",X"40",X"42",X"55",X"54",
		X"54",X"4F",X"4E",X"20",X"54",X"4F",X"20",X"47",X"45",X"54",X"20",X"41",X"57",X"41",X"59",X"20",
		X"46",X"52",X"4F",X"4D",X"00",X"CF",X"60",X"50",X"41",X"20",X"52",X"4F",X"42",X"42",X"45",X"52",
		X"00",X"CD",X"D3",X"26",X"CD",X"E3",X"46",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",
		X"90",X"3E",X"07",X"32",X"42",X"90",X"3E",X"93",X"32",X"43",X"90",X"32",X"47",X"90",X"DD",X"21",
		X"40",X"90",X"3E",X"0C",X"32",X"45",X"90",X"3E",X"03",X"32",X"46",X"90",X"06",X"25",X"0E",X"01",
		X"3E",X"07",X"CD",X"0C",X"08",X"DD",X"70",X"00",X"DD",X"71",X"04",X"C5",X"DD",X"E5",X"3E",X"01",
		X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"0C",X"3E",X"78",X"B8",X"30",X"06",X"04",X"3E",X"08",
		X"CD",X"0C",X"08",X"3E",X"F0",X"B8",X"30",X"07",X"06",X"F1",X"3E",X"00",X"CD",X"0C",X"08",X"3E",
		X"F1",X"B9",X"20",X"D1",X"3E",X"00",X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"CD",X"83",
		X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",
		X"DF",X"13",X"E7",X"09",X"06",X"05",X"CF",X"18",X"30",X"50",X"49",X"43",X"4B",X"49",X"4E",X"47",
		X"20",X"55",X"50",X"20",X"54",X"48",X"45",X"20",X"4D",X"4F",X"4E",X"45",X"59",X"20",X"47",X"49",
		X"56",X"45",X"53",X"00",X"CF",X"48",X"40",X"59",X"4F",X"55",X"20",X"31",X"30",X"30",X"20",X"50",
		X"4F",X"49",X"4E",X"54",X"53",X"00",X"CF",X"38",X"50",X"45",X"56",X"45",X"52",X"59",X"20",X"46",
		X"4F",X"55",X"52",X"20",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"53",X"00",X"CF",X"30",X"60",X"59",
		X"4F",X"55",X"20",X"47",X"45",X"54",X"20",X"54",X"4F",X"20",X"54",X"48",X"45",X"20",X"42",X"41",
		X"4E",X"4B",X"00",X"CF",X"28",X"70",X"47",X"49",X"56",X"45",X"53",X"20",X"59",X"4F",X"55",X"20",
		X"4F",X"4E",X"45",X"20",X"53",X"41",X"57",X"48",X"4F",X"52",X"53",X"45",X"00",X"CD",X"D3",X"26",
		X"CD",X"E3",X"46",X"3E",X"4F",X"32",X"D3",X"8A",X"32",X"53",X"8A",X"32",X"D3",X"89",X"32",X"53",
		X"89",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",X"32",X"42",X"90",
		X"3E",X"93",X"32",X"43",X"90",X"DD",X"21",X"40",X"90",X"06",X"01",X"3E",X"07",X"CD",X"0C",X"08",
		X"DD",X"70",X"00",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"3E",
		X"46",X"B8",X"20",X"0A",X"3E",X"04",X"CD",X"0C",X"08",X"3E",X"10",X"32",X"D3",X"8A",X"3E",X"66",
		X"B8",X"20",X"0A",X"3E",X"04",X"CD",X"0C",X"08",X"3E",X"10",X"32",X"53",X"8A",X"3E",X"86",X"B8",
		X"20",X"0A",X"3E",X"04",X"CD",X"0C",X"08",X"3E",X"10",X"32",X"D3",X"89",X"3E",X"A6",X"B8",X"20",
		X"0A",X"3E",X"04",X"CD",X"0C",X"08",X"3E",X"10",X"32",X"53",X"89",X"3E",X"F1",X"B8",X"C2",X"10",
		X"1F",X"3E",X"00",X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",
		X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",
		X"09",X"06",X"06",X"CF",X"28",X"30",X"54",X"48",X"45",X"20",X"53",X"54",X"45",X"41",X"4D",X"20",
		X"52",X"4F",X"4C",X"4C",X"45",X"52",X"20",X"57",X"49",X"4C",X"4C",X"00",X"CF",X"18",X"40",X"43",
		X"48",X"41",X"4E",X"47",X"45",X"20",X"41",X"52",X"52",X"4F",X"57",X"20",X"49",X"4E",X"54",X"45",
		X"52",X"53",X"45",X"43",X"54",X"49",X"4F",X"4E",X"53",X"00",X"CF",X"18",X"50",X"54",X"4F",X"20",
		X"53",X"41",X"57",X"48",X"4F",X"52",X"53",X"45",X"53",X"20",X"20",X"59",X"4F",X"55",X"20",X"43",
		X"41",X"4E",X"20",X"50",X"41",X"53",X"53",X"00",X"CF",X"38",X"60",X"54",X"48",X"52",X"55",X"20",
		X"54",X"48",X"45",X"20",X"53",X"41",X"57",X"48",X"4F",X"52",X"53",X"45",X"53",X"00",X"CF",X"30",
		X"70",X"42",X"55",X"54",X"20",X"54",X"48",X"45",X"20",X"52",X"4F",X"42",X"42",X"45",X"52",X"53",
		X"20",X"43",X"41",X"4E",X"54",X"00",X"CD",X"D3",X"26",X"CD",X"E3",X"46",X"3E",X"4C",X"32",X"53",
		X"8A",X"3C",X"32",X"D3",X"89",X"3E",X"4F",X"32",X"53",X"89",X"3E",X"06",X"CD",X"A4",X"14",X"3E",
		X"2B",X"32",X"41",X"90",X"3E",X"02",X"32",X"42",X"90",X"3E",X"93",X"32",X"43",X"90",X"DD",X"21",
		X"40",X"90",X"06",X"F1",X"0E",X"2B",X"DD",X"70",X"00",X"DD",X"71",X"01",X"C5",X"DD",X"E5",X"3E",
		X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"05",X"0D",X"3E",X"27",X"B9",X"20",X"02",X"0E",X"2B",
		X"3E",X"86",X"B8",X"20",X"05",X"3E",X"2F",X"32",X"D3",X"89",X"3E",X"66",X"B8",X"20",X"05",X"3E",
		X"2F",X"32",X"53",X"8A",X"3E",X"00",X"B8",X"20",X"CD",X"3E",X"00",X"CD",X"0C",X"08",X"3E",X"01",
		X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",
		X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",X"07",X"CF",X"20",X"30",X"54",X"48",
		X"45",X"20",X"53",X"54",X"52",X"45",X"45",X"54",X"20",X"53",X"57",X"45",X"45",X"50",X"45",X"52",
		X"20",X"57",X"49",X"4C",X"4C",X"00",X"CF",X"30",X"40",X"53",X"57",X"45",X"45",X"50",X"20",X"55",
		X"50",X"20",X"41",X"52",X"52",X"4F",X"57",X"53",X"20",X"41",X"4E",X"44",X"00",X"CF",X"58",X"50",
		X"53",X"41",X"57",X"48",X"4F",X"52",X"53",X"45",X"53",X"00",X"CD",X"D3",X"26",X"CD",X"E3",X"46",
		X"3E",X"4C",X"32",X"D3",X"8A",X"3C",X"32",X"53",X"8A",X"3E",X"4F",X"32",X"D3",X"89",X"3E",X"2F",
		X"32",X"53",X"89",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"AC",X"32",X"41",X"90",X"3E",X"07",X"32",
		X"42",X"90",X"3E",X"93",X"32",X"43",X"90",X"DD",X"21",X"40",X"90",X"06",X"F1",X"0E",X"AC",X"DD",
		X"70",X"00",X"DD",X"71",X"01",X"C5",X"DD",X"E5",X"3E",X"02",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",
		X"05",X"0C",X"3E",X"AE",X"B9",X"20",X"02",X"0E",X"B0",X"3E",X"B2",X"B9",X"20",X"02",X"0E",X"AC",
		X"3E",X"A6",X"B8",X"20",X"05",X"3E",X"10",X"32",X"53",X"89",X"3E",X"66",X"B8",X"20",X"05",X"3E",
		X"10",X"32",X"53",X"8A",X"3E",X"46",X"B8",X"20",X"05",X"3E",X"10",X"32",X"D3",X"8A",X"3E",X"00",
		X"B8",X"20",X"BC",X"3E",X"00",X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"CD",X"83",X"05",
		X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"DF",
		X"13",X"E7",X"09",X"06",X"03",X"CF",X"20",X"30",X"4B",X"45",X"45",X"50",X"20",X"41",X"4E",X"20",
		X"45",X"59",X"45",X"20",X"4F",X"4E",X"20",X"54",X"48",X"45",X"20",X"46",X"55",X"45",X"4C",X"00",
		X"CF",X"28",X"40",X"54",X"48",X"45",X"52",X"45",X"20",X"41",X"52",X"45",X"20",X"54",X"57",X"4F",
		X"20",X"46",X"55",X"45",X"4C",X"49",X"4E",X"47",X"00",X"CF",X"28",X"50",X"53",X"54",X"41",X"54",
		X"49",X"4F",X"4E",X"53",X"20",X"42",X"45",X"54",X"57",X"45",X"45",X"4E",X"20",X"45",X"41",X"43",
		X"48",X"00",X"CF",X"28",X"60",X"42",X"41",X"4E",X"4B",X"20",X"20",X"55",X"53",X"45",X"20",X"54",
		X"48",X"45",X"4D",X"20",X"57",X"49",X"53",X"45",X"4C",X"59",X"00",X"CD",X"E8",X"27",X"CD",X"D3",
		X"26",X"CD",X"E3",X"46",X"3E",X"CD",X"32",X"B2",X"89",X"3E",X"CE",X"32",X"B3",X"89",X"3E",X"CF",
		X"32",X"B4",X"89",X"3E",X"CC",X"32",X"D2",X"89",X"3E",X"D0",X"32",X"D3",X"89",X"3E",X"D1",X"32",
		X"D4",X"89",X"3E",X"CB",X"32",X"F2",X"89",X"3E",X"D2",X"32",X"F3",X"89",X"3E",X"D3",X"32",X"F4",
		X"89",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",X"32",X"42",X"90",
		X"3E",X"93",X"32",X"43",X"90",X"DD",X"21",X"40",X"90",X"06",X"01",X"3E",X"07",X"CD",X"0C",X"08",
		X"DD",X"70",X"00",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"3E",
		X"86",X"B8",X"20",X"10",X"3E",X"09",X"CD",X"0C",X"08",X"21",X"D3",X"89",X"CD",X"68",X"2D",X"C5",
		X"CD",X"C8",X"27",X"C1",X"3E",X"F1",X"B8",X"C2",X"20",X"22",X"3E",X"00",X"CD",X"0C",X"08",X"3E",
		X"01",X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",
		X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",X"01",X"CF",X"20",X"30",X"59",
		X"4F",X"55",X"20",X"47",X"45",X"54",X"20",X"41",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"41",
		X"52",X"4D",X"4F",X"52",X"45",X"44",X"00",X"CF",X"40",X"40",X"43",X"41",X"52",X"20",X"41",X"54",
		X"20",X"42",X"41",X"4E",X"4B",X"20",X"46",X"4F",X"55",X"52",X"00",X"CF",X"48",X"50",X"41",X"4E",
		X"44",X"20",X"42",X"41",X"4E",X"4B",X"20",X"45",X"49",X"47",X"48",X"54",X"00",X"E7",X"0A",X"0E",
		X"05",X"CD",X"6F",X"06",X"CD",X"4D",X"06",X"21",X"B0",X"89",X"11",X"1A",X"00",X"36",X"62",X"23",
		X"36",X"65",X"23",X"36",X"65",X"23",X"36",X"65",X"23",X"36",X"65",X"23",X"36",X"65",X"23",X"36",
		X"6E",X"19",X"36",X"61",X"23",X"36",X"64",X"23",X"36",X"64",X"23",X"36",X"6D",X"23",X"36",X"66",
		X"23",X"36",X"66",X"23",X"36",X"68",X"19",X"36",X"61",X"23",X"36",X"64",X"23",X"36",X"64",X"23",
		X"36",X"6C",X"23",X"36",X"66",X"23",X"36",X"66",X"23",X"36",X"68",X"19",X"36",X"61",X"23",X"36",
		X"64",X"23",X"36",X"64",X"23",X"36",X"6B",X"23",X"36",X"66",X"23",X"36",X"66",X"23",X"36",X"68",
		X"19",X"36",X"61",X"23",X"36",X"64",X"23",X"36",X"64",X"23",X"36",X"6A",X"23",X"36",X"66",X"23",
		X"36",X"66",X"23",X"36",X"68",X"19",X"36",X"61",X"23",X"36",X"64",X"23",X"36",X"64",X"23",X"36",
		X"69",X"23",X"36",X"66",X"23",X"36",X"66",X"23",X"36",X"68",X"19",X"36",X"60",X"23",X"36",X"63",
		X"23",X"36",X"63",X"23",X"36",X"63",X"23",X"36",X"63",X"23",X"36",X"63",X"23",X"36",X"67",X"3E",
		X"04",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",X"32",X"42",X"90",X"3E",X"93",
		X"32",X"43",X"90",X"DD",X"21",X"40",X"90",X"06",X"01",X"DD",X"70",X"00",X"C5",X"DD",X"E5",X"3E",
		X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"3E",X"76",X"B8",X"20",X"EC",X"3E",X"00",X"DD",
		X"77",X"00",X"06",X"05",X"C5",X"E7",X"0A",X"0E",X"01",X"3E",X"03",X"CD",X"CF",X"14",X"E7",X"0A",
		X"0E",X"02",X"3E",X"03",X"CD",X"CF",X"14",X"E7",X"0A",X"0E",X"03",X"3E",X"03",X"CD",X"CF",X"14",
		X"E7",X"0A",X"0E",X"04",X"3E",X"03",X"CD",X"CF",X"14",X"E7",X"0A",X"0E",X"06",X"3E",X"03",X"CD",
		X"CF",X"14",X"E7",X"0A",X"0E",X"05",X"3E",X"03",X"CD",X"CF",X"14",X"C1",X"10",X"C6",X"3E",X"01",
		X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",X"45",X"44",
		X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",X"04",X"CF",X"38",X"30",X"57",X"41",
		X"54",X"43",X"48",X"20",X"4F",X"55",X"54",X"20",X"46",X"4F",X"52",X"20",X"54",X"48",X"45",X"00",
		X"CF",X"28",X"40",X"41",X"4D",X"42",X"55",X"4C",X"41",X"4E",X"43",X"45",X"20",X"20",X"49",X"46",
		X"20",X"49",X"54",X"20",X"43",X"4F",X"4D",X"45",X"53",X"00",X"CF",X"28",X"50",X"4F",X"55",X"54",
		X"20",X"4F",X"4E",X"20",X"59",X"4F",X"55",X"52",X"20",X"53",X"54",X"52",X"45",X"45",X"54",X"20",
		X"47",X"45",X"54",X"00",X"CF",X"30",X"60",X"4F",X"46",X"46",X"20",X"54",X"48",X"41",X"54",X"20",
		X"53",X"54",X"52",X"45",X"45",X"54",X"20",X"46",X"41",X"53",X"54",X"00",X"CD",X"D3",X"26",X"3E",
		X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",X"32",X"42",X"90",X"3E",X"93",
		X"32",X"43",X"90",X"32",X"47",X"90",X"DD",X"21",X"40",X"90",X"3E",X"AF",X"32",X"45",X"90",X"3E",
		X"02",X"32",X"46",X"90",X"06",X"01",X"0E",X"02",X"DD",X"70",X"00",X"C5",X"DD",X"E5",X"3E",X"01",
		X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"3E",X"56",X"B8",X"20",X"EC",X"3E",X"10",X"CD",X"0C",
		X"08",X"0C",X"0C",X"04",X"DD",X"70",X"00",X"DD",X"71",X"04",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",
		X"CF",X"14",X"DD",X"E1",X"C1",X"3E",X"86",X"B8",X"20",X"E7",X"3E",X"F9",X"32",X"41",X"90",X"06",
		X"93",X"DD",X"71",X"04",X"DD",X"70",X"03",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",
		X"E1",X"C1",X"0C",X"0C",X"3E",X"D6",X"B8",X"38",X"01",X"04",X"3E",X"F0",X"B9",X"30",X"E2",X"3E",
		X"00",X"CD",X"0C",X"08",X"3E",X"01",X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",
		X"52",X"4D",X"4F",X"52",X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",
		X"01",X"CF",X"30",X"30",X"50",X"49",X"43",X"4B",X"20",X"55",X"50",X"20",X"54",X"48",X"45",X"20",
		X"4B",X"45",X"59",X"20",X"41",X"4E",X"44",X"00",X"CF",X"40",X"40",X"42",X"52",X"49",X"4E",X"47",
		X"20",X"49",X"54",X"20",X"54",X"4F",X"20",X"54",X"48",X"45",X"00",X"CF",X"48",X"50",X"4C",X"4F",
		X"43",X"4B",X"20",X"46",X"4F",X"52",X"20",X"20",X"31",X"30",X"30",X"30",X"00",X"CF",X"50",X"60",
		X"42",X"4F",X"4E",X"55",X"53",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"CD",X"D3",X"26",
		X"3E",X"CA",X"32",X"52",X"8A",X"3E",X"C9",X"32",X"53",X"8A",X"3E",X"4E",X"32",X"52",X"89",X"3E",
		X"2D",X"32",X"53",X"89",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",
		X"32",X"42",X"90",X"3E",X"93",X"32",X"43",X"90",X"DD",X"21",X"40",X"90",X"06",X"25",X"3E",X"07",
		X"CD",X"0C",X"08",X"DD",X"70",X"00",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",X"E1",
		X"C1",X"04",X"3E",X"66",X"B8",X"20",X"0D",X"3E",X"10",X"32",X"52",X"8A",X"32",X"53",X"8A",X"3E",
		X"13",X"CD",X"0C",X"08",X"3E",X"A6",X"B8",X"20",X"0D",X"3E",X"10",X"32",X"52",X"89",X"32",X"53",
		X"89",X"3E",X"13",X"CD",X"0C",X"08",X"3E",X"F1",X"B8",X"20",X"C8",X"3E",X"00",X"CD",X"0C",X"08",
		X"3E",X"01",X"CD",X"A4",X"14",X"CD",X"83",X"05",X"CF",X"50",X"10",X"41",X"52",X"4D",X"4F",X"52",
		X"45",X"44",X"20",X"43",X"41",X"52",X"00",X"DF",X"13",X"E7",X"09",X"06",X"04",X"CF",X"30",X"30",
		X"43",X"52",X"41",X"53",X"48",X"20",X"54",X"48",X"45",X"20",X"54",X"4E",X"54",X"20",X"54",X"52",
		X"55",X"43",X"4B",X"00",X"CF",X"38",X"40",X"49",X"4E",X"54",X"4F",X"20",X"54",X"48",X"45",X"20",
		X"57",X"41",X"4C",X"4C",X"20",X"46",X"4F",X"52",X"00",X"CF",X"38",X"50",X"31",X"30",X"30",X"30",
		X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"CD",X"D3",
		X"26",X"3E",X"06",X"CD",X"A4",X"14",X"3E",X"3C",X"32",X"41",X"90",X"3E",X"07",X"32",X"42",X"90",
		X"3E",X"93",X"32",X"43",X"90",X"32",X"47",X"90",X"DD",X"21",X"40",X"90",X"3E",X"27",X"32",X"45",
		X"90",X"3E",X"05",X"32",X"46",X"90",X"06",X"01",X"0E",X"F0",X"3E",X"07",X"CD",X"0C",X"08",X"DD",
		X"70",X"00",X"DD",X"71",X"04",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",
		X"04",X"0D",X"3E",X"46",X"B8",X"20",X"E8",X"3E",X"F9",X"32",X"41",X"90",X"06",X"93",X"DD",X"71",
		X"04",X"DD",X"70",X"03",X"C5",X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"0D",
		X"3E",X"B6",X"B8",X"38",X"01",X"04",X"3E",X"46",X"B9",X"20",X"E3",X"3E",X"3C",X"32",X"41",X"90",
		X"3E",X"66",X"32",X"45",X"90",X"06",X"46",X"0E",X"93",X"DD",X"71",X"07",X"DD",X"70",X"00",X"C5",
		X"DD",X"E5",X"3E",X"01",X"CD",X"CF",X"14",X"DD",X"E1",X"C1",X"04",X"0C",X"3E",X"C0",X"B9",X"20",
		X"E8",X"3E",X"38",X"32",X"45",X"90",X"3E",X"0E",X"CD",X"0C",X"08",X"3E",X"06",X"CD",X"CF",X"14",
		X"3E",X"37",X"32",X"45",X"90",X"3E",X"06",X"CD",X"CF",X"14",X"3E",X"36",X"32",X"45",X"90",X"3E",
		X"06",X"CD",X"CF",X"14",X"3E",X"38",X"32",X"45",X"90",X"3E",X"06",X"CD",X"CF",X"14",X"3E",X"37",
		X"32",X"45",X"90",X"3E",X"00",X"CD",X"0C",X"08",X"3E",X"14",X"CD",X"CF",X"14",X"3E",X"00",X"32",
		X"9A",X"86",X"C9",X"E7",X"03",X"10",X"05",X"E7",X"04",X"14",X"05",X"DF",X"9C",X"CD",X"6F",X"06",
		X"CD",X"4D",X"06",X"21",X"5F",X"27",X"11",X"F0",X"88",X"01",X"07",X"00",X"ED",X"B0",X"11",X"10",
		X"89",X"01",X"07",X"00",X"ED",X"B0",X"11",X"30",X"89",X"01",X"07",X"00",X"ED",X"B0",X"11",X"70",
		X"89",X"01",X"07",X"00",X"ED",X"B0",X"11",X"90",X"89",X"01",X"07",X"00",X"ED",X"B0",X"11",X"B0",
		X"89",X"01",X"07",X"00",X"ED",X"B0",X"11",X"F0",X"89",X"01",X"07",X"00",X"ED",X"B0",X"11",X"10",
		X"8A",X"01",X"07",X"00",X"ED",X"B0",X"11",X"30",X"8A",X"01",X"07",X"00",X"ED",X"B0",X"11",X"70",
		X"8A",X"01",X"07",X"00",X"ED",X"B0",X"11",X"90",X"8A",X"01",X"07",X"00",X"ED",X"B0",X"11",X"B0",
		X"8A",X"01",X"07",X"00",X"ED",X"B0",X"11",X"F0",X"8A",X"01",X"07",X"00",X"ED",X"B0",X"11",X"10",
		X"8B",X"01",X"07",X"00",X"ED",X"B0",X"11",X"30",X"8B",X"01",X"07",X"00",X"ED",X"B0",X"C9",X"58",
		X"52",X"5E",X"10",X"46",X"5B",X"55",X"40",X"49",X"45",X"10",X"50",X"41",X"45",X"42",X"59",X"44",
		X"10",X"4A",X"4B",X"53",X"51",X"47",X"48",X"10",X"46",X"47",X"5E",X"57",X"49",X"54",X"10",X"57",
		X"41",X"5D",X"4A",X"43",X"44",X"10",X"56",X"4B",X"44",X"46",X"47",X"5E",X"10",X"58",X"52",X"48",
		X"57",X"41",X"45",X"10",X"57",X"41",X"5D",X"4A",X"59",X"5C",X"10",X"42",X"43",X"53",X"58",X"52",
		X"5E",X"10",X"46",X"5B",X"55",X"40",X"49",X"45",X"10",X"50",X"41",X"45",X"42",X"59",X"44",X"10",
		X"4A",X"4B",X"53",X"51",X"47",X"48",X"10",X"46",X"47",X"5E",X"57",X"49",X"54",X"10",X"57",X"41",
		X"5D",X"4A",X"43",X"44",X"10",X"56",X"4B",X"44",X"3E",X"FF",X"06",X"18",X"21",X"59",X"88",X"11",
		X"20",X"00",X"77",X"19",X"10",X"FC",X"3E",X"1C",X"77",X"19",X"3E",X"15",X"77",X"19",X"3E",X"25",
		X"77",X"19",X"3E",X"16",X"77",X"DF",X"CF",X"C9",X"3E",X"F7",X"06",X"17",X"21",X"59",X"88",X"11",
		X"20",X"00",X"77",X"19",X"10",X"FC",X"3E",X"FF",X"77",X"19",X"3E",X"1C",X"77",X"19",X"3E",X"15",
		X"77",X"19",X"3E",X"25",X"77",X"19",X"3E",X"16",X"77",X"DF",X"7F",X"CD",X"6F",X"06",X"CD",X"4D",
		X"06",X"C9",X"DD",X"CB",X"00",X"6E",X"CA",X"37",X"28",X"DD",X"7E",X"03",X"FE",X"28",X"C2",X"6E",
		X"28",X"DF",X"1F",X"DF",X"3F",X"DF",X"5F",X"DF",X"7F",X"DF",X"9F",X"DF",X"BF",X"DF",X"DF",X"3E",
		X"06",X"CD",X"0C",X"08",X"C3",X"6E",X"28",X"DF",X"1C",X"DF",X"3C",X"DF",X"5C",X"DF",X"7C",X"DF",
		X"9C",X"DF",X"BC",X"DF",X"DC",X"3E",X"FF",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"21",X"6F",
		X"28",X"06",X"38",X"0E",X"4B",X"5E",X"23",X"56",X"23",X"1A",X"FE",X"4C",X"28",X"06",X"FE",X"4D",
		X"28",X"02",X"18",X"07",X"3D",X"B9",X"C2",X"6B",X"28",X"3E",X"4D",X"12",X"10",X"E7",X"C9",X"63",
		X"88",X"67",X"88",X"6B",X"88",X"6F",X"88",X"73",X"88",X"77",X"88",X"7B",X"88",X"E3",X"88",X"E7",
		X"88",X"EB",X"88",X"EF",X"88",X"F3",X"88",X"F7",X"88",X"FB",X"88",X"63",X"89",X"67",X"89",X"6B",
		X"89",X"6F",X"89",X"73",X"89",X"77",X"89",X"7B",X"89",X"E3",X"89",X"E7",X"89",X"EB",X"89",X"EF",
		X"89",X"F3",X"89",X"F7",X"89",X"FB",X"89",X"63",X"8A",X"67",X"8A",X"6B",X"8A",X"6F",X"8A",X"73",
		X"8A",X"77",X"8A",X"7B",X"8A",X"E3",X"8A",X"E7",X"8A",X"EB",X"8A",X"EF",X"8A",X"F3",X"8A",X"F7",
		X"8A",X"FB",X"8A",X"63",X"8B",X"67",X"8B",X"6B",X"8B",X"6F",X"8B",X"73",X"8B",X"77",X"8B",X"7B",
		X"8B",X"E3",X"8B",X"E7",X"8B",X"EB",X"8B",X"EF",X"8B",X"F3",X"8B",X"F7",X"8B",X"FB",X"8B",X"E0",
		X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"04",X"8D",X"02",X"10",X"08",X"04",X"8C",X"02",X"00",
		X"01",X"E5",X"28",X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"04",X"0D",X"02",X"10",X"08",X"04",
		X"0C",X"02",X"00",X"01",X"F8",X"28",X"00",X"00",X"01",X"00",X"00",X"08",X"10",X"04",X"0F",X"02",
		X"08",X"10",X"04",X"0E",X"02",X"00",X"01",X"0B",X"29",X"00",X"00",X"01",X"00",X"00",X"08",X"10",
		X"04",X"4F",X"02",X"08",X"10",X"04",X"4E",X"02",X"00",X"01",X"1E",X"29",X"00",X"00",X"01",X"00",
		X"00",X"10",X"08",X"04",X"8D",X"03",X"10",X"08",X"04",X"8C",X"03",X"00",X"01",X"31",X"29",X"00",
		X"00",X"01",X"00",X"00",X"10",X"08",X"04",X"0D",X"03",X"10",X"08",X"04",X"0C",X"03",X"00",X"01",
		X"44",X"29",X"00",X"00",X"01",X"00",X"00",X"08",X"10",X"04",X"0F",X"03",X"08",X"10",X"04",X"0E",
		X"03",X"00",X"01",X"57",X"29",X"00",X"00",X"01",X"00",X"00",X"08",X"10",X"04",X"4F",X"03",X"08",
		X"10",X"04",X"4E",X"03",X"00",X"01",X"6A",X"29",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"04",
		X"38",X"01",X"01",X"00",X"04",X"B8",X"02",X"01",X"00",X"04",X"F8",X"03",X"01",X"00",X"04",X"38",
		X"02",X"01",X"00",X"04",X"B8",X"03",X"01",X"00",X"04",X"F8",X"01",X"01",X"00",X"04",X"38",X"03",
		X"01",X"00",X"04",X"B8",X"01",X"01",X"00",X"04",X"F8",X"02",X"01",X"00",X"05",X"37",X"01",X"01",
		X"00",X"05",X"B7",X"02",X"01",X"00",X"05",X"F7",X"03",X"01",X"00",X"05",X"37",X"02",X"01",X"00",
		X"05",X"B7",X"01",X"01",X"00",X"05",X"F7",X"03",X"01",X"00",X"05",X"36",X"01",X"01",X"00",X"05",
		X"B6",X"02",X"01",X"00",X"05",X"F6",X"03",X"00",X"00",X"00",X"00",X"CD",X"C5",X"08",X"D2",X"7F",
		X"09",X"CD",X"9F",X"08",X"D2",X"7F",X"2C",X"FD",X"2A",X"DA",X"80",X"FD",X"66",X"02",X"FD",X"6E",
		X"01",X"E5",X"DD",X"E1",X"CD",X"87",X"2C",X"CD",X"AD",X"2C",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",
		X"0C",X"D6",X"FD",X"CB",X"00",X"D6",X"DD",X"E5",X"CD",X"5B",X"09",X"FD",X"E1",X"FD",X"CB",X"00",
		X"76",X"C2",X"78",X"2C",X"FD",X"CB",X"00",X"4E",X"CC",X"22",X"2A",X"FD",X"E5",X"CD",X"5B",X"09",
		X"18",X"E9",X"FD",X"CB",X"00",X"DE",X"DD",X"7E",X"0A",X"E6",X"0E",X"FE",X"02",X"C2",X"34",X"2B",
		X"DD",X"7E",X"0A",X"CB",X"67",X"CA",X"34",X"2B",X"3A",X"E5",X"80",X"47",X"DD",X"7E",X"08",X"90",
		X"47",X"E6",X"0E",X"FE",X"0C",X"C2",X"34",X"2B",X"78",X"CB",X"67",X"CA",X"34",X"2B",X"CB",X"47",
		X"28",X"03",X"DD",X"35",X"08",X"FD",X"36",X"01",X"07",X"FD",X"CB",X"00",X"CE",X"DD",X"7E",X"08",
		X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"DF",X"04",X"7E",X"FE",X"2F",X"CA",
		X"D3",X"2B",X"FE",X"4F",X"20",X"02",X"36",X"10",X"DD",X"CB",X"00",X"A6",X"CD",X"3D",X"2B",X"32",
		X"9C",X"86",X"FE",X"00",X"20",X"2A",X"2A",X"2E",X"86",X"CD",X"BF",X"2C",X"FD",X"75",X"03",X"FD",
		X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"E0",X"28",X"DD",X"CB",X"0B",
		X"5E",X"28",X"03",X"21",X"2C",X"29",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",
		X"FE",X"01",X"20",X"27",X"2A",X"2E",X"86",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",
		X"00",X"FD",X"36",X"0A",X"00",X"21",X"F3",X"28",X"DD",X"CB",X"0B",X"5E",X"28",X"03",X"21",X"3F",
		X"29",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FE",X"02",X"20",X"2A",X"2A",
		X"2E",X"86",X"CD",X"BF",X"2C",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"FD",X"36",X"03",X"00",X"FD",
		X"36",X"04",X"00",X"21",X"06",X"29",X"DD",X"CB",X"0B",X"5E",X"28",X"03",X"21",X"52",X"29",X"DD",
		X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FE",X"03",X"20",X"27",X"2A",X"2E",X"86",
		X"FD",X"75",X"09",X"FD",X"74",X"0A",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"19",
		X"29",X"DD",X"CB",X"0B",X"5E",X"28",X"03",X"21",X"65",X"29",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"9E",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"CB",X"0B",
		X"DE",X"FD",X"7E",X"06",X"E6",X"F8",X"FE",X"68",X"20",X"0E",X"3A",X"61",X"81",X"FD",X"BE",X"0C",
		X"38",X"03",X"3E",X"03",X"C9",X"3E",X"02",X"C9",X"3A",X"61",X"81",X"E6",X"F8",X"47",X"FD",X"7E",
		X"0C",X"E6",X"F8",X"B8",X"20",X"0D",X"3E",X"6D",X"FD",X"BE",X"06",X"38",X"03",X"3E",X"01",X"C9",
		X"3E",X"00",X"C9",X"CD",X"3D",X"08",X"DD",X"CB",X"0B",X"9E",X"E6",X"03",X"CD",X"98",X"2B",X"47",
		X"DD",X"7E",X"0A",X"FE",X"16",X"38",X"0A",X"FE",X"D0",X"78",X"D8",X"FE",X"03",X"C0",X"3E",X"02",
		X"C9",X"78",X"FE",X"02",X"C0",X"3E",X"03",X"C9",X"FE",X"00",X"20",X"0B",X"3A",X"9C",X"86",X"FE",
		X"01",X"3E",X"00",X"C0",X"3E",X"01",X"C9",X"FE",X"01",X"20",X"0B",X"3A",X"9C",X"86",X"FE",X"00",
		X"3E",X"01",X"C0",X"3E",X"00",X"C9",X"FE",X"02",X"20",X"0B",X"3A",X"9C",X"86",X"FE",X"03",X"3E",
		X"02",X"C0",X"3E",X"03",X"C9",X"FE",X"03",X"C0",X"3A",X"9C",X"86",X"FE",X"02",X"3E",X"03",X"C0",
		X"3E",X"02",X"C9",X"AF",X"FD",X"77",X"04",X"FD",X"77",X"03",X"FD",X"77",X"0A",X"FD",X"77",X"09",
		X"FD",X"CB",X"00",X"9E",X"C1",X"E5",X"3E",X"0E",X"CD",X"0C",X"08",X"01",X"02",X"02",X"CD",X"73",
		X"17",X"DD",X"CB",X"0C",X"96",X"DD",X"CB",X"00",X"A6",X"21",X"78",X"29",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"66",X"28",X"39",
		X"DD",X"66",X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"CB",X"00",X"76",X"20",X"2A",X"3E",
		X"FF",X"32",X"05",X"A8",X"3E",X"03",X"CD",X"AF",X"09",X"3E",X"00",X"32",X"05",X"A8",X"3E",X"04",
		X"CD",X"AF",X"09",X"3E",X"FF",X"32",X"03",X"A8",X"3E",X"02",X"CD",X"AF",X"09",X"3E",X"00",X"32",
		X"03",X"A8",X"3E",X"04",X"CD",X"AF",X"09",X"18",X"C1",X"E1",X"36",X"10",X"3E",X"00",X"32",X"03",
		X"A8",X"3E",X"00",X"32",X"05",X"A8",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"08",X"00",X"DD",X"66",
		X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"36",X"06",X"00",X"FD",X"36",X"0C",X"00",X"DD",
		X"CB",X"00",X"96",X"3E",X"FF",X"CD",X"AF",X"09",X"FD",X"CB",X"00",X"B6",X"C3",X"E7",X"29",X"CD",
		X"D5",X"09",X"CD",X"5B",X"09",X"18",X"FB",X"FD",X"36",X"08",X"EB",X"CD",X"3D",X"08",X"E6",X"E0",
		X"F6",X"13",X"FD",X"77",X"0A",X"2A",X"2E",X"86",X"CD",X"BF",X"2C",X"DD",X"74",X"04",X"DD",X"75",
		X"03",X"3E",X"00",X"32",X"9C",X"86",X"DD",X"77",X"0A",X"DD",X"77",X"09",X"C9",X"21",X"E0",X"28",
		X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"7C",
		X"2F",X"67",X"7D",X"2F",X"6F",X"23",X"C9",X"3E",X"FF",X"06",X"18",X"21",X"5F",X"88",X"11",X"20",
		X"00",X"77",X"19",X"10",X"FC",X"3E",X"1C",X"77",X"19",X"3E",X"15",X"77",X"19",X"3E",X"25",X"77",
		X"19",X"3E",X"16",X"77",X"21",X"5F",X"88",X"22",X"8F",X"86",X"3A",X"8E",X"86",X"FD",X"77",X"01",
		X"FD",X"CB",X"00",X"CE",X"DD",X"CB",X"0D",X"9E",X"DF",X"FF",X"C9",X"FD",X"7E",X"01",X"B7",X"20",
		X"66",X"3A",X"8E",X"86",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"2A",X"8F",X"86",X"E5",X"3E",
		X"8A",X"BC",X"20",X"0C",X"3E",X"9F",X"BD",X"30",X"07",X"3E",X"01",X"CD",X"0C",X"08",X"DF",X"FA",
		X"E1",X"3E",X"8B",X"BC",X"20",X"34",X"3E",X"5F",X"BD",X"20",X"2F",X"DD",X"CB",X"0D",X"DE",X"CF",
		X"10",X"F8",X"46",X"55",X"45",X"4C",X"20",X"20",X"20",X"20",X"20",X"20",X"4F",X"55",X"54",X"20",
		X"20",X"20",X"4F",X"46",X"20",X"20",X"20",X"47",X"41",X"53",X"20",X"20",X"20",X"20",X"00",X"21",
		X"3F",X"90",X"34",X"3E",X"07",X"32",X"8E",X"86",X"18",X"0D",X"35",X"7E",X"FE",X"F7",X"20",X"07",
		X"11",X"20",X"00",X"19",X"22",X"8F",X"86",X"C9",X"E5",X"D5",X"23",X"11",X"20",X"00",X"ED",X"52",
		X"3E",X"4A",X"77",X"3E",X"10",X"2B",X"77",X"3E",X"44",X"2B",X"77",X"19",X"3E",X"10",X"77",X"23",
		X"77",X"23",X"77",X"19",X"3E",X"46",X"77",X"2B",X"3E",X"10",X"77",X"2B",X"3E",X"5E",X"77",X"D1",
		X"E1",X"C9",X"CF",X"10",X"E8",X"53",X"41",X"57",X"48",X"4F",X"52",X"53",X"45",X"53",X"00",X"21",
		X"9D",X"8A",X"22",X"95",X"86",X"3A",X"30",X"86",X"B7",X"C8",X"47",X"3E",X"00",X"32",X"30",X"86",
		X"CD",X"B6",X"2D",X"10",X"FB",X"C9",X"21",X"30",X"86",X"34",X"11",X"20",X"00",X"3E",X"13",X"BE",
		X"D8",X"2A",X"95",X"86",X"B7",X"ED",X"52",X"22",X"95",X"86",X"3E",X"2F",X"18",X"1E",X"3A",X"30",
		X"86",X"B7",X"C8",X"21",X"30",X"86",X"35",X"3E",X"13",X"BE",X"D8",X"3E",X"10",X"CD",X"EC",X"2D",
		X"2A",X"95",X"86",X"11",X"20",X"00",X"19",X"22",X"95",X"86",X"3F",X"C9",X"2A",X"95",X"86",X"77",
		X"C9",X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"02",X"2B",X"02",X"10",X"08",X"02",X"2A",X"02",
		X"10",X"08",X"02",X"29",X"02",X"10",X"08",X"02",X"28",X"02",X"00",X"01",X"F6",X"2D",X"00",X"00",
		X"01",X"00",X"00",X"10",X"10",X"04",X"38",X"03",X"10",X"10",X"04",X"78",X"03",X"10",X"10",X"04",
		X"39",X"03",X"10",X"10",X"04",X"79",X"03",X"10",X"10",X"04",X"3A",X"03",X"10",X"10",X"04",X"7A",
		X"03",X"10",X"10",X"04",X"3B",X"00",X"10",X"10",X"04",X"7B",X"00",X"10",X"10",X"04",X"3A",X"00",
		X"10",X"10",X"04",X"39",X"00",X"10",X"10",X"04",X"38",X"00",X"00",X"00",X"00",X"00",X"CD",X"C5",
		X"08",X"D2",X"7F",X"09",X"DD",X"E5",X"CD",X"9F",X"08",X"D2",X"05",X"2F",X"DD",X"E5",X"3E",X"FE",
		X"CD",X"AF",X"09",X"3E",X"32",X"CD",X"AF",X"09",X"DD",X"E1",X"FD",X"E1",X"CD",X"2E",X"2F",X"CD",
		X"45",X"2F",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"FD",X"CB",X"00",X"D6",X"FD",X"36",
		X"03",X"0F",X"DD",X"E5",X"CD",X"5B",X"09",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"05",X"2F",
		X"DD",X"7E",X"0D",X"B7",X"FD",X"CB",X"00",X"76",X"C2",X"05",X"2F",X"FD",X"CB",X"00",X"4E",X"CC",
		X"A9",X"2E",X"FD",X"E5",X"CD",X"5B",X"09",X"18",X"DE",X"FD",X"CB",X"00",X"DE",X"DD",X"7E",X"0A",
		X"E6",X"0E",X"FE",X"02",X"C2",X"FC",X"2E",X"DD",X"7E",X"0A",X"CB",X"67",X"CA",X"FC",X"2E",X"3A",
		X"E5",X"80",X"47",X"DD",X"7E",X"08",X"90",X"47",X"E6",X"0E",X"FE",X"0C",X"C2",X"FC",X"2E",X"78",
		X"CB",X"67",X"CA",X"FC",X"2E",X"FD",X"36",X"01",X"05",X"FD",X"CB",X"00",X"CE",X"DD",X"7E",X"08",
		X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"DF",X"04",X"7E",X"FE",X"4C",X"28",
		X"04",X"FE",X"4D",X"20",X"07",X"36",X"2F",X"DD",X"35",X"03",X"28",X"09",X"FD",X"CB",X"00",X"9E",
		X"DD",X"CB",X"00",X"E6",X"C9",X"CD",X"D5",X"09",X"3A",X"2A",X"86",X"FE",X"04",X"38",X"07",X"CD",
		X"3D",X"08",X"CB",X"47",X"28",X"0C",X"FD",X"21",X"4E",X"2E",X"CD",X"43",X"09",X"CD",X"5B",X"09",
		X"18",X"FB",X"FD",X"21",X"CB",X"11",X"CD",X"43",X"09",X"CD",X"5B",X"09",X"18",X"FB",X"FD",X"36",
		X"08",X"EB",X"CD",X"3D",X"08",X"E6",X"E0",X"F6",X"13",X"FD",X"77",X"0A",X"DD",X"36",X"04",X"FE",
		X"DD",X"36",X"03",X"9C",X"C9",X"21",X"F1",X"2D",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",
		X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"3A",X"12",X"81",X"B7",X"C8",X"06",X"80",X"FE",X"01",
		X"28",X"02",X"06",X"C0",X"3A",X"01",X"98",X"2F",X"A0",X"C8",X"CD",X"87",X"14",X"21",X"00",X"00",
		X"22",X"4F",X"81",X"22",X"51",X"81",X"22",X"53",X"81",X"22",X"0A",X"81",X"08",X"AF",X"32",X"27",
		X"86",X"32",X"39",X"86",X"08",X"21",X"22",X"86",X"06",X"01",X"70",X"CB",X"77",X"CA",X"AB",X"2F",
		X"34",X"CD",X"99",X"0E",X"21",X"39",X"86",X"36",X"02",X"23",X"CD",X"4B",X"30",X"23",X"36",X"00",
		X"23",X"36",X"01",X"23",X"23",X"23",X"23",X"23",X"23",X"36",X"04",X"CD",X"99",X"0E",X"21",X"27",
		X"86",X"36",X"01",X"23",X"CD",X"4B",X"30",X"23",X"36",X"00",X"23",X"36",X"01",X"3E",X"00",X"32",
		X"92",X"86",X"21",X"9D",X"8A",X"22",X"95",X"86",X"3E",X"04",X"32",X"30",X"86",X"AF",X"32",X"A2",
		X"86",X"32",X"A3",X"86",X"32",X"A4",X"86",X"AF",X"32",X"1F",X"86",X"CD",X"81",X"0A",X"CD",X"AD",
		X"30",X"3E",X"3C",X"CD",X"AF",X"09",X"CD",X"08",X"0A",X"CD",X"FA",X"05",X"AF",X"CD",X"0C",X"08",
		X"3A",X"28",X"86",X"C6",X"99",X"27",X"32",X"28",X"86",X"B7",X"CC",X"59",X"30",X"CD",X"36",X"30",
		X"3A",X"28",X"86",X"B7",X"C2",X"D7",X"2F",X"CD",X"36",X"30",X"3A",X"28",X"86",X"B7",X"20",X"C7",
		X"2A",X"A3",X"86",X"ED",X"4B",X"A5",X"86",X"09",X"22",X"A5",X"86",X"2A",X"A7",X"86",X"23",X"3A",
		X"22",X"86",X"FE",X"02",X"20",X"01",X"23",X"22",X"A7",X"86",X"CD",X"C3",X"15",X"CD",X"36",X"30",
		X"CD",X"C3",X"15",X"C3",X"61",X"14",X"E5",X"21",X"27",X"86",X"11",X"39",X"86",X"06",X"12",X"1A",
		X"4E",X"EB",X"12",X"71",X"EB",X"23",X"13",X"10",X"F6",X"E1",X"C9",X"3A",X"01",X"98",X"2F",X"E6",
		X"01",X"28",X"03",X"36",X"05",X"C9",X"36",X"03",X"C9",X"DF",X"18",X"3A",X"22",X"86",X"FE",X"01",
		X"28",X"2E",X"CF",X"28",X"78",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"00",X"21",X"78",
		X"68",X"11",X"27",X"86",X"06",X"01",X"CD",X"28",X"05",X"CF",X"78",X"78",X"20",X"47",X"41",X"4D",
		X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"00",X"3E",X"02",X"3E",X"78",X"CD",X"AF",X"09",X"C9",
		X"CF",X"38",X"78",X"20",X"20",X"20",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",
		X"20",X"20",X"20",X"20",X"00",X"3E",X"02",X"3E",X"78",X"CD",X"AF",X"09",X"C9",X"CD",X"83",X"05",
		X"CD",X"FA",X"05",X"CD",X"A7",X"06",X"CD",X"8E",X"10",X"3E",X"00",X"32",X"9A",X"86",X"CD",X"36",
		X"31",X"21",X"E3",X"80",X"36",X"00",X"FD",X"21",X"53",X"34",X"CD",X"43",X"09",X"FD",X"21",X"46",
		X"38",X"CD",X"43",X"09",X"3E",X"50",X"CD",X"AF",X"09",X"21",X"23",X"86",X"34",X"FD",X"21",X"DB",
		X"29",X"CD",X"43",X"09",X"FD",X"21",X"E2",X"43",X"CD",X"43",X"09",X"3A",X"2A",X"86",X"FE",X"01",
		X"28",X"12",X"FD",X"21",X"4E",X"2E",X"CD",X"43",X"09",X"21",X"23",X"86",X"34",X"FD",X"21",X"DB",
		X"29",X"CD",X"43",X"09",X"FD",X"21",X"46",X"10",X"CD",X"43",X"09",X"FD",X"21",X"7F",X"09",X"CD",
		X"43",X"09",X"DD",X"21",X"18",X"82",X"DD",X"7E",X"00",X"B7",X"C8",X"3A",X"1F",X"86",X"B7",X"C4",
		X"57",X"2F",X"3A",X"1D",X"86",X"B7",X"C4",X"A7",X"06",X"3A",X"92",X"86",X"B7",X"C2",X"67",X"39",
		X"CD",X"5B",X"09",X"C3",X"12",X"31",X"3E",X"FF",X"32",X"9D",X"86",X"3A",X"2A",X"86",X"E6",X"03",
		X"FE",X"01",X"CA",X"52",X"31",X"FE",X"02",X"CA",X"7B",X"31",X"FE",X"03",X"CA",X"A4",X"31",X"C3",
		X"CD",X"31",X"DF",X"1C",X"E7",X"03",X"04",X"05",X"DF",X"3C",X"E7",X"03",X"08",X"05",X"DF",X"5C",
		X"E7",X"03",X"0C",X"05",X"DF",X"7C",X"E7",X"03",X"10",X"05",X"DF",X"9C",X"E7",X"03",X"14",X"05",
		X"DF",X"BC",X"E7",X"03",X"18",X"05",X"DF",X"DC",X"C3",X"F6",X"31",X"DF",X"1C",X"E7",X"03",X"04",
		X"04",X"DF",X"3C",X"E7",X"03",X"08",X"04",X"DF",X"5C",X"E7",X"03",X"0C",X"04",X"DF",X"7C",X"E7",
		X"03",X"10",X"04",X"DF",X"9C",X"E7",X"03",X"14",X"04",X"DF",X"BC",X"E7",X"03",X"18",X"04",X"DF",
		X"DC",X"C3",X"F6",X"31",X"DF",X"1C",X"E7",X"03",X"04",X"00",X"DF",X"3C",X"E7",X"03",X"08",X"00",
		X"DF",X"5C",X"E7",X"03",X"0C",X"00",X"DF",X"7C",X"E7",X"03",X"10",X"00",X"DF",X"9C",X"E7",X"03",
		X"14",X"00",X"DF",X"BC",X"E7",X"03",X"18",X"00",X"DF",X"DC",X"C3",X"F6",X"31",X"DF",X"1C",X"E7",
		X"03",X"04",X"06",X"DF",X"3C",X"E7",X"03",X"08",X"06",X"DF",X"5C",X"E7",X"03",X"0C",X"06",X"DF",
		X"7C",X"E7",X"03",X"10",X"06",X"DF",X"9C",X"E7",X"03",X"14",X"06",X"DF",X"BC",X"E7",X"03",X"18",
		X"06",X"DF",X"DC",X"C3",X"F6",X"31",X"21",X"85",X"42",X"3A",X"2A",X"86",X"4F",X"06",X"00",X"09",
		X"7E",X"32",X"32",X"86",X"3E",X"21",X"3D",X"F5",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"6F",X"3A",
		X"32",X"86",X"3D",X"67",X"CD",X"83",X"32",X"F1",X"20",X"EC",X"3E",X"00",X"32",X"9D",X"86",X"C9",
		X"3A",X"31",X"86",X"47",X"3A",X"E5",X"80",X"90",X"06",X"00",X"F2",X"2E",X"32",X"05",X"4F",X"2A",
		X"31",X"86",X"55",X"09",X"22",X"31",X"86",X"7D",X"AA",X"CB",X"5F",X"C8",X"78",X"B7",X"28",X"2A",
		X"FD",X"21",X"18",X"82",X"FD",X"CB",X"0B",X"CE",X"3A",X"32",X"86",X"67",X"3A",X"31",X"86",X"F6",
		X"07",X"6F",X"01",X"FF",X"00",X"37",X"3F",X"ED",X"42",X"CD",X"70",X"33",X"F5",X"21",X"4C",X"86",
		X"09",X"73",X"23",X"72",X"CD",X"95",X"33",X"C3",X"91",X"32",X"FD",X"21",X"18",X"82",X"FD",X"CB",
		X"0B",X"D6",X"3A",X"32",X"86",X"67",X"3A",X"31",X"86",X"E6",X"F8",X"6F",X"01",X"01",X"00",X"37",
		X"3F",X"ED",X"42",X"CD",X"70",X"33",X"F5",X"21",X"4C",X"86",X"09",X"73",X"23",X"72",X"CD",X"95",
		X"33",X"E5",X"EB",X"01",X"1B",X"00",X"ED",X"B0",X"E1",X"C1",X"3E",X"13",X"B8",X"CA",X"FA",X"32",
		X"3C",X"B8",X"CA",X"0F",X"33",X"3C",X"B8",X"28",X"77",X"3C",X"B8",X"CA",X"35",X"33",X"3C",X"B8",
		X"CA",X"4A",X"33",X"3C",X"B8",X"CA",X"5B",X"33",X"3E",X"00",X"B8",X"C2",X"F9",X"32",X"11",X"04",
		X"00",X"06",X"07",X"3A",X"2D",X"86",X"4F",X"23",X"3A",X"E3",X"80",X"CB",X"7F",X"20",X"10",X"3A",
		X"9D",X"86",X"B7",X"20",X"0A",X"CD",X"3D",X"08",X"1F",X"1F",X"1F",X"E6",X"01",X"18",X"14",X"CD",
		X"3D",X"08",X"FE",X"20",X"D2",X"EB",X"32",X"3E",X"03",X"18",X"08",X"B9",X"30",X"08",X"1F",X"1F",
		X"1F",X"E6",X"01",X"C6",X"4C",X"77",X"19",X"10",X"CF",X"C9",X"21",X"23",X"82",X"CB",X"76",X"C8",
		X"3E",X"46",X"21",X"90",X"88",X"77",X"2B",X"3E",X"10",X"77",X"2B",X"3E",X"5E",X"77",X"C9",X"21",
		X"23",X"82",X"CB",X"76",X"C8",X"3E",X"10",X"21",X"70",X"88",X"77",X"2B",X"77",X"2B",X"77",X"C9",
		X"21",X"23",X"82",X"CB",X"76",X"C8",X"3E",X"4A",X"21",X"50",X"88",X"77",X"2B",X"3E",X"10",X"77",
		X"2B",X"3E",X"44",X"77",X"C9",X"21",X"23",X"82",X"CB",X"7E",X"C8",X"3E",X"46",X"21",X"90",X"8B",
		X"77",X"2B",X"3E",X"10",X"77",X"2B",X"3E",X"55",X"77",X"C9",X"21",X"23",X"82",X"CB",X"7E",X"C8",
		X"3E",X"10",X"21",X"70",X"8B",X"77",X"2B",X"77",X"2B",X"77",X"C9",X"21",X"23",X"82",X"CB",X"7E",
		X"C8",X"3E",X"56",X"21",X"50",X"8B",X"77",X"2B",X"3E",X"10",X"77",X"2B",X"3E",X"53",X"77",X"C9",
		X"EB",X"06",X"00",X"4A",X"21",X"DF",X"42",X"09",X"09",X"7E",X"23",X"66",X"6F",X"7B",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"06",X"00",X"4F",X"09",X"5E",X"16",X"00",X"7B",X"21",X"61",X"3B",X"19",
		X"19",X"5E",X"23",X"56",X"C9",X"69",X"60",X"06",X"05",X"CB",X"25",X"CB",X"14",X"10",X"FA",X"01",
		X"02",X"88",X"09",X"C9",X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"04",X"BC",X"07",X"10",X"08",
		X"04",X"BB",X"07",X"00",X"01",X"A9",X"33",X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"04",X"3C",
		X"07",X"10",X"08",X"04",X"3B",X"07",X"00",X"01",X"BC",X"33",X"00",X"00",X"01",X"00",X"00",X"08",
		X"10",X"04",X"3A",X"07",X"08",X"10",X"04",X"39",X"07",X"00",X"01",X"CF",X"33",X"00",X"00",X"01",
		X"00",X"00",X"08",X"10",X"04",X"7A",X"07",X"08",X"10",X"04",X"79",X"07",X"00",X"01",X"E2",X"33",
		X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"04",X"38",X"01",X"01",X"00",X"04",X"B8",X"02",X"01",
		X"00",X"04",X"F8",X"03",X"01",X"00",X"04",X"38",X"02",X"01",X"00",X"04",X"B8",X"03",X"01",X"00",
		X"04",X"F8",X"01",X"01",X"00",X"04",X"38",X"03",X"01",X"00",X"04",X"B8",X"01",X"01",X"00",X"04",
		X"F8",X"02",X"01",X"00",X"05",X"37",X"01",X"01",X"00",X"05",X"B7",X"02",X"01",X"00",X"05",X"F7",
		X"03",X"01",X"00",X"05",X"37",X"02",X"01",X"00",X"05",X"B7",X"01",X"01",X"00",X"05",X"F7",X"03",
		X"01",X"00",X"05",X"36",X"01",X"01",X"00",X"05",X"B6",X"02",X"01",X"00",X"05",X"F6",X"03",X"00",
		X"00",X"00",X"00",X"CD",X"7B",X"08",X"DD",X"21",X"18",X"82",X"FD",X"21",X"55",X"81",X"DD",X"36",
		X"08",X"6D",X"DD",X"36",X"0A",X"73",X"CD",X"A1",X"37",X"DD",X"CB",X"00",X"D6",X"DD",X"36",X"03",
		X"FF",X"DD",X"CB",X"00",X"EE",X"CD",X"C7",X"2C",X"CD",X"92",X"2D",X"DD",X"CB",X"00",X"F6",X"DD",
		X"CB",X"0C",X"C6",X"CD",X"5B",X"09",X"3A",X"17",X"86",X"47",X"3E",X"04",X"32",X"26",X"86",X"AF",
		X"4F",X"3E",X"00",X"32",X"9B",X"86",X"3E",X"07",X"CD",X"0C",X"08",X"FD",X"21",X"55",X"81",X"DD",
		X"7E",X"0D",X"CB",X"57",X"C2",X"21",X"37",X"CD",X"C8",X"36",X"CD",X"F3",X"36",X"DD",X"CB",X"00",
		X"96",X"FD",X"CB",X"00",X"B6",X"DD",X"7E",X"0A",X"E6",X"1E",X"FE",X"12",X"C2",X"E4",X"35",X"3A",
		X"E5",X"80",X"E6",X"1E",X"FE",X"0E",X"C2",X"E4",X"35",X"DD",X"CB",X"0B",X"5E",X"CA",X"DA",X"34",
		X"01",X"01",X"01",X"CD",X"73",X"17",X"DD",X"CB",X"0B",X"9E",X"21",X"00",X"00",X"22",X"E2",X"80",
		X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",
		X"0A",X"C6",X"08",X"6F",X"CD",X"DF",X"04",X"E5",X"7E",X"CD",X"2A",X"35",X"E1",X"7E",X"FE",X"2F",
		X"28",X"1A",X"FE",X"7C",X"28",X"16",X"3A",X"0F",X"86",X"DD",X"CB",X"0B",X"6E",X"28",X"0D",X"DD",
		X"CB",X"0B",X"AE",X"E5",X"CD",X"CE",X"2D",X"E1",X"30",X"02",X"36",X"2F",X"FD",X"CB",X"00",X"6E",
		X"CA",X"E8",X"35",X"FD",X"CB",X"00",X"AE",X"C3",X"B8",X"36",X"FE",X"4C",X"20",X"17",X"CD",X"5C",
		X"36",X"FD",X"CB",X"00",X"EE",X"3A",X"0F",X"86",X"CB",X"6F",X"20",X"03",X"CB",X"67",X"C8",X"3E",
		X"13",X"CD",X"0C",X"08",X"C9",X"FE",X"D0",X"20",X"25",X"CD",X"68",X"2D",X"3E",X"88",X"BC",X"20",
		X"06",X"DD",X"CB",X"0B",X"F6",X"18",X"04",X"DD",X"CB",X"0B",X"FE",X"CD",X"C7",X"2C",X"01",X"05",
		X"01",X"CD",X"73",X"17",X"3E",X"09",X"CD",X"0C",X"08",X"21",X"94",X"86",X"34",X"C9",X"FE",X"4D",
		X"20",X"17",X"CD",X"F4",X"35",X"FD",X"CB",X"00",X"EE",X"3A",X"11",X"86",X"CB",X"67",X"20",X"03",
		X"CB",X"77",X"C8",X"3E",X"13",X"CD",X"0C",X"08",X"C9",X"FE",X"4F",X"C2",X"A0",X"35",X"36",X"10",
		X"01",X"01",X"02",X"CD",X"73",X"17",X"3E",X"04",X"CD",X"0C",X"08",X"21",X"93",X"86",X"34",X"C9",
		X"DD",X"CB",X"0B",X"76",X"20",X"06",X"DD",X"CB",X"0B",X"7E",X"28",X"1B",X"FE",X"D4",X"28",X"0C",
		X"FE",X"D5",X"28",X"08",X"FE",X"D6",X"28",X"04",X"FE",X"D7",X"20",X"0B",X"3E",X"01",X"32",X"92",
		X"86",X"3E",X"0A",X"CD",X"0C",X"08",X"C9",X"FE",X"C9",X"CA",X"E9",X"13",X"FE",X"2D",X"CA",X"FB",
		X"13",X"FE",X"7C",X"20",X"0E",X"CD",X"5C",X"36",X"3A",X"0F",X"86",X"CD",X"24",X"36",X"FD",X"CB",
		X"00",X"EE",X"C9",X"C9",X"DD",X"CB",X"0B",X"DE",X"DD",X"7E",X"0A",X"E6",X"1E",X"FE",X"12",X"CC",
		X"F4",X"35",X"18",X"5C",X"3A",X"0F",X"86",X"CB",X"6F",X"28",X"29",X"3A",X"E3",X"80",X"B8",X"20",
		X"05",X"3A",X"E2",X"80",X"B9",X"C8",X"ED",X"43",X"E2",X"80",X"FD",X"36",X"0A",X"00",X"FD",X"36",
		X"09",X"00",X"DD",X"CB",X"00",X"A6",X"21",X"A4",X"33",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",
		X"CB",X"00",X"E6",X"C9",X"CB",X"67",X"C8",X"3A",X"E3",X"80",X"BA",X"20",X"05",X"3A",X"E2",X"80",
		X"BB",X"C8",X"ED",X"53",X"E2",X"80",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"DD",X"CB",
		X"00",X"A6",X"21",X"B7",X"33",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"CB",X"00",X"E6",X"C9",
		X"3A",X"E5",X"80",X"E6",X"1E",X"FE",X"0E",X"CC",X"5C",X"36",X"18",X"5C",X"3A",X"11",X"86",X"CB",
		X"67",X"28",X"29",X"FD",X"7E",X"0A",X"BA",X"20",X"05",X"FD",X"7E",X"09",X"BB",X"C8",X"FD",X"72",
		X"0A",X"FD",X"73",X"09",X"21",X"00",X"00",X"22",X"E2",X"80",X"DD",X"CB",X"00",X"A6",X"21",X"CA",
		X"33",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"CB",X"00",X"E6",X"C9",X"CB",X"77",X"C8",X"FD",
		X"7E",X"0A",X"B8",X"20",X"05",X"FD",X"7E",X"09",X"B9",X"C8",X"FD",X"70",X"0A",X"FD",X"71",X"09",
		X"21",X"00",X"00",X"22",X"E2",X"80",X"DD",X"CB",X"00",X"A6",X"21",X"DD",X"33",X"DD",X"75",X"05",
		X"DD",X"74",X"06",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"CB",X"00",X"D6",X"CD",X"12",X"28",X"CD",
		X"FB",X"2C",X"CD",X"5B",X"09",X"C3",X"9B",X"34",X"3A",X"0F",X"86",X"CB",X"5F",X"28",X"1F",X"DD",
		X"CB",X"0B",X"66",X"C0",X"DD",X"CB",X"0B",X"E6",X"DD",X"CB",X"0B",X"EE",X"3A",X"30",X"86",X"B7",
		X"28",X"06",X"3E",X"02",X"CD",X"0C",X"08",X"C9",X"3E",X"0B",X"CD",X"0C",X"08",X"C9",X"DD",X"CB",
		X"0B",X"A6",X"C9",X"01",X"80",X"00",X"11",X"80",X"FF",X"DD",X"7E",X"0D",X"CB",X"5F",X"C0",X"01",
		X"00",X"01",X"11",X"00",X"FF",X"3E",X"08",X"32",X"8E",X"86",X"3A",X"0F",X"86",X"CB",X"4F",X"C8",
		X"3E",X"04",X"32",X"8E",X"86",X"3E",X"08",X"CD",X"0C",X"08",X"01",X"00",X"02",X"11",X"00",X"FE",
		X"C9",X"3E",X"0E",X"CD",X"0C",X"08",X"21",X"00",X"00",X"22",X"E2",X"80",X"FD",X"36",X"0A",X"00",
		X"FD",X"36",X"09",X"00",X"DD",X"21",X"18",X"82",X"DD",X"CB",X"00",X"A6",X"21",X"F0",X"33",X"DD",
		X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",
		X"66",X"28",X"2A",X"3E",X"FF",X"32",X"05",X"A8",X"3E",X"03",X"CD",X"AF",X"09",X"3E",X"00",X"32",
		X"05",X"A8",X"3E",X"04",X"CD",X"AF",X"09",X"3E",X"FF",X"32",X"03",X"A8",X"3E",X"02",X"CD",X"AF",
		X"09",X"3E",X"00",X"32",X"03",X"A8",X"3E",X"04",X"CD",X"AF",X"09",X"18",X"D0",X"3E",X"00",X"32",
		X"03",X"A8",X"32",X"05",X"A8",X"3E",X"00",X"32",X"93",X"86",X"32",X"94",X"86",X"3A",X"30",X"86",
		X"FE",X"04",X"30",X"05",X"3E",X"04",X"32",X"30",X"86",X"CD",X"D5",X"09",X"CD",X"5B",X"09",X"18",
		X"FB",X"DD",X"CB",X"0B",X"46",X"C0",X"DD",X"CB",X"0B",X"C6",X"DD",X"CB",X"00",X"A6",X"21",X"B7",
		X"33",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"3E",X"04",X"32",X"20",X"86",
		X"32",X"21",X"86",X"DD",X"CB",X"00",X"E6",X"C9",X"0D",X"2C",X"F7",X"F7",X"2E",X"F7",X"F7",X"2E",
		X"F7",X"F7",X"2E",X"F7",X"F7",X"2C",X"F7",X"F7",X"2E",X"F7",X"F7",X"2E",X"F7",X"F7",X"2E",X"F7",
		X"F7",X"10",X"20",X"11",X"1D",X"00",X"28",X"40",X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",
		X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",
		X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",
		X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",
		X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",
		X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",X"58",X"70",X"88",X"A0",X"B8",X"D0",X"28",X"40",
		X"58",X"70",X"88",X"A0",X"B8",X"D0",X"DF",X"F6",X"06",X"1C",X"DD",X"21",X"5E",X"88",X"11",X"20",
		X"00",X"21",X"C9",X"37",X"7E",X"DD",X"77",X"00",X"DD",X"19",X"23",X"10",X"F7",X"CD",X"DD",X"08",
		X"DD",X"E5",X"CD",X"B0",X"08",X"FD",X"E1",X"3E",X"EA",X"DD",X"77",X"0C",X"21",X"23",X"82",X"CB",
		X"8E",X"CB",X"96",X"21",X"E5",X"37",X"3A",X"2A",X"86",X"4F",X"06",X"00",X"09",X"7E",X"32",X"97",
		X"86",X"3E",X"01",X"32",X"98",X"86",X"3E",X"02",X"FD",X"77",X"03",X"FD",X"CB",X"00",X"EE",X"DD",
		X"E5",X"FD",X"E5",X"DD",X"E1",X"FD",X"E1",X"21",X"23",X"82",X"CB",X"4E",X"28",X"18",X"CB",X"8E",
		X"21",X"98",X"86",X"34",X"3A",X"98",X"86",X"FE",X"0C",X"20",X"24",X"3E",X"01",X"32",X"98",X"86",
		X"21",X"97",X"86",X"34",X"18",X"19",X"CB",X"56",X"28",X"15",X"CB",X"96",X"21",X"98",X"86",X"35",
		X"3A",X"98",X"86",X"B7",X"20",X"09",X"3E",X"0B",X"32",X"98",X"86",X"21",X"97",X"86",X"35",X"DD",
		X"7E",X"03",X"B7",X"20",X"18",X"3E",X"02",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"FD",X"34",
		X"0C",X"FD",X"7E",X"0C",X"FE",X"EC",X"20",X"05",X"3E",X"E9",X"FD",X"77",X"0C",X"3A",X"97",X"86",
		X"FE",X"29",X"30",X"02",X"3E",X"29",X"FD",X"77",X"06",X"FD",X"E5",X"DD",X"E5",X"CD",X"5B",X"09",
		X"C3",X"93",X"38",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"10",X"11",X"12",
		X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",
		X"29",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"40",X"41",X"42",X"43",X"44",
		X"45",X"46",X"47",X"48",X"49",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"60",
		X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"70",X"71",X"72",X"73",X"74",X"75",X"76",
		X"77",X"78",X"79",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"90",X"91",X"92",
		X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"CD",X"08",X"0A",X"3E",X"00",X"32",X"03",X"A8",X"32",
		X"05",X"A8",X"21",X"00",X"00",X"22",X"E2",X"80",X"06",X"03",X"C5",X"D7",X"01",X"3E",X"04",X"CD",
		X"AF",X"09",X"D7",X"02",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"03",X"3E",X"04",X"CD",X"AF",X"09",
		X"D7",X"04",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"05",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"06",
		X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"07",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"08",X"3E",X"04",
		X"CD",X"AF",X"09",X"C1",X"10",X"C4",X"CD",X"FA",X"05",X"CD",X"83",X"05",X"D7",X"00",X"CD",X"A7",
		X"06",X"CD",X"F1",X"06",X"3A",X"2A",X"86",X"4F",X"06",X"00",X"21",X"03",X"39",X"09",X"7E",X"32",
		X"99",X"86",X"DF",X"25",X"CF",X"38",X"20",X"4D",X"41",X"44",X"45",X"20",X"49",X"54",X"20",X"54",
		X"4F",X"20",X"42",X"41",X"4E",X"4B",X"20",X"20",X"20",X"00",X"21",X"20",X"B8",X"11",X"99",X"86",
		X"06",X"02",X"CD",X"28",X"05",X"3E",X"0A",X"CD",X"AF",X"09",X"E7",X"03",X"06",X"03",X"CF",X"28",
		X"30",X"4D",X"4F",X"4E",X"45",X"59",X"20",X"43",X"4F",X"4C",X"4C",X"45",X"43",X"54",X"45",X"44",
		X"20",X"42",X"4F",X"4E",X"55",X"53",X"00",X"CF",X"58",X"40",X"31",X"30",X"30",X"20",X"50",X"4F",
		X"49",X"4E",X"54",X"53",X"00",X"3E",X"14",X"CD",X"AF",X"09",X"3A",X"93",X"86",X"B7",X"28",X"32",
		X"FE",X"4E",X"38",X"02",X"3E",X"4E",X"21",X"50",X"18",X"F5",X"E5",X"CD",X"DA",X"04",X"36",X"4F",
		X"01",X"01",X"02",X"CD",X"73",X"17",X"CD",X"A7",X"06",X"3E",X"0C",X"CD",X"0C",X"08",X"E1",X"CD",
		X"53",X"3B",X"E5",X"3E",X"05",X"CD",X"AF",X"09",X"E1",X"F1",X"3D",X"20",X"DC",X"3E",X"0A",X"CD",
		X"AF",X"09",X"E7",X"03",X"12",X"01",X"CF",X"40",X"90",X"42",X"4F",X"4E",X"55",X"53",X"20",X"53",
		X"41",X"57",X"48",X"4F",X"52",X"53",X"45",X"53",X"00",X"CF",X"20",X"A0",X"31",X"20",X"53",X"41",
		X"57",X"48",X"4F",X"52",X"53",X"45",X"20",X"50",X"45",X"52",X"20",X"34",X"20",X"4D",X"4F",X"4E",
		X"45",X"59",X"53",X"00",X"3E",X"14",X"CD",X"AF",X"09",X"3A",X"93",X"86",X"CB",X"3F",X"CB",X"3F",
		X"28",X"2D",X"FE",X"48",X"38",X"02",X"3E",X"48",X"21",X"B0",X"18",X"F5",X"E5",X"CD",X"DA",X"04",
		X"36",X"2F",X"21",X"30",X"86",X"34",X"3E",X"0D",X"CD",X"0C",X"08",X"E1",X"CD",X"53",X"3B",X"E5",
		X"3E",X"0A",X"CD",X"AF",X"09",X"E1",X"F1",X"3D",X"20",X"E1",X"3E",X"14",X"CD",X"AF",X"09",X"AF",
		X"32",X"93",X"86",X"32",X"94",X"86",X"3E",X"FF",X"3E",X"00",X"32",X"92",X"86",X"21",X"2A",X"86",
		X"34",X"06",X"05",X"C5",X"D7",X"01",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"02",X"3E",X"04",X"CD",
		X"AF",X"09",X"D7",X"03",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"04",X"3E",X"04",X"CD",X"AF",X"09",
		X"D7",X"05",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"06",X"3E",X"04",X"CD",X"AF",X"09",X"D7",X"00",
		X"3E",X"04",X"CD",X"AF",X"09",X"C1",X"10",X"CB",X"3A",X"2A",X"86",X"3D",X"FE",X"04",X"28",X"04",
		X"FE",X"08",X"20",X"18",X"FD",X"21",X"55",X"45",X"CD",X"43",X"09",X"3E",X"FE",X"CD",X"AF",X"09",
		X"21",X"28",X"86",X"34",X"CD",X"F1",X"06",X"3E",X"FA",X"CD",X"AF",X"09",X"CD",X"08",X"0A",X"CD",
		X"83",X"05",X"C3",X"AD",X"30",X"7C",X"C6",X"08",X"67",X"FE",X"E0",X"C0",X"26",X"18",X"7D",X"C6",
		X"08",X"6F",X"C9",X"7C",X"C6",X"10",X"67",X"FE",X"E0",X"D8",X"26",X"18",X"7D",X"C6",X"08",X"6F",
		X"C9",X"C9",X"3B",X"E4",X"3B",X"FF",X"3B",X"1A",X"3C",X"35",X"3C",X"50",X"3C",X"6B",X"3C",X"86",
		X"3C",X"A1",X"3C",X"BC",X"3C",X"D7",X"3C",X"F2",X"3C",X"0D",X"3D",X"28",X"3D",X"43",X"3D",X"5E",
		X"3D",X"79",X"3D",X"94",X"3D",X"AF",X"3D",X"CA",X"3D",X"E5",X"3D",X"00",X"3E",X"1B",X"3E",X"36",
		X"3E",X"51",X"3E",X"6C",X"3E",X"87",X"3E",X"A2",X"3E",X"BD",X"3E",X"D8",X"3E",X"F3",X"3E",X"0E",
		X"3F",X"29",X"3F",X"44",X"3F",X"5F",X"3F",X"7A",X"3F",X"95",X"3F",X"B0",X"3F",X"CB",X"3F",X"E6",
		X"3F",X"01",X"40",X"1C",X"40",X"37",X"40",X"52",X"40",X"6D",X"40",X"88",X"40",X"A3",X"40",X"BE",
		X"40",X"D9",X"40",X"F4",X"40",X"0F",X"41",X"2A",X"41",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",X"10",X"56",X"59",
		X"5C",X"10",X"4A",X"43",X"44",X"10",X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",X"10",X"5F",X"5F",
		X"10",X"4A",X"43",X"5C",X"10",X"42",X"43",X"44",X"10",X"42",X"43",X"44",X"10",X"56",X"4B",X"53",
		X"10",X"42",X"4B",X"44",X"10",X"56",X"59",X"53",X"10",X"5F",X"5F",X"10",X"56",X"4B",X"5C",X"10",
		X"4A",X"59",X"5C",X"10",X"42",X"4B",X"44",X"10",X"42",X"59",X"5C",X"10",X"42",X"43",X"53",X"10",
		X"4A",X"4B",X"44",X"10",X"5F",X"5F",X"10",X"40",X"49",X"45",X"10",X"50",X"41",X"45",X"10",X"40",
		X"5A",X"45",X"10",X"40",X"49",X"54",X"10",X"50",X"5A",X"5D",X"10",X"57",X"5A",X"45",X"10",X"5F",
		X"5F",X"10",X"50",X"49",X"54",X"10",X"57",X"49",X"54",X"10",X"50",X"41",X"5D",X"10",X"57",X"41",
		X"5D",X"10",X"40",X"41",X"45",X"10",X"40",X"41",X"5D",X"10",X"5F",X"5F",X"10",X"57",X"5A",X"5D",
		X"10",X"40",X"5A",X"5D",X"10",X"57",X"49",X"54",X"10",X"50",X"49",X"45",X"10",X"57",X"49",X"54",
		X"10",X"50",X"49",X"54",X"10",X"5F",X"5F",X"10",X"58",X"52",X"5E",X"10",X"46",X"5B",X"55",X"10",
		X"58",X"52",X"5E",X"10",X"51",X"5B",X"48",X"10",X"51",X"47",X"5E",X"10",X"58",X"47",X"55",X"10",
		X"5F",X"5F",X"10",X"46",X"5B",X"48",X"10",X"51",X"47",X"48",X"10",X"51",X"47",X"48",X"10",X"46",
		X"47",X"5E",X"10",X"58",X"52",X"55",X"10",X"46",X"5B",X"5E",X"10",X"5F",X"5F",X"10",X"51",X"47",
		X"55",X"10",X"58",X"52",X"5E",X"10",X"46",X"5B",X"55",X"10",X"58",X"52",X"55",X"10",X"46",X"5B",
		X"5E",X"10",X"51",X"52",X"48",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"D4",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",X"10",X"60",X"63",X"63",X"63",
		X"63",X"63",X"67",X"10",X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",X"10",X"5F",X"5F",X"10",X"40",
		X"49",X"45",X"10",X"50",X"41",X"45",X"10",X"61",X"64",X"64",X"69",X"66",X"66",X"68",X"10",X"50",
		X"5A",X"5D",X"10",X"57",X"5A",X"45",X"10",X"5F",X"5F",X"10",X"51",X"47",X"55",X"10",X"58",X"52",
		X"5E",X"10",X"61",X"64",X"64",X"6A",X"66",X"66",X"68",X"10",X"46",X"5B",X"5E",X"10",X"51",X"52",
		X"48",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"D7",X"61",X"64",X"64",
		X"6B",X"66",X"66",X"68",X"D6",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",
		X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",X"10",X"61",X"64",X"64",X"6C",X"66",X"66",X"68",X"10",
		X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",X"10",X"5F",X"5F",X"10",X"57",X"5A",X"5D",X"10",X"40",
		X"5A",X"5D",X"10",X"61",X"64",X"64",X"6D",X"66",X"66",X"68",X"10",X"57",X"49",X"54",X"10",X"50",
		X"49",X"54",X"10",X"5F",X"5F",X"10",X"58",X"52",X"5E",X"10",X"46",X"5B",X"55",X"10",X"62",X"65",
		X"65",X"65",X"65",X"65",X"6E",X"10",X"51",X"47",X"5E",X"10",X"58",X"47",X"55",X"10",X"5F",X"5F",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"D5",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",X"51",X"47",X"5E",X"10",
		X"46",X"5B",X"55",X"10",X"51",X"52",X"CB",X"D2",X"D3",X"52",X"5E",X"10",X"46",X"5B",X"55",X"10",
		X"51",X"52",X"55",X"10",X"5F",X"5F",X"4C",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"CC",X"D0",X"D1",X"10",X"10",X"4C",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",
		X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"44",X"10",X"4A",X"43",X"CD",X"CE",X"CF",X"43",
		X"44",X"10",X"42",X"59",X"5C",X"10",X"42",X"4B",X"5C",X"10",X"5F",X"5F",X"10",X"51",X"52",X"55",
		X"10",X"46",X"52",X"5E",X"10",X"51",X"52",X"CB",X"D2",X"D3",X"52",X"48",X"10",X"46",X"5B",X"55",
		X"10",X"51",X"47",X"48",X"10",X"5F",X"5F",X"4C",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"CC",X"D0",X"D1",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"5F",X"5F",X"10",X"42",X"59",X"53",X"10",X"56",X"43",X"5C",X"10",X"4A",X"43",X"CD",X"CE",X"CF",
		X"43",X"44",X"10",X"42",X"4B",X"5C",X"10",X"42",X"4B",X"44",X"10",X"5F",X"5F",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"D4",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",
		X"10",X"60",X"63",X"63",X"63",X"63",X"63",X"67",X"10",X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",
		X"10",X"5F",X"5F",X"10",X"40",X"49",X"45",X"10",X"50",X"41",X"45",X"10",X"61",X"64",X"6F",X"74",
		X"66",X"66",X"68",X"10",X"50",X"5A",X"5D",X"10",X"57",X"5A",X"45",X"10",X"5F",X"5F",X"10",X"51",
		X"47",X"55",X"10",X"58",X"52",X"5E",X"10",X"61",X"64",X"70",X"75",X"66",X"66",X"68",X"10",X"46",
		X"5B",X"5E",X"10",X"51",X"52",X"48",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"D7",X"61",X"64",X"71",X"76",X"66",X"66",X"68",X"D6",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",X"10",X"61",X"64",X"72",
		X"77",X"66",X"66",X"68",X"10",X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",X"10",X"5F",X"5F",X"10",
		X"57",X"5A",X"5D",X"10",X"40",X"5A",X"5D",X"10",X"61",X"64",X"73",X"78",X"66",X"66",X"68",X"10",
		X"57",X"49",X"54",X"10",X"50",X"49",X"54",X"10",X"5F",X"5F",X"10",X"58",X"52",X"5E",X"10",X"46",
		X"5B",X"55",X"10",X"62",X"65",X"65",X"65",X"65",X"65",X"6E",X"10",X"51",X"47",X"5E",X"10",X"58",
		X"47",X"55",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"D5",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"D4",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",
		X"4A",X"4B",X"53",X"10",X"60",X"63",X"16",X"22",X"63",X"63",X"67",X"10",X"4A",X"59",X"5C",X"10",
		X"42",X"43",X"5C",X"10",X"5F",X"5F",X"10",X"40",X"49",X"45",X"10",X"50",X"41",X"45",X"10",X"61",
		X"64",X"15",X"15",X"66",X"66",X"68",X"10",X"50",X"5A",X"5D",X"10",X"57",X"5A",X"45",X"10",X"5F",
		X"5F",X"10",X"51",X"47",X"55",X"10",X"58",X"52",X"5E",X"10",X"61",X"64",X"14",X"23",X"66",X"66",
		X"68",X"10",X"46",X"5B",X"5E",X"10",X"51",X"52",X"48",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"D7",X"61",X"64",X"15",X"15",X"66",X"66",X"68",X"D6",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",X"10",
		X"61",X"64",X"22",X"22",X"66",X"66",X"68",X"10",X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",X"10",
		X"5F",X"5F",X"10",X"57",X"5A",X"5D",X"10",X"40",X"5A",X"5D",X"10",X"61",X"64",X"11",X"26",X"66",
		X"66",X"68",X"10",X"57",X"49",X"54",X"10",X"50",X"49",X"54",X"10",X"5F",X"5F",X"10",X"58",X"52",
		X"5E",X"10",X"46",X"5B",X"55",X"10",X"62",X"65",X"1C",X"15",X"65",X"65",X"6E",X"10",X"51",X"47",
		X"5E",X"10",X"58",X"47",X"55",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"D5",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"5F",X"5F",X"10",X"42",X"59",X"44",X"10",X"4A",X"4B",X"53",X"10",X"8E",X"8F",X"87",X"10",
		X"8E",X"8F",X"87",X"10",X"4A",X"59",X"5C",X"10",X"42",X"43",X"5C",X"10",X"5F",X"5F",X"10",X"40",
		X"49",X"45",X"10",X"50",X"41",X"45",X"10",X"8C",X"8D",X"88",X"10",X"8C",X"8D",X"88",X"10",X"50",
		X"5A",X"5D",X"10",X"57",X"5A",X"45",X"10",X"5F",X"5F",X"10",X"58",X"52",X"5E",X"10",X"46",X"5B",
		X"55",X"10",X"8A",X"8B",X"89",X"10",X"8A",X"8B",X"89",X"10",X"51",X"47",X"5E",X"10",X"58",X"47",
		X"55",X"10",X"5F",X"5F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"CA",X"C9",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",
		X"10",X"10",X"4E",X"2D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"5F",X"10",X"8E",X"8F",X"87",X"10",X"8E",
		X"8F",X"87",X"10",X"8E",X"8F",X"87",X"10",X"8E",X"8F",X"87",X"10",X"8E",X"8F",X"87",X"10",X"8E",
		X"8F",X"87",X"10",X"5F",X"5F",X"10",X"8C",X"8D",X"88",X"10",X"8C",X"8D",X"88",X"10",X"8C",X"8D",
		X"88",X"10",X"8C",X"8D",X"88",X"10",X"8C",X"8D",X"88",X"10",X"8C",X"8D",X"88",X"10",X"5F",X"5F",
		X"10",X"8A",X"8B",X"89",X"10",X"8A",X"8B",X"89",X"10",X"8A",X"8B",X"89",X"10",X"8A",X"8B",X"89",
		X"10",X"8A",X"8B",X"89",X"10",X"8A",X"8B",X"89",X"10",X"5F",X"5F",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"5F",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"2D",X"2C",X"2B",
		X"00",X"07",X"05",X"01",X"00",X"09",X"06",X"03",X"00",X"08",X"05",X"02",X"00",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"00",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"09",X"05",X"02",
		X"00",X"07",X"05",X"01",X"12",X"11",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"00",X"08",X"04",X"15",X"14",X"13",X"06",X"03",X"00",X"09",X"05",X"02",
		X"00",X"07",X"05",X"03",X"00",X"09",X"06",X"03",X"00",X"08",X"05",X"02",X"00",X"07",X"04",X"01",
		X"00",X"07",X"04",X"03",X"00",X"08",X"04",X"01",X"00",X"09",X"06",X"03",X"00",X"09",X"05",X"02",
		X"00",X"07",X"05",X"03",X"00",X"09",X"06",X"03",X"00",X"08",X"05",X"02",X"00",X"07",X"04",X"18",
		X"17",X"16",X"04",X"03",X"00",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"09",X"05",X"02",
		X"00",X"07",X"05",X"01",X"21",X"20",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"00",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"09",X"05",X"02",
		X"00",X"07",X"05",X"01",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",X"23",X"22",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"00",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"2D",X"2C",X"2B",
		X"00",X"07",X"05",X"01",X"00",X"09",X"06",X"03",X"00",X"08",X"05",X"02",X"2E",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"00",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"2D",X"2C",X"2B",
		X"00",X"07",X"05",X"01",X"00",X"09",X"06",X"03",X"00",X"08",X"05",X"02",X"2F",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"00",X"32",X"31",X"30",X"00",X"32",X"31",X"30",X"00",X"32",X"31",X"30",
		X"00",X"32",X"31",X"30",X"00",X"32",X"31",X"30",X"00",X"32",X"31",X"30",X"00",X"32",X"31",X"30",
		X"00",X"32",X"31",X"30",X"00",X"08",X"04",X"01",X"00",X"07",X"06",X"03",X"00",X"2D",X"2C",X"2B",
		X"00",X"07",X"05",X"01",X"00",X"09",X"06",X"03",X"00",X"08",X"05",X"02",X"00",X"07",X"04",X"03",
		X"00",X"09",X"04",X"03",X"33",X"00",X"48",X"41",X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",
		X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",
		X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",
		X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",
		X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",
		X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"41",X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"45",
		X"41",X"45",X"41",X"45",X"41",X"45",X"41",X"45",X"41",X"45",X"41",X"45",X"41",X"45",X"41",X"65",
		X"41",X"45",X"41",X"A5",X"41",X"25",X"42",X"45",X"41",X"85",X"41",X"05",X"42",X"E5",X"41",X"45",
		X"41",X"A5",X"41",X"25",X"42",X"45",X"41",X"85",X"41",X"05",X"42",X"65",X"41",X"45",X"41",X"A5",
		X"41",X"25",X"42",X"45",X"41",X"85",X"41",X"05",X"42",X"65",X"41",X"45",X"41",X"A5",X"41",X"25",
		X"42",X"45",X"41",X"85",X"41",X"05",X"42",X"65",X"41",X"45",X"41",X"A5",X"41",X"25",X"42",X"45",
		X"41",X"85",X"41",X"05",X"42",X"C5",X"41",X"45",X"41",X"A5",X"41",X"25",X"42",X"45",X"41",X"85",
		X"41",X"05",X"42",X"65",X"41",X"45",X"41",X"A5",X"41",X"25",X"42",X"45",X"41",X"85",X"41",X"05",
		X"42",X"65",X"41",X"45",X"41",X"A5",X"41",X"25",X"42",X"45",X"41",X"85",X"41",X"05",X"42",X"65",
		X"41",X"45",X"41",X"A5",X"41",X"25",X"42",X"45",X"41",X"85",X"41",X"05",X"42",X"65",X"42",X"45",
		X"42",X"45",X"42",X"45",X"42",X"45",X"42",X"45",X"42",X"45",X"42",X"45",X"42",X"45",X"42",X"45",
		X"42",X"45",X"42",X"45",X"42",X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"03",X"B0",X"07",X"10",
		X"08",X"03",X"B1",X"07",X"10",X"08",X"03",X"AC",X"07",X"10",X"08",X"03",X"AD",X"07",X"00",X"01",
		X"8A",X"43",X"00",X"00",X"01",X"00",X"00",X"10",X"10",X"04",X"38",X"03",X"10",X"10",X"04",X"78",
		X"03",X"10",X"10",X"04",X"39",X"03",X"10",X"10",X"04",X"79",X"03",X"10",X"10",X"04",X"3A",X"03",
		X"10",X"10",X"04",X"7A",X"03",X"10",X"10",X"04",X"3B",X"00",X"10",X"10",X"04",X"7B",X"00",X"10",
		X"10",X"04",X"3A",X"00",X"10",X"10",X"04",X"39",X"00",X"10",X"10",X"04",X"38",X"00",X"00",X"00",
		X"00",X"00",X"CD",X"C5",X"08",X"D2",X"7F",X"09",X"DD",X"E5",X"CD",X"9F",X"08",X"D2",X"B7",X"44",
		X"FD",X"E1",X"CD",X"E0",X"44",X"CD",X"F7",X"44",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",
		X"FD",X"CB",X"00",X"D6",X"DD",X"E5",X"CD",X"5B",X"09",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",
		X"B7",X"44",X"DD",X"7E",X"0D",X"B7",X"FD",X"CB",X"00",X"76",X"C2",X"B7",X"44",X"FD",X"CB",X"00",
		X"4E",X"CC",X"2B",X"44",X"FD",X"E5",X"CD",X"5B",X"09",X"18",X"DE",X"FD",X"CB",X"00",X"DE",X"DD",
		X"7E",X"0A",X"E6",X"0E",X"FE",X"02",X"C2",X"7D",X"44",X"DD",X"7E",X"0A",X"CB",X"67",X"CA",X"7D",
		X"44",X"3A",X"E5",X"80",X"47",X"DD",X"7E",X"08",X"90",X"47",X"E6",X"0E",X"FE",X"0C",X"C2",X"7D",
		X"44",X"78",X"CB",X"67",X"CA",X"7D",X"44",X"FD",X"36",X"01",X"07",X"FD",X"CB",X"00",X"CE",X"DD",
		X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"DF",X"04",X"7E",X"FE",
		X"2F",X"28",X"08",X"FE",X"4C",X"28",X"04",X"FE",X"4D",X"20",X"02",X"36",X"10",X"FD",X"CB",X"00",
		X"9E",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"19",X"AF",X"06",X"04",
		X"77",X"23",X"10",X"FC",X"23",X"06",X"04",X"77",X"23",X"10",X"FC",X"DD",X"CB",X"0C",X"96",X"DD",
		X"CB",X"00",X"A6",X"21",X"A2",X"43",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",
		X"DD",X"CB",X"00",X"E6",X"CD",X"AF",X"09",X"CD",X"D5",X"09",X"3A",X"2A",X"86",X"FE",X"03",X"38",
		X"07",X"CD",X"3D",X"08",X"CB",X"47",X"28",X"0C",X"FD",X"21",X"E2",X"43",X"CD",X"43",X"09",X"CD",
		X"5B",X"09",X"18",X"FB",X"FD",X"21",X"14",X"46",X"CD",X"43",X"09",X"CD",X"5B",X"09",X"18",X"FB",
		X"FD",X"36",X"08",X"EB",X"CD",X"3D",X"08",X"E6",X"E0",X"F6",X"13",X"FD",X"77",X"0A",X"DD",X"36",
		X"04",X"FF",X"DD",X"36",X"03",X"6A",X"C9",X"21",X"85",X"43",X"FD",X"75",X"05",X"FD",X"74",X"06",
		X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",X"00",X"01",X"00",X"00",X"10",X"08",
		X"04",X"BC",X"05",X"10",X"08",X"04",X"BB",X"05",X"00",X"01",X"0E",X"45",X"00",X"00",X"01",X"00",
		X"00",X"10",X"08",X"04",X"3C",X"05",X"10",X"08",X"04",X"3B",X"05",X"00",X"01",X"21",X"45",X"00",
		X"00",X"01",X"00",X"00",X"08",X"10",X"04",X"3A",X"05",X"08",X"10",X"04",X"39",X"05",X"00",X"01",
		X"34",X"45",X"00",X"00",X"01",X"00",X"00",X"08",X"10",X"04",X"7A",X"05",X"08",X"10",X"04",X"79",
		X"05",X"00",X"01",X"47",X"45",X"CD",X"C5",X"08",X"D2",X"7F",X"09",X"DD",X"E5",X"CD",X"9F",X"08",
		X"D2",X"B6",X"45",X"FD",X"E1",X"CD",X"DE",X"45",X"CD",X"EF",X"45",X"FD",X"CB",X"00",X"F6",X"FD",
		X"CB",X"0C",X"D6",X"FD",X"CB",X"00",X"D6",X"3E",X"12",X"CD",X"0C",X"08",X"DD",X"E5",X"CD",X"5B",
		X"09",X"FD",X"E1",X"DD",X"7E",X"0A",X"FE",X"D3",X"20",X"1D",X"FD",X"36",X"0A",X"00",X"FD",X"36",
		X"09",X"00",X"FD",X"36",X"04",X"FE",X"21",X"09",X"45",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",
		X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"DD",X"7E",X"08",X"FE",X"78",X"CA",X"B6",X"45",X"FD",
		X"E5",X"CD",X"5B",X"09",X"18",X"CB",X"FD",X"36",X"04",X"00",X"21",X"42",X"45",X"DD",X"75",X"05",
		X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"32",X"CD",X"AF",X"09",
		X"CD",X"D5",X"09",X"3E",X"0E",X"CD",X"0C",X"08",X"CD",X"5B",X"09",X"C3",X"DB",X"45",X"FD",X"36",
		X"08",X"D2",X"FD",X"36",X"0A",X"32",X"DD",X"36",X"0A",X"01",X"DD",X"36",X"09",X"64",X"C9",X"21",
		X"42",X"45",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",
		X"C9",X"00",X"00",X"01",X"00",X"00",X"10",X"08",X"06",X"AE",X"02",X"10",X"08",X"06",X"AF",X"02",
		X"00",X"01",X"06",X"46",X"CD",X"C5",X"08",X"D2",X"7F",X"09",X"DD",X"E5",X"CD",X"9F",X"08",X"D2",
		X"57",X"46",X"FD",X"E1",X"3E",X"10",X"CD",X"0C",X"08",X"CD",X"7E",X"46",X"CD",X"95",X"46",X"FD",
		X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"FD",X"CB",X"00",X"D6",X"DD",X"E5",X"CD",X"5B",X"09",
		X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"57",X"46",X"FD",X"CB",X"00",X"76",X"C2",X"57",X"46",
		X"FD",X"E5",X"CD",X"5B",X"09",X"18",X"E9",X"3E",X"07",X"CD",X"0C",X"08",X"CD",X"D5",X"09",X"CD",
		X"3D",X"08",X"CB",X"47",X"28",X"0C",X"FD",X"21",X"E2",X"43",X"CD",X"43",X"09",X"CD",X"5B",X"09",
		X"18",X"FB",X"FD",X"21",X"14",X"46",X"CD",X"43",X"09",X"CD",X"5B",X"09",X"18",X"FB",X"FD",X"36",
		X"08",X"09",X"CD",X"3D",X"08",X"E6",X"E0",X"F6",X"13",X"FD",X"77",X"0A",X"DD",X"36",X"04",X"02",
		X"DD",X"36",X"03",X"00",X"C9",X"21",X"01",X"46",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",
		X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"AD",X"21",X"6B",X"47",X"7E",X"32",X"0F",X"86",X"23",
		X"7E",X"32",X"11",X"86",X"23",X"7E",X"32",X"A0",X"86",X"23",X"22",X"9E",X"86",X"3E",X"FF",X"32",
		X"1F",X"86",X"C9",X"21",X"A0",X"86",X"35",X"20",X"19",X"2A",X"9E",X"86",X"7E",X"FE",X"FF",X"28",
		X"D7",X"32",X"0F",X"86",X"23",X"7E",X"32",X"11",X"86",X"23",X"7E",X"32",X"A0",X"86",X"23",X"22",
		X"9E",X"86",X"C9",X"3A",X"0F",X"86",X"E6",X"1A",X"FE",X"1A",X"C0",X"21",X"80",X"88",X"11",X"20",
		X"00",X"3A",X"A5",X"86",X"E6",X"0F",X"CD",X"50",X"47",X"3A",X"A5",X"86",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CD",X"50",X"47",X"3A",X"A6",X"86",X"E6",X"0F",X"CD",X"50",X"47",X"3A",
		X"A6",X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"50",X"47",X"21",X"00",X"8B",
		X"11",X"20",X"00",X"3A",X"A7",X"86",X"E6",X"0F",X"CD",X"50",X"47",X"3A",X"A7",X"86",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"50",X"47",X"3A",X"A8",X"86",X"E6",X"0F",X"CD",X"50",
		X"47",X"3A",X"A8",X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"50",X"47",X"C9",
		X"01",X"59",X"47",X"81",X"4F",X"0A",X"77",X"19",X"C9",X"00",X"01",X"02",X"03",X"04",X"05",X"06",
		X"07",X"08",X"09",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"00",X"00",X"20",X"10",X"00",
		X"40",X"00",X"40",X"20",X"10",X"00",X"30",X"00",X"10",X"90",X"12",X"00",X"20",X"08",X"40",X"10",
		X"00",X"40",X"50",X"10",X"00",X"20",X"12",X"00",X"10",X"00",X"40",X"20",X"10",X"00",X"30",X"00",
		X"10",X"70",X"12",X"00",X"20",X"08",X"40",X"20",X"00",X"40",X"40",X"10",X"00",X"20",X"12",X"00",
		X"10",X"00",X"40",X"20",X"10",X"00",X"30",X"00",X"10",X"80",X"12",X"00",X"20",X"08",X"40",X"10",
		X"00",X"40",X"50",X"10",X"00",X"20",X"12",X"00",X"10",X"00",X"40",X"20",X"10",X"00",X"30",X"00",
		X"10",X"80",X"12",X"00",X"20",X"08",X"40",X"20",X"00",X"40",X"40",X"10",X"00",X"20",X"12",X"00",
		X"10",X"00",X"40",X"20",X"10",X"00",X"30",X"00",X"10",X"70",X"12",X"00",X"20",X"08",X"40",X"10",
		X"00",X"40",X"50",X"10",X"00",X"20",X"12",X"00",X"10",X"00",X"40",X"20",X"10",X"00",X"30",X"00",
		X"10",X"50",X"12",X"00",X"20",X"08",X"40",X"20",X"00",X"40",X"40",X"10",X"00",X"20",X"FF",X"FF",
		X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
