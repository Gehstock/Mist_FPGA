library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity timber_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of timber_bg_bits_2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"80",X"71",X"40",X"30",X"00",X"10",X"04",X"05",X"50",X"04",X"10",X"28",X"28",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"A9",
		X"80",X"AA",X"0A",X"AA",X"00",X"00",X"AA",X"AA",X"59",X"55",X"59",X"55",X"AA",X"AA",X"55",X"95",
		X"A8",X"AA",X"A2",X"AA",X"0A",X"AA",X"AA",X"AA",X"88",X"AA",X"8A",X"AA",X"AA",X"AA",X"5A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"A8",X"01",X"A0",X"02",X"A0",X"31",X"80",X"01",X"80",X"02",X"03",X"01",X"00",X"01",X"AA",X"AA",
		X"55",X"95",X"AA",X"AA",X"59",X"55",X"59",X"55",X"AA",X"AA",X"55",X"95",X"55",X"95",X"AA",X"AA",
		X"5A",X"80",X"AA",X"80",X"9A",X"00",X"9A",X"00",X"A8",X"00",X"58",X"00",X"50",X"00",X"AA",X"AA",
		X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"03",X"AA",X"00",X"A8",X"AA",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"A0",X"30",X"A0",X"00",X"80",X"00",X"80",X"00",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"51",X"14",X"11",X"10",X"05",X"40",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"15",X"05",X"50",X"00",X"40",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"AA",X"A2",
		X"80",X"00",X"15",X"55",X"03",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"45",X"55",X"03",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"55",X"55",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"55",X"55",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"55",X"55",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"C0",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"03",X"AA",X"00",X"A8",X"00",X"A8",X"AA",
		X"A0",X"00",X"A0",X"30",X"A0",X"00",X"80",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",X"00",X"00",
		X"0A",X"A0",X"28",X"A8",X"00",X"28",X"00",X"A0",X"02",X"80",X"0A",X"00",X"2A",X"A8",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"00",X"28",X"02",X"A0",X"00",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"02",X"28",X"0A",X"28",X"08",X"28",X"28",X"28",X"2A",X"A8",X"00",X"28",X"00",X"28",X"00",X"00",
		X"2A",X"A8",X"28",X"00",X"2A",X"A0",X"00",X"28",X"00",X"28",X"2A",X"A8",X"2A",X"A0",X"00",X"00",
		X"02",X"A0",X"0A",X"08",X"28",X"00",X"2A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"2A",X"A8",X"20",X"28",X"00",X"A0",X"02",X"80",X"0A",X"80",X"0A",X"00",X"0A",X"00",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A8",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"00",
		X"2A",X"A0",X"80",X"08",X"8A",X"88",X"88",X"08",X"8A",X"88",X"80",X"08",X"2A",X"A0",X"00",X"00",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"00",X"00",X"00",X"00",X"02",X"2A",X"8A",X"20",X"22",X"2A",X"02",X"20",X"02",X"2A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"82",X"02",X"08",X"02",X"08",X"02",X"08",X"02",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"82",X"82",X"22",X"82",X"82",X"82",X"22",X"02",X"82",X"00",X"00",
		X"00",X"00",X"00",X"00",X"82",X"2A",X"08",X"88",X"8A",X"88",X"08",X"88",X"88",X"88",X"00",X"00",
		X"02",X"80",X"71",X"40",X"30",X"00",X"10",X"04",X"01",X"40",X"04",X"10",X"28",X"28",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A0",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"08",X"0A",X"A0",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"08",X"28",X"08",X"28",X"08",X"28",X"28",X"2A",X"A0",X"00",X"00",
		X"2A",X"A8",X"28",X"00",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",X"2A",X"A8",X"00",X"00",
		X"2A",X"A8",X"28",X"00",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",X"28",X"00",X"00",X"00",
		X"0A",X"A8",X"28",X"00",X"28",X"00",X"28",X"A8",X"28",X"08",X"2A",X"A8",X"0A",X"88",X"00",X"00",
		X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",
		X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",X"00",X"00",
		X"0A",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A0",X"2A",X"A0",X"0A",X"80",X"00",X"00",
		X"28",X"08",X"28",X"28",X"28",X"A0",X"2A",X"A0",X"28",X"28",X"28",X"08",X"28",X"08",X"00",X"00",
		X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"2A",X"A8",X"00",X"00",
		X"28",X"28",X"28",X"28",X"22",X"88",X"22",X"88",X"20",X"08",X"20",X"08",X"20",X"08",X"00",X"00",
		X"28",X"08",X"2A",X"08",X"2A",X"08",X"22",X"88",X"20",X"88",X"20",X"A8",X"20",X"28",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"08",X"2A",X"A8",X"28",X"00",X"28",X"00",X"28",X"00",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"20",X"08",X"20",X"08",X"20",X"88",X"28",X"A0",X"0A",X"A8",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"08",X"2A",X"A8",X"28",X"20",X"28",X"28",X"28",X"08",X"00",X"00",
		X"0A",X"A8",X"28",X"08",X"28",X"00",X"2A",X"A8",X"00",X"28",X"20",X"28",X"2A",X"A0",X"00",X"00",
		X"2A",X"A8",X"2A",X"A8",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"00",X"00",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"20",X"08",X"20",X"08",X"28",X"28",X"08",X"20",X"0A",X"A0",X"02",X"80",X"02",X"80",X"00",X"00",
		X"20",X"08",X"20",X"08",X"20",X"08",X"22",X"88",X"22",X"88",X"2A",X"A8",X"08",X"20",X"00",X"00",
		X"20",X"08",X"28",X"28",X"0A",X"A0",X"02",X"80",X"0A",X"A0",X"28",X"28",X"20",X"08",X"00",X"00",
		X"20",X"08",X"20",X"08",X"28",X"28",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",X"00",X"00",
		X"2A",X"A8",X"20",X"28",X"00",X"A0",X"02",X"80",X"0A",X"00",X"28",X"08",X"2A",X"A8",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"50",X"01",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"41",X"55",X"55",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"45",X"55",X"55",
		X"AA",X"AA",X"80",X"02",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"80",X"AA",X"00",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"A5",
		X"AA",X"AA",X"AA",X"A5",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"0A",X"95",X"00",X"25",
		X"AA",X"AA",X"55",X"55",X"55",X"6A",X"55",X"6B",X"55",X"6A",X"55",X"50",X"55",X"5A",X"55",X"5A",
		X"AA",X"AA",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"55",X"55",X"A9",X"55",X"E9",X"55",X"A9",X"55",X"55",X"55",X"A5",X"55",X"A5",X"55",
		X"AA",X"AA",X"55",X"55",X"54",X"00",X"54",X"00",X"54",X"30",X"54",X"00",X"55",X"54",X"55",X"02",
		X"AA",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",
		X"AA",X"AA",X"A5",X"55",X"A5",X"55",X"A5",X"15",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"AA",X"AA",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",
		X"00",X"2A",X"00",X"25",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"25",
		X"00",X"2A",X"00",X"25",X"00",X"95",X"00",X"95",X"40",X"95",X"50",X"95",X"58",X"95",X"54",X"25",
		X"AA",X"02",X"55",X"02",X"55",X"02",X"51",X"02",X"55",X"06",X"55",X"15",X"55",X"14",X"55",X"10",
		X"AA",X"10",X"55",X"10",X"55",X"00",X"54",X"00",X"40",X"14",X"01",X"50",X"15",X"13",X"55",X"13",
		X"AA",X"50",X"54",X"50",X"54",X"50",X"54",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"55",X"13",X"AA",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"00",X"A0",X"00",
		X"54",X"50",X"AA",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"AA",X"50",
		X"55",X"55",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"AA",X"96",X"55",X"55",X"45",X"54",X"55",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"55",X"50",X"AA",X"50",X"15",X"50",X"15",X"50",X"15",X"50",X"15",X"50",X"15",X"50",X"AA",X"50",
		X"55",X"55",X"AA",X"AA",X"55",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"54",X"16",X"14",X"55",X"58",X"54",X"48",X"50",X"48",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"14",X"50",X"56",X"50",X"54",X"50",X"40",X"50",X"55",X"50",X"55",X"50",X"45",X"50",X"55",X"50",
		X"95",X"55",X"94",X"54",X"59",X"55",X"55",X"45",X"56",X"51",X"65",X"95",X"55",X"54",X"55",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"96",X"56",X"00",X"00",X"00",X"00",X"55",X"55",
		X"58",X"54",X"65",X"55",X"95",X"55",X"55",X"54",X"95",X"65",X"55",X"55",X"56",X"55",X"55",X"96",
		X"01",X"00",X"41",X"50",X"45",X"50",X"55",X"40",X"59",X"50",X"55",X"44",X"55",X"54",X"55",X"50",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"84",X"50",X"55",X"50",X"55",X"50",X"59",X"50",X"55",X"50",X"65",X"50",X"55",X"50",X"55",X"50",
		X"55",X"55",X"59",X"55",X"55",X"54",X"95",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"55",X"59",X"55",X"55",X"55",X"55",X"56",X"55",X"5A",X"55",X"65",X"55",X"51",X"69",X"55",X"55",
		X"04",X"11",X"04",X"45",X"41",X"59",X"50",X"59",X"16",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"AA",X"AA",X"02",X"AA",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"40",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"44",X"01",X"45",
		X"00",X"59",X"00",X"56",X"15",X"55",X"45",X"54",X"55",X"69",X"59",X"95",X"66",X"55",X"95",X"55",
		X"55",X"15",X"55",X"56",X"55",X"56",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"55",X"56",X"45",X"55",X"59",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"56",X"5A",X"55",X"95",
		X"14",X"50",X"55",X"50",X"15",X"50",X"01",X"50",X"46",X"50",X"59",X"50",X"55",X"50",X"55",X"50",
		X"01",X"55",X"01",X"55",X"00",X"54",X"05",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"01",
		X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",
		X"00",X"14",X"00",X"55",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"AA",X"A8",X"0A",X"AA",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"54",X"14",X"55",X"55",X"55",X"54",X"54",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",
		X"50",X"50",X"54",X"50",X"55",X"50",X"55",X"50",X"54",X"50",X"55",X"50",X"68",X"50",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"56",X"55",X"55",X"55",X"5A",X"55",X"55",X"55",X"41",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",X"05",X"00",X"14",X"00",X"40",X"00",X"54",X"00",
		X"44",X"54",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"59",X"55",X"59",X"55",
		X"51",X"54",X"55",X"50",X"54",X"50",X"55",X"44",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"50",
		X"45",X"6A",X"54",X"AA",X"55",X"1A",X"55",X"56",X"51",X"5A",X"55",X"6A",X"15",X"1A",X"54",X"46",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"06",X"AA",X"52",X"AA",X"5A",X"AA",
		X"AA",X"AA",X"A8",X"2A",X"A8",X"2A",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A8",X"2A",X"AA",X"AA",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"00",X"00",X"AA",X"AA",X"A8",X"08",X"AA",X"28",X"AA",X"28",X"AA",X"28",X"AA",X"28",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"28",X"20",X"88",X"A2",X"28",X"20",X"88",X"A2",X"88",X"20",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"A0",X"AA",X"8A",X"AA",X"A2",X"AA",X"A8",X"AA",X"80",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"8A",X"08",X"8A",X"28",X"8A",X"08",X"8A",X"28",X"82",X"08",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"20",X"2A",X"A8",X"AA",X"28",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"AA",X"80",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"88",X"20",X"88",X"00",X"88",X"88",X"88",X"A8",X"88",X"A8",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"82",X"AA",X"8A",X"AA",X"82",X"AA",X"8A",X"AA",X"82",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"28",X"20",X"28",X"A2",X"28",X"20",X"28",X"A2",X"08",X"22",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"80",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"41",X"55",X"84",X"54",X"00",X"00",X"00",X"00",
		X"01",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"45",X"50",X"51",X"50",X"14",X"50",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"55",X"50",X"05",X"50",X"00",X"50",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"15",X"55",X"55",X"95",X"00",X"54",X"00",X"00",
		X"00",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"54",X"50",X"00",X"50",X"00",X"50",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"59",X"15",X"14",X"05",X"00",X"00",X"00",X"00",
		X"0A",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"54",X"50",X"50",X"50",X"00",X"50",X"00",X"10",
		X"00",X"00",X"31",X"44",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"10",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"50",X"00",X"50",X"00",X"50",X"55",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"10",
		X"80",X"14",X"01",X"50",X"15",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"92",X"AA",X"56",X"AA",X"52",X"AA",X"52",X"80",X"52",X"00",X"52",X"00",X"52",X"55",X"52",
		X"AA",X"52",X"00",X"50",X"00",X"50",X"55",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"10",
		X"AA",X"52",X"AA",X"52",X"AA",X"7F",X"AA",X"7F",X"AA",X"52",X"AA",X"52",X"AA",X"52",X"AA",X"52",
		X"00",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"55",X"56",X"AA",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"02",X"55",X"02",X"55",X"02",X"51",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"02",X"A0",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"55",X"5A",X"55",X"50",X"55",X"6A",X"55",X"6B",X"55",X"6A",X"55",X"50",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"55",X"55",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"A9",X"55",X"E9",X"55",X"A9",X"55",X"05",X"55",X"55",X"55",
		X"AA",X"AA",X"A1",X"55",X"A1",X"55",X"A1",X"55",X"A1",X"55",X"A1",X"55",X"A1",X"41",X"A1",X"00",
		X"00",X"03",X"00",X"0F",X"00",X"3B",X"00",X"EB",X"03",X"AB",X"03",X"AB",X"03",X"AB",X"0E",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"C0",X"00",X"B0",X"00",X"B0",X"00",X"AC",X"00",X"AB",X"00",X"AA",X"C0",X"AA",X"B0",X"AA",X"AC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"AA",X"0E",X"AA",X"0E",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"00",X"EA",
		X"00",X"00",X"00",X"3F",X"03",X"FA",X"0F",X"AA",X"0E",X"AA",X"3E",X"AA",X"3A",X"AA",X"3A",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"AA",X"AA",X"A0",X"0A",X"80",X"00",X"82",X"A8",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"82",X"AA",X"80",X"A0",X"A0",X"02",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"28",X"82",X"00",X"8A",X"88",X"0A",X"88",X"82",X"08",X"A0",X"28",
		X"AA",X"AA",X"AA",X"AA",X"82",X"A0",X"20",X"82",X"28",X"8A",X"28",X"8A",X"28",X"A2",X"28",X"08",
		X"AA",X"AA",X"AA",X"AA",X"28",X"82",X"08",X"28",X"88",X"AA",X"88",X"2A",X"00",X"2A",X"08",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"AA",X"A8",X"82",X"28",X"08",X"28",X"2A",X"28",X"2A",X"28",X"08",X"28",X"80",X"82",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A2",X"82",X"A2",X"82",X"A2",X"82",X"A2",X"82",X"A2",X"82",X"08",X"20",
		X"22",X"AA",X"22",X"AA",X"22",X"82",X"22",X"08",X"22",X"2A",X"22",X"2A",X"82",X"08",X"08",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"8A",X"AA",X"22",X"AA",X"22",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"40",X"A1",X"50",X"00",X"50",X"A8",X"50",X"E8",X"50",X"A8",X"50",X"01",X"50",X"54",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"80",X"0A",
		X"A8",X"A2",X"A8",X"AA",X"28",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"A2",X"02",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"80",X"A2",X"08",X"00",X"2A",X"20",X"2A",X"20",X"08",X"20",X"80",X"A0",
		X"AA",X"AA",X"AA",X"80",X"0A",X"2A",X"82",X"2A",X"A2",X"82",X"A2",X"A8",X"A2",X"A8",X"A0",X"02",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"A2",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"AB",X"8A",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"20",X"02",X"80",X"A0",X"82",X"A8",X"82",X"A8",X"82",X"A8",X"82",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A2",X"A2",X"82",X"A2",X"8A",X"88",X"8A",X"88",X"A0",
		X"8A",X"AA",X"0A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"80",X"02",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"00",X"A0",
		X"88",X"AA",X"88",X"AA",X"88",X"A0",X"88",X"82",X"88",X"8A",X"88",X"8A",X"A0",X"82",X"02",X"20",
		X"AA",X"AA",X"AA",X"AA",X"88",X"A2",X"08",X"A2",X"88",X"A2",X"88",X"A2",X"08",X"A2",X"22",X"00",
		X"AA",X"AA",X"AA",X"AA",X"80",X"A2",X"2A",X"20",X"28",X"A2",X"02",X"A0",X"2A",X"80",X"80",X"20",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"A8",X"A8",X"A0",X"AA",X"A2",X"0A",X"82",X"A0",X"82",X"AA",
		X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"A2",X"AA",X"A8",X"A8",X"AA",X"02",
		X"0A",X"AA",X"0A",X"AA",X"08",X"82",X"08",X"28",X"08",X"A8",X"28",X"A8",X"A8",X"A8",X"A8",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"22",X"AA",X"0A",X"AA",X"8A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"8A",X"8A",X"8A",X"2A",X"80",X"A8",X"8A",X"A2",X"20",X"0A",
		X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"82",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",
		X"AA",X"A2",X"AA",X"82",X"AA",X"22",X"A8",X"A2",X"A8",X"A2",X"A8",X"A2",X"AA",X"0A",X"AA",X"AA",
		X"A0",X"20",X"A8",X"A8",X"A8",X"20",X"AA",X"02",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"02",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"08",X"28",X"8A",X"28",X"8A",X"28",X"8A",X"82",X"A0",
		X"AA",X"A8",X"AA",X"A0",X"AA",X"A2",X"2A",X"A2",X"2A",X"A2",X"2A",X"A2",X"2A",X"A0",X"AA",X"A8",
		X"08",X"2A",X"A2",X"2A",X"A2",X"2A",X"AA",X"02",X"AA",X"28",X"AA",X"28",X"A2",X"28",X"0A",X"28",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"88",X"8A",X"22",X"8A",X"22",X"8A",X"22",X"A0",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"22",X"0A",X"88",X"A2",X"88",X"A2",X"88",X"A2",X"28",X"0A",
		X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"82",X"A0",X"28",X"8A",X"00",X"8A",X"2A",X"8A",X"80",X"A0",
		X"2A",X"A0",X"2A",X"A2",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"8A",X"AA",
		X"00",X"22",X"8A",X"22",X"8A",X"A2",X"8A",X"A0",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"02",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"0A",X"88",X"A2",X"88",X"02",X"88",X"AA",X"8A",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"82",X"82",X"0A",X"88",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"82",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",
		X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"AA",X"AA",X"AA",X"00",X"02",X"28",X"A2",X"A8",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"88",X"8A",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"0A",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"0A",X"02",X"A2",X"2A",X"A2",X"0A",X"A2",X"A2",X"0A",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"A8",X"A8",X"A2",X"A8",X"A2",X"A8",X"A2",X"A0",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"20",X"A8",X"8A",X"22",X"80",X"20",X"8A",X"A2",X"A0",X"28",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"28",X"0A",X"88",X"AA",X"08",X"0A",X"AA",X"8A",X"08",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"0A",X"0A",X"82",X"0A",X"A2",
		X"00",X"00",X"00",X"00",X"05",X"00",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"54",
		X"00",X"00",X"00",X"00",X"01",X"40",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"54",
		X"00",X"00",X"00",X"00",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"40",X"55",X"40",X"55",
		X"00",X"00",X"00",X"00",X"55",X"00",X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"01",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"50",X"01",X"54",X"05",X"55",X"55",X"54",X"15",X"54",X"05",X"50",X"01",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"50",
		X"00",X"00",X"00",X"00",X"40",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"15",X"50",X"05",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"40",X"05",X"50",X"55",X"54",X"55",X"54",X"15",X"54",X"05",X"54",X"01",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"51",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",
		X"54",X"2A",X"54",X"AA",X"54",X"AA",X"54",X"AA",X"54",X"2A",X"14",X"0A",X"15",X"02",X"15",X"00",
		X"55",X"55",X"50",X"05",X"52",X"A1",X"52",X"A1",X"52",X"A8",X"52",X"AA",X"52",X"AA",X"52",X"AA",
		X"05",X"55",X"01",X"55",X"29",X"55",X"29",X"55",X"29",X"55",X"29",X"55",X"29",X"55",X"09",X"55",
		X"85",X"54",X"81",X"54",X"A1",X"54",X"A1",X"55",X"A1",X"55",X"A1",X"55",X"A1",X"55",X"21",X"55",
		X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"60",X"55",X"40",
		X"58",X"01",X"5A",X"21",X"5A",X"A1",X"5A",X"A1",X"5A",X"A1",X"58",X"A1",X"50",X"21",X"50",X"01",
		X"08",X"55",X"28",X"55",X"28",X"55",X"20",X"55",X"21",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"55",X"80",X"55",X"A0",X"55",X"A0",X"55",X"60",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"50",
		X"00",X"15",X"0A",X"15",X"AA",X"15",X"AA",X"15",X"AA",X"15",X"82",X"15",X"80",X"15",X"00",X"55",
		X"15",X"55",X"05",X"55",X"85",X"56",X"85",X"56",X"85",X"56",X"85",X"56",X"85",X"56",X"85",X"56",
		X"01",X"54",X"A1",X"54",X"A0",X"56",X"A8",X"56",X"A8",X"16",X"AA",X"16",X"AA",X"06",X"AA",X"86",
		X"15",X"54",X"15",X"56",X"15",X"56",X"15",X"56",X"15",X"56",X"15",X"56",X"15",X"56",X"15",X"56",
		X"15",X"50",X"15",X"6A",X"15",X"6A",X"15",X"AA",X"15",X"AA",X"16",X"AA",X"16",X"AA",X"1A",X"AA",
		X"AA",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",
		X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",
		X"2A",X"A8",X"0A",X"A8",X"0A",X"A8",X"02",X"A8",X"02",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"28",
		X"85",X"56",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"50",X"01",X"50",X"01",X"50",X"01",X"50",X"01",X"54",X"01",X"54",X"01",X"54",X"01",X"54",X"01",
		X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",
		X"21",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"54",X"55",X"54",
		X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"52",X"AA",X"50",X"0A",X"50",X"0A",X"50",X"02",X"50",X"00",X"50",X"00",X"50",X"04",X"50",X"04",
		X"85",X"00",X"85",X"00",X"A1",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"2A",X"80",
		X"55",X"4A",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"50",
		X"2A",X"80",X"0A",X"80",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"50",X"00",
		X"50",X"04",X"54",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"95",
		X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"41",X"55",
		X"55",X"50",X"55",X"50",X"15",X"50",X"05",X"50",X"85",X"54",X"81",X"55",X"A1",X"55",X"A0",X"55",
		X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",
		X"54",X"01",X"54",X"01",X"54",X"01",X"54",X"01",X"54",X"01",X"54",X"01",X"55",X"01",X"55",X"01",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",
		X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"05",X"55",
		X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"05",X"54",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"85",X"55",X"85",X"55",X"81",X"55",X"A1",X"55",X"A0",X"55",X"A8",X"55",X"A8",X"55",X"28",X"15",
		X"55",X"85",X"55",X"85",X"55",X"85",X"56",X"85",X"56",X"85",X"5A",X"85",X"5A",X"85",X"5A",X"05",
		X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"41",X"55",X"41",X"55",X"41",X"55",X"41",X"55",X"41",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"A8",X"55",X"A8",X"55",X"A8",X"55",X"A8",X"55",X"A8",X"55",X"28",X"55",X"20",X"55",X"01",X"55",
		X"41",X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"52",X"A5",X"52",X"AA",X"52",X"AA",X"52",X"AA",X"52",X"AA",X"50",X"2A",X"50",X"0A",X"50",X"00",
		X"50",X"00",X"50",X"00",X"94",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"10",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"41",X"55",X"49",
		X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"42",X"55",X"40",
		X"28",X"10",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"01",X"50",X"01",X"50",X"55",X"50",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"55",X"40",X"55",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"A9",X"55",X"AA",X"95",
		X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"15",X"5A",X"02",X"AA",X"0A",X"AA",X"AA",X"AA",
		X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",
		X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"5A",X"5A",X"8A",X"AA",X"8A",X"AA",X"AA",
		X"6A",X"05",X"6A",X"05",X"68",X"05",X"A0",X"15",X"A0",X"55",X"A0",X"55",X"81",X"2A",X"80",X"2A",
		X"2A",X"15",X"2A",X"15",X"0A",X"05",X"0A",X"85",X"02",X"81",X"02",X"A2",X"02",X"AA",X"00",X"AA",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"54",X"05",X"54",X"05",X"54",X"15",X"54",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"5A",X"55",X"6A",X"96",X"AA",X"AA",X"AA",
		X"40",X"AA",X"54",X"AA",X"50",X"2A",X"00",X"2A",X"00",X"08",X"00",X"00",X"00",X"00",X"80",X"00",
		X"80",X"2A",X"80",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A9",X"AA",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"02",X"AA",X"00",X"2A",X"00",X"02",
		X"55",X"55",X"95",X"55",X"AA",X"55",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"A5",X"58",X"A9",X"54",X"AA",X"95",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"55",X"50",X"55",X"54",X"55",X"54",X"95",X"54",X"A5",X"54",X"A9",X"54",X"AA",X"54",X"AA",X"A5",
		X"AA",X"A5",X"AA",X"A9",X"AA",X"A8",X"AA",X"A8",X"0A",X"A0",X"02",X"A8",X"00",X"2A",X"00",X"0A",
		X"2A",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",
		X"80",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"80",X"28",X"00",X"00",X"00",X"00",X"00",
		X"55",X"58",X"55",X"68",X"55",X"AA",X"56",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"16",X"00",X"1A",
		X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"56",X"55",X"56",
		X"00",X"0A",X"54",X"2A",X"50",X"2A",X"40",X"AA",X"40",X"AA",X"00",X"A8",X"00",X"A0",X"A8",X"00",
		X"AA",X"80",X"AA",X"00",X"A8",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",
		X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"20",X"00",X"20",X"20",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A9",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",
		X"28",X"02",X"28",X"02",X"28",X"02",X"08",X"02",X"08",X"02",X"08",X"02",X"08",X"02",X"08",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"A8",X"00",X"A8",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"02",X"28",X"02",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"80",X"2A",X"80",X"2A",X"A0",X"AA",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"A8",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5A",X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"AA",X"56",X"A8",X"56",X"A8",X"5A",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"2A",X"00",X"2A",
		X"5A",X"A0",X"6A",X"80",X"6A",X"80",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"A8",X"02",X"A0",X"0A",X"80",X"2A",X"80",X"AA",X"00",
		X"AA",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"A0",X"02",X"A0",X"02",
		X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"00",X"02",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"2A",X"00",X"2A",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",
		X"AA",X"A0",X"2A",X"80",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"A8",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"02",
		X"A0",X"0A",X"A0",X"0A",X"80",X"0A",X"80",X"2A",X"80",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"02",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",
		X"2A",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"AA",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"AA",X"AA",X"02",X"8A",X"02",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"A0",X"02",X"A8",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"AA",X"00",X"AA",X"02",X"AA",X"02",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"0A",X"02",X"0A",X"02",
		X"08",X"02",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",X"0A",X"20",X"0A",
		X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"80",X"0A",X"80",X"02",X"00",X"00",X"00",X"02",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"AA",X"80",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",
		X"00",X"0A",X"00",X"0A",X"00",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A0",X"0A",X"A0",X"02",X"80",X"00",X"80",X"00",X"A0",X"02",X"A8",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"AA",X"02",X"AA",
		X"02",X"80",X"02",X"80",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A8",X"02",X"A8",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",
		X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",
		X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",
		X"80",X"02",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"80",X"02",X"80",X"02",X"80",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"A0",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A5",X"2A",X"A9",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"0A",
		X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"09",X"00",X"02",X"00",X"02",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",
		X"55",X"50",X"55",X"50",X"95",X"50",X"A5",X"54",X"A9",X"54",X"AA",X"54",X"AA",X"95",X"AA",X"A5",
		X"55",X"00",X"55",X"00",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",
		X"00",X"95",X"00",X"A5",X"00",X"A9",X"00",X"A9",X"00",X"55",X"80",X"55",X"80",X"15",X"80",X"25",
		X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"00",
		X"01",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"95",X"02",X"95",X"02",X"95",
		X"29",X"55",X"29",X"55",X"29",X"55",X"29",X"55",X"09",X"55",X"09",X"55",X"09",X"55",X"01",X"55",
		X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"42",X"95",X"52",X"95",X"50",X"95",X"54",X"95",X"54",X"A5",X"54",X"A5",X"54",X"25",X"55",
		X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"42",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",
		X"28",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"48",X"00",X"08",X"00",X"28",X"00",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"A9",X"55",X"A9",X"55",X"29",X"55",X"09",X"55",X"09",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",
		X"55",X"50",X"55",X"54",X"55",X"54",X"95",X"54",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A9",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"55",X"50",
		X"6A",X"AA",X"6A",X"9A",X"6A",X"96",X"59",X"D6",X"55",X"D6",X"55",X"D5",X"57",X"55",X"57",X"55",
		X"A9",X"AA",X"A9",X"A6",X"A5",X"A6",X"95",X"65",X"55",X"55",X"55",X"55",X"D1",X"55",X"54",X"55",
		X"AA",X"AA",X"AA",X"A6",X"AA",X"A5",X"AA",X"95",X"AA",X"95",X"69",X"95",X"59",X"75",X"59",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"9A",X"69",X"99",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"6A",X"AA",X"5A",X"A6",X"5A",X"A5",X"5A",X"95",X"56",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"9A",X"AA",X"9A",X"9A",X"96",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"A9",X"AA",X"A6",X"69",X"A5",X"55",X"55",X"55",X"55",X"55",X"71",X"55",X"D5",X"55",X"D5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"46",X"AA",
		X"55",X"55",X"57",X"55",X"D5",X"D7",X"D5",X"75",X"55",X"5D",X"5D",X"5F",X"55",X"57",X"57",X"57",
		X"55",X"55",X"D5",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"54",X"D5",X"55",X"55",X"15",X"55",
		X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"7D",X"57",X"55",X"5D",X"55",X"55",X"57",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"54",X"55",X"D5",X"57",X"55",X"55",X"54",X"5D",X"55",X"55",X"51",X"55",X"54",
		X"55",X"A9",X"56",X"A9",X"55",X"A5",X"55",X"95",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A6",X"A6",X"57",X"D6",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"9A",X"AA",X"56",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"A9",X"A9",X"6A",X"A5",X"6A",X"55",X"69",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"9A",X"5A",X"9A",X"5A",X"5A",X"55",X"56",X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"AA",X"AA",X"AA",X"AA",X"A9",X"A9",X"99",X"95",X"75",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",
		X"AA",X"AA",X"6A",X"9A",X"5A",X"5A",X"55",X"59",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"69",X"66",X"69",X"55",X"69",X"55",X"59",X"55",X"55",X"55",X"55",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"99",X"6A",X"59",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"D5",
		X"55",X"D4",X"55",X"55",X"55",X"55",X"55",X"45",X"5D",X"45",X"57",X"55",X"55",X"D5",X"55",X"55",
		X"55",X"55",X"57",X"55",X"57",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"57",X"55",
		X"D5",X"55",X"55",X"55",X"75",X"55",X"75",X"55",X"55",X"D5",X"57",X"55",X"57",X"55",X"55",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"75",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",
		X"55",X"55",X"45",X"D5",X"55",X"55",X"45",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"54",X"51",
		X"55",X"15",X"55",X"51",X"55",X"15",X"41",X"55",X"55",X"50",X"55",X"55",X"45",X"41",X"55",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"D5",X"57",X"55",X"55",X"55",X"D5",X"55",X"75",X"75",X"D5",X"55",X"55",X"55",X"D5",X"5D",
		X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"54",X"55",X"55",X"55",X"51",X"55",X"D5",X"75",
		X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",
		X"5D",X"55",X"55",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",X"5D",X"55",X"57",X"55",X"55",X"55",
		X"95",X"55",X"E5",X"55",X"F9",X"55",X"FE",X"55",X"FE",X"55",X"AA",X"95",X"AA",X"95",X"AA",X"A5",
		X"55",X"5D",X"55",X"75",X"5D",X"75",X"55",X"55",X"5D",X"57",X"57",X"55",X"55",X"55",X"15",X"D5",
		X"55",X"57",X"5D",X"55",X"D5",X"55",X"75",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",
		X"55",X"57",X"D5",X"55",X"D5",X"55",X"75",X"57",X"5D",X"55",X"55",X"57",X"75",X"55",X"D5",X"55",
		X"55",X"55",X"D5",X"57",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",
		X"D5",X"55",X"51",X"55",X"54",X"D5",X"D5",X"54",X"71",X"55",X"D5",X"45",X"55",X"54",X"54",X"45",
		X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"51",X"45",X"55",X"55",X"55",X"54",X"55",X"55",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5D",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"75",X"55",X"D5",X"57",X"55",X"55",X"D5",X"55",X"75",X"55",X"DD",X"55",X"75",X"55",X"55",
		X"55",X"D5",X"55",X"D5",X"55",X"75",X"55",X"75",X"55",X"DD",X"55",X"75",X"55",X"57",X"55",X"5D",
		X"55",X"51",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"41",X"55",X"51",X"55",X"15",X"55",X"45",
		X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"57",X"55",X"55",
		X"55",X"55",X"55",X"D5",X"55",X"75",X"55",X"D5",X"57",X"55",X"5D",X"55",X"77",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5C",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",X"15",X"51",X"55",X"55",X"55",X"45",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"5D",X"55",X"75",X"55",X"75",X"55",X"5D",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"51",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",
		X"FF",X"E5",X"FF",X"E5",X"FF",X"F9",X"FF",X"F9",X"FF",X"F9",X"FF",X"F9",X"FF",X"F9",X"AA",X"AA",
		X"D5",X"55",X"75",X"55",X"5D",X"54",X"5D",X"55",X"57",X"55",X"55",X"D5",X"55",X"51",X"55",X"55",
		X"55",X"55",X"F5",X"55",X"75",X"55",X"D5",X"55",X"75",X"55",X"75",X"55",X"5D",X"55",X"57",X"55",
		X"D5",X"57",X"55",X"D5",X"55",X"55",X"57",X"55",X"55",X"55",X"75",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"57",X"55",X"55",X"55",X"75",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",
		X"5D",X"15",X"55",X"51",X"55",X"55",X"54",X"51",X"55",X"55",X"75",X"11",X"5C",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"45",X"5D",X"55",X"55",X"55",X"55",X"51",X"75",X"55",X"55",X"14",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"07",X"55",X"00",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"54",X"55",X"51",X"55",X"55",X"55",X"75",X"55",X"55",X"15",X"5D",X"00",X"00",X"00",X"00",
		X"55",X"75",X"55",X"5D",X"55",X"17",X"54",X"55",X"55",X"57",X"55",X"55",X"00",X"07",X"00",X"00",
		X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"57",X"55",X"55",X"40",X"50",X"00",X"00",X"00",
		X"D5",X"D5",X"55",X"75",X"55",X"75",X"55",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"05",X"00",X"15",X"00",X"00",X"00",X"00",
		X"54",X"51",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"11",X"51",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"51",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"D5",X"55",X"55",X"55",X"75",X"55",X"D5",X"00",X"3D",X"00",X"03",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"00",X"00",
		X"75",X"55",X"75",X"55",X"75",X"55",X"5D",X"55",X"75",X"40",X"75",X"00",X"50",X"01",X"00",X"00",
		X"55",X"55",X"54",X"55",X"55",X"55",X"45",X"15",X"15",X"55",X"51",X"45",X"55",X"51",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"01",X"54",X"00",X"00",X"00",
		X"95",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"AA",X"01",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"AA",X"55",X"00",X"AA",X"00",X"00",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A5",X"00",X"0A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"45",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A5",
		X"55",X"55",X"55",X"55",X"50",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"01",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"45",X"55",X"55",X"55",X"55",
		X"00",X"09",X"02",X"A5",X"09",X"55",X"25",X"55",X"95",X"69",X"95",X"55",X"A5",X"55",X"0A",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"BF",X"FF",X"AB",X"FF",X"AE",X"FF",X"AF",X"BF",X"AF",X"EA",X"BB",X"EA",X"BE",X"FA",
		X"55",X"AA",X"56",X"AA",X"5B",X"FE",X"5B",X"FE",X"6F",X"AA",X"6E",X"FE",X"AE",X"FE",X"AB",X"EA",
		X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"55",X"25",X"55",X"0A",X"95",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"6A",X"5A",X"55",X"55",X"A9",X"55",X"02",X"A9",X"00",X"02",X"00",X"00",X"00",X"0A",
		X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",
		X"BE",X"FB",X"EF",X"BB",X"EF",X"BE",X"FB",X"BE",X"BB",X"BE",X"BB",X"BE",X"AB",X"EE",X"AA",X"EF",
		X"AA",X"BE",X"AA",X"BE",X"AA",X"AA",X"EA",X"A0",X"EE",X"A0",X"EE",X"E0",X"BE",X"E0",X"BB",X"E0",
		X"00",X"A5",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"55",X"55",X"55",X"A9",X"55",X"02",X"95",X"00",X"25",X"00",X"09",X"00",X"A9",X"00",X"95",
		X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"55",X"02",X"95",X"00",X"25",X"00",X"29",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"95",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"95",X"55",X"25",X"59",X"09",X"55",
		X"55",X"15",X"54",X"55",X"51",X"50",X"45",X"45",X"15",X"15",X"54",X"55",X"51",X"55",X"51",X"55",
		X"14",X"55",X"45",X"15",X"51",X"45",X"51",X"51",X"54",X"54",X"55",X"15",X"55",X"45",X"55",X"50",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"75",X"55",X"7D",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",
		X"50",X"55",X"05",X"56",X"55",X"56",X"55",X"02",X"50",X"02",X"40",X"5B",X"05",X"5B",X"40",X"57",
		X"50",X"05",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"05",X"55",X"50",X"55",X"55",X"05",
		X"55",X"75",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"5D",X"55",X"D5",X"55",X"55",X"57",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"41",X"55",X"55",X"55",X"55",X"00",
		X"55",X"5D",X"55",X"75",X"D5",X"75",X"FD",X"57",X"55",X"55",X"55",X"75",X"55",X"57",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"57",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5D",X"DD",X"55",X"DD",X"55",X"75",X"55",X"57",X"55",X"D5",X"55",X"75",X"55",X"51",X"D5",
		X"55",X"5D",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"A0",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"9A",
		X"55",X"55",X"55",X"55",X"55",X"50",X"50",X"55",X"55",X"55",X"55",X"55",X"5A",X"9A",X"60",X"00",
		X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"5A",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A6",X"9A",X"00",X"00",X"00",X"03",X"FF",X"0C",X"00",
		X"55",X"55",X"55",X"55",X"5A",X"AA",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"55",X"56",X"69",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",X"00",X"00",
		X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"15",X"3F",X"55",X"C3",X"D5",X"00",X"37",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5D",X"55",X"53",X"F5",X"50",X"0D",X"70",X"0F",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"73",X"55",X"C3",X"55",X"0D",X"55",X"0D",X"55",X"0D",X"F5",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"FD",X"55",X"03",X"DD",X"03",X"55",X"03",X"55",
		X"00",X"D5",X"00",X"37",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"FC",X"03",X"F0",
		X"55",X"55",X"69",X"A8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"56",X"9A",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"6A",X"9A",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"15",X"15",X"55",X"55",X"55",X"55",X"55",X"56",X"69",X"68",X"80",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"56",X"96",X"58",X"00",
		X"55",X"5A",X"55",X"6E",X"55",X"6E",X"55",X"BE",X"55",X"BA",X"56",X"F8",X"02",X"A8",X"02",X"A0",
		X"AA",X"AA",X"AA",X"FF",X"BE",X"BF",X"AF",X"BF",X"0B",X"EF",X"02",X"AA",X"02",X"AA",X"02",X"FA",
		X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"41",X"00",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"AA",X"AA",
		X"80",X"BE",X"20",X"BE",X"20",X"BE",X"20",X"AA",X"20",X"AA",X"20",X"BE",X"20",X"BE",X"20",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"55",X"54",X"55",X"40",X"54",X"01",X"41",X"05",X"15",X"15",X"45",X"41",X"51",X"54",X"54",X"15",
		X"10",X"55",X"05",X"50",X"55",X"44",X"54",X"10",X"55",X"05",X"55",X"50",X"15",X"55",X"45",X"55",
		X"56",X"E2",X"02",X"E2",X"02",X"A2",X"55",X"A2",X"05",X"62",X"10",X"56",X"41",X"05",X"54",X"10",
		X"7B",X"AA",X"57",X"AB",X"05",X"6B",X"00",X"57",X"50",X"05",X"55",X"00",X"55",X"50",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"55",X"55",X"05",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"04",X"00",X"55",X"55",
		X"41",X"55",X"04",X"00",X"50",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"40",X"55",X"55",X"15",X"55",X"41",X"55",X"54",X"05",X"15",X"50",X"40",X"55",X"55",X"05",
		X"50",X"55",X"55",X"01",X"05",X"54",X"54",X"15",X"55",X"41",X"55",X"54",X"55",X"55",X"55",X"55",
		X"55",X"41",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"14",X"10",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"10",X"00",X"55",X"55",
		X"55",X"55",X"00",X"04",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"01",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"50",X"55",X"55",
		X"55",X"55",X"00",X"50",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"00",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"10",X"55",X"55",
		X"55",X"55",X"00",X"14",X"40",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"54",X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"01",X"55",X"55",
		X"01",X"44",X"05",X"51",X"55",X"45",X"54",X"14",X"41",X"51",X"15",X"05",X"50",X"55",X"05",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"41",X"55",X"14",X"15",X"41",X"45",X"14",X"11",
		X"41",X"55",X"14",X"15",X"41",X"41",X"14",X"14",X"01",X"41",X"40",X"14",X"54",X"01",X"55",X"40",
		X"BA",X"AF",X"EE",X"AA",X"EE",X"AA",X"EE",X"EA",X"6E",X"EA",X"56",X"EE",X"05",X"6F",X"00",X"57",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",
		X"A9",X"55",X"FE",X"55",X"FF",X"95",X"FF",X"95",X"FF",X"E5",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",
		X"55",X"55",X"55",X"55",X"55",X"95",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"10",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"59",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A0",X"02",X"A0",X"02",X"80",X"02",X"80",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"0A",
		X"00",X"2A",X"00",X"2A",X"80",X"2A",X"80",X"0A",X"80",X"0A",X"80",X"02",X"00",X"02",X"00",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",
		X"15",X"50",X"41",X"55",X"54",X"55",X"55",X"15",X"55",X"41",X"55",X"54",X"55",X"55",X"55",X"55",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"0A",X"A0",X"0A",X"A0",X"0A",X"80",X"0A",X"00",X"0A",X"00",X"28",X"00",X"20",X"00",X"20",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"0A",
		X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"2A",X"A8",X"2A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"28",
		X"AA",X"0A",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"00",X"28",X"00",X"28",X"00",X"2A",X"80",X"0A",X"80",X"0A",X"A0",X"0A",X"A8",X"0A",X"A8",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"AA",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"80",X"2A",X"80",X"0A",X"80",X"0A",X"80",X"0A",
		X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",
		X"55",X"55",X"05",X"55",X"50",X"55",X"55",X"05",X"55",X"50",X"15",X"55",X"40",X"55",X"55",X"05",
		X"50",X"05",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"05",X"55",X"50",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"04",X"00",X"55",X"55",
		X"00",X"00",X"2A",X"80",X"AA",X"A8",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"2A",X"80",X"AA",X"A0",X"2A",X"80",X"AA",X"80",X"AA",X"82",X"AA",X"82",X"AA",X"82",
		X"00",X"00",X"20",X"2A",X"A8",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"8A",X"AA",X"8A",X"AA",X"82",
		X"00",X"00",X"80",X"AA",X"A2",X"AA",X"80",X"AA",X"A2",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"8A",
		X"00",X"00",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A0",X"8A",
		X"00",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"20",X"A0",X"20",X"A0",X"20",X"A0",X"20",X"A0",X"20",X"20",X"20",X"00",
		X"AA",X"82",X"AA",X"8A",X"20",X"88",X"20",X"88",X"20",X"88",X"20",X"88",X"20",X"88",X"A0",X"88",
		X"AA",X"A2",X"AA",X"A0",X"08",X"20",X"28",X"20",X"22",X"08",X"28",X"08",X"20",X"08",X"02",X"08",
		X"AA",X"8A",X"AA",X"0A",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"08",
		X"A8",X"0A",X"AA",X"0A",X"00",X"88",X"00",X"88",X"20",X"88",X"28",X"88",X"22",X"08",X"20",X"88",
		X"A2",X"AA",X"A2",X"AA",X"08",X"08",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"28",X"08",
		X"2A",X"AA",X"2A",X"A8",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",
		X"2A",X"8A",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"A8",X"2A",X"A0",X"2A",X"80",
		X"AA",X"AA",X"A2",X"AA",X"A0",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"00",X"2A",
		X"AA",X"A8",X"AA",X"A8",X"A2",X"A8",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A8",X"AA",X"A8",X"AA",
		X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"A0",X"2A",X"A8",X"2A",X"A8",X"2A",X"A0",
		X"AA",X"00",X"28",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"A0",X"2A",X"A0",X"20",X"20",X"20",X"20",
		X"00",X"00",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"82",X"80",X"82",
		X"00",X"00",X"02",X"AA",X"8A",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"28",X"00",X"28",
		X"00",X"82",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"00",X"80",X"00",X"80",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"0A",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",
		X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"2A",X"A0",X"2A",X"A0",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"80",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"00",X"00",X"00",
		X"80",X"28",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",X"8A",X"AA",X"02",X"8A",X"00",X"00",X"00",X"00",
		X"28",X"80",X"A2",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"AA",X"00",X"2A",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"80",X"AA",X"A8",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"2A",X"80",X"AA",X"A0",X"2A",X"80",X"AA",X"80",X"AA",X"82",X"AA",X"82",X"AA",X"82",
		X"00",X"00",X"20",X"2A",X"A8",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"8A",X"AA",X"8A",X"AA",X"82",
		X"00",X"00",X"80",X"AA",X"A2",X"AA",X"80",X"AA",X"A2",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"8A",
		X"00",X"00",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A0",X"8A",
		X"00",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"20",X"A0",X"20",X"A0",X"20",X"A0",X"20",X"A0",X"20",X"20",X"20",X"00",
		X"AA",X"82",X"AA",X"8A",X"20",X"88",X"20",X"88",X"20",X"88",X"20",X"88",X"20",X"88",X"A0",X"88",
		X"AA",X"A2",X"AA",X"A0",X"08",X"20",X"28",X"20",X"22",X"08",X"28",X"08",X"20",X"08",X"02",X"08",
		X"AA",X"8A",X"AA",X"0A",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"08",
		X"A8",X"0A",X"AA",X"0A",X"00",X"88",X"00",X"88",X"20",X"88",X"28",X"88",X"22",X"08",X"20",X"88",
		X"A2",X"AA",X"A2",X"AA",X"08",X"08",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"28",X"08",
		X"2A",X"AA",X"2A",X"A8",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",
		X"2A",X"8A",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"A8",X"2A",X"A0",X"2A",X"80",
		X"AA",X"AA",X"A2",X"AA",X"A0",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"00",X"2A",
		X"AA",X"A8",X"AA",X"A8",X"A2",X"A8",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A8",X"AA",X"A8",X"AA",
		X"2A",X"80",X"2A",X"80",X"2A",X"82",X"2A",X"82",X"2A",X"A2",X"2A",X"A8",X"2A",X"A8",X"2A",X"A0",
		X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"A8",X"02",X"08",X"02",X"08",
		X"80",X"00",X"AA",X"A0",X"AA",X"A8",X"AA",X"A2",X"AA",X"AA",X"AA",X"A2",X"08",X"0A",X"02",X"08",
		X"00",X"00",X"02",X"A8",X"0A",X"AA",X"A2",X"AA",X"AA",X"AA",X"A2",X"AA",X"28",X"08",X"08",X"28",
		X"00",X"02",X"2A",X"A8",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A8",X"2A",X"08",X"20",X"08",X"20",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"82",X"AA",X"80",X"AA",X"A0",X"2A",X"20",X"2A",X"20",X"0A",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",
		X"A8",X"00",X"AA",X"00",X"2A",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"20",X"A8",X"2A",X"A8",X"2A",X"AA",X"AA",X"AA",X"AA",X"2A",X"A8",X"00",X"00",X"00",X"00",
		X"20",X"02",X"A0",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"28",X"AA",X"AA",X"2A",X"A2",X"2A",X"82",X"0A",X"80",X"02",X"00",X"00",X"00",X"00",X"00",
		X"02",X"08",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"20",X"00",X"00",X"00",X"00",
		X"02",X"08",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"0A",X"AA",X"02",X"A8",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"A8",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"02",X"AA",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"A0",X"02",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"0A",X"80",X"0A",X"80",X"2A",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",
		X"00",X"AA",X"00",X"AA",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"02",X"80",X"02",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"2A",
		X"AA",X"AA",X"AA",X"82",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"02",X"A0",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",
		X"A8",X"02",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"0A",X"A0",X"0A",
		X"AA",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"A8",X"00",X"A8",X"02",X"AA",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A0",X"2A",X"A0",X"AA",X"A8",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"A8",X"2A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"0A",X"A8",X"0A",X"A0",X"0A",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"80",X"00",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"AA",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"AA",X"80",X"AA",X"00",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"80",
		X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",
		X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"00",X"00",X"00",X"A0",X"2A",X"A8",
		X"00",X"2A",X"A0",X"0A",X"A0",X"0A",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"00",X"02",X"28",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"AA",
		X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",X"AA",X"82",X"AA",X"02",X"AA",X"02",X"A8",X"02",X"A0",X"02",
		X"A0",X"00",X"A0",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",
		X"AA",X"02",X"AA",X"02",X"AA",X"02",X"2A",X"02",X"2A",X"00",X"02",X"00",X"02",X"00",X"02",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"02",X"AA",X"0A",X"AA",
		X"00",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",
		X"AA",X"AA",X"2A",X"A8",X"2A",X"A0",X"2A",X"A0",X"2A",X"A8",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"2A",X"00",X"2A",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"8A",X"0A",X"0A",X"00",X"28",X"00",X"A8",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"2A",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"80",X"80",X"80",X"80",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"28",X"00",X"0A",X"00",X"0A",
		X"2A",X"AA",X"0A",X"A8",X"0A",X"A8",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"00",X"80",X"00",X"80",
		X"80",X"00",X"00",X"00",X"2A",X"80",X"2A",X"80",X"2A",X"A0",X"2A",X"A0",X"2A",X"80",X"28",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",
		X"00",X"0A",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"00",X"80",X"00",
		X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"82",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"A2",
		X"00",X"00",X"A8",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",X"0A",X"80",X"00",X"00",X"80",X"02",
		X"00",X"00",X"2A",X"00",X"AA",X"A0",X"AA",X"A8",X"0A",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"82",
		X"AA",X"80",X"AA",X"00",X"A8",X"0A",X"28",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"A8",X"00",
		X"00",X"AA",X"00",X"2A",X"A0",X"2A",X"A8",X"2A",X"A0",X"2A",X"80",X"0A",X"00",X"0A",X"00",X"0A",
		X"20",X"02",X"20",X"0A",X"20",X"0A",X"20",X"0A",X"20",X"00",X"28",X"00",X"A8",X"00",X"AA",X"00",
		X"A0",X"0A",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"00",X"00",X"00",X"08",X"00",X"AA",X"00",
		X"AA",X"A0",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"8A",X"00",X"0A",X"00",X"2A",X"00",X"A0",X"00",
		X"0A",X"A2",X"00",X"02",X"0A",X"8A",X"0A",X"8A",X"0A",X"A2",X"0A",X"A2",X"0A",X"82",X"00",X"0A",
		X"80",X"28",X"0A",X"08",X"2A",X"88",X"2A",X"88",X"2A",X"88",X"2A",X"88",X"0A",X"08",X"80",X"28",
		X"20",X"A0",X"08",X"28",X"2A",X"28",X"2A",X"28",X"2A",X"28",X"2A",X"28",X"2A",X"28",X"2A",X"2A",
		X"A8",X"28",X"A8",X"20",X"A8",X"20",X"A8",X"28",X"A8",X"2A",X"A8",X"2A",X"28",X"22",X"00",X"A8",
		X"0A",X"AA",X"A2",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"82",X"AA",X"A2",X"AA",X"0A",X"AA",
		X"AA",X"AA",X"8A",X"AA",X"80",X"00",X"82",X"82",X"8A",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",
		X"AA",X"AA",X"A2",X"AA",X"02",X"AA",X"82",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"82",X"A2",X"82",X"A0",X"82",X"22",X"82",X"22",X"82",X"22",X"A0",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"80",X"A2",X"08",X"0A",X"2A",X"2A",X"2A",X"2A",X"08",X"2A",X"80",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A2",X"AA",X"82",X"AA",X"8A",X"AA",X"8A",X"AA",X"A0",
		X"AA",X"AA",X"80",X"AA",X"08",X"22",X"2A",X"0A",X"2A",X"2A",X"2A",X"2A",X"08",X"2A",X"80",X"AA",
		X"AA",X"AA",X"A8",X"0A",X"A0",X"82",X"A2",X"A0",X"A2",X"A2",X"A2",X"A2",X"A0",X"82",X"A8",X"0A",
		X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"00",
		X"AA",X"AA",X"2A",X"AA",X"00",X"00",X"0A",X"82",X"2A",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",
		X"AA",X"AA",X"A8",X"AA",X"00",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"8A",X"AA",X"0A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",X"AA",X"88",X"AA",X"88",X"AA",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"AA",X"88",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"00",X"0A",X"2A",X"82",X"2A",X"A0",X"2A",X"A8",X"2A",X"A8",X"00",X"00",X"2A",X"82",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"00",X"2A",X"2A",X"0A",X"2A",X"82",X"2A",X"A2",X"2A",X"A2",X"2A",X"8A",
		X"AA",X"AA",X"A0",X"8A",X"82",X"08",X"8A",X"88",X"8A",X"88",X"0A",X"88",X"82",X"00",X"A0",X"8A",
		X"A8",X"AA",X"08",X"AA",X"20",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"20",X"8A",X"08",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",
		X"80",X"82",X"2A",X"22",X"2A",X"22",X"2A",X"A0",X"2A",X"A2",X"2A",X"A2",X"2A",X"22",X"80",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"08",X"88",X"A2",X"88",X"A2",X"88",X"A2",X"8A",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"A0",X"A0",X"A2",X"A0",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"A0",X"A8",X"8A",X"22",X"80",X"22",X"8A",X"A2",X"80",X"22",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"28",X"08",X"88",X"A8",X"08",X"08",X"8A",X"88",X"00",X"08",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"28",X"AA",X"28",X"AA",X"28",X"AA",X"02",X"AA",
		X"A0",X"02",X"A8",X"A2",X"A8",X"AA",X"A8",X"08",X"A8",X"AA",X"A8",X"A0",X"A8",X"A2",X"A0",X"28",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",X"AA",X"80",X"AA",
		X"A2",X"22",X"A2",X"22",X"A2",X"82",X"A2",X"82",X"82",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"82",X"08",X"28",X"88",X"00",X"A2",X"2A",X"88",X"80",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"22",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"00",X"8A",X"28",X"AA",X"2A",
		X"AA",X"28",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"A8",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"28",X"22",X"28",X"88",X"28",X"88",X"28",X"88",X"08",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"A0",X"A2",X"8A",X"22",X"80",X"22",X"8A",X"AA",X"80",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",
		X"AA",X"80",X"AA",X"A2",X"AA",X"A2",X"2A",X"A0",X"2A",X"A2",X"2A",X"A2",X"2A",X"A2",X"AA",X"80",
		X"0A",X"AA",X"88",X"AA",X"AA",X"AA",X"20",X"80",X"A8",X"8A",X"A8",X"8A",X"A8",X"8A",X"A0",X"0A",
		X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"A0",X"80",X"28",X"8A",X"28",X"A2",X"28",X"A8",X"20",X"00",
		X"0A",X"AA",X"8A",X"AA",X"8A",X"AA",X"80",X"A8",X"8A",X"22",X"8A",X"20",X"8A",X"22",X"8A",X"28",
		X"AA",X"82",X"AA",X"A2",X"AA",X"A2",X"2A",X"02",X"88",X"A2",X"08",X"A2",X"A8",X"A2",X"0A",X"08",
		X"AA",X"02",X"AA",X"8A",X"AA",X"8A",X"AA",X"A2",X"AA",X"A2",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"A0",X"2A",X"A8",X"8A",X"A8",X"A8",X"22",X"0A",X"22",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"02",
		X"20",X"AA",X"28",X"AA",X"08",X"AA",X"28",X"0A",X"28",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"A2",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"2A",X"8A",X"22",X"8A",X"AA",
		X"8A",X"82",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"02",X"80",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"08",X"A8",X"22",X"22",X"22",X"20",X"2A",X"22",X"2A",X"28",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"2A",X"AA",X"8A",X"AA",X"0A",X"AA",X"AA",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"0A",X"A2",X"8A",X"A2",X"AA",
		X"A2",X"A0",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"80",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"00",X"A0",X"8A",X"A8",X"8A",X"A8",X"8A",X"02",X"80",X"AA",X"8A",X"AA",X"8A",X"AA",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"A8",X"AA",X"AA",X"AA",
		X"A0",X"2A",X"2A",X"88",X"28",X"08",X"22",X"88",X"A0",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"08",X"28",X"A2",X"88",X"A0",X"08",X"A2",X"AA",X"A8",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"80",X"0A",X"00",X"02",X"00",X"00",X"28",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"28",X"00",X"20",X"00",
		X"80",X"0A",X"00",X"0A",X"00",X"02",X"00",X"00",X"28",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",X"2A",X"A0",X"0A",X"80",
		X"AA",X"A8",X"AA",X"A0",X"AA",X"80",X"AA",X"02",X"AA",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",
		X"28",X"00",X"28",X"00",X"28",X"02",X"08",X"00",X"08",X"00",X"0A",X"00",X"02",X"00",X"00",X"A0",
		X"0A",X"AA",X"00",X"AA",X"A0",X"2A",X"A8",X"0A",X"AA",X"02",X"A8",X"02",X"A0",X"0A",X"00",X"2A",
		X"02",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A0",X"0A",X"82",X"00",X"02",X"00",X"0A",
		X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"80",
		X"A0",X"00",X"A0",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",X"AA",X"82",X"AA",X"02",X"AA",X"02",X"A8",X"02",
		X"FF",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"AA",X"00",X"A8",X"AA",X"80",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"8A",X"AA",X"8A",X"AA",
		X"88",X"20",X"8A",X"28",X"8A",X"28",X"8A",X"28",X"2A",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",
		X"80",X"8A",X"8A",X"8A",X"A2",X"8A",X"A8",X"8A",X"80",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"8A",X"AA",X"02",
		X"AA",X"28",X"AA",X"28",X"AA",X"28",X"AA",X"28",X"A8",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"0A",X"AA",X"2A",X"AA",X"2A",
		X"0A",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"A8",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"28",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"28",X"A2",X"A8",X"AA",
		X"28",X"00",X"28",X"88",X"28",X"88",X"28",X"88",X"08",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"A0",X"A8",X"8A",X"28",X"80",X"28",X"8A",X"AA",X"A0",X"28",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"AB",X"55",X"AB",X"55",X"AD",X"55",X"AD",X"55",X"B5",X"55",X"B5",X"55",X"D5",X"55",X"D5",X"55",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AD",X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",X"AA",X"D5",X"AA",X"D5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"A8",X"A8",X"A0",X"A0",X"02",X"A0",X"0A",X"80",
		X"0A",X"A0",X"0A",X"80",X"0A",X"00",X"0A",X"00",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",
		X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"02",X"A0",X"02",X"80",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"02",X"A0",X"00",X"80",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"02",X"A0",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"02",X"A0",X"02",X"A8",X"02",X"A8",X"02",X"A8",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"28",
		X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"A8",X"02",X"A8",X"02",X"A0",X"02",X"A0",X"00",X"A0",
		X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"20",X"80",X"28",X"80",X"28",X"00",X"0A",X"00",X"02",
		X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"A8",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"02",X"A0",X"02",X"A0",X"0A",X"A0",X"0A",X"A0",X"2A",X"A0",X"2A",X"A0",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"0A",X"80",X"2A",X"80",X"2A",X"00",X"2A",X"00",X"2A",
		X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"0A",X"80",X"0A",X"80",X"00",X"80",X"00",X"80",X"00",
		X"0A",X"A8",X"02",X"A8",X"00",X"AA",X"80",X"2A",X"80",X"0A",X"A0",X"02",X"A0",X"02",X"A8",X"00",
		X"AA",X"00",X"AA",X"00",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",
		X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",
		X"80",X"02",X"80",X"0A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",
		X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"0A",X"00",X"02",X"00",X"02",
		X"80",X"AA",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"A0",X"2A",X"A0",X"0A",
		X"A0",X"0A",X"A0",X"0A",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"80",X"00",X"80",X"00",
		X"A8",X"02",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"00",X"2A",X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",
		X"80",X"2A",X"80",X"2A",X"80",X"0A",X"80",X"0A",X"A0",X"0A",X"A0",X"02",X"A0",X"02",X"A8",X"02",
		X"80",X"0A",X"80",X"0A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"80",X"2A",X"80",X"AA",
		X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A8",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"0A",
		X"AA",X"00",X"A8",X"00",X"A0",X"08",X"A0",X"2A",X"80",X"2A",X"80",X"AA",X"00",X"AA",X"00",X"AA",
		X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"2A",X"80",X"2A",X"80",X"0A",X"80",X"0A",
		X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"A0",X"0A",X"A0",X"02",X"A0",X"02",X"A0",X"02",
		X"80",X"02",X"80",X"0A",X"80",X"0A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"AA",
		X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"80",X"00",X"80",X"00",X"A0",X"00",X"A8",X"00",
		X"80",X"0A",X"A0",X"02",X"A0",X"02",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",
		X"00",X"02",X"00",X"02",X"A0",X"02",X"A8",X"02",X"A8",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"80",
		X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",
		X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",
		X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"28",X"00",X"28",X"00",X"A8",X"00",X"A8",X"00",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"28",X"00",X"20",X"00",X"A0",X"00",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"02",X"00",X"02",X"20",X"02",X"A8",X"02",X"AA",X"00",X"AA",X"80",X"AA",X"A0",
		X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"28",X"0A",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",
		X"A8",X"00",X"A8",X"00",X"28",X"00",X"28",X"02",X"28",X"02",X"28",X"02",X"28",X"0A",X"08",X"0A",
		X"08",X"2A",X"20",X"2A",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"28",X"80",X"28",X"80",X"2A",X"80",X"2A",X"80",X"2A",
		X"02",X"00",X"02",X"00",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"82",X"80",
		X"80",X"80",X"80",X"80",X"A0",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"80",X"2A",X"00",X"0A",X"00",X"02",X"00",X"02",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"2A",X"00",X"2A",X"00",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"02",X"A0",X"02",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
