library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity egs0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of egs0 is
	type rom is array(0 to  1023) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"00",X"32",X"2B",X"22",X"C3",X"00",X"08",X"3E",X"01",X"32",X"2A",X"22",X"C3",X"15",X"00",
		X"3E",X"02",X"32",X"2A",X"22",X"F3",X"F1",X"CD",X"10",X"1A",X"C9",X"3E",X"01",X"32",X"2B",X"22",
		X"C3",X"38",X"00",X"3E",X"02",X"C3",X"1D",X"00",X"3A",X"2B",X"22",X"FE",X"00",X"CA",X"3C",X"00",
		X"47",X"3A",X"2A",X"22",X"B8",X"CA",X"3C",X"00",X"FB",X"C3",X"38",X"00",X"3E",X"00",X"32",X"2B",
		X"22",X"C9",X"78",X"F5",X"1A",X"77",X"13",X"23",X"05",X"CA",X"4F",X"00",X"C3",X"44",X"00",X"F1",
		X"F5",X"47",X"D5",X"3E",X"20",X"90",X"5F",X"97",X"57",X"19",X"D1",X"0D",X"CA",X"63",X"00",X"F1",
		X"C3",X"42",X"00",X"F1",X"C9",X"06",X"40",X"21",X"00",X"23",X"97",X"77",X"BE",X"C2",X"6B",X"00",
		X"23",X"7C",X"B8",X"C2",X"6A",X"00",X"C9",X"1A",X"47",X"13",X"1A",X"4F",X"13",X"C9",X"21",X"02",
		X"24",X"22",X"10",X"20",X"CD",X"60",X"01",X"21",X"04",X"24",X"22",X"12",X"20",X"CD",X"60",X"01",
		X"21",X"06",X"24",X"22",X"14",X"20",X"CD",X"60",X"01",X"21",X"18",X"28",X"22",X"16",X"20",X"11",
		X"10",X"1C",X"CD",X"63",X"01",X"21",X"1A",X"28",X"22",X"18",X"20",X"11",X"10",X"1C",X"CD",X"63",
		X"01",X"21",X"1C",X"28",X"22",X"1A",X"20",X"11",X"10",X"1C",X"CD",X"63",X"01",X"21",X"C2",X"25",
		X"22",X"1C",X"20",X"CD",X"6A",X"01",X"21",X"C4",X"25",X"22",X"1E",X"20",X"CD",X"6A",X"01",X"21",
		X"C6",X"25",X"22",X"20",X"20",X"CD",X"6A",X"01",X"21",X"D8",X"29",X"22",X"22",X"20",X"11",X"4C",
		X"1C",X"CD",X"63",X"01",X"21",X"DA",X"29",X"22",X"24",X"20",X"11",X"4C",X"1C",X"CD",X"63",X"01",
		X"21",X"DC",X"29",X"22",X"26",X"20",X"11",X"4C",X"1C",X"CD",X"63",X"01",X"21",X"82",X"27",X"22",
		X"28",X"20",X"CD",X"74",X"01",X"21",X"84",X"27",X"22",X"2A",X"20",X"CD",X"74",X"01",X"21",X"86",
		X"27",X"22",X"2C",X"20",X"CD",X"74",X"01",X"21",X"98",X"2B",X"22",X"2E",X"20",X"11",X"2E",X"1C",
		X"CD",X"63",X"01",X"21",X"9A",X"2B",X"22",X"30",X"20",X"11",X"2E",X"1C",X"CD",X"63",X"01",X"21",
		X"9C",X"2B",X"22",X"32",X"20",X"11",X"2E",X"1C",X"CD",X"63",X"01",X"21",X"D6",X"25",X"CD",X"7E",
		X"01",X"21",X"C3",X"29",X"CD",X"7E",X"01",X"21",X"D7",X"2D",X"CD",X"7E",X"01",X"21",X"C2",X"31",
		X"CD",X"7E",X"01",X"21",X"D8",X"35",X"CD",X"7E",X"01",X"21",X"C2",X"39",X"CD",X"7E",X"01",X"C9",
		X"11",X"6A",X"1C",X"CD",X"77",X"00",X"CD",X"42",X"00",X"C9",X"11",X"A6",X"1C",X"CD",X"77",X"00",
		X"CD",X"42",X"00",X"C9",X"11",X"88",X"1C",X"CD",X"77",X"00",X"CD",X"42",X"00",X"C9",X"11",X"C4",
		X"1C",X"CD",X"77",X"00",X"CD",X"42",X"00",X"C9",X"1A",X"00",X"00",X"00",X"00",X"B6",X"77",X"23",
		X"13",X"1A",X"00",X"00",X"00",X"00",X"B6",X"77",X"23",X"13",X"1A",X"00",X"00",X"00",X"00",X"B6",
		X"77",X"23",X"13",X"1A",X"00",X"00",X"00",X"00",X"B6",X"77",X"23",X"13",X"AF",X"00",X"00",X"00",
		X"00",X"B6",X"77",X"C9",X"1A",X"00",X"00",X"00",X"00",X"2F",X"A6",X"77",X"23",X"13",X"1A",X"00",
		X"00",X"00",X"00",X"2F",X"A6",X"77",X"23",X"13",X"1A",X"00",X"00",X"00",X"00",X"2F",X"A6",X"77",
		X"23",X"13",X"1A",X"00",X"00",X"00",X"00",X"2F",X"A6",X"77",X"23",X"13",X"AF",X"00",X"00",X"00",
		X"00",X"2F",X"A6",X"77",X"C9",X"21",X"4E",X"3D",X"11",X"1A",X"1D",X"CD",X"63",X"01",X"21",X"02",
		X"3C",X"11",X"8A",X"1D",X"CD",X"63",X"01",X"21",X"04",X"3C",X"11",X"6C",X"1D",X"CD",X"63",X"01",
		X"21",X"19",X"3C",X"11",X"6C",X"1D",X"CD",X"63",X"01",X"C9",X"21",X"2C",X"25",X"11",X"9A",X"1D",
		X"CD",X"63",X"01",X"21",X"8C",X"26",X"11",X"CD",X"1D",X"CD",X"63",X"01",X"C9",X"2A",X"0A",X"20",
		X"EB",X"CD",X"77",X"00",X"3A",X"08",X"20",X"D3",X"05",X"2A",X"06",X"20",X"CD",X"88",X"01",X"CD",
		X"72",X"02",X"C2",X"2C",X"02",X"C9",X"2A",X"06",X"20",X"7D",X"E6",X"1F",X"6F",X"3E",X"EB",X"85",
		X"D8",X"3A",X"08",X"20",X"D3",X"05",X"2A",X"0A",X"20",X"EB",X"CD",X"77",X"00",X"2A",X"06",X"20",
		X"CD",X"B4",X"01",X"CD",X"72",X"02",X"C2",X"50",X"02",X"3A",X"08",X"20",X"3C",X"E6",X"07",X"CA",
		X"66",X"02",X"32",X"08",X"20",X"C9",X"AF",X"32",X"08",X"20",X"2A",X"06",X"20",X"23",X"22",X"06",
		X"20",X"C9",X"D5",X"11",X"1C",X"00",X"19",X"D1",X"0D",X"C9",X"2A",X"0A",X"20",X"EB",X"CD",X"77",
		X"00",X"3A",X"08",X"20",X"D3",X"05",X"2A",X"06",X"20",X"CD",X"88",X"01",X"CD",X"72",X"02",X"C2",
		X"89",X"02",X"C9",X"2A",X"06",X"20",X"7D",X"E6",X"1F",X"6F",X"3E",X"F7",X"85",X"D0",X"3A",X"08",
		X"20",X"D3",X"07",X"2A",X"0A",X"20",X"EB",X"CD",X"77",X"00",X"2A",X"06",X"20",X"CD",X"B4",X"01",
		X"CD",X"72",X"02",X"C2",X"AD",X"02",X"3A",X"08",X"20",X"B7",X"CA",X"C2",X"02",X"3D",X"32",X"08",
		X"20",X"C9",X"3E",X"07",X"32",X"08",X"20",X"2A",X"06",X"20",X"2B",X"22",X"06",X"20",X"C9",X"2A",
		X"04",X"20",X"EB",X"CD",X"77",X"00",X"3A",X"02",X"20",X"D3",X"05",X"2A",X"00",X"20",X"CD",X"9A",
		X"01",X"CD",X"41",X"03",X"C2",X"DE",X"02",X"C9",X"2A",X"04",X"20",X"EB",X"CD",X"77",X"00",X"3A",
		X"02",X"20",X"D3",X"05",X"2A",X"00",X"20",X"CD",X"C8",X"01",X"CD",X"41",X"03",X"C2",X"F7",X"02",
		X"3A",X"02",X"20",X"3C",X"E6",X"07",X"CA",X"12",X"03",X"FE",X"04",X"32",X"02",X"20",X"CA",X"2A",
		X"03",X"C9",X"AF",X"32",X"02",X"20",X"2A",X"00",X"20",X"23",X"22",X"00",X"20",X"3A",X"03",X"20",
		X"3C",X"FE",X"17",X"C2",X"27",X"03",X"AF",X"32",X"03",X"20",X"7D",X"E6",X"1F",X"6F",X"3E",X"F8",
		X"85",X"D0",X"3E",X"E8",X"85",X"D8",X"11",X"20",X"00",X"2A",X"00",X"20",X"19",X"22",X"00",X"20",
		X"C9",X"D5",X"11",X"1E",X"00",X"19",X"D1",X"0D",X"C9",X"2A",X"04",X"20",X"EB",X"CD",X"77",X"00",
		X"3A",X"02",X"20",X"D3",X"05",X"2A",X"00",X"20",X"CD",X"9A",X"01",X"CD",X"41",X"03",X"C2",X"58",
		X"03",X"C9",X"2A",X"04",X"20",X"EB",X"CD",X"77",X"00",X"3A",X"02",X"20",X"D3",X"05",X"2A",X"00",
		X"20",X"CD",X"C8",X"01",X"CD",X"41",X"03",X"C2",X"71",X"03",X"3A",X"02",X"20",X"B7",X"CA",X"8B",
		X"03",X"3D",X"32",X"02",X"20",X"FE",X"04",X"CA",X"A4",X"03",X"C9",X"3E",X"07",X"32",X"02",X"20",
		X"2A",X"00",X"20",X"2B",X"22",X"00",X"20",X"3A",X"03",X"20",X"3C",X"FE",X"18",X"C2",X"A1",X"03",
		X"AF",X"32",X"03",X"20",X"7D",X"E6",X"1F",X"6F",X"3E",X"F8",X"85",X"D0",X"3E",X"E8",X"85",X"D8",
		X"11",X"20",X"00",X"2A",X"00",X"20",X"19",X"22",X"00",X"20",X"C9",X"3E",X"01",X"32",X"34",X"20",
		X"0E",X"05",X"3E",X"07",X"47",X"32",X"35",X"20",X"11",X"36",X"20",X"21",X"48",X"3D",X"7E",X"B7",
		X"C2",X"D7",X"03",X"23",X"C3",X"40",X"0C",X"22",X"3D",X"20",X"7E",X"12",X"C5",X"01",X"20",X"00",
		X"09",X"C1",X"13",X"05",X"0D",X"C2",X"DA",X"03",X"AF",X"12",X"05",X"C8",X"13",X"C3",X"E8",X"03",
		X"11",X"36",X"20",X"2A",X"3D",X"20",X"0E",X"05",X"CD",X"26",X"04",X"CD",X"1F",X"04",X"0D",X"C2");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
