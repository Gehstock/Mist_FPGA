`define BUILD_DATE "190307"
`define BUILD_TIME "160242"
