library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"02",X"32",X"22",X"4E",X"C9",X"06",X"01",X"0E",X"0A",X"CD",X"A4",X"80",X"3A",X"E3",X"4D",
		X"A7",X"C0",X"0E",X"02",X"16",X"00",X"1E",X"00",X"CD",X"CA",X"80",X"C9",X"06",X"06",X"0E",X"0A",
		X"CD",X"A4",X"80",X"3A",X"E3",X"4D",X"A7",X"C0",X"0E",X"02",X"16",X"00",X"1E",X"00",X"CD",X"CA",
		X"80",X"C9",X"06",X"00",X"18",X"12",X"06",X"02",X"18",X"0E",X"06",X"03",X"18",X"0A",X"06",X"04",
		X"18",X"06",X"06",X"05",X"18",X"02",X"06",X"07",X"0E",X"0A",X"CD",X"A4",X"80",X"3A",X"E3",X"4D",
		X"A7",X"C0",X"21",X"22",X"4E",X"34",X"C9",X"06",X"00",X"0E",X"01",X"CD",X"A4",X"80",X"3A",X"E3",
		X"4D",X"A7",X"C0",X"0E",X"02",X"16",X"01",X"1E",X"00",X"CD",X"CA",X"80",X"C9",X"06",X"05",X"0E",
		X"01",X"CD",X"A4",X"80",X"3A",X"E3",X"4D",X"A7",X"C0",X"0E",X"01",X"16",X"01",X"1E",X"00",X"CD",
		X"CA",X"80",X"C9",X"06",X"01",X"18",X"0E",X"06",X"02",X"18",X"0A",X"06",X"03",X"18",X"06",X"06",
		X"04",X"18",X"02",X"06",X"06",X"0E",X"01",X"CD",X"A4",X"80",X"3A",X"E3",X"4D",X"A7",X"C0",X"21",
		X"22",X"4E",X"34",X"C9",X"21",X"E3",X"4D",X"AF",X"86",X"20",X"04",X"71",X"79",X"23",X"70",X"E7",
		X"44",X"B0",X"DF",X"80",X"37",X"81",X"4E",X"81",X"62",X"81",X"76",X"81",X"A6",X"81",X"B2",X"81",
		X"44",X"B0",X"44",X"B0",X"DC",X"81",X"0C",X"82",X"23",X"82",X"3A",X"13",X"4E",X"A7",X"47",X"79",
		X"28",X"06",X"7A",X"CB",X"08",X"38",X"01",X"7B",X"21",X"22",X"4E",X"86",X"3C",X"77",X"C9",X"21",
		X"E4",X"4D",X"7E",X"87",X"86",X"87",X"21",X"26",X"0A",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"11",
		X"E5",X"4D",X"01",X"06",X"00",X"ED",X"B0",X"AF",X"12",X"1E",X"F0",X"16",X"00",X"CD",X"31",X"82",
		X"16",X"03",X"1E",X"01",X"21",X"0A",X"4C",X"3A",X"EA",X"4D",X"4F",X"82",X"77",X"23",X"3A",X"E9",
		X"4D",X"47",X"77",X"23",X"79",X"83",X"77",X"23",X"70",X"CD",X"20",X"81",X"CD",X"32",X"81",X"C9",
		X"CD",X"B8",X"90",X"C8",X"21",X"0A",X"4C",X"3E",X"C0",X"47",X"AE",X"77",X"23",X"23",X"78",X"AE",
		X"77",X"C9",X"21",X"E3",X"4D",X"34",X"C9",X"11",X"70",X"0A",X"06",X"01",X"CD",X"45",X"82",X"C0",
		X"1E",X"F4",X"16",X"00",X"CD",X"31",X"82",X"16",X"05",X"1E",X"04",X"C3",X"04",X"81",X"11",X"70",
		X"0A",X"06",X"02",X"CD",X"45",X"82",X"C0",X"1E",X"F8",X"16",X"08",X"CD",X"31",X"82",X"CD",X"32",
		X"81",X"C9",X"11",X"70",X"0A",X"06",X"03",X"CD",X"45",X"82",X"C0",X"1E",X"FC",X"16",X"0C",X"CD",
		X"31",X"82",X"CD",X"32",X"81",X"C9",X"11",X"70",X"0A",X"06",X"04",X"CD",X"45",X"82",X"C0",X"3E",
		X"04",X"32",X"EC",X"4E",X"AF",X"32",X"BC",X"4E",X"1E",X"00",X"16",X"10",X"CD",X"31",X"82",X"16",
		X"07",X"1E",X"06",X"CD",X"04",X"81",X"2A",X"E7",X"4D",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",
		X"23",X"EB",X"CD",X"C3",X"81",X"C9",X"11",X"70",X"0A",X"06",X"05",X"CD",X"45",X"82",X"C0",X"C3",
		X"F9",X"80",X"11",X"70",X"0A",X"06",X"06",X"CD",X"45",X"82",X"C0",X"CD",X"55",X"82",X"AF",X"32",
		X"E3",X"4D",X"C9",X"D5",X"DD",X"E1",X"11",X"20",X"00",X"7B",X"91",X"5F",X"C5",X"DD",X"7E",X"00",
		X"77",X"23",X"DD",X"23",X"0D",X"20",X"F6",X"C1",X"19",X"10",X"F1",X"C9",X"21",X"E4",X"4D",X"7E",
		X"87",X"87",X"21",X"50",X"0A",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"5E",X"23",X"56",X"ED",X"53",
		X"E5",X"4D",X"23",X"5E",X"23",X"56",X"ED",X"53",X"E9",X"4D",X"AF",X"32",X"EB",X"4D",X"1E",X"00",
		X"16",X"08",X"CD",X"31",X"82",X"16",X"11",X"1E",X"10",X"C3",X"04",X"81",X"11",X"78",X"0A",X"06",
		X"01",X"CD",X"45",X"82",X"C0",X"3A",X"E4",X"4D",X"47",X"CD",X"F6",X"08",X"CD",X"55",X"82",X"CD",
		X"32",X"81",X"C9",X"11",X"78",X"0A",X"06",X"02",X"CD",X"45",X"82",X"C0",X"AF",X"32",X"E3",X"4D",
		X"C9",X"2A",X"E5",X"4D",X"22",X"08",X"4D",X"3A",X"EA",X"4D",X"A7",X"28",X"03",X"AF",X"92",X"57",
		X"19",X"22",X"0A",X"4D",X"C9",X"21",X"EB",X"4D",X"34",X"4E",X"EB",X"AF",X"86",X"23",X"10",X"FC",
		X"91",X"C8",X"D0",X"AF",X"C9",X"21",X"00",X"00",X"22",X"0A",X"4C",X"22",X"0C",X"4C",X"22",X"08",
		X"4D",X"22",X"0A",X"4D",X"C9",X"21",X"E4",X"F8",X"22",X"08",X"4D",X"2E",X"34",X"26",X"1C",X"22",
		X"0A",X"4C",X"21",X"0C",X"AC",X"22",X"0A",X"4D",X"2E",X"00",X"26",X"1C",X"22",X"0C",X"4C",X"AF",
		X"32",X"EB",X"4D",X"CD",X"DA",X"01",X"CD",X"20",X"81",X"C9",X"3E",X"02",X"32",X"CC",X"4E",X"CD",
		X"DA",X"01",X"C9",X"21",X"EB",X"4D",X"34",X"7E",X"E6",X"07",X"C0",X"DD",X"21",X"08",X"4D",X"FD",
		X"21",X"0A",X"03",X"CD",X"47",X"91",X"22",X"08",X"4D",X"AF",X"11",X"E4",X"DC",X"ED",X"52",X"28",
		X"0B",X"DD",X"21",X"00",X"4C",X"CD",X"63",X"89",X"CD",X"C4",X"82",X"C9",X"CD",X"DA",X"01",X"AF",
		X"32",X"EB",X"4D",X"C9",X"CD",X"B8",X"90",X"C8",X"21",X"0A",X"4C",X"3E",X"C0",X"AE",X"77",X"C9",
		X"CD",X"BD",X"93",X"EF",X"04",X"00",X"CD",X"DA",X"01",X"C9",X"21",X"EB",X"4D",X"34",X"7E",X"FE",
		X"1E",X"28",X"12",X"FE",X"2A",X"D8",X"21",X"0C",X"AC",X"22",X"0A",X"4D",X"3E",X"01",X"32",X"CC",
		X"4E",X"32",X"22",X"4E",X"C9",X"3E",X"01",X"32",X"0C",X"4C",X"21",X"08",X"B4",X"22",X"0A",X"4D",
		X"21",X"AC",X"4E",X"36",X"04",X"CD",X"09",X"83",X"C9",X"CD",X"B8",X"90",X"C8",X"21",X"0C",X"4C",
		X"3E",X"C0",X"AE",X"77",X"C9",X"AF",X"32",X"DE",X"4D",X"21",X"00",X"00",X"22",X"0A",X"4D",X"C9",
		X"EF",X"1C",X"A2",X"C9",X"57",X"21",X"B7",X"4D",X"86",X"C8",X"5F",X"72",X"19",X"14",X"72",X"C9",
		X"21",X"E2",X"4D",X"7E",X"A7",X"C8",X"36",X"00",X"07",X"07",X"07",X"E6",X"07",X"47",X"CD",X"E3",
		X"08",X"C9",X"3A",X"B0",X"4D",X"4F",X"3A",X"DD",X"4D",X"B1",X"C0",X"3A",X"B8",X"4D",X"E7",X"44",
		X"B0",X"5B",X"83",X"6F",X"83",X"7E",X"83",X"44",X"B0",X"44",X"B0",X"21",X"00",X"00",X"22",X"0C",
		X"4D",X"22",X"3C",X"4D",X"22",X"00",X"4D",X"CD",X"71",X"85",X"22",X"EC",X"4D",X"18",X"0A",X"2A",
		X"EC",X"4D",X"2B",X"22",X"EC",X"4D",X"7C",X"B5",X"C0",X"21",X"B8",X"4D",X"34",X"C9",X"0E",X"00",
		X"CD",X"DA",X"84",X"22",X"0C",X"4D",X"22",X"3C",X"4D",X"D9",X"22",X"00",X"4D",X"EB",X"22",X"18",
		X"4D",X"22",X"24",X"4D",X"79",X"32",X"30",X"4D",X"32",X"36",X"4D",X"3E",X"02",X"32",X"03",X"4C",
		X"AF",X"32",X"B8",X"4D",X"32",X"AC",X"4D",X"C9",X"3A",X"B0",X"4D",X"4F",X"3A",X"DD",X"4D",X"B1",
		X"C0",X"3A",X"B9",X"4D",X"E7",X"44",X"B0",X"C1",X"83",X"D5",X"83",X"E4",X"83",X"44",X"B0",X"44",
		X"B0",X"21",X"00",X"00",X"22",X"0E",X"4D",X"22",X"3E",X"4D",X"22",X"02",X"4D",X"CD",X"71",X"85",
		X"22",X"EE",X"4D",X"18",X"0A",X"2A",X"EE",X"4D",X"2B",X"22",X"EE",X"4D",X"7C",X"B5",X"C0",X"21",
		X"B9",X"4D",X"34",X"C9",X"0E",X"01",X"CD",X"DA",X"84",X"22",X"0E",X"4D",X"22",X"3E",X"4D",X"D9",
		X"22",X"02",X"4D",X"EB",X"22",X"1A",X"4D",X"22",X"26",X"4D",X"79",X"32",X"31",X"4D",X"32",X"37",
		X"4D",X"3E",X"04",X"32",X"05",X"4C",X"AF",X"32",X"B9",X"4D",X"32",X"AD",X"4D",X"C9",X"3A",X"B0",
		X"4D",X"4F",X"3A",X"DD",X"4D",X"B1",X"C0",X"3A",X"BA",X"4D",X"E7",X"44",X"B0",X"27",X"84",X"3B",
		X"84",X"4A",X"84",X"44",X"B0",X"44",X"B0",X"21",X"00",X"00",X"22",X"10",X"4D",X"22",X"40",X"4D",
		X"22",X"04",X"4D",X"CD",X"71",X"85",X"22",X"F0",X"4D",X"18",X"0A",X"2A",X"F0",X"4D",X"2B",X"22",
		X"F0",X"4D",X"7C",X"B5",X"C0",X"21",X"BA",X"4D",X"34",X"C9",X"0E",X"02",X"CD",X"DA",X"84",X"22",
		X"10",X"4D",X"22",X"40",X"4D",X"D9",X"22",X"04",X"4D",X"EB",X"22",X"1C",X"4D",X"22",X"28",X"4D",
		X"79",X"32",X"32",X"4D",X"32",X"38",X"4D",X"3E",X"06",X"32",X"07",X"4C",X"AF",X"32",X"BA",X"4D",
		X"32",X"AE",X"4D",X"C9",X"3A",X"B0",X"4D",X"4F",X"3A",X"DD",X"4D",X"B1",X"C0",X"3A",X"BB",X"4D",
		X"E7",X"44",X"B0",X"8D",X"84",X"A1",X"84",X"B0",X"84",X"44",X"B0",X"44",X"B0",X"21",X"00",X"00",
		X"22",X"12",X"4D",X"22",X"42",X"4D",X"22",X"06",X"4D",X"CD",X"71",X"85",X"22",X"F2",X"4D",X"18",
		X"0A",X"2A",X"F2",X"4D",X"2B",X"22",X"F2",X"4D",X"7C",X"B5",X"C0",X"21",X"BB",X"4D",X"34",X"C9",
		X"0E",X"03",X"CD",X"DA",X"84",X"22",X"12",X"4D",X"22",X"42",X"4D",X"D9",X"22",X"06",X"4D",X"EB",
		X"22",X"1E",X"4D",X"22",X"2A",X"4D",X"79",X"32",X"33",X"4D",X"32",X"39",X"4D",X"3E",X"08",X"32",
		X"09",X"4C",X"AF",X"32",X"BB",X"4D",X"32",X"AF",X"4D",X"C9",X"06",X"00",X"3A",X"8B",X"4C",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"07",X"0F",X"CE",X"00",X"4F",X"21",X"16",X"4E",X"09",X"06",X"08",X"3E",
		X"07",X"B9",X"30",X"04",X"21",X"1D",X"4E",X"4F",X"7E",X"A7",X"28",X"04",X"FE",X"05",X"38",X"06",
		X"2B",X"0D",X"10",X"EB",X"0E",X"00",X"3E",X"07",X"B9",X"79",X"20",X"04",X"3A",X"0D",X"4E",X"81",
		X"07",X"07",X"07",X"4F",X"06",X"00",X"21",X"29",X"85",X"09",X"06",X"04",X"5E",X"23",X"56",X"23",
		X"D5",X"10",X"F9",X"C1",X"D1",X"E1",X"D9",X"E1",X"C9",X"24",X"22",X"24",X"24",X"00",X"01",X"02",
		X"02",X"27",X"39",X"3C",X"DC",X"00",X"FF",X"00",X"00",X"2E",X"22",X"74",X"24",X"00",X"01",X"02",
		X"02",X"33",X"39",X"9C",X"DC",X"00",X"FF",X"00",X"00",X"3C",X"22",X"E4",X"24",X"00",X"01",X"02",
		X"02",X"2A",X"22",X"54",X"24",X"00",X"01",X"02",X"02",X"2E",X"39",X"74",X"DC",X"00",X"FF",X"00",
		X"00",X"33",X"22",X"9C",X"24",X"00",X"01",X"02",X"02",X"3C",X"39",X"E4",X"DC",X"00",X"FF",X"00",
		X"00",X"2A",X"8B",X"4C",X"3E",X"03",X"A4",X"FE",X"03",X"20",X"01",X"3D",X"67",X"C9",X"CD",X"8B",
		X"85",X"C0",X"3A",X"DD",X"4D",X"4F",X"3A",X"B0",X"4D",X"B1",X"C9",X"21",X"16",X"4E",X"06",X"07",
		X"7E",X"23",X"B6",X"10",X"FC",X"A7",X"C9",X"3E",X"40",X"32",X"CC",X"4E",X"3E",X"1C",X"CD",X"FF",
		X"B0",X"F7",X"43",X"07",X"00",X"C3",X"BB",X"91",X"3E",X"00",X"CD",X"FF",X"B0",X"F7",X"42",X"07",
		X"00",X"C3",X"BB",X"91",X"3E",X"0C",X"18",X"E6",X"3E",X"02",X"18",X"E2",X"3A",X"CC",X"4E",X"A7",
		X"C0",X"C3",X"BB",X"91",X"AF",X"32",X"06",X"4E",X"3E",X"0C",X"32",X"04",X"4E",X"C9",X"AF",X"32",
		X"CC",X"4E",X"32",X"DC",X"4E",X"32",X"EC",X"4E",X"32",X"9C",X"4E",X"32",X"AC",X"4E",X"32",X"BC",
		X"4E",X"21",X"02",X"4C",X"06",X"08",X"CF",X"32",X"0C",X"4C",X"32",X"0D",X"4C",X"3E",X"06",X"18",
		X"AD",X"3A",X"B0",X"4D",X"A7",X"C8",X"E1",X"3A",X"DD",X"4D",X"E7",X"44",X"B0",X"0F",X"86",X"15",
		X"86",X"1B",X"86",X"21",X"86",X"44",X"B0",X"42",X"86",X"50",X"86",X"44",X"B0",X"48",X"86",X"AF",
		X"32",X"03",X"4C",X"18",X"10",X"AF",X"32",X"05",X"4C",X"18",X"0A",X"AF",X"32",X"07",X"4C",X"18",
		X"04",X"AF",X"32",X"09",X"4C",X"3A",X"DC",X"4D",X"C6",X"18",X"4F",X"06",X"1C",X"CD",X"42",X"00",
		X"3E",X"05",X"32",X"DD",X"4D",X"CD",X"6D",X"86",X"F7",X"42",X"03",X"00",X"3E",X"60",X"CD",X"73",
		X"86",X"C9",X"3A",X"B0",X"4D",X"32",X"B7",X"4D",X"AF",X"32",X"B0",X"4D",X"32",X"DD",X"4D",X"C9",
		X"CD",X"C1",X"90",X"CD",X"30",X"83",X"3E",X"08",X"32",X"DD",X"4D",X"CD",X"6D",X"86",X"F7",X"42",
		X"03",X"00",X"0E",X"60",X"CD",X"73",X"86",X"C9",X"21",X"DD",X"4D",X"34",X"C9",X"3E",X"20",X"32",
		X"AC",X"4E",X"C9",X"3A",X"39",X"4F",X"A7",X"3E",X"03",X"32",X"39",X"4F",X"28",X"1A",X"21",X"91",
		X"4C",X"06",X"10",X"11",X"03",X"00",X"3E",X"0A",X"BE",X"20",X"09",X"2B",X"AF",X"BE",X"28",X"03",
		X"71",X"0E",X"00",X"23",X"19",X"10",X"EF",X"C9",X"F7",X"60",X"0A",X"00",X"C9",X"3A",X"B1",X"4D",
		X"E7",X"C7",X"86",X"D1",X"86",X"D1",X"86",X"D1",X"86",X"D1",X"86",X"EB",X"86",X"19",X"87",X"25",
		X"87",X"2C",X"87",X"33",X"87",X"3A",X"87",X"41",X"87",X"48",X"87",X"7A",X"87",X"84",X"87",X"A0",
		X"87",X"EB",X"86",X"19",X"87",X"CD",X"86",X"3E",X"00",X"32",X"B1",X"4D",X"C9",X"3E",X"07",X"18",
		X"15",X"2A",X"D1",X"4D",X"23",X"22",X"D1",X"4D",X"11",X"78",X"00",X"A7",X"ED",X"52",X"20",X"09",
		X"AF",X"32",X"AC",X"4E",X"3E",X"05",X"32",X"B1",X"4D",X"E1",X"C9",X"21",X"00",X"00",X"22",X"0A",
		X"4D",X"CD",X"72",X"95",X"3E",X"34",X"11",X"B4",X"00",X"4F",X"CD",X"B8",X"90",X"28",X"04",X"3E",
		X"C0",X"A9",X"4F",X"79",X"32",X"0A",X"4C",X"2A",X"D1",X"4D",X"23",X"22",X"D1",X"4D",X"A7",X"ED",
		X"52",X"20",X"D6",X"21",X"B1",X"4D",X"34",X"E1",X"C9",X"21",X"CC",X"4E",X"36",X"04",X"3E",X"35",
		X"11",X"C8",X"00",X"18",X"D4",X"3E",X"37",X"11",X"D3",X"00",X"18",X"CD",X"3E",X"39",X"11",X"E3",
		X"00",X"18",X"C6",X"3E",X"3B",X"11",X"F3",X"00",X"18",X"BF",X"3E",X"3D",X"11",X"03",X"01",X"18",
		X"B8",X"3E",X"75",X"11",X"23",X"01",X"18",X"B1",X"3E",X"F5",X"4F",X"CD",X"B8",X"90",X"28",X"04",
		X"3E",X"C0",X"A9",X"4F",X"79",X"32",X"0A",X"4C",X"2A",X"D1",X"4D",X"23",X"22",X"D1",X"4D",X"11",
		X"63",X"01",X"A7",X"ED",X"52",X"28",X"02",X"E1",X"C9",X"21",X"14",X"4E",X"35",X"21",X"15",X"4E",
		X"35",X"CD",X"69",X"95",X"21",X"04",X"4E",X"34",X"E1",X"C9",X"AF",X"32",X"AC",X"4E",X"CD",X"06",
		X"09",X"C3",X"13",X"87",X"21",X"CC",X"4E",X"36",X"20",X"11",X"A8",X"00",X"2A",X"D1",X"4D",X"23",
		X"22",X"D1",X"4D",X"A7",X"ED",X"52",X"28",X"02",X"E1",X"C9",X"CD",X"06",X"09",X"C3",X"13",X"87",
		X"11",X"48",X"01",X"2A",X"D1",X"4D",X"23",X"22",X"D1",X"4D",X"A7",X"ED",X"52",X"28",X"02",X"E1",
		X"C9",X"21",X"78",X"00",X"22",X"D1",X"4D",X"C3",X"13",X"87",X"3A",X"04",X"4E",X"FE",X"03",X"C8",
		X"E1",X"C9",X"06",X"06",X"1A",X"2F",X"DD",X"86",X"00",X"77",X"23",X"23",X"13",X"13",X"DD",X"23",
		X"10",X"F2",X"C9",X"06",X"06",X"1A",X"DD",X"86",X"00",X"77",X"23",X"23",X"13",X"13",X"DD",X"23",
		X"10",X"F3",X"C9",X"08",X"08",X"08",X"08",X"08",X"08",X"07",X"07",X"08",X"08",X"08",X"08",X"21",
		X"13",X"4C",X"11",X"00",X"4D",X"DD",X"21",X"E3",X"87",X"CD",X"D3",X"87",X"21",X"12",X"4C",X"11",
		X"01",X"4D",X"CD",X"C2",X"87",X"18",X"28",X"09",X"09",X"09",X"09",X"09",X"09",X"06",X"06",X"07",
		X"07",X"07",X"07",X"CD",X"B8",X"90",X"4F",X"20",X"D6",X"21",X"13",X"4C",X"11",X"00",X"4D",X"DD",
		X"21",X"07",X"88",X"CD",X"C2",X"87",X"21",X"12",X"4C",X"11",X"01",X"4D",X"CD",X"D3",X"87",X"3A",
		X"22",X"4E",X"FE",X"01",X"28",X"03",X"FE",X"14",X"D8",X"41",X"DD",X"21",X"00",X"4C",X"CD",X"C5",
		X"BD",X"A7",X"C2",X"5A",X"88",X"3A",X"B0",X"4D",X"A7",X"C0",X"21",X"5A",X"88",X"E5",X"3A",X"3A",
		X"4D",X"E7",X"63",X"89",X"7B",X"89",X"76",X"89",X"83",X"89",X"21",X"CC",X"4D",X"56",X"3E",X"20",
		X"82",X"4F",X"3A",X"2D",X"4F",X"A7",X"20",X"05",X"3A",X"36",X"4D",X"87",X"81",X"DD",X"77",X"02",
		X"3A",X"2E",X"4F",X"A7",X"20",X"05",X"3A",X"37",X"4D",X"87",X"81",X"DD",X"77",X"04",X"3A",X"2F",
		X"4F",X"A7",X"20",X"05",X"3A",X"38",X"4D",X"87",X"81",X"DD",X"77",X"06",X"3A",X"30",X"4F",X"A7",
		X"20",X"05",X"3A",X"39",X"4D",X"87",X"81",X"DD",X"77",X"08",X"3A",X"32",X"4F",X"A7",X"20",X"0F",
		X"3A",X"1A",X"4F",X"A7",X"3A",X"1C",X"4F",X"28",X"04",X"C6",X"14",X"18",X"02",X"C6",X"00",X"DD",
		X"77",X"0C",X"78",X"A7",X"C8",X"DD",X"56",X"02",X"3A",X"36",X"4D",X"CD",X"88",X"89",X"DD",X"72",
		X"02",X"DD",X"56",X"04",X"3A",X"37",X"4D",X"CD",X"88",X"89",X"DD",X"72",X"04",X"DD",X"56",X"06",
		X"3A",X"38",X"4D",X"CD",X"88",X"89",X"DD",X"72",X"06",X"DD",X"56",X"08",X"3A",X"39",X"4D",X"CD",
		X"88",X"89",X"DD",X"72",X"08",X"3A",X"1A",X"4F",X"A7",X"28",X"1E",X"DD",X"56",X"0C",X"3A",X"3B",
		X"4D",X"CD",X"88",X"89",X"DD",X"72",X"0C",X"3A",X"B1",X"4D",X"A7",X"C0",X"DD",X"56",X"0A",X"3A",
		X"3A",X"4D",X"CD",X"88",X"89",X"DD",X"72",X"0A",X"C9",X"DD",X"7E",X"0C",X"EE",X"C0",X"DD",X"77",
		X"0C",X"18",X"E4",X"34",X"34",X"35",X"35",X"36",X"36",X"37",X"37",X"38",X"38",X"35",X"35",X"39",
		X"39",X"3A",X"3A",X"B4",X"B4",X"B5",X"B5",X"B6",X"B6",X"B7",X"B7",X"B8",X"B8",X"B5",X"B5",X"B9",
		X"B9",X"BA",X"BA",X"3B",X"3B",X"3B",X"3B",X"3C",X"3C",X"3C",X"3C",X"3D",X"3D",X"3D",X"3D",X"3C",
		X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"3C",X"3F",X"3F",X"3F",X"3F",X"3C",
		X"3C",X"3C",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"21",X"13",X"89",X"3A",X"09",X"4D",X"E6",X"0F",X"D5",X"5F",X"16",X"00",X"19",
		X"7E",X"DD",X"77",X"0A",X"D1",X"C9",X"21",X"23",X"89",X"18",X"EB",X"21",X"33",X"89",X"3A",X"08",
		X"4D",X"18",X"E6",X"21",X"43",X"89",X"18",X"F6",X"5F",X"0E",X"C0",X"7A",X"A1",X"20",X"04",X"7A",
		X"B1",X"57",X"C9",X"7B",X"FE",X"02",X"20",X"05",X"CB",X"7A",X"C8",X"18",X"06",X"FE",X"03",X"C0",
		X"CB",X"72",X"C8",X"7A",X"A9",X"57",X"C9",X"06",X"05",X"ED",X"5B",X"44",X"4D",X"3A",X"2C",X"4F",
		X"A7",X"20",X"13",X"3A",X"1A",X"4F",X"FE",X"01",X"38",X"0C",X"FE",X"08",X"30",X"08",X"2A",X"46",
		X"4D",X"A7",X"ED",X"52",X"28",X"4B",X"05",X"3A",X"13",X"4E",X"FE",X"02",X"38",X"0E",X"3A",X"BB",
		X"4D",X"A7",X"20",X"08",X"2A",X"42",X"4D",X"A7",X"ED",X"52",X"28",X"35",X"05",X"3A",X"13",X"4E",
		X"FE",X"01",X"38",X"0E",X"3A",X"BA",X"4D",X"A7",X"20",X"08",X"2A",X"40",X"4D",X"A7",X"ED",X"52",
		X"28",X"1F",X"05",X"3A",X"B9",X"4D",X"A7",X"20",X"08",X"2A",X"3E",X"4D",X"A7",X"ED",X"52",X"28",
		X"10",X"05",X"3A",X"B8",X"4D",X"A7",X"20",X"08",X"2A",X"3C",X"4D",X"A7",X"ED",X"52",X"28",X"01",
		X"05",X"78",X"FE",X"05",X"20",X"06",X"3E",X"08",X"32",X"1A",X"4F",X"C9",X"32",X"B0",X"4D",X"32",
		X"DD",X"4D",X"32",X"B1",X"4D",X"A7",X"C8",X"3A",X"33",X"4E",X"A7",X"C8",X"AF",X"32",X"B1",X"4D",
		X"21",X"DC",X"4D",X"7E",X"3C",X"FE",X"0E",X"38",X"02",X"3E",X"0D",X"77",X"C6",X"04",X"47",X"CD",
		X"C5",X"98",X"C9",X"3A",X"B0",X"4D",X"A7",X"C0",X"3A",X"B2",X"4D",X"A7",X"C8",X"01",X"04",X"05",
		X"DD",X"21",X"08",X"4D",X"3A",X"2C",X"4F",X"A7",X"20",X"1D",X"3A",X"1A",X"4F",X"FE",X"01",X"38",
		X"16",X"FE",X"08",X"30",X"12",X"3A",X"0A",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"09",X"3A",X"0B",
		X"4D",X"DD",X"96",X"01",X"B9",X"38",X"9A",X"05",X"3A",X"13",X"4E",X"FE",X"02",X"38",X"19",X"3A",
		X"BB",X"4D",X"A7",X"20",X"13",X"3A",X"06",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"07",
		X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"11",X"8A",X"05",X"3A",X"13",X"4E",X"FE",X"01",X"38",X"19",
		X"3A",X"BA",X"4D",X"A7",X"20",X"13",X"3A",X"04",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",
		X"05",X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"11",X"8A",X"05",X"3A",X"B9",X"4D",X"A7",X"20",X"13",
		X"3A",X"02",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"03",X"4D",X"DD",X"96",X"01",X"B9",
		X"DA",X"11",X"8A",X"05",X"3A",X"B8",X"4D",X"A7",X"20",X"13",X"3A",X"00",X"4D",X"DD",X"96",X"00",
		X"B9",X"30",X"0A",X"3A",X"01",X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"11",X"8A",X"05",X"C3",X"11",
		X"8A",X"3A",X"1A",X"4F",X"FE",X"08",X"D0",X"3A",X"B0",X"4D",X"A7",X"28",X"02",X"E1",X"C9",X"21",
		X"A9",X"4D",X"3E",X"FF",X"BE",X"28",X"02",X"35",X"C9",X"2A",X"54",X"4D",X"29",X"22",X"54",X"4D",
		X"2A",X"52",X"4D",X"ED",X"6A",X"22",X"52",X"4D",X"D0",X"21",X"54",X"4D",X"34",X"3A",X"0E",X"4E",
		X"32",X"AA",X"4D",X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"4F",X"21",X"45",X"4D",X"7E",
		X"06",X"21",X"90",X"38",X"09",X"7E",X"06",X"3B",X"90",X"30",X"03",X"C3",X"82",X"8B",X"3E",X"01",
		X"32",X"CB",X"4D",X"3A",X"00",X"4E",X"FE",X"01",X"CA",X"CA",X"91",X"3A",X"04",X"4E",X"FE",X"10",
		X"D2",X"CA",X"91",X"79",X"A7",X"3A",X"40",X"50",X"20",X"03",X"3A",X"00",X"50",X"CB",X"4F",X"C2",
		X"70",X"8B",X"2A",X"0E",X"03",X"3E",X"02",X"32",X"3A",X"4D",X"22",X"20",X"4D",X"C3",X"31",X"8C",
		X"CB",X"57",X"C2",X"31",X"8C",X"2A",X"0A",X"03",X"AF",X"32",X"3A",X"4D",X"22",X"20",X"4D",X"C3",
		X"31",X"8C",X"3A",X"00",X"4E",X"FE",X"01",X"CA",X"CA",X"91",X"3A",X"04",X"4E",X"FE",X"10",X"D2",
		X"CA",X"91",X"79",X"A7",X"3A",X"40",X"50",X"20",X"03",X"3A",X"00",X"50",X"C3",X"01",X"0C",X"00",
		X"00",X"CB",X"57",X"CA",X"06",X"8D",X"CB",X"47",X"CA",X"0D",X"8D",X"CB",X"5F",X"CA",X"14",X"8D",
		X"2A",X"20",X"4D",X"22",X"2C",X"4D",X"06",X"01",X"DD",X"21",X"2C",X"4D",X"FD",X"21",X"44",X"4D",
		X"CD",X"56",X"91",X"FE",X"E0",X"28",X"5B",X"FE",X"E1",X"28",X"57",X"E6",X"C0",X"D6",X"C0",X"20",
		X"51",X"21",X"EC",X"4E",X"CB",X"86",X"05",X"20",X"1A",X"3A",X"3A",X"4D",X"0F",X"38",X"0A",X"3A",
		X"09",X"4D",X"E6",X"07",X"FE",X"04",X"C8",X"18",X"39",X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"04",
		X"C8",X"18",X"2F",X"DD",X"21",X"20",X"4D",X"CD",X"56",X"91",X"FE",X"E0",X"28",X"33",X"FE",X"E1",
		X"28",X"2F",X"E6",X"C0",X"D6",X"C0",X"20",X"29",X"3A",X"3A",X"4D",X"0F",X"38",X"0A",X"3A",X"09",
		X"4D",X"CD",X"72",X"0C",X"00",X"C8",X"18",X"19",X"3A",X"08",X"4D",X"CD",X"72",X"0C",X"00",X"C8",
		X"18",X"0F",X"2A",X"2C",X"4D",X"22",X"20",X"4D",X"05",X"28",X"06",X"3A",X"34",X"4D",X"32",X"3A",
		X"4D",X"3A",X"BC",X"4E",X"A7",X"20",X"05",X"21",X"EC",X"4E",X"CB",X"C6",X"DD",X"21",X"20",X"4D",
		X"FD",X"21",X"08",X"4D",X"CD",X"47",X"91",X"3A",X"3A",X"4D",X"0F",X"38",X"0F",X"7D",X"E6",X"07",
		X"FE",X"04",X"28",X"15",X"38",X"03",X"2D",X"18",X"10",X"2C",X"18",X"0D",X"7C",X"E6",X"07",X"FE",
		X"04",X"28",X"06",X"38",X"03",X"25",X"18",X"01",X"24",X"22",X"08",X"4D",X"CD",X"5F",X"91",X"22",
		X"44",X"4D",X"DD",X"21",X"CB",X"4D",X"DD",X"7E",X"00",X"DD",X"36",X"00",X"00",X"A7",X"C0",X"21",
		X"CC",X"8C",X"E5",X"2A",X"44",X"4D",X"CD",X"22",X"91",X"7E",X"FE",X"20",X"30",X"48",X"DD",X"21",
		X"0E",X"4E",X"DD",X"34",X"00",X"FE",X"1A",X"28",X"40",X"FE",X"1C",X"30",X"33",X"FE",X"18",X"00",
		X"00",X"00",X"FE",X"10",X"D8",X"3E",X"01",X"32",X"0C",X"4F",X"11",X"00",X"04",X"19",X"7E",X"32",
		X"E2",X"4D",X"21",X"30",X"4E",X"22",X"2E",X"4E",X"2A",X"2C",X"4E",X"CD",X"80",X"0A",X"EF",X"19",
		X"00",X"3E",X"07",X"32",X"B0",X"4D",X"32",X"DD",X"4D",X"3E",X"06",X"C9",X"32",X"A9",X"4D",X"C9",
		X"C6",X"C0",X"77",X"3E",X"01",X"C9",X"3E",X"FF",X"C9",X"36",X"40",X"11",X"0A",X"43",X"ED",X"52",
		X"21",X"1E",X"4E",X"28",X"03",X"21",X"1F",X"4E",X"36",X"00",X"2A",X"C9",X"4D",X"CD",X"26",X"0B",
		X"3E",X"01",X"32",X"33",X"4E",X"AF",X"32",X"DC",X"4D",X"32",X"D4",X"4D",X"3E",X"06",X"C9",X"21",
		X"00",X"01",X"3E",X"02",X"18",X"13",X"21",X"00",X"FF",X"3E",X"00",X"18",X"0C",X"21",X"FF",X"00",
		X"3E",X"03",X"18",X"05",X"21",X"01",X"00",X"3E",X"01",X"32",X"34",X"4D",X"22",X"2C",X"4D",X"06",
		X"00",X"C3",X"B8",X"8B",X"CD",X"E9",X"B4",X"3A",X"B8",X"4D",X"A7",X"C0",X"CD",X"8B",X"91",X"2A",
		X"3C",X"4D",X"01",X"A5",X"4D",X"CD",X"7C",X"91",X"3A",X"A5",X"4D",X"A7",X"28",X"17",X"2A",X"6C",
		X"4D",X"29",X"22",X"6C",X"4D",X"2A",X"6A",X"4D",X"ED",X"6A",X"22",X"6A",X"4D",X"D0",X"21",X"6C",
		X"4D",X"34",X"C3",X"A3",X"8D",X"3A",X"C3",X"4D",X"A7",X"28",X"17",X"2A",X"5C",X"4D",X"29",X"22",
		X"5C",X"4D",X"2A",X"5A",X"4D",X"ED",X"6A",X"22",X"5A",X"4D",X"D0",X"21",X"5C",X"4D",X"34",X"C3",
		X"A3",X"8D",X"3A",X"C2",X"4D",X"A7",X"28",X"17",X"2A",X"60",X"4D",X"29",X"22",X"60",X"4D",X"2A",
		X"5E",X"4D",X"ED",X"6A",X"22",X"5E",X"4D",X"D0",X"21",X"60",X"4D",X"34",X"C3",X"A3",X"8D",X"2A",
		X"64",X"4D",X"29",X"22",X"64",X"4D",X"2A",X"62",X"4D",X"ED",X"6A",X"22",X"62",X"4D",X"D0",X"21",
		X"64",X"4D",X"34",X"21",X"18",X"4D",X"7E",X"A7",X"28",X"0C",X"3A",X"00",X"4D",X"E6",X"07",X"FE",
		X"04",X"28",X"0C",X"C3",X"FC",X"8D",X"3A",X"01",X"4D",X"E6",X"07",X"FE",X"04",X"20",X"3D",X"3E",
		X"01",X"CD",X"28",X"90",X"38",X"19",X"3A",X"33",X"4E",X"A7",X"28",X"05",X"EF",X"0C",X"00",X"18",
		X"0E",X"2A",X"0C",X"4D",X"CD",X"74",X"91",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"08",X"00",X"CD",
		X"50",X"90",X"DD",X"21",X"24",X"4D",X"FD",X"21",X"0C",X"4D",X"CD",X"47",X"91",X"22",X"0C",X"4D",
		X"2A",X"24",X"4D",X"22",X"18",X"4D",X"3A",X"36",X"4D",X"32",X"30",X"4D",X"DD",X"21",X"18",X"4D",
		X"FD",X"21",X"00",X"4D",X"CD",X"47",X"91",X"22",X"00",X"4D",X"CD",X"5F",X"91",X"22",X"3C",X"4D",
		X"C9",X"CD",X"F8",X"B4",X"3A",X"B9",X"4D",X"A7",X"C0",X"2A",X"3E",X"4D",X"01",X"A6",X"4D",X"CD",
		X"7C",X"91",X"3A",X"A6",X"4D",X"A7",X"28",X"17",X"2A",X"78",X"4D",X"29",X"22",X"78",X"4D",X"2A",
		X"76",X"4D",X"ED",X"6A",X"22",X"76",X"4D",X"D0",X"21",X"78",X"4D",X"34",X"C3",X"53",X"8E",X"2A",
		X"70",X"4D",X"29",X"22",X"70",X"4D",X"2A",X"6E",X"4D",X"ED",X"6A",X"22",X"6E",X"4D",X"D0",X"21",
		X"70",X"4D",X"34",X"21",X"1A",X"4D",X"7E",X"A7",X"28",X"0B",X"3A",X"02",X"4D",X"E6",X"07",X"FE",
		X"04",X"28",X"0B",X"18",X"46",X"3A",X"03",X"4D",X"E6",X"07",X"FE",X"04",X"20",X"3D",X"3E",X"02",
		X"CD",X"28",X"90",X"38",X"19",X"3A",X"33",X"4E",X"A7",X"28",X"05",X"EF",X"0D",X"00",X"18",X"0E",
		X"2A",X"0E",X"4D",X"CD",X"74",X"91",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"09",X"00",X"CD",X"6A",
		X"90",X"DD",X"21",X"26",X"4D",X"FD",X"21",X"0E",X"4D",X"CD",X"47",X"91",X"22",X"0E",X"4D",X"2A",
		X"26",X"4D",X"22",X"1A",X"4D",X"3A",X"37",X"4D",X"32",X"31",X"4D",X"DD",X"21",X"1A",X"4D",X"FD",
		X"21",X"02",X"4D",X"CD",X"47",X"91",X"22",X"02",X"4D",X"CD",X"5F",X"91",X"22",X"3E",X"4D",X"C9",
		X"3A",X"13",X"4E",X"FE",X"01",X"D8",X"CD",X"07",X"B5",X"3A",X"BA",X"4D",X"A7",X"C0",X"2A",X"40",
		X"4D",X"01",X"A7",X"4D",X"CD",X"7C",X"91",X"3A",X"A7",X"4D",X"A7",X"28",X"16",X"2A",X"84",X"4D",
		X"29",X"22",X"84",X"4D",X"2A",X"82",X"4D",X"ED",X"6A",X"22",X"82",X"4D",X"D0",X"21",X"84",X"4D",
		X"34",X"18",X"14",X"2A",X"7C",X"4D",X"29",X"22",X"7C",X"4D",X"2A",X"7A",X"4D",X"ED",X"6A",X"22",
		X"7A",X"4D",X"D0",X"21",X"7C",X"4D",X"34",X"21",X"1C",X"4D",X"7E",X"A7",X"28",X"0B",X"3A",X"04",
		X"4D",X"E6",X"07",X"FE",X"04",X"28",X"0B",X"18",X"46",X"3A",X"05",X"4D",X"E6",X"07",X"FE",X"04",
		X"20",X"3D",X"3E",X"03",X"CD",X"28",X"90",X"38",X"19",X"3A",X"33",X"4E",X"A7",X"28",X"05",X"EF",
		X"0E",X"00",X"18",X"0E",X"2A",X"10",X"4D",X"CD",X"74",X"91",X"7E",X"FE",X"1A",X"28",X"03",X"EF",
		X"0A",X"00",X"CD",X"84",X"90",X"DD",X"21",X"28",X"4D",X"FD",X"21",X"10",X"4D",X"CD",X"47",X"91",
		X"22",X"10",X"4D",X"2A",X"28",X"4D",X"22",X"1C",X"4D",X"3A",X"38",X"4D",X"32",X"32",X"4D",X"DD",
		X"21",X"1C",X"4D",X"FD",X"21",X"04",X"4D",X"CD",X"47",X"91",X"22",X"04",X"4D",X"CD",X"5F",X"91",
		X"22",X"40",X"4D",X"C9",X"3A",X"13",X"4E",X"FE",X"02",X"D8",X"CD",X"16",X"B5",X"3A",X"BB",X"4D",
		X"A7",X"C0",X"2A",X"42",X"4D",X"01",X"A8",X"4D",X"CD",X"7C",X"91",X"3A",X"A8",X"4D",X"A7",X"28",
		X"16",X"2A",X"90",X"4D",X"29",X"22",X"90",X"4D",X"2A",X"8E",X"4D",X"ED",X"6A",X"22",X"8E",X"4D",
		X"D0",X"21",X"90",X"4D",X"34",X"18",X"14",X"2A",X"88",X"4D",X"29",X"22",X"88",X"4D",X"2A",X"86",
		X"4D",X"ED",X"6A",X"22",X"86",X"4D",X"D0",X"21",X"88",X"4D",X"34",X"21",X"1E",X"4D",X"7E",X"A7",
		X"28",X"0B",X"3A",X"06",X"4D",X"E6",X"07",X"FE",X"04",X"28",X"0B",X"18",X"46",X"3A",X"07",X"4D",
		X"E6",X"07",X"FE",X"04",X"20",X"3D",X"3E",X"04",X"CD",X"28",X"90",X"38",X"19",X"3A",X"33",X"4E",
		X"A7",X"28",X"05",X"EF",X"0F",X"00",X"18",X"0E",X"2A",X"12",X"4D",X"CD",X"74",X"91",X"7E",X"FE",
		X"1A",X"28",X"03",X"EF",X"0B",X"00",X"CD",X"9E",X"90",X"DD",X"21",X"2A",X"4D",X"FD",X"21",X"12",
		X"4D",X"CD",X"47",X"91",X"22",X"12",X"4D",X"2A",X"2A",X"4D",X"22",X"1E",X"4D",X"3A",X"39",X"4D",
		X"32",X"33",X"4D",X"DD",X"21",X"1E",X"4D",X"FD",X"21",X"06",X"4D",X"CD",X"47",X"91",X"22",X"06",
		X"4D",X"CD",X"5F",X"91",X"22",X"42",X"4D",X"C9",X"87",X"4F",X"06",X"00",X"21",X"0B",X"4D",X"09",
		X"7E",X"FE",X"1D",X"20",X"04",X"36",X"3D",X"18",X"15",X"FE",X"3E",X"20",X"04",X"36",X"1E",X"18",
		X"0D",X"06",X"21",X"90",X"38",X"08",X"7E",X"06",X"3B",X"90",X"30",X"02",X"A7",X"C9",X"37",X"C9",
		X"3A",X"BD",X"4D",X"A7",X"C8",X"AF",X"32",X"BD",X"4D",X"21",X"0A",X"03",X"3A",X"30",X"4D",X"EE",
		X"02",X"32",X"36",X"4D",X"47",X"DF",X"22",X"24",X"4D",X"C9",X"3A",X"BE",X"4D",X"A7",X"C8",X"AF",
		X"32",X"BE",X"4D",X"21",X"0A",X"03",X"3A",X"31",X"4D",X"EE",X"02",X"32",X"37",X"4D",X"47",X"DF",
		X"22",X"26",X"4D",X"C9",X"3A",X"BF",X"4D",X"A7",X"C8",X"AF",X"32",X"BF",X"4D",X"21",X"0A",X"03",
		X"3A",X"32",X"4D",X"EE",X"02",X"32",X"38",X"4D",X"47",X"DF",X"22",X"28",X"4D",X"C9",X"3A",X"C0",
		X"4D",X"A7",X"C8",X"AF",X"32",X"C0",X"4D",X"21",X"0A",X"03",X"3A",X"33",X"4D",X"EE",X"02",X"32",
		X"39",X"4D",X"47",X"DF",X"22",X"2A",X"4D",X"C9",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",
		X"C9",X"CD",X"06",X"91",X"21",X"C1",X"40",X"11",X"31",X"4E",X"01",X"03",X"02",X"1A",X"0F",X"0F",
		X"0F",X"0F",X"CD",X"DD",X"90",X"1A",X"CD",X"DD",X"90",X"1B",X"10",X"F1",X"C9",X"E6",X"0F",X"28",
		X"04",X"0E",X"00",X"18",X"03",X"B9",X"20",X"0A",X"C6",X"30",X"77",X"D5",X"11",X"E0",X"FF",X"19",
		X"D1",X"C9",X"0D",X"36",X"40",X"18",X"F4",X"3E",X"0D",X"0E",X"02",X"06",X"03",X"18",X"10",X"21",
		X"01",X"47",X"3E",X"06",X"18",X"05",X"21",X"61",X"44",X"3E",X"04",X"0E",X"01",X"06",X"04",X"11",
		X"20",X"00",X"F5",X"7B",X"91",X"5F",X"F1",X"C5",X"77",X"23",X"0D",X"20",X"FB",X"C1",X"19",X"10",
		X"F6",X"C9",X"F5",X"C5",X"7D",X"D6",X"20",X"6F",X"7C",X"D6",X"20",X"67",X"06",X"00",X"CB",X"24",
		X"CB",X"24",X"CB",X"24",X"CB",X"24",X"CB",X"10",X"CB",X"24",X"CB",X"10",X"4C",X"26",X"00",X"09",
		X"01",X"40",X"40",X"09",X"C1",X"F1",X"C9",X"FD",X"7E",X"00",X"DD",X"86",X"00",X"6F",X"FD",X"7E",
		X"01",X"DD",X"86",X"01",X"67",X"C9",X"CD",X"47",X"91",X"CD",X"22",X"91",X"7E",X"A7",X"C9",X"7D",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"20",X"6F",X"7C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"C6",X"1E",X"67",X"C9",X"CD",X"22",X"91",X"11",X"00",X"04",X"19",X"C9",X"CD",X"74",X"91",X"7E",
		X"FE",X"1B",X"20",X"04",X"3E",X"01",X"02",X"C9",X"AF",X"02",X"C9",X"3A",X"AF",X"4D",X"A7",X"C8",
		X"21",X"0E",X"4E",X"3A",X"C2",X"4D",X"A7",X"20",X"0E",X"3E",X"F4",X"96",X"47",X"3A",X"C7",X"4D",
		X"90",X"D8",X"3E",X"01",X"32",X"C2",X"4D",X"3A",X"C3",X"4D",X"A7",X"C0",X"3E",X"F4",X"96",X"47",
		X"3A",X"C8",X"4D",X"90",X"D8",X"3E",X"01",X"32",X"C3",X"4D",X"C9",X"21",X"06",X"4E",X"34",X"C9",
		X"21",X"07",X"4E",X"34",X"C9",X"21",X"08",X"4E",X"34",X"C9",X"3A",X"07",X"4E",X"E7",X"E4",X"91",
		X"EF",X"91",X"FD",X"91",X"08",X"92",X"1A",X"92",X"CD",X"C0",X"91",X"C3",X"FF",X"8C",X"CD",X"C0",
		X"91",X"C3",X"0D",X"8D",X"3A",X"45",X"4D",X"FE",X"2D",X"C2",X"06",X"8D",X"C3",X"DE",X"91",X"3A",
		X"44",X"4D",X"FE",X"2E",X"C2",X"0D",X"8D",X"CD",X"C0",X"91",X"C3",X"06",X"8D",X"3A",X"45",X"4D",
		X"FE",X"22",X"C2",X"06",X"8D",X"C3",X"D8",X"91",X"3A",X"45",X"4D",X"FE",X"2D",X"20",X"05",X"CD",
		X"C3",X"B7",X"18",X"CA",X"DA",X"FF",X"8C",X"C3",X"06",X"8D",X"3A",X"44",X"4D",X"FE",X"22",X"28",
		X"B7",X"C3",X"0D",X"8D",X"21",X"00",X"50",X"06",X"08",X"AF",X"77",X"2C",X"10",X"FC",X"21",X"00",
		X"40",X"06",X"04",X"32",X"C0",X"50",X"32",X"07",X"50",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",
		X"10",X"F1",X"06",X"04",X"32",X"C0",X"50",X"AF",X"32",X"07",X"50",X"3E",X"0D",X"77",X"2C",X"20",
		X"FC",X"24",X"10",X"F0",X"ED",X"56",X"AF",X"32",X"07",X"50",X"3C",X"32",X"00",X"50",X"FB",X"76",
		X"32",X"C0",X"50",X"31",X"C0",X"4F",X"AF",X"21",X"00",X"50",X"06",X"08",X"CF",X"21",X"00",X"4C",
		X"06",X"BE",X"CF",X"CF",X"CF",X"CF",X"21",X"40",X"50",X"06",X"40",X"CF",X"32",X"C0",X"50",X"CD",
		X"21",X"93",X"32",X"C0",X"50",X"06",X"00",X"CD",X"01",X"93",X"32",X"C0",X"50",X"21",X"C0",X"4C",
		X"22",X"80",X"4C",X"22",X"82",X"4C",X"3E",X"FF",X"06",X"40",X"CF",X"3E",X"01",X"32",X"00",X"50",
		X"FB",X"2A",X"82",X"4C",X"7E",X"A7",X"FA",X"A1",X"92",X"36",X"FF",X"2C",X"46",X"36",X"FF",X"2C",
		X"20",X"02",X"2E",X"C0",X"22",X"82",X"4C",X"21",X"A1",X"92",X"E5",X"E7",X"01",X"93",X"16",X"94",
		X"2D",X"93",X"6B",X"93",X"88",X"94",X"7F",X"95",X"21",X"93",X"90",X"95",X"20",X"96",X"5C",X"96",
		X"99",X"96",X"E1",X"96",X"35",X"96",X"6B",X"96",X"A8",X"96",X"F0",X"96",X"12",X"03",X"9A",X"95",
		X"0D",X"94",X"B3",X"98",X"D6",X"95",X"44",X"B0",X"FC",X"92",X"2B",X"97",X"7E",X"99",X"C5",X"98",
		X"EC",X"99",X"98",X"9A",X"F2",X"9A",X"27",X"9A",X"69",X"95",X"B8",X"95",X"21",X"04",X"4E",X"34",
		X"C9",X"78",X"E7",X"07",X"93",X"14",X"93",X"3E",X"40",X"01",X"04",X"00",X"21",X"00",X"40",X"CF",
		X"0D",X"20",X"FC",X"C9",X"3E",X"40",X"21",X"40",X"40",X"01",X"04",X"80",X"CF",X"0D",X"20",X"FC",
		X"C9",X"AF",X"01",X"04",X"00",X"21",X"00",X"44",X"CF",X"0D",X"20",X"FC",X"C9",X"CD",X"E5",X"0B",
		X"CD",X"4F",X"93",X"3A",X"00",X"4E",X"3D",X"C8",X"CD",X"D8",X"B0",X"3E",X"9B",X"C3",X"FF",X"B0",
		X"21",X"3F",X"40",X"01",X"D0",X"A0",X"0A",X"FE",X"27",X"C8",X"23",X"77",X"03",X"18",X"F7",X"3A",
		X"13",X"4E",X"A7",X"C8",X"CD",X"64",X"93",X"0F",X"D8",X"21",X"1C",X"1D",X"22",X"EB",X"42",X"7C",
		X"32",X"ED",X"42",X"C9",X"21",X"60",X"61",X"22",X"E5",X"41",X"C9",X"21",X"16",X"4E",X"06",X"08",
		X"AF",X"BE",X"28",X"02",X"36",X"01",X"23",X"10",X"F8",X"CD",X"1C",X"09",X"AF",X"32",X"BC",X"4E",
		X"3E",X"04",X"32",X"EC",X"4E",X"3A",X"1D",X"4E",X"A7",X"28",X"2A",X"3A",X"0D",X"4E",X"A7",X"F5",
		X"CC",X"BD",X"93",X"F1",X"C4",X"C4",X"93",X"CD",X"DF",X"93",X"3A",X"13",X"4E",X"A7",X"C8",X"0F",
		X"38",X"06",X"CD",X"FD",X"93",X"CD",X"E9",X"93",X"CD",X"F8",X"93",X"CD",X"F3",X"93",X"CD",X"EE",
		X"93",X"CD",X"E4",X"93",X"C9",X"CD",X"CB",X"93",X"CD",X"DA",X"93",X"18",X"DA",X"CD",X"CB",X"93",
		X"CD",X"D0",X"93",X"C9",X"CD",X"D5",X"93",X"CD",X"DA",X"93",X"C9",X"21",X"6C",X"09",X"18",X"30",
		X"21",X"76",X"09",X"18",X"2B",X"21",X"80",X"09",X"18",X"26",X"21",X"8A",X"09",X"18",X"21",X"21",
		X"94",X"09",X"18",X"1C",X"21",X"AA",X"09",X"18",X"17",X"21",X"B7",X"09",X"18",X"12",X"21",X"C7",
		X"09",X"18",X"0D",X"21",X"D4",X"09",X"18",X"08",X"21",X"E1",X"09",X"18",X"03",X"21",X"F1",X"09",
		X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"EB",X"CD",X"C3",X"81",X"C9",X"21",X"16",X"4E",
		X"3E",X"01",X"06",X"0A",X"CF",X"C9",X"C5",X"78",X"FE",X"02",X"3E",X"1E",X"28",X"17",X"3A",X"13",
		X"4E",X"FE",X"0F",X"38",X"02",X"3E",X"0F",X"4F",X"06",X"00",X"21",X"78",X"94",X"09",X"7E",X"32",
		X"20",X"4E",X"32",X"21",X"4E",X"21",X"40",X"44",X"01",X"04",X"80",X"CF",X"0D",X"20",X"FC",X"3E",
		X"0D",X"06",X"40",X"21",X"C0",X"47",X"CF",X"C1",X"05",X"C0",X"06",X"00",X"0E",X"0A",X"21",X"23",
		X"07",X"C5",X"DF",X"11",X"00",X"04",X"19",X"78",X"0F",X"0F",X"0F",X"E6",X"E0",X"C6",X"0D",X"06",
		X"03",X"0E",X"02",X"CD",X"0F",X"91",X"C1",X"04",X"0D",X"20",X"E3",X"21",X"5B",X"47",X"3E",X"ED",
		X"06",X"03",X"0E",X"02",X"CD",X"F3",X"0B",X"C9",X"0C",X"9B",X"1D",X"9A",X"18",X"13",X"1D",X"9B",
		X"1D",X"9A",X"18",X"0C",X"0C",X"0C",X"0C",X"0C",X"78",X"FE",X"01",X"20",X"09",X"21",X"02",X"4C",
		X"06",X"0C",X"AF",X"CF",X"18",X"0B",X"21",X"EF",X"94",X"11",X"02",X"4C",X"01",X"0C",X"00",X"ED",
		X"B0",X"21",X"FB",X"94",X"11",X"00",X"4D",X"01",X"48",X"00",X"ED",X"B0",X"CD",X"43",X"95",X"3A",
		X"13",X"4E",X"FE",X"01",X"30",X"19",X"22",X"06",X"4C",X"22",X"04",X"4D",X"22",X"10",X"4D",X"22",
		X"40",X"4D",X"22",X"1C",X"4D",X"22",X"28",X"4D",X"AF",X"32",X"32",X"4D",X"32",X"38",X"4D",X"3A",
		X"13",X"4E",X"FE",X"02",X"D0",X"22",X"08",X"4C",X"22",X"06",X"4D",X"22",X"12",X"4D",X"22",X"42",
		X"4D",X"22",X"1E",X"4D",X"22",X"2A",X"4D",X"AF",X"32",X"33",X"4D",X"32",X"39",X"4D",X"C9",X"20",
		X"02",X"20",X"04",X"20",X"06",X"20",X"08",X"34",X"1C",X"00",X"1C",X"24",X"24",X"3C",X"DC",X"74",
		X"24",X"9C",X"DC",X"E4",X"DC",X"0C",X"AC",X"24",X"22",X"27",X"39",X"2E",X"22",X"33",X"39",X"3C",
		X"38",X"21",X"33",X"00",X"01",X"00",X"FF",X"00",X"01",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"01",X"00",X"FF",X"00",X"01",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"02",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"24",X"22",X"27",X"39",X"2E",X"22",X"33",X"39",X"3C",
		X"38",X"21",X"33",X"3A",X"0D",X"4E",X"A7",X"C8",X"21",X"9C",X"24",X"22",X"08",X"4D",X"21",X"33",
		X"22",X"22",X"14",X"4D",X"22",X"44",X"4D",X"21",X"00",X"01",X"22",X"20",X"4D",X"22",X"2C",X"4D",
		X"3E",X"02",X"32",X"3A",X"4D",X"32",X"34",X"4D",X"C9",X"21",X"00",X"00",X"22",X"0A",X"4D",X"22",
		X"08",X"4D",X"22",X"00",X"4D",X"22",X"02",X"4D",X"22",X"04",X"4D",X"22",X"06",X"4D",X"C9",X"21",
		X"28",X"4E",X"06",X"0C",X"AF",X"CF",X"21",X"00",X"01",X"22",X"29",X"4E",X"CD",X"D0",X"06",X"C9",
		X"3E",X"01",X"32",X"00",X"4E",X"AF",X"32",X"01",X"4E",X"C9",X"AF",X"11",X"00",X"4D",X"21",X"00",
		X"4E",X"12",X"13",X"A7",X"ED",X"52",X"C2",X"9E",X"95",X"21",X"00",X"4F",X"06",X"80",X"AF",X"CF",
		X"21",X"40",X"4C",X"06",X"40",X"AF",X"CF",X"C9",X"DD",X"21",X"56",X"41",X"3A",X"71",X"4E",X"E6",
		X"0F",X"C6",X"30",X"DD",X"77",X"00",X"3A",X"71",X"4E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C8",
		X"C6",X"30",X"DD",X"77",X"20",X"C9",X"3A",X"80",X"50",X"47",X"E6",X"03",X"20",X"05",X"21",X"6E",
		X"4E",X"36",X"FF",X"4F",X"1F",X"CE",X"00",X"32",X"6B",X"4E",X"E6",X"02",X"A9",X"32",X"6D",X"4E",
		X"78",X"0F",X"0F",X"E6",X"03",X"3C",X"FE",X"04",X"20",X"01",X"3C",X"32",X"6F",X"4E",X"78",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"03",X"21",X"1C",X"96",X"D7",X"32",X"71",X"4E",X"21",X"B5",X"05",X"22",
		X"73",X"4E",X"78",X"07",X"07",X"2F",X"E6",X"01",X"32",X"72",X"4E",X"C9",X"05",X"10",X"15",X"FF",
		X"3A",X"CD",X"4D",X"CB",X"47",X"C2",X"48",X"96",X"3A",X"C2",X"4D",X"A7",X"20",X"1A",X"3A",X"04",
		X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0C",X"4D",X"3A",X"36",X"4D",X"11",X"32",X"39",X"CD",X"D4",
		X"97",X"22",X"24",X"4D",X"32",X"36",X"4D",X"C9",X"2A",X"0C",X"4D",X"ED",X"5B",X"44",X"4D",X"3A",
		X"36",X"4D",X"CD",X"D4",X"97",X"22",X"24",X"4D",X"32",X"36",X"4D",X"C9",X"3A",X"CD",X"4D",X"CB",
		X"47",X"C2",X"7E",X"96",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0E",X"4D",X"3A",X"37",
		X"4D",X"11",X"2D",X"22",X"CD",X"D4",X"97",X"22",X"26",X"4D",X"32",X"37",X"4D",X"C9",X"ED",X"5B",
		X"44",X"4D",X"2A",X"2C",X"4D",X"29",X"29",X"19",X"EB",X"2A",X"0E",X"4D",X"3A",X"37",X"4D",X"CD",
		X"D4",X"97",X"22",X"26",X"4D",X"32",X"37",X"4D",X"C9",X"3A",X"CD",X"4D",X"CB",X"47",X"C2",X"BB",
		X"96",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"10",X"4D",X"3A",X"38",X"4D",X"11",X"26",
		X"39",X"CD",X"D4",X"97",X"22",X"28",X"4D",X"32",X"38",X"4D",X"C9",X"ED",X"4B",X"0C",X"4D",X"ED",
		X"5B",X"44",X"4D",X"2A",X"20",X"4D",X"29",X"19",X"7D",X"87",X"91",X"6F",X"7C",X"87",X"90",X"67",
		X"EB",X"2A",X"10",X"4D",X"3A",X"38",X"4D",X"CD",X"D4",X"97",X"22",X"28",X"4D",X"32",X"38",X"4D",
		X"C9",X"3A",X"CD",X"4D",X"CB",X"47",X"C2",X"03",X"97",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",
		X"2A",X"12",X"4D",X"3A",X"39",X"4D",X"11",X"23",X"22",X"CD",X"D4",X"97",X"22",X"2A",X"4D",X"32",
		X"39",X"4D",X"C9",X"DD",X"21",X"44",X"4D",X"FD",X"21",X"12",X"4D",X"CD",X"6C",X"98",X"11",X"40",
		X"00",X"A7",X"ED",X"52",X"DA",X"F0",X"96",X"2A",X"12",X"4D",X"ED",X"5B",X"44",X"4D",X"3A",X"39",
		X"4D",X"CD",X"D4",X"97",X"22",X"2A",X"4D",X"32",X"39",X"4D",X"C9",X"78",X"E7",X"35",X"97",X"52",
		X"97",X"58",X"97",X"70",X"97",X"ED",X"5B",X"44",X"4D",X"3E",X"03",X"32",X"10",X"4F",X"2A",X"16",
		X"4D",X"3A",X"3B",X"4D",X"CD",X"D4",X"97",X"22",X"2E",X"4D",X"32",X"3B",X"4D",X"AF",X"32",X"10",
		X"4F",X"C9",X"ED",X"5B",X"12",X"4F",X"18",X"E1",X"AF",X"32",X"10",X"4F",X"ED",X"5B",X"12",X"4F",
		X"2A",X"14",X"4D",X"3A",X"34",X"4D",X"CD",X"D4",X"97",X"22",X"2C",X"4D",X"32",X"34",X"4D",X"C9",
		X"3A",X"11",X"4F",X"32",X"10",X"4F",X"ED",X"5B",X"12",X"4F",X"2A",X"14",X"4F",X"3A",X"16",X"4F",
		X"CD",X"D4",X"97",X"22",X"17",X"4F",X"32",X"19",X"4F",X"AF",X"32",X"10",X"4F",X"C9",X"22",X"4A",
		X"4D",X"EE",X"02",X"32",X"49",X"4D",X"CD",X"A1",X"98",X"E6",X"03",X"21",X"48",X"4D",X"77",X"87",
		X"5F",X"16",X"00",X"DD",X"21",X"0A",X"03",X"DD",X"19",X"FD",X"21",X"4A",X"4D",X"3A",X"49",X"4D",
		X"BE",X"28",X"13",X"CD",X"56",X"91",X"E6",X"C0",X"D6",X"C0",X"28",X"0A",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"3A",X"48",X"4D",X"C9",X"DD",X"23",X"DD",X"23",X"21",X"48",X"4D",X"7E",X"3C",X"E6",
		X"03",X"77",X"18",X"D9",X"22",X"4A",X"4D",X"ED",X"53",X"4C",X"4D",X"32",X"48",X"4D",X"EE",X"02",
		X"32",X"49",X"4D",X"21",X"FF",X"FF",X"22",X"50",X"4D",X"DD",X"21",X"0A",X"03",X"FD",X"21",X"4A",
		X"4D",X"AF",X"32",X"E1",X"4D",X"21",X"D3",X"4D",X"36",X"00",X"3A",X"49",X"4D",X"BE",X"28",X"40",
		X"CD",X"47",X"91",X"22",X"4E",X"4D",X"3A",X"10",X"4F",X"A7",X"20",X"0A",X"CD",X"22",X"91",X"7E",
		X"E6",X"C0",X"D6",X"C0",X"28",X"2A",X"21",X"E1",X"4D",X"34",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",
		X"4C",X"4D",X"FD",X"21",X"4E",X"4D",X"CD",X"6C",X"98",X"FD",X"E1",X"DD",X"E1",X"EB",X"2A",X"50",
		X"4D",X"A7",X"ED",X"52",X"38",X"0A",X"ED",X"53",X"50",X"4D",X"3A",X"D3",X"4D",X"32",X"48",X"4D",
		X"DD",X"23",X"DD",X"23",X"21",X"D3",X"4D",X"34",X"3E",X"04",X"BE",X"20",X"AD",X"3A",X"E1",X"4D",
		X"A7",X"3A",X"49",X"4D",X"28",X"03",X"3A",X"48",X"4D",X"87",X"5F",X"16",X"00",X"DD",X"21",X"0A",
		X"03",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CB",X"3F",X"C9",X"DD",X"7E",X"00",X"FD",
		X"46",X"00",X"90",X"30",X"05",X"78",X"DD",X"46",X"00",X"90",X"CD",X"92",X"98",X"E5",X"DD",X"7E",
		X"01",X"FD",X"46",X"01",X"90",X"30",X"05",X"78",X"DD",X"46",X"01",X"90",X"CD",X"92",X"98",X"C1",
		X"09",X"C9",X"67",X"5F",X"2E",X"00",X"55",X"0E",X"08",X"29",X"30",X"01",X"19",X"0D",X"20",X"F9",
		X"C9",X"2A",X"D5",X"4D",X"54",X"5D",X"29",X"29",X"19",X"23",X"7C",X"E6",X"1F",X"67",X"7E",X"22",
		X"D5",X"4D",X"C9",X"06",X"0A",X"C5",X"05",X"21",X"23",X"07",X"DF",X"11",X"F9",X"06",X"CD",X"3D",
		X"09",X"C1",X"10",X"F1",X"C9",X"3A",X"00",X"4E",X"FE",X"01",X"C8",X"78",X"A7",X"21",X"5E",X"99",
		X"20",X"03",X"2A",X"2E",X"4E",X"DF",X"EB",X"CD",X"A9",X"99",X"7B",X"86",X"27",X"77",X"23",X"7A",
		X"8E",X"27",X"77",X"5F",X"23",X"3E",X"00",X"8E",X"27",X"77",X"57",X"EB",X"29",X"29",X"29",X"29",
		X"3A",X"71",X"4E",X"3D",X"BC",X"DC",X"B5",X"99",X"CD",X"21",X"99",X"13",X"13",X"13",X"21",X"8A",
		X"4E",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"CD",X"A9",X"99",
		X"11",X"88",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"1B",X"01",X"04",X"03",X"21",X"F2",X"43",X"18",
		X"0F",X"3A",X"09",X"4E",X"01",X"04",X"03",X"21",X"FC",X"43",X"A7",X"28",X"03",X"21",X"E9",X"43",
		X"1A",X"0F",X"0F",X"0F",X"0F",X"CD",X"40",X"99",X"1A",X"CD",X"40",X"99",X"1B",X"10",X"F1",X"C9",
		X"E6",X"0F",X"28",X"07",X"0E",X"00",X"CD",X"55",X"99",X"18",X"07",X"79",X"A7",X"28",X"F7",X"3E",
		X"40",X"0D",X"77",X"2B",X"C9",X"E6",X"0F",X"C6",X"90",X"27",X"CE",X"40",X"27",X"C9",X"10",X"00",
		X"50",X"00",X"30",X"00",X"50",X"00",X"70",X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"05",
		X"00",X"07",X"00",X"10",X"00",X"20",X"00",X"30",X"00",X"50",X"00",X"70",X"00",X"90",X"06",X"00",
		X"CD",X"F2",X"9A",X"AF",X"21",X"80",X"4E",X"06",X"08",X"CF",X"01",X"04",X"03",X"11",X"82",X"4E",
		X"21",X"FC",X"43",X"CD",X"30",X"99",X"01",X"04",X"03",X"11",X"86",X"4E",X"21",X"E9",X"43",X"3A",
		X"70",X"4E",X"A7",X"20",X"8B",X"0E",X"06",X"18",X"87",X"3A",X"09",X"4E",X"21",X"80",X"4E",X"A7",
		X"C8",X"21",X"84",X"4E",X"C9",X"13",X"6B",X"62",X"1B",X"CB",X"46",X"C0",X"CB",X"C6",X"21",X"EC",
		X"4E",X"36",X"02",X"21",X"14",X"4E",X"34",X"21",X"15",X"4E",X"34",X"46",X"21",X"1C",X"40",X"0E",
		X"05",X"78",X"A7",X"28",X"0E",X"FE",X"06",X"30",X"0A",X"3E",X"7C",X"CD",X"11",X"9A",X"2B",X"2B",
		X"0D",X"10",X"F6",X"0D",X"F8",X"CD",X"00",X"9A",X"2B",X"2B",X"18",X"F7",X"3A",X"00",X"4E",X"FE",
		X"01",X"C8",X"CD",X"53",X"9A",X"14",X"44",X"1C",X"05",X"02",X"21",X"15",X"4E",X"46",X"18",X"CC",
		X"3E",X"40",X"E5",X"D5",X"77",X"23",X"77",X"11",X"1F",X"00",X"19",X"77",X"23",X"77",X"D1",X"E1",
		X"C9",X"E5",X"CD",X"17",X"9A",X"E1",X"C9",X"D5",X"11",X"1F",X"00",X"77",X"3C",X"23",X"77",X"3C",
		X"19",X"77",X"3C",X"23",X"77",X"D1",X"C9",X"3A",X"6E",X"4E",X"FE",X"FF",X"20",X"05",X"06",X"02",
		X"C3",X"F2",X"9A",X"06",X"01",X"CD",X"F2",X"9A",X"3A",X"6E",X"4E",X"E6",X"F0",X"28",X"09",X"0F",
		X"0F",X"0F",X"0F",X"C6",X"30",X"32",X"36",X"40",X"3A",X"6E",X"4E",X"E6",X"0F",X"C6",X"30",X"32",
		X"35",X"40",X"C9",X"E1",X"5E",X"23",X"56",X"23",X"4E",X"23",X"7E",X"87",X"47",X"23",X"7E",X"23",
		X"E5",X"EB",X"11",X"16",X"00",X"C5",X"71",X"23",X"10",X"FC",X"C1",X"19",X"3D",X"20",X"F6",X"C9",
		X"80",X"13",X"80",X"9B",X"80",X"1D",X"80",X"9A",X"80",X"18",X"80",X"0C",X"80",X"13",X"80",X"9B",
		X"80",X"1D",X"80",X"9A",X"80",X"0C",X"80",X"0C",X"80",X"0C",X"80",X"0C",X"80",X"0C",X"80",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"00",X"4E",X"FE",X"01",X"C8",X"3A",X"13",
		X"4E",X"3C",X"FE",X"06",X"D2",X"DC",X"9A",X"11",X"70",X"9A",X"47",X"0E",X"05",X"21",X"02",X"40",
		X"1A",X"CD",X"11",X"9A",X"3E",X"04",X"84",X"67",X"13",X"1A",X"CD",X"02",X"9A",X"3E",X"FC",X"84",
		X"67",X"13",X"23",X"23",X"0D",X"10",X"E9",X"0D",X"F8",X"CD",X"00",X"9A",X"3E",X"04",X"84",X"67",
		X"AF",X"CD",X"02",X"9A",X"3E",X"FC",X"84",X"67",X"23",X"23",X"18",X"EB",X"FE",X"0F",X"38",X"02",
		X"3E",X"0F",X"D6",X"05",X"4F",X"06",X"00",X"21",X"70",X"9A",X"09",X"09",X"EB",X"06",X"05",X"C3",
		X"AB",X"9A",X"21",X"72",X"A0",X"DF",X"5E",X"23",X"3E",X"7F",X"A6",X"57",X"DD",X"21",X"00",X"44",
		X"DD",X"19",X"DD",X"E5",X"11",X"00",X"FC",X"DD",X"19",X"11",X"FF",X"FF",X"CB",X"7E",X"20",X"03",
		X"11",X"E0",X"FF",X"23",X"78",X"01",X"00",X"00",X"87",X"38",X"28",X"7E",X"FE",X"27",X"28",X"09",
		X"DD",X"77",X"00",X"23",X"DD",X"19",X"04",X"18",X"F2",X"23",X"DD",X"E1",X"7E",X"A7",X"FA",X"3B",
		X"9B",X"7E",X"DD",X"77",X"00",X"23",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"77",X"00",X"DD",X"19",
		X"10",X"F9",X"C9",X"7E",X"FE",X"27",X"28",X"0A",X"DD",X"36",X"00",X"40",X"23",X"DD",X"19",X"04",
		X"18",X"F1",X"23",X"04",X"ED",X"B1",X"18",X"D2",X"21",X"55",X"9C",X"DD",X"21",X"CC",X"4E",X"FD",
		X"21",X"8C",X"4E",X"CD",X"DB",X"9B",X"47",X"3A",X"CC",X"4E",X"A7",X"28",X"04",X"78",X"32",X"91",
		X"4E",X"21",X"65",X"9C",X"DD",X"21",X"DC",X"4E",X"FD",X"21",X"92",X"4E",X"CD",X"DB",X"9B",X"47",
		X"3A",X"DC",X"4E",X"A7",X"28",X"04",X"78",X"32",X"96",X"4E",X"21",X"75",X"9C",X"DD",X"21",X"EC",
		X"4E",X"FD",X"21",X"97",X"4E",X"CD",X"DB",X"9B",X"47",X"3A",X"EC",X"4E",X"A7",X"C8",X"78",X"32",
		X"9B",X"4E",X"C9",X"21",X"85",X"9C",X"DD",X"21",X"9C",X"4E",X"FD",X"21",X"8C",X"4E",X"CD",X"8E",
		X"9D",X"32",X"91",X"4E",X"21",X"C5",X"9C",X"DD",X"21",X"AC",X"4E",X"FD",X"21",X"92",X"4E",X"CD",
		X"8E",X"9D",X"32",X"96",X"4E",X"21",X"05",X"9D",X"DD",X"21",X"BC",X"4E",X"FD",X"21",X"97",X"4E",
		X"CD",X"8E",X"9D",X"32",X"9B",X"4E",X"AF",X"32",X"90",X"4E",X"C9",X"DD",X"7E",X"00",X"A7",X"CA",
		X"94",X"9D",X"4F",X"06",X"08",X"1E",X"80",X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",
		X"DD",X"7E",X"02",X"A3",X"20",X"07",X"DD",X"73",X"02",X"05",X"DF",X"18",X"0C",X"DD",X"35",X"0C",
		X"C2",X"77",X"9D",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",
		X"07",X"FE",X"F0",X"DA",X"45",X"9D",X"21",X"03",X"9C",X"E5",X"E6",X"0F",X"E7",X"EA",X"9E",X"FA",
		X"9E",X"0C",X"9F",X"1E",X"9F",X"30",X"9F",X"EF",X"9B",X"EF",X"9B",X"EF",X"9B",X"EF",X"9B",X"EF",
		X"9B",X"EF",X"9B",X"EF",X"9B",X"EF",X"9B",X"EF",X"9B",X"EF",X"9B",X"42",X"9F",X"00",X"57",X"5C",
		X"61",X"67",X"6D",X"74",X"7B",X"82",X"8A",X"92",X"9A",X"A3",X"AD",X"B8",X"C3",X"01",X"02",X"04",
		X"08",X"10",X"20",X"40",X"80",X"51",X"A4",X"A8",X"A4",X"EF",X"A4",X"FF",X"FF",X"11",X"A5",X"2E",
		X"A5",X"46",X"A5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"A4",X"DC",X"A4",X"FE",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"76",X"10",X"02",X"8E",X"00",X"01",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"37",X"10",X"02",X"8E",X"00",X"01",X"0F",X"00",X"12",X"10",X"02",
		X"8E",X"00",X"01",X"0F",X"00",X"24",X"20",X"00",X"0E",X"00",X"01",X"1F",X"00",X"14",X"20",X"00",
		X"12",X"00",X"01",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"42",X"00",X"02",
		X"20",X"00",X"01",X"0C",X"00",X"40",X"00",X"06",X"08",X"00",X"00",X"0A",X"00",X"56",X"10",X"02",
		X"8C",X"00",X"00",X"0A",X"00",X"40",X"40",X"08",X"88",X"00",X"01",X"15",X"00",X"41",X"40",X"08",
		X"88",X"00",X"01",X"15",X"00",X"32",X"40",X"08",X"88",X"00",X"01",X"15",X"00",X"43",X"40",X"08",
		X"88",X"00",X"01",X"15",X"00",X"24",X"40",X"08",X"88",X"00",X"01",X"15",X"00",X"15",X"40",X"08",
		X"88",X"00",X"01",X"15",X"00",X"46",X"40",X"08",X"88",X"00",X"01",X"15",X"00",X"37",X"40",X"08",
		X"88",X"00",X"01",X"15",X"00",X"47",X"E6",X"1F",X"28",X"03",X"DD",X"70",X"0D",X"DD",X"4E",X"09",
		X"DD",X"7E",X"0B",X"E6",X"08",X"28",X"02",X"0E",X"00",X"DD",X"71",X"0F",X"78",X"07",X"07",X"07",
		X"E6",X"07",X"21",X"4D",X"9C",X"D7",X"DD",X"77",X"0C",X"78",X"E6",X"1F",X"28",X"09",X"E6",X"0F",
		X"21",X"3D",X"9C",X"D7",X"DD",X"77",X"0E",X"DD",X"6E",X"0E",X"26",X"00",X"DD",X"7E",X"0D",X"E6",
		X"10",X"28",X"02",X"3E",X"01",X"DD",X"86",X"04",X"CA",X"88",X"9E",X"C3",X"84",X"9E",X"DD",X"7E",
		X"00",X"A7",X"20",X"27",X"DD",X"7E",X"02",X"A7",X"C8",X"DD",X"36",X"02",X"00",X"DD",X"36",X"0D",
		X"00",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"00",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",
		X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",X"00",X"AF",X"C9",X"4F",X"06",X"08",X"1E",X"80",
		X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",X"DD",X"7E",X"02",X"A3",X"20",X"3F",X"DD",
		X"73",X"02",X"05",X"78",X"07",X"07",X"07",X"4F",X"06",X"00",X"E5",X"09",X"DD",X"E5",X"D1",X"13",
		X"13",X"13",X"01",X"08",X"00",X"ED",X"B0",X"E1",X"DD",X"7E",X"06",X"E6",X"7F",X"DD",X"77",X"0C",
		X"DD",X"7E",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"DD",X"77",X"0B",X"E6",X"08",X"20",X"07",X"DD",X"70",X"0F",X"DD",X"36",X"0D",X"00",X"DD",X"35",
		X"0C",X"20",X"5A",X"DD",X"7E",X"08",X"A7",X"28",X"10",X"DD",X"35",X"08",X"20",X"0B",X"7B",X"2F",
		X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"8E",X"9D",X"DD",X"7E",X"06",X"E6",X"7F",X"DD",X"77",
		X"0C",X"DD",X"CB",X"06",X"7E",X"28",X"16",X"DD",X"7E",X"05",X"ED",X"44",X"DD",X"77",X"05",X"DD",
		X"CB",X"0D",X"46",X"DD",X"CB",X"0D",X"C6",X"28",X"24",X"DD",X"CB",X"0D",X"86",X"DD",X"7E",X"04",
		X"DD",X"86",X"07",X"DD",X"77",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",X"DD",X"86",X"0A",X"DD",
		X"77",X"09",X"47",X"DD",X"7E",X"0B",X"E6",X"08",X"20",X"03",X"DD",X"70",X"0F",X"DD",X"7E",X"0E",
		X"DD",X"86",X"05",X"DD",X"77",X"0E",X"6F",X"26",X"00",X"DD",X"7E",X"03",X"E6",X"70",X"28",X"08",
		X"0F",X"0F",X"0F",X"0F",X"47",X"29",X"10",X"FD",X"FD",X"75",X"00",X"7D",X"0F",X"0F",X"0F",X"0F",
		X"FD",X"77",X"01",X"FD",X"74",X"02",X"7C",X"0F",X"0F",X"0F",X"0F",X"FD",X"77",X"03",X"DD",X"7E",
		X"0B",X"E7",X"C2",X"9E",X"C6",X"9E",X"CB",X"9E",X"DC",X"9E",X"E3",X"9E",X"C5",X"9E",X"C5",X"9E",
		X"C5",X"9E",X"C5",X"9E",X"C5",X"9E",X"C5",X"9E",X"C5",X"9E",X"C5",X"9E",X"C5",X"9E",X"C5",X"9E",
		X"C5",X"9E",X"DD",X"7E",X"0F",X"C9",X"DD",X"7E",X"0F",X"18",X"09",X"3A",X"84",X"4C",X"E6",X"01",
		X"DD",X"7E",X"0F",X"C0",X"E6",X"0F",X"C8",X"3D",X"DD",X"77",X"0F",X"C9",X"3A",X"84",X"4C",X"E6",
		X"03",X"18",X"ED",X"3A",X"84",X"4C",X"E6",X"07",X"18",X"E6",X"DD",X"6E",X"06",X"DD",X"66",X"07",
		X"7E",X"DD",X"77",X"06",X"23",X"7E",X"DD",X"77",X"07",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",
		X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"03",X"C9",X"DD",X"6E",X"06",X"DD",
		X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"04",X"C9",X"DD",X"6E",
		X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"09",X"C9",
		X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",
		X"0B",X"C9",X"DD",X"7E",X"02",X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"94",X"9D",X"31",
		X"C0",X"4F",X"21",X"00",X"4C",X"06",X"04",X"32",X"C0",X"50",X"36",X"00",X"2C",X"20",X"FB",X"24",
		X"10",X"F5",X"21",X"00",X"40",X"06",X"04",X"32",X"C0",X"50",X"3E",X"40",X"77",X"2C",X"20",X"FC",
		X"24",X"10",X"F4",X"06",X"04",X"32",X"C0",X"50",X"3E",X"0D",X"77",X"2C",X"20",X"FC",X"24",X"10",
		X"F4",X"21",X"06",X"50",X"3E",X"01",X"77",X"2D",X"20",X"FC",X"AF",X"32",X"03",X"50",X"3E",X"01",
		X"ED",X"47",X"31",X"C0",X"4F",X"32",X"C0",X"50",X"AF",X"32",X"00",X"4E",X"3C",X"32",X"01",X"4E",
		X"32",X"00",X"50",X"FB",X"3A",X"80",X"50",X"E6",X"03",X"C6",X"25",X"47",X"CD",X"F2",X"9A",X"3A",
		X"80",X"50",X"0F",X"0F",X"0F",X"0F",X"E6",X"03",X"FE",X"03",X"20",X"0E",X"06",X"2A",X"CD",X"F2",
		X"9A",X"C3",X"E7",X"9F",X"35",X"40",X"30",X"31",X"35",X"31",X"07",X"5F",X"D5",X"06",X"2B",X"CD",
		X"F2",X"9A",X"06",X"2E",X"CD",X"F2",X"9A",X"D1",X"16",X"00",X"21",X"C4",X"9F",X"19",X"7E",X"32",
		X"2A",X"42",X"23",X"7E",X"32",X"4A",X"42",X"3A",X"80",X"50",X"0F",X"0F",X"E6",X"03",X"C6",X"31",
		X"FE",X"34",X"20",X"01",X"3C",X"32",X"0C",X"42",X"06",X"29",X"CD",X"F2",X"9A",X"3A",X"80",X"50",
		X"07",X"07",X"E6",X"01",X"C6",X"2C",X"47",X"CD",X"F2",X"9A",X"3A",X"80",X"50",X"07",X"D2",X"95",
		X"9F",X"AF",X"32",X"00",X"50",X"F3",X"21",X"07",X"50",X"AF",X"77",X"2D",X"20",X"FC",X"31",X"54",
		X"A0",X"06",X"03",X"D9",X"E1",X"D1",X"32",X"C0",X"50",X"C1",X"3E",X"3C",X"77",X"23",X"72",X"23",
		X"10",X"F8",X"3B",X"3B",X"C1",X"71",X"23",X"3E",X"3F",X"77",X"23",X"10",X"F8",X"3B",X"3B",X"1D",
		X"C2",X"26",X"A0",X"F1",X"D9",X"10",X"DC",X"31",X"C0",X"4F",X"06",X"08",X"CD",X"66",X"A0",X"10",
		X"FB",X"C3",X"60",X"92",X"02",X"40",X"01",X"3E",X"3D",X"10",X"40",X"40",X"0E",X"3D",X"3E",X"10",
		X"C2",X"43",X"01",X"3E",X"3D",X"10",X"32",X"C0",X"50",X"21",X"00",X"28",X"2B",X"7C",X"B5",X"20",
		X"FB",X"C9",X"5D",X"A5",X"6D",X"A5",X"7C",X"A5",X"85",X"A7",X"85",X"A7",X"8B",X"A5",X"9A",X"A5",
		X"A6",X"A5",X"BD",X"A5",X"D1",X"A5",X"E5",X"A5",X"04",X"A6",X"85",X"A7",X"85",X"A7",X"85",X"A7",
		X"85",X"A7",X"85",X"A7",X"85",X"A7",X"85",X"A7",X"12",X"A6",X"28",X"A6",X"32",X"A6",X"3C",X"A6",
		X"46",X"A6",X"50",X"A6",X"5A",X"A6",X"64",X"A6",X"6E",X"A6",X"78",X"A6",X"82",X"A6",X"8C",X"A6",
		X"96",X"A6",X"A0",X"A6",X"AA",X"A6",X"B4",X"A6",X"BE",X"A6",X"CE",X"A6",X"DE",X"A6",X"F5",X"A6",
		X"0C",X"A7",X"23",X"A7",X"3A",X"A7",X"45",X"A7",X"56",X"A7",X"62",X"A7",X"6F",X"A7",X"7C",X"A7",
		X"E4",X"E8",X"E5",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"D0",X"D0",X"D0",X"40",X"C4",X"C5",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",
		X"E6",X"D0",X"E7",X"74",X"E1",X"D6",X"C7",X"D0",X"D0",X"74",X"E1",X"D6",X"C7",X"74",X"E1",X"D6",
		X"C7",X"D0",X"74",X"E1",X"D5",X"C0",X"40",X"C6",X"C7",X"D0",X"D0",X"74",X"E1",X"D6",X"C7",X"00",
		X"E6",X"D0",X"E7",X"73",X"75",X"D3",X"C0",X"D0",X"D0",X"73",X"75",X"D3",X"C0",X"73",X"75",X"D3",
		X"C0",X"D0",X"73",X"75",X"D3",X"C5",X"40",X"C2",X"C0",X"D0",X"D0",X"73",X"75",X"D3",X"C0",X"00",
		X"E6",X"D0",X"E7",X"72",X"E0",X"D4",X"C5",X"D0",X"D0",X"72",X"E0",X"D4",X"C5",X"72",X"E0",X"D4",
		X"C5",X"D0",X"72",X"E0",X"D4",X"C0",X"40",X"C4",X"C5",X"D0",X"D0",X"72",X"E0",X"D4",X"C5",X"00",
		X"E6",X"D0",X"E7",X"D0",X"40",X"C2",X"C0",X"D0",X"D0",X"D0",X"40",X"C2",X"C0",X"D0",X"40",X"C2",
		X"C0",X"D0",X"D0",X"40",X"CC",X"CD",X"63",X"C9",X"C0",X"40",X"C6",X"C7",X"40",X"C2",X"C0",X"00",
		X"E2",X"E8",X"E3",X"D0",X"40",X"C4",X"C5",X"40",X"DB",X"DE",X"63",X"C9",X"C5",X"D0",X"40",X"C4",
		X"C5",X"D0",X"D0",X"40",X"60",X"61",X"61",X"C4",X"C5",X"40",X"CC",X"CD",X"63",X"C9",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"C2",X"C0",X"40",X"60",X"61",X"61",X"C2",X"C0",X"D0",X"40",X"C2",
		X"C0",X"D0",X"D0",X"40",X"CA",X"CB",X"62",X"C8",X"C0",X"40",X"60",X"61",X"61",X"C2",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"C4",X"C5",X"40",X"CA",X"CB",X"62",X"C8",X"C5",X"D0",X"40",X"C4",
		X"C5",X"D0",X"D0",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"40",X"CA",X"CB",X"62",X"C8",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"CC",X"CD",X"63",X"C9",X"C5",X"40",X"CC",X"CD",X"CF",X"63",X"C9",
		X"C0",X"E9",X"D0",X"40",X"C4",X"C5",X"40",X"CC",X"CD",X"63",X"C9",X"C5",X"40",X"C2",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"60",X"61",X"61",X"C2",X"C0",X"40",X"60",X"61",X"61",X"61",X"C4",
		X"C5",X"D0",X"40",X"40",X"C2",X"C0",X"40",X"1C",X"1D",X"61",X"C2",X"C0",X"40",X"C4",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"CA",X"CB",X"62",X"C8",X"C5",X"40",X"CA",X"CB",X"CE",X"62",X"C8",
		X"C0",X"40",X"40",X"C6",X"F3",X"C5",X"40",X"CA",X"CB",X"62",X"C8",X"C5",X"40",X"C2",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"C2",X"C0",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"D0",X"40",X"C4",
		X"C5",X"40",X"C6",X"F3",X"F7",X"C0",X"40",X"C4",X"C5",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"CC",X"CD",X"63",X"F1",X"CD",X"63",X"F1",X"CD",X"CF",X"63",X"F1",
		X"CD",X"63",X"F1",X"F5",X"F5",X"CD",X"63",X"F1",X"CD",X"63",X"F1",X"CD",X"63",X"C9",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"1C",X"1D",X"61",X"60",X"61",X"61",X"1C",X"1D",X"1D",X"61",X"60",
		X"61",X"61",X"1C",X"1D",X"1D",X"1D",X"61",X"60",X"61",X"61",X"1C",X"1D",X"61",X"C4",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"CA",X"CB",X"62",X"F0",X"CB",X"62",X"F0",X"CB",X"CE",X"62",X"F0",
		X"CB",X"62",X"F0",X"F4",X"F4",X"CB",X"62",X"F0",X"CB",X"62",X"F0",X"CB",X"62",X"C8",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"C2",X"C0",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"D0",X"40",X"C2",
		X"C5",X"40",X"C1",X"F2",X"F6",X"C5",X"40",X"C4",X"C5",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"C4",X"C5",X"40",X"C4",X"C5",X"40",X"CC",X"CD",X"CF",X"63",X"C9",
		X"C0",X"40",X"40",X"C1",X"F2",X"C0",X"40",X"C2",X"C0",X"40",X"C4",X"C5",X"40",X"C2",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"CC",X"CD",X"63",X"C9",X"C0",X"40",X"60",X"61",X"61",X"61",X"C2",
		X"C5",X"D0",X"40",X"40",X"CC",X"CD",X"63",X"C9",X"C5",X"40",X"CC",X"CD",X"63",X"C9",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"60",X"61",X"61",X"C4",X"C5",X"40",X"CA",X"CB",X"CE",X"62",X"C8",
		X"C0",X"D0",X"D0",X"40",X"60",X"61",X"61",X"C2",X"C0",X"40",X"60",X"61",X"61",X"C2",X"C0",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"CA",X"CB",X"62",X"C8",X"C0",X"40",X"C4",X"C5",X"D0",X"40",X"C4",
		X"C5",X"DF",X"D0",X"40",X"CA",X"CB",X"62",X"C8",X"C5",X"40",X"CA",X"CB",X"62",X"C8",X"C5",X"00",
		X"D0",X"D0",X"D0",X"E7",X"40",X"C4",X"C5",X"40",X"C4",X"C5",X"40",X"CC",X"CD",X"CF",X"63",X"C9",
		X"C0",X"D0",X"D0",X"40",X"C2",X"C0",X"40",X"CC",X"CD",X"63",X"C9",X"C5",X"40",X"C2",X"C0",X"00",
		X"E4",X"E8",X"E5",X"74",X"E1",X"D5",X"C0",X"40",X"C2",X"C0",X"40",X"60",X"61",X"61",X"61",X"C4",
		X"C5",X"D0",X"D0",X"40",X"C4",X"C5",X"40",X"60",X"61",X"61",X"C2",X"C0",X"40",X"C4",X"C5",X"00",
		X"E6",X"D0",X"E7",X"73",X"75",X"D2",X"C5",X"40",X"C4",X"C5",X"40",X"D9",X"DA",X"CE",X"62",X"C8",
		X"C0",X"D0",X"D0",X"40",X"C2",X"C0",X"40",X"D9",X"DA",X"62",X"C8",X"C5",X"40",X"C2",X"C0",X"00",
		X"E6",X"D0",X"E7",X"72",X"E0",X"D1",X"C3",X"40",X"C2",X"C0",X"D0",X"D0",X"D0",X"D0",X"40",X"C4",
		X"C5",X"D0",X"D0",X"40",X"C4",X"C5",X"D0",X"D0",X"D0",X"D0",X"C1",X"C3",X"40",X"C4",X"C5",X"00",
		X"E6",X"D0",X"E7",X"D0",X"D0",X"D0",X"74",X"E1",X"D5",X"C0",X"D0",X"D0",X"D0",X"74",X"E1",X"D5",
		X"C0",X"D0",X"74",X"E1",X"D5",X"C0",X"D0",X"D0",X"D0",X"D0",X"D0",X"74",X"E1",X"D5",X"C0",X"00",
		X"E6",X"D0",X"E7",X"D0",X"D0",X"D0",X"73",X"75",X"D2",X"C5",X"D0",X"D0",X"D0",X"73",X"75",X"D2",
		X"C5",X"D0",X"73",X"75",X"D2",X"C5",X"D0",X"D0",X"D0",X"D0",X"D0",X"73",X"75",X"D2",X"C5",X"00",
		X"E2",X"E8",X"E3",X"D0",X"D0",X"D0",X"72",X"E0",X"D1",X"C3",X"D0",X"D0",X"D0",X"72",X"E0",X"D1",
		X"C3",X"D0",X"72",X"E0",X"D1",X"C3",X"D0",X"D0",X"D0",X"D0",X"D0",X"72",X"E0",X"D4",X"C0",X"00",
		X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"40",X"C2",X"C0",X"00",
		X"27",X"F1",X"07",X"F2",X"03",X"F3",X"08",X"F4",X"01",X"82",X"86",X"8B",X"69",X"8B",X"84",X"87",
		X"8D",X"6B",X"8D",X"86",X"89",X"F2",X"04",X"84",X"62",X"64",X"62",X"62",X"82",X"84",X"82",X"F2",
		X"03",X"6D",X"6B",X"69",X"67",X"67",X"87",X"F2",X"04",X"82",X"F2",X"03",X"8D",X"6B",X"69",X"67",
		X"66",X"66",X"86",X"62",X"62",X"66",X"66",X"64",X"64",X"67",X"67",X"66",X"66",X"69",X"69",X"67",
		X"67",X"6B",X"6B",X"69",X"69",X"6D",X"6D",X"6B",X"6B",X"6D",X"6D",X"F2",X"04",X"64",X"62",X"F3",
		X"00",X"60",X"F3",X"0F",X"82",X"FF",X"FF",X"FF",X"F1",X"07",X"F2",X"03",X"F3",X"0F",X"F4",X"01",
		X"82",X"86",X"8B",X"69",X"8B",X"84",X"87",X"8D",X"6B",X"8D",X"86",X"89",X"F2",X"04",X"84",X"62",
		X"64",X"62",X"62",X"82",X"FF",X"FF",X"FF",X"F1",X"05",X"F2",X"01",X"F3",X"0F",X"F4",X"03",X"46",
		X"F3",X"00",X"40",X"F3",X"0F",X"42",X"F3",X"00",X"40",X"FF",X"FF",X"FF",X"F1",X"04",X"F2",X"01",
		X"F3",X"0F",X"F4",X"00",X"49",X"47",X"46",X"44",X"42",X"49",X"47",X"46",X"44",X"42",X"FF",X"F1",
		X"06",X"F2",X"03",X"F3",X"0F",X"F4",X"01",X"67",X"6B",X"6E",X"F2",X"04",X"A7",X"FF",X"F1",X"06",
		X"F2",X"03",X"F3",X"0F",X"F4",X"02",X"29",X"27",X"26",X"24",X"22",X"29",X"27",X"26",X"24",X"22",
		X"FF",X"F1",X"06",X"F2",X"06",X"F3",X"0F",X"F4",X"01",X"89",X"89",X"89",X"89",X"89",X"89",X"8D",
		X"89",X"86",X"86",X"84",X"86",X"88",X"89",X"8B",X"8B",X"8D",X"8D",X"89",X"89",X"FF",X"F1",X"06",
		X"F2",X"05",X"F3",X"0F",X"F4",X"02",X"89",X"66",X"82",X"89",X"66",X"82",X"89",X"66",X"8E",X"F3",
		X"00",X"60",X"F3",X"0F",X"AE",X"FF",X"F1",X"06",X"F2",X"05",X"F3",X"0F",X"F4",X"02",X"82",X"F2",
		X"04",X"69",X"F2",X"05",X"62",X"86",X"62",X"66",X"89",X"89",X"69",X"89",X"FF",X"D4",X"83",X"48",
		X"49",X"47",X"48",X"40",X"53",X"43",X"4F",X"52",X"45",X"27",X"8D",X"27",X"80",X"3D",X"80",X"43",
		X"52",X"45",X"44",X"49",X"54",X"40",X"40",X"40",X"27",X"8D",X"27",X"80",X"3D",X"80",X"46",X"52",
		X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"27",X"8D",X"27",X"80",X"1D",X"80",X"47",X"41",X"4D",
		X"45",X"40",X"4F",X"56",X"45",X"52",X"27",X"9C",X"27",X"80",X"12",X"80",X"53",X"54",X"41",X"52",
		X"54",X"5B",X"27",X"9C",X"27",X"93",X"EE",X"02",X"50",X"55",X"53",X"48",X"40",X"53",X"54",X"41",
		X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"27",X"88",X"27",X"80",X"B2",X"02",X"31",
		X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"4C",X"59",X"40",X"27",X"86",X"27",
		X"80",X"B2",X"02",X"31",X"40",X"4F",X"52",X"40",X"32",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"53",X"27",X"86",X"27",X"80",X"76",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"4D",X"4F",X"55",
		X"53",X"45",X"40",X"46",X"4F",X"52",X"40",X"40",X"40",X"30",X"30",X"30",X"40",X"5D",X"5E",X"5F",
		X"27",X"8B",X"27",X"80",X"33",X"80",X"40",X"51",X"40",X"52",X"49",X"56",X"45",X"52",X"27",X"84",
		X"27",X"80",X"FA",X"02",X"40",X"40",X"40",X"51",X"55",X"45",X"45",X"4E",X"40",X"52",X"49",X"56",
		X"45",X"52",X"40",X"40",X"27",X"84",X"27",X"80",X"C1",X"00",X"40",X"40",X"40",X"40",X"27",X"84",
		X"27",X"80",X"C1",X"00",X"40",X"40",X"40",X"40",X"27",X"93",X"27",X"80",X"C1",X"00",X"40",X"40",
		X"33",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",X"40",X"40",X"35",X"30",X"27",X"84",X"27",X"80",
		X"C1",X"00",X"40",X"40",X"37",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",X"40",X"31",X"30",X"30",
		X"27",X"84",X"27",X"80",X"C1",X"00",X"40",X"32",X"30",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",
		X"40",X"33",X"30",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",X"40",X"35",X"30",X"30",X"27",X"84",
		X"27",X"80",X"C1",X"00",X"40",X"37",X"30",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",X"31",X"30",
		X"30",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",X"32",X"30",X"30",X"30",X"27",X"84",X"27",X"80",
		X"C1",X"00",X"33",X"30",X"30",X"30",X"27",X"84",X"27",X"80",X"C1",X"00",X"35",X"30",X"30",X"30",
		X"27",X"84",X"27",X"80",X"C1",X"00",X"37",X"30",X"30",X"30",X"27",X"84",X"27",X"80",X"04",X"03",
		X"4D",X"45",X"4D",X"4F",X"52",X"59",X"40",X"40",X"4F",X"4B",X"27",X"8D",X"27",X"80",X"04",X"03",
		X"42",X"41",X"44",X"40",X"40",X"40",X"40",X"52",X"40",X"4D",X"27",X"8D",X"27",X"80",X"08",X"03",
		X"46",X"52",X"45",X"45",X"40",X"40",X"50",X"4C",X"41",X"59",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"27",X"8D",X"27",X"80",X"08",X"03",X"31",X"40",X"43",X"4F",X"49",X"4E",X"40",X"40",X"31",
		X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"27",X"8D",X"27",X"80",X"08",X"03",X"31",X"40",
		X"43",X"4F",X"49",X"4E",X"40",X"40",X"32",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"27",
		X"8D",X"27",X"80",X"08",X"03",X"32",X"40",X"43",X"4F",X"49",X"4E",X"53",X"40",X"31",X"40",X"43",
		X"52",X"45",X"44",X"49",X"54",X"40",X"27",X"8D",X"27",X"80",X"0C",X"03",X"4D",X"4F",X"55",X"53",
		X"45",X"27",X"8D",X"27",X"80",X"0A",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"4E",X"4F",
		X"4E",X"45",X"27",X"8D",X"27",X"80",X"0A",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"27",X"8D",
		X"27",X"80",X"0E",X"03",X"54",X"41",X"42",X"4C",X"45",X"40",X"40",X"27",X"8D",X"27",X"80",X"0E",
		X"03",X"55",X"50",X"52",X"49",X"47",X"48",X"54",X"27",X"8D",X"27",X"80",X"0A",X"02",X"30",X"30",
		X"30",X"27",X"8D",X"27",X"80",X"52",X"02",X"4E",X"4F",X"40",X"45",X"4E",X"54",X"52",X"59",X"40",
		X"44",X"41",X"54",X"41",X"27",X"82",X"27",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"00",X"4E",X"E7",X"0C",X"B0",X"30",X"B0",X"52",X"B1",X"28",X"B2",X"3A",X"01",X"4E",X"E7",
		X"14",X"B0",X"44",X"B0",X"EF",X"00",X"00",X"EF",X"06",X"00",X"EF",X"01",X"00",X"EF",X"14",X"00",
		X"EF",X"18",X"00",X"EF",X"07",X"00",X"21",X"01",X"4E",X"34",X"21",X"01",X"50",X"36",X"01",X"C9",
		X"CD",X"27",X"9A",X"3A",X"6E",X"4E",X"A7",X"28",X"0C",X"AF",X"32",X"04",X"4E",X"32",X"02",X"4E",
		X"21",X"00",X"4E",X"34",X"C9",X"3A",X"02",X"4E",X"E7",X"77",X"B0",X"44",X"B0",X"91",X"B0",X"44",
		X"B0",X"AA",X"B0",X"44",X"B0",X"9F",X"B0",X"44",X"B0",X"AA",X"B0",X"44",X"B0",X"9F",X"B0",X"44",
		X"B0",X"AA",X"B0",X"44",X"B0",X"9F",X"B0",X"44",X"B0",X"AA",X"B0",X"44",X"B0",X"9F",X"B0",X"44",
		X"B0",X"B6",X"B0",X"44",X"B0",X"D4",X"B0",X"EF",X"00",X"01",X"EF",X"06",X"00",X"EF",X"02",X"00",
		X"EF",X"01",X"01",X"EF",X"11",X"00",X"EF",X"1C",X"05",X"CD",X"62",X"B2",X"0E",X"0B",X"C3",X"1E",
		X"B1",X"AF",X"CD",X"FF",X"B0",X"CD",X"D8",X"B0",X"F7",X"45",X"02",X"00",X"C3",X"27",X"B1",X"AF",
		X"CD",X"FF",X"B0",X"F7",X"45",X"02",X"00",X"C3",X"27",X"B1",X"3E",X"9A",X"CD",X"FF",X"B0",X"F7",
		X"45",X"02",X"00",X"C3",X"27",X"B1",X"3E",X"9B",X"CD",X"FF",X"B0",X"F7",X"45",X"02",X"00",X"AF",
		X"32",X"15",X"4E",X"32",X"70",X"4E",X"3C",X"32",X"14",X"4E",X"AF",X"32",X"07",X"4E",X"32",X"08",
		X"4E",X"C3",X"27",X"B1",X"CD",X"28",X"B2",X"C9",X"06",X"07",X"21",X"01",X"41",X"11",X"1F",X"00",
		X"3E",X"9E",X"CD",X"17",X"9A",X"19",X"3C",X"10",X"F9",X"77",X"23",X"3C",X"77",X"21",X"60",X"42",
		X"11",X"20",X"00",X"3C",X"77",X"19",X"3C",X"77",X"19",X"3C",X"77",X"19",X"3C",X"77",X"C9",X"21",
		X"01",X"45",X"11",X"40",X"00",X"06",X"07",X"CD",X"02",X"9A",X"19",X"10",X"FA",X"77",X"23",X"77",
		X"21",X"60",X"46",X"11",X"20",X"00",X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"C9",X"06",X"1C",
		X"CD",X"42",X"00",X"F7",X"4A",X"02",X"00",X"21",X"02",X"4E",X"34",X"C9",X"06",X"1C",X"CD",X"42",
		X"00",X"F7",X"45",X"02",X"00",X"C3",X"27",X"B1",X"3A",X"C1",X"4D",X"A7",X"C8",X"AF",X"32",X"C1",
		X"4D",X"3A",X"3A",X"4D",X"EE",X"02",X"32",X"34",X"4D",X"47",X"21",X"0A",X"03",X"DF",X"22",X"2C",
		X"4D",X"C9",X"3A",X"03",X"4E",X"E7",X"60",X"B1",X"8A",X"B1",X"DF",X"B1",X"44",X"B0",X"12",X"B2",
		X"CD",X"27",X"9A",X"EF",X"1C",X"85",X"EF",X"00",X"01",X"EF",X"1C",X"07",X"EF",X"1C",X"8B",X"EF",
		X"1C",X"13",X"EF",X"1E",X"00",X"CD",X"0D",X"B2",X"3E",X"01",X"32",X"E0",X"4D",X"3A",X"71",X"4E",
		X"FE",X"FF",X"C8",X"EF",X"1C",X"0A",X"EF",X"1F",X"00",X"C9",X"CD",X"27",X"9A",X"3A",X"6E",X"4E",
		X"FE",X"01",X"06",X"09",X"20",X"02",X"06",X"08",X"CD",X"F2",X"9A",X"3A",X"6E",X"4E",X"FE",X"01",
		X"3A",X"40",X"50",X"28",X"0B",X"CB",X"77",X"20",X"07",X"3E",X"01",X"32",X"70",X"4E",X"18",X"07",
		X"CB",X"6F",X"C0",X"AF",X"32",X"70",X"4E",X"3A",X"6B",X"4E",X"A7",X"28",X"15",X"3A",X"70",X"4E",
		X"A7",X"3A",X"6E",X"4E",X"28",X"03",X"C6",X"99",X"27",X"C6",X"99",X"27",X"32",X"6E",X"4E",X"CD",
		X"27",X"9A",X"CD",X"0D",X"B2",X"AF",X"32",X"E0",X"4D",X"3E",X"02",X"32",X"CC",X"4E",X"C9",X"EF",
		X"00",X"01",X"EF",X"01",X"01",X"EF",X"02",X"00",X"EF",X"12",X"00",X"EF",X"1C",X"06",X"EF",X"18",
		X"00",X"EF",X"1B",X"00",X"AF",X"32",X"13",X"4E",X"3A",X"6F",X"4E",X"32",X"14",X"4E",X"32",X"15",
		X"4E",X"C6",X"02",X"32",X"23",X"4E",X"EF",X"1A",X"00",X"F7",X"4A",X"01",X"00",X"21",X"03",X"4E",
		X"34",X"C9",X"21",X"15",X"4E",X"35",X"CD",X"EC",X"99",X"AF",X"32",X"03",X"4E",X"32",X"02",X"4E",
		X"32",X"04",X"4E",X"21",X"00",X"4E",X"34",X"C9",X"3A",X"04",X"4E",X"E7",X"86",X"B2",X"8B",X"B2",
		X"44",X"B0",X"CF",X"B2",X"4C",X"B3",X"44",X"B0",X"71",X"B3",X"44",X"B0",X"AD",X"B3",X"C3",X"B3",
		X"44",X"B0",X"2E",X"B4",X"34",X"B4",X"44",X"B0",X"40",X"B4",X"44",X"B0",X"59",X"B4",X"7D",X"B4",
		X"44",X"B0",X"2E",X"B4",X"44",X"B0",X"44",X"B0",X"44",X"B0",X"44",X"B0",X"06",X"B4",X"44",X"B0",
		X"2E",X"B4",X"21",X"09",X"4E",X"AF",X"06",X"0B",X"CF",X"32",X"22",X"4E",X"CD",X"0D",X"94",X"2A",
		X"73",X"4E",X"22",X"0A",X"4E",X"21",X"0A",X"4E",X"11",X"38",X"4E",X"01",X"1E",X"00",X"ED",X"B0",
		X"C9",X"21",X"04",X"4E",X"34",X"C9",X"CD",X"62",X"B2",X"18",X"F6",X"3A",X"00",X"4E",X"3D",X"20",
		X"06",X"3E",X"18",X"32",X"04",X"4E",X"C9",X"EF",X"11",X"00",X"EF",X"05",X"00",X"EF",X"10",X"00",
		X"EF",X"1A",X"00",X"F7",X"54",X"00",X"00",X"F7",X"54",X"06",X"00",X"3A",X"72",X"4E",X"47",X"3A",
		X"09",X"4E",X"A0",X"32",X"03",X"50",X"18",X"C9",X"3A",X"00",X"50",X"CB",X"67",X"20",X"09",X"21",
		X"04",X"4E",X"36",X"0E",X"EF",X"13",X"00",X"C9",X"CD",X"7E",X"85",X"28",X"36",X"18",X"64",X"3A",
		X"22",X"4E",X"E7",X"00",X"80",X"B8",X"B2",X"46",X"80",X"3E",X"80",X"57",X"80",X"87",X"80",X"83",
		X"80",X"3A",X"80",X"36",X"80",X"1C",X"80",X"8B",X"80",X"8F",X"80",X"42",X"80",X"06",X"80",X"6D",
		X"80",X"93",X"80",X"32",X"80",X"65",X"82",X"8A",X"82",X"93",X"82",X"D0",X"82",X"DA",X"82",X"FF",
		X"FF",X"FF",X"FF",X"3A",X"06",X"4E",X"E7",X"CE",X"85",X"44",X"B0",X"97",X"85",X"44",X"B0",X"A8",
		X"85",X"44",X"B0",X"B4",X"85",X"44",X"B0",X"A8",X"85",X"44",X"B0",X"B8",X"85",X"44",X"B0",X"A8",
		X"85",X"44",X"B0",X"9C",X"85",X"44",X"B0",X"A8",X"85",X"44",X"B0",X"B8",X"85",X"44",X"B0",X"BC",
		X"85",X"C4",X"85",X"CD",X"96",X"06",X"CD",X"B1",X"B4",X"CD",X"B1",X"B4",X"CD",X"44",X"06",X"CD",
		X"60",X"06",X"CD",X"FA",X"05",X"CD",X"CD",X"05",X"CD",X"85",X"B7",X"C9",X"3E",X"01",X"32",X"12",
		X"4E",X"CD",X"81",X"B2",X"3A",X"14",X"4E",X"A7",X"C2",X"81",X"B2",X"3A",X"70",X"4E",X"A7",X"CA",
		X"81",X"B2",X"3A",X"42",X"4E",X"A7",X"CA",X"81",X"B2",X"EF",X"1C",X"05",X"F7",X"54",X"00",X"00",
		X"C9",X"3A",X"70",X"4E",X"A7",X"28",X"06",X"3A",X"42",X"4E",X"A7",X"20",X"13",X"3A",X"14",X"4E",
		X"A7",X"20",X"24",X"CD",X"27",X"9A",X"EF",X"1C",X"05",X"F7",X"54",X"00",X"00",X"C3",X"81",X"B2",
		X"CD",X"DD",X"05",X"3A",X"09",X"4E",X"EE",X"01",X"32",X"09",X"4E",X"3A",X"22",X"4E",X"A7",X"3E",
		X"11",X"20",X"04",X"32",X"04",X"4E",X"C9",X"3E",X"09",X"32",X"04",X"4E",X"C9",X"AF",X"32",X"02",
		X"4E",X"32",X"04",X"4E",X"32",X"70",X"4E",X"32",X"09",X"4E",X"32",X"03",X"50",X"3E",X"01",X"32",
		X"00",X"4E",X"C9",X"EF",X"00",X"01",X"EF",X"01",X"01",X"EF",X"02",X"00",X"EF",X"11",X"00",X"EF",
		X"13",X"00",X"EF",X"04",X"00",X"EF",X"05",X"00",X"EF",X"10",X"00",X"EF",X"03",X"00",X"EF",X"1A",
		X"00",X"EF",X"1C",X"06",X"F7",X"54",X"00",X"00",X"F7",X"54",X"06",X"00",X"3A",X"72",X"4E",X"47",
		X"3A",X"09",X"4E",X"A0",X"32",X"03",X"50",X"3E",X"01",X"32",X"22",X"4E",X"21",X"0D",X"4E",X"3E",
		X"01",X"AE",X"77",X"C3",X"81",X"B2",X"EF",X"11",X"00",X"EF",X"13",X"00",X"EF",X"05",X"00",X"EF",
		X"10",X"00",X"EF",X"1A",X"00",X"EF",X"1C",X"05",X"EF",X"1D",X"00",X"F7",X"54",X"00",X"00",X"AF",
		X"32",X"03",X"50",X"32",X"22",X"4E",X"3E",X"02",X"32",X"13",X"4E",X"C3",X"81",X"B2",X"3E",X"03",
		X"32",X"04",X"4E",X"C9",X"F7",X"45",X"00",X"00",X"CD",X"81",X"B2",X"AF",X"32",X"CC",X"4E",X"C9",
		X"EF",X"00",X"01",X"EF",X"06",X"00",X"EF",X"11",X"00",X"EF",X"13",X"00",X"EF",X"05",X"00",X"EF",
		X"10",X"13",X"F7",X"43",X"00",X"00",X"C3",X"81",X"B2",X"AF",X"32",X"CC",X"4E",X"06",X"06",X"21",
		X"0C",X"4E",X"CF",X"CD",X"0D",X"94",X"CD",X"81",X"B2",X"21",X"23",X"4E",X"34",X"21",X"13",X"4E",
		X"34",X"2A",X"0A",X"4E",X"7E",X"FE",X"14",X"C8",X"23",X"22",X"0A",X"4E",X"C9",X"EF",X"00",X"01",
		X"EF",X"01",X"01",X"EF",X"02",X"00",X"EF",X"11",X"00",X"EF",X"05",X"00",X"EF",X"10",X"00",X"EF",
		X"1A",X"00",X"EF",X"1C",X"06",X"F7",X"54",X"00",X"00",X"F7",X"54",X"06",X"00",X"3A",X"72",X"4E",
		X"47",X"3A",X"09",X"4E",X"A0",X"32",X"03",X"50",X"AF",X"32",X"22",X"4E",X"21",X"04",X"4E",X"34",
		X"C9",X"CD",X"9D",X"86",X"CD",X"24",X"83",X"CD",X"42",X"83",X"CD",X"A8",X"83",X"CD",X"0E",X"84",
		X"CD",X"74",X"84",X"CD",X"F1",X"85",X"CD",X"A7",X"89",X"CD",X"43",X"8A",X"3A",X"1A",X"4F",X"FE",
		X"08",X"30",X"03",X"CD",X"F1",X"8A",X"CD",X"24",X"8D",X"CD",X"11",X"8E",X"CD",X"C0",X"8E",X"CD",
		X"74",X"8F",X"CD",X"04",X"B8",X"CD",X"BA",X"87",X"C9",X"3A",X"28",X"4F",X"A7",X"C8",X"E1",X"E7",
		X"44",X"B0",X"25",X"B5",X"6A",X"B5",X"AB",X"B5",X"3A",X"29",X"4F",X"A7",X"C8",X"E1",X"E7",X"44",
		X"B0",X"BD",X"B5",X"02",X"B6",X"43",X"B6",X"3A",X"2A",X"4F",X"A7",X"C8",X"E1",X"E7",X"44",X"B0",
		X"55",X"B6",X"9A",X"B6",X"DB",X"B6",X"3A",X"2B",X"4F",X"A7",X"C8",X"E1",X"E7",X"44",X"B0",X"ED",
		X"B6",X"32",X"B7",X"73",X"B7",X"DD",X"21",X"00",X"4D",X"FD",X"21",X"40",X"4C",X"CD",X"BE",X"BB",
		X"DD",X"21",X"3C",X"4D",X"FD",X"21",X"44",X"4D",X"CD",X"6C",X"98",X"CD",X"F9",X"BC",X"30",X"21",
		X"21",X"46",X"4C",X"CD",X"94",X"BC",X"DD",X"21",X"40",X"4C",X"ED",X"5B",X"3C",X"4D",X"CD",X"B0",
		X"BC",X"2A",X"44",X"4C",X"22",X"42",X"4C",X"21",X"33",X"4F",X"36",X"00",X"21",X"28",X"4F",X"34",
		X"C9",X"DD",X"21",X"40",X"4C",X"CD",X"9C",X"BC",X"18",X"DC",X"DD",X"21",X"40",X"4C",X"FD",X"21",
		X"00",X"4D",X"21",X"42",X"4C",X"01",X"00",X"00",X"78",X"ED",X"5B",X"44",X"4C",X"BB",X"28",X"18",
		X"CD",X"6B",X"BC",X"2A",X"00",X"4D",X"CD",X"E5",X"BC",X"38",X"15",X"3A",X"33",X"4F",X"0F",X"0F",
		X"E6",X"C0",X"C6",X"00",X"32",X"2D",X"4F",X"C9",X"BA",X"28",X"05",X"CD",X"75",X"BC",X"18",X"E3",
		X"AF",X"32",X"03",X"4C",X"32",X"2D",X"4F",X"CD",X"5C",X"B5",X"C9",X"3A",X"B7",X"4D",X"A7",X"C0",
		X"3E",X"01",X"32",X"B7",X"4D",X"AF",X"32",X"28",X"4F",X"CD",X"C3",X"BC",X"C9",X"DD",X"21",X"02",
		X"4D",X"FD",X"21",X"48",X"4C",X"CD",X"BE",X"BB",X"DD",X"21",X"3E",X"4D",X"FD",X"21",X"44",X"4D",
		X"CD",X"6C",X"98",X"CD",X"F9",X"BC",X"30",X"21",X"21",X"4E",X"4C",X"CD",X"94",X"BC",X"DD",X"21",
		X"48",X"4C",X"ED",X"5B",X"3E",X"4D",X"CD",X"B0",X"BC",X"2A",X"4C",X"4C",X"22",X"4A",X"4C",X"21",
		X"34",X"4F",X"36",X"00",X"21",X"29",X"4F",X"34",X"C9",X"DD",X"21",X"48",X"4C",X"CD",X"9C",X"BC",
		X"18",X"DC",X"DD",X"21",X"48",X"4C",X"FD",X"21",X"02",X"4D",X"21",X"4A",X"4C",X"01",X"00",X"00",
		X"78",X"ED",X"5B",X"4C",X"4C",X"BB",X"28",X"18",X"CD",X"6B",X"BC",X"2A",X"02",X"4D",X"CD",X"E5",
		X"BC",X"38",X"15",X"3A",X"34",X"4F",X"0F",X"0F",X"E6",X"C0",X"C6",X"00",X"32",X"2E",X"4F",X"C9",
		X"BA",X"28",X"05",X"CD",X"75",X"BC",X"18",X"E3",X"AF",X"32",X"05",X"4C",X"32",X"2E",X"4F",X"CD",
		X"F4",X"B5",X"C9",X"3A",X"B7",X"4D",X"A7",X"C0",X"3E",X"02",X"32",X"B7",X"4D",X"AF",X"32",X"29",
		X"4F",X"CD",X"C3",X"BC",X"C9",X"DD",X"21",X"04",X"4D",X"FD",X"21",X"50",X"4C",X"CD",X"BE",X"BB",
		X"DD",X"21",X"40",X"4D",X"FD",X"21",X"44",X"4D",X"CD",X"6C",X"98",X"CD",X"F9",X"BC",X"30",X"21",
		X"21",X"56",X"4C",X"CD",X"94",X"BC",X"DD",X"21",X"50",X"4C",X"ED",X"5B",X"40",X"4D",X"CD",X"B0",
		X"BC",X"2A",X"54",X"4C",X"22",X"52",X"4C",X"21",X"35",X"4F",X"36",X"00",X"21",X"2A",X"4F",X"34",
		X"C9",X"DD",X"21",X"50",X"4C",X"CD",X"9C",X"BC",X"18",X"DC",X"DD",X"21",X"50",X"4C",X"FD",X"21",
		X"04",X"4D",X"21",X"52",X"4C",X"01",X"00",X"00",X"78",X"ED",X"5B",X"54",X"4C",X"BB",X"28",X"18",
		X"CD",X"6B",X"BC",X"2A",X"04",X"4D",X"CD",X"E5",X"BC",X"38",X"15",X"3A",X"35",X"4F",X"0F",X"0F",
		X"E6",X"C0",X"C6",X"00",X"32",X"2F",X"4F",X"C9",X"BA",X"28",X"05",X"CD",X"75",X"BC",X"18",X"E3",
		X"AF",X"32",X"07",X"4C",X"32",X"2F",X"4F",X"CD",X"8C",X"B6",X"C9",X"3A",X"B7",X"4D",X"A7",X"C0",
		X"3E",X"03",X"32",X"B7",X"4D",X"AF",X"32",X"2A",X"4F",X"CD",X"C3",X"BC",X"C9",X"DD",X"21",X"06",
		X"4D",X"FD",X"21",X"58",X"4C",X"CD",X"BE",X"BB",X"DD",X"21",X"42",X"4D",X"FD",X"21",X"44",X"4D",
		X"CD",X"6C",X"98",X"CD",X"F9",X"BC",X"30",X"21",X"21",X"5E",X"4C",X"CD",X"94",X"BC",X"DD",X"21",
		X"58",X"4C",X"ED",X"5B",X"42",X"4D",X"CD",X"B0",X"BC",X"2A",X"5C",X"4C",X"22",X"5A",X"4C",X"21",
		X"36",X"4F",X"36",X"00",X"21",X"2B",X"4F",X"34",X"C9",X"DD",X"21",X"58",X"4C",X"CD",X"9C",X"BC",
		X"18",X"DC",X"DD",X"21",X"58",X"4C",X"FD",X"21",X"06",X"4D",X"21",X"5A",X"4C",X"01",X"00",X"00",
		X"78",X"ED",X"5B",X"5C",X"4C",X"BB",X"28",X"18",X"CD",X"6B",X"BC",X"2A",X"06",X"4D",X"CD",X"E5",
		X"BC",X"38",X"15",X"3A",X"36",X"4F",X"0F",X"0F",X"E6",X"C0",X"C6",X"00",X"32",X"30",X"4F",X"C9",
		X"BA",X"28",X"05",X"CD",X"75",X"BC",X"18",X"E3",X"AF",X"32",X"09",X"4C",X"32",X"30",X"4F",X"CD",
		X"24",X"B7",X"C9",X"3A",X"B7",X"4D",X"A7",X"C0",X"3E",X"04",X"32",X"B7",X"4D",X"AF",X"32",X"2B",
		X"4F",X"CD",X"C3",X"BC",X"C9",X"3A",X"26",X"4F",X"47",X"3A",X"B1",X"4D",X"B0",X"47",X"3A",X"1A",
		X"4F",X"D6",X"08",X"3E",X"00",X"38",X"02",X"3E",X"01",X"B0",X"C0",X"CD",X"8D",X"0B",X"4F",X"3A",
		X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"20",X"4B",X"CB",X"61",X"28",X"01",X"37",X"3A",X"76",
		X"4E",X"17",X"E6",X"0F",X"32",X"76",X"4E",X"D6",X"0C",X"C0",X"CD",X"D5",X"BD",X"18",X"04",X"3D",
		X"32",X"23",X"4E",X"3E",X"0F",X"32",X"26",X"4F",X"3E",X"40",X"32",X"AC",X"4E",X"21",X"27",X"4F",
		X"06",X"06",X"3E",X"01",X"CF",X"21",X"B8",X"4D",X"06",X"04",X"3E",X"04",X"CF",X"3A",X"13",X"4E",
		X"A7",X"20",X"0D",X"32",X"2A",X"4F",X"32",X"BA",X"4D",X"32",X"2B",X"4F",X"32",X"BB",X"4D",X"C9",
		X"3D",X"28",X"F6",X"C9",X"79",X"17",X"3A",X"77",X"4E",X"17",X"E6",X"0F",X"32",X"77",X"4E",X"D6",
		X"0C",X"28",X"B7",X"C9",X"3A",X"2C",X"4F",X"A7",X"C2",X"DC",X"BA",X"3A",X"1A",X"4F",X"E7",X"25",
		X"B8",X"BE",X"B8",X"0C",X"B9",X"3C",X"BA",X"66",X"BA",X"78",X"BA",X"0A",X"BD",X"0E",X"BD",X"46",
		X"BD",X"7A",X"BD",X"BF",X"BD",X"3A",X"0C",X"4F",X"20",X"26",X"2A",X"0A",X"4F",X"29",X"22",X"0A",
		X"4F",X"2A",X"08",X"4F",X"ED",X"6A",X"22",X"08",X"4F",X"D0",X"21",X"0A",X"4F",X"34",X"21",X"1E",
		X"4F",X"35",X"20",X"22",X"CD",X"D9",X"BC",X"AF",X"32",X"0C",X"4F",X"21",X"1A",X"4F",X"34",X"C9",
		X"2A",X"02",X"4F",X"29",X"22",X"02",X"4F",X"2A",X"00",X"4F",X"ED",X"6A",X"22",X"00",X"4F",X"D0",
		X"21",X"02",X"4F",X"34",X"18",X"D8",X"ED",X"4B",X"44",X"4D",X"3A",X"47",X"4D",X"B8",X"28",X"D4",
		X"3A",X"0B",X"4D",X"E6",X"07",X"FE",X"04",X"20",X"1C",X"3A",X"47",X"4D",X"FE",X"27",X"38",X"37",
		X"FE",X"34",X"30",X"33",X"3A",X"3B",X"4D",X"32",X"3B",X"4D",X"47",X"21",X"0A",X"03",X"DF",X"22",
		X"2E",X"4D",X"CD",X"9E",X"BA",X"CD",X"B9",X"BA",X"21",X"1B",X"4F",X"34",X"3E",X"08",X"BE",X"D0",
		X"36",X"00",X"23",X"3A",X"3B",X"4D",X"A7",X"06",X"80",X"28",X"02",X"06",X"00",X"7E",X"3C",X"E6",
		X"01",X"80",X"77",X"CD",X"09",X"83",X"C9",X"3A",X"35",X"4D",X"EE",X"02",X"18",X"C9",X"2E",X"14",
		X"26",X"18",X"22",X"0C",X"4C",X"21",X"01",X"00",X"06",X"01",X"CD",X"CE",X"BA",X"3E",X"01",X"32",
		X"23",X"4F",X"2A",X"46",X"4D",X"22",X"1F",X"4F",X"2A",X"0A",X"4D",X"22",X"21",X"4F",X"3A",X"1D",
		X"4F",X"47",X"AF",X"CB",X"40",X"28",X"02",X"3E",X"02",X"32",X"24",X"4F",X"78",X"32",X"1E",X"4F",
		X"06",X"00",X"FE",X"10",X"30",X"02",X"06",X"80",X"78",X"32",X"25",X"4F",X"AF",X"32",X"1B",X"4F",
		X"32",X"1C",X"4F",X"3E",X"80",X"32",X"AC",X"4E",X"CD",X"4B",X"B8",X"C9",X"21",X"23",X"4F",X"3A",
		X"25",X"4F",X"CB",X"7F",X"20",X"07",X"7E",X"A7",X"CA",X"60",X"B9",X"3D",X"77",X"21",X"01",X"00",
		X"06",X"01",X"CD",X"CE",X"BA",X"3A",X"0A",X"4D",X"E6",X"07",X"FE",X"04",X"20",X"1E",X"3A",X"46",
		X"4D",X"47",X"3A",X"44",X"4D",X"90",X"38",X"20",X"FE",X"08",X"30",X"0D",X"3A",X"46",X"4D",X"FE",
		X"25",X"38",X"06",X"EF",X"17",X"00",X"CD",X"4B",X"B8",X"CD",X"9E",X"BA",X"CD",X"B9",X"BA",X"3A",
		X"37",X"4F",X"E6",X"03",X"32",X"1C",X"4F",X"C9",X"3E",X"04",X"32",X"1A",X"4F",X"C3",X"8A",X"BA",
		X"3A",X"25",X"4F",X"A7",X"20",X"75",X"34",X"21",X"00",X"FF",X"06",X"00",X"3A",X"24",X"4F",X"A7",
		X"28",X"09",X"FE",X"03",X"28",X"05",X"21",X"00",X"01",X"06",X"02",X"CD",X"CE",X"BA",X"3A",X"24",
		X"4F",X"0F",X"30",X"27",X"3A",X"0B",X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"4C",X"B9",X"3A",X"47",
		X"4D",X"47",X"3A",X"20",X"4F",X"90",X"C2",X"49",X"B9",X"3A",X"1D",X"4F",X"32",X"1E",X"4F",X"3A",
		X"24",X"4F",X"3C",X"E6",X"03",X"32",X"24",X"4F",X"C3",X"49",X"B9",X"21",X"1E",X"4F",X"35",X"3E",
		X"08",X"BE",X"30",X"10",X"3A",X"47",X"4D",X"FE",X"25",X"38",X"04",X"FE",X"37",X"38",X"0F",X"3E",
		X"08",X"32",X"1E",X"4F",X"3E",X"01",X"32",X"25",X"4F",X"3E",X"02",X"32",X"23",X"4F",X"3A",X"0B",
		X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"4C",X"B9",X"C3",X"49",X"B9",X"CB",X"77",X"20",X"35",X"3C",
		X"32",X"25",X"4F",X"3C",X"E6",X"1F",X"32",X"23",X"4F",X"FE",X"08",X"38",X"0E",X"CB",X"F7",X"32",
		X"25",X"4F",X"3A",X"24",X"4F",X"3C",X"E6",X"03",X"32",X"24",X"4F",X"21",X"00",X"FF",X"06",X"00",
		X"3A",X"24",X"4F",X"A7",X"28",X"09",X"FE",X"03",X"28",X"05",X"21",X"00",X"01",X"06",X"02",X"CD",
		X"CE",X"BA",X"18",X"BA",X"21",X"25",X"4F",X"3E",X"1F",X"A6",X"32",X"23",X"4F",X"35",X"3D",X"20",
		X"01",X"77",X"21",X"00",X"FF",X"06",X"00",X"3A",X"24",X"4F",X"A7",X"28",X"09",X"FE",X"03",X"28",
		X"05",X"21",X"00",X"01",X"06",X"02",X"CD",X"CE",X"BA",X"C3",X"84",X"B9",X"3A",X"0A",X"4D",X"E6",
		X"07",X"FE",X"04",X"C2",X"4C",X"B9",X"3A",X"46",X"4D",X"47",X"3A",X"44",X"4D",X"90",X"30",X"03",
		X"CD",X"4B",X"B8",X"3A",X"47",X"4D",X"FE",X"25",X"38",X"05",X"FE",X"37",X"DA",X"49",X"B9",X"3E",
		X"05",X"32",X"1A",X"4F",X"18",X"12",X"3A",X"25",X"4F",X"CB",X"7F",X"20",X"0B",X"A7",X"CA",X"60",
		X"B9",X"3A",X"23",X"4F",X"3D",X"32",X"23",X"4F",X"21",X"01",X"00",X"06",X"01",X"CD",X"CE",X"BA",
		X"3A",X"0A",X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"4C",X"B9",X"3A",X"46",X"4D",X"FE",X"3E",X"30",
		X"03",X"C3",X"49",X"B9",X"3E",X"06",X"32",X"1A",X"4F",X"AF",X"32",X"EB",X"4D",X"C9",X"DD",X"21",
		X"2E",X"4D",X"FD",X"21",X"16",X"4D",X"CD",X"47",X"91",X"22",X"16",X"4D",X"2A",X"2E",X"4D",X"22",
		X"22",X"4D",X"3A",X"3B",X"4D",X"32",X"35",X"4D",X"C9",X"DD",X"21",X"22",X"4D",X"FD",X"21",X"0A",
		X"4D",X"CD",X"47",X"91",X"22",X"0A",X"4D",X"CD",X"5F",X"91",X"22",X"46",X"4D",X"C9",X"22",X"22",
		X"4D",X"22",X"2E",X"4D",X"78",X"32",X"35",X"4D",X"32",X"3B",X"4D",X"C9",X"E7",X"44",X"B0",X"E5",
		X"BA",X"2A",X"BB",X"94",X"BB",X"DD",X"21",X"0A",X"4D",X"FD",X"21",X"60",X"4C",X"CD",X"BE",X"BB",
		X"DD",X"21",X"46",X"4D",X"FD",X"21",X"44",X"4D",X"CD",X"6C",X"98",X"CD",X"F9",X"BC",X"30",X"21",
		X"21",X"66",X"4C",X"CD",X"94",X"BC",X"DD",X"21",X"60",X"4C",X"ED",X"5B",X"46",X"4D",X"CD",X"B0",
		X"BC",X"2A",X"64",X"4C",X"22",X"62",X"4C",X"21",X"37",X"4F",X"36",X"00",X"21",X"2C",X"4F",X"34",
		X"C9",X"DD",X"21",X"60",X"4C",X"CD",X"9C",X"BC",X"18",X"DC",X"DD",X"21",X"60",X"4C",X"FD",X"21",
		X"0A",X"4D",X"21",X"62",X"4C",X"01",X"00",X"00",X"78",X"ED",X"5B",X"64",X"4C",X"BB",X"28",X"18",
		X"CD",X"6B",X"BC",X"2A",X"0A",X"4D",X"CD",X"E5",X"BC",X"38",X"15",X"3A",X"37",X"4F",X"0F",X"0F",
		X"E6",X"C0",X"C6",X"14",X"32",X"32",X"4F",X"C9",X"BA",X"28",X"05",X"CD",X"75",X"BC",X"18",X"E3",
		X"21",X"00",X"00",X"22",X"0C",X"4C",X"21",X"0C",X"AC",X"22",X"0A",X"4D",X"21",X"21",X"33",X"22",
		X"16",X"4D",X"22",X"46",X"4D",X"21",X"00",X"FF",X"22",X"22",X"4D",X"22",X"2E",X"4D",X"3E",X"00",
		X"32",X"35",X"4D",X"32",X"3B",X"4D",X"AF",X"32",X"32",X"4F",X"32",X"1B",X"4F",X"32",X"1C",X"4F",
		X"CD",X"1C",X"BB",X"C9",X"21",X"1B",X"4F",X"34",X"3E",X"08",X"BE",X"D8",X"36",X"00",X"CD",X"D9",
		X"BC",X"2E",X"80",X"26",X"1C",X"22",X"0C",X"4C",X"CD",X"09",X"83",X"AF",X"32",X"1A",X"4F",X"32",
		X"2C",X"4F",X"CD",X"C3",X"BC",X"C9",X"01",X"01",X"01",X"FF",X"FF",X"01",X"FF",X"FF",X"21",X"08",
		X"4D",X"DD",X"7E",X"00",X"96",X"FD",X"36",X"00",X"00",X"30",X"08",X"7E",X"DD",X"96",X"00",X"FD",
		X"36",X"00",X"01",X"FD",X"77",X"02",X"23",X"DD",X"7E",X"01",X"96",X"FD",X"36",X"01",X"00",X"30",
		X"08",X"7E",X"DD",X"96",X"01",X"FD",X"36",X"01",X"01",X"FD",X"77",X"03",X"FD",X"7E",X"01",X"1F",
		X"FD",X"7E",X"00",X"17",X"FD",X"77",X"00",X"21",X"B6",X"BB",X"47",X"DF",X"FD",X"75",X"06",X"FD",
		X"74",X"07",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"7D",X"2C",X"A7",X"28",X"01",X"6F",X"7C",X"24",
		X"A7",X"28",X"01",X"67",X"7D",X"94",X"20",X"09",X"FD",X"36",X"04",X"01",X"FD",X"36",X"05",X"01",
		X"C9",X"38",X"10",X"7C",X"65",X"6F",X"CD",X"52",X"BC",X"7D",X"A7",X"20",X"15",X"FD",X"6E",X"02",
		X"FD",X"66",X"03",X"CD",X"52",X"BC",X"7D",X"A7",X"20",X"10",X"FD",X"66",X"02",X"FD",X"6E",X"03",
		X"18",X"E4",X"FD",X"36",X"04",X"01",X"FD",X"75",X"05",X"C9",X"FD",X"75",X"04",X"FD",X"36",X"05",
		X"01",X"C9",X"F5",X"C5",X"7D",X"6C",X"ED",X"44",X"4F",X"26",X"00",X"06",X"09",X"7C",X"81",X"30",
		X"01",X"67",X"ED",X"6A",X"10",X"F7",X"CB",X"3C",X"C1",X"F1",X"C9",X"35",X"20",X"03",X"73",X"06",
		X"01",X"23",X"BA",X"28",X"06",X"35",X"20",X"03",X"72",X"0E",X"01",X"B8",X"28",X"09",X"DD",X"7E",
		X"06",X"FD",X"86",X"00",X"FD",X"77",X"00",X"79",X"A7",X"C8",X"DD",X"7E",X"07",X"FD",X"86",X"01",
		X"FD",X"77",X"01",X"C9",X"7E",X"87",X"77",X"23",X"7E",X"87",X"77",X"C9",X"78",X"A7",X"C8",X"DD",
		X"7E",X"04",X"87",X"DD",X"77",X"04",X"DD",X"7E",X"05",X"87",X"DD",X"77",X"05",X"10",X"F0",X"C9",
		X"2A",X"44",X"4D",X"7D",X"BB",X"20",X"04",X"DD",X"36",X"04",X"00",X"7C",X"BA",X"C0",X"DD",X"36",
		X"05",X"00",X"C9",X"21",X"28",X"4F",X"06",X"04",X"7E",X"23",X"B6",X"10",X"FC",X"A7",X"C0",X"21",
		X"AC",X"4E",X"CB",X"B6",X"F7",X"02",X"0C",X"00",X"C9",X"3A",X"8E",X"4C",X"E6",X"3F",X"32",X"1D",
		X"4F",X"32",X"1E",X"4F",X"C9",X"7D",X"FE",X"11",X"D8",X"FE",X"F0",X"30",X"0A",X"7C",X"FE",X"11",
		X"D8",X"FE",X"F0",X"30",X"02",X"AF",X"C9",X"37",X"C9",X"06",X"03",X"7C",X"A7",X"C0",X"7D",X"05",
		X"FE",X"40",X"D0",X"05",X"FE",X"10",X"D0",X"FE",X"08",X"C9",X"CD",X"4B",X"B8",X"C9",X"2E",X"00",
		X"26",X"1C",X"22",X"0C",X"4C",X"3A",X"3B",X"4D",X"E6",X"02",X"21",X"00",X"FF",X"06",X"00",X"28",
		X"05",X"21",X"00",X"01",X"06",X"02",X"CD",X"CE",X"BA",X"2A",X"1F",X"4F",X"22",X"16",X"4D",X"22",
		X"46",X"4D",X"2A",X"21",X"4F",X"22",X"0A",X"4D",X"CD",X"D9",X"BC",X"AF",X"32",X"1A",X"4F",X"32",
		X"1B",X"4F",X"32",X"1C",X"4F",X"C9",X"3A",X"33",X"4E",X"A7",X"28",X"0E",X"AF",X"32",X"33",X"4E",
		X"CD",X"6E",X"0B",X"21",X"EC",X"4E",X"CB",X"8E",X"18",X"B4",X"32",X"CC",X"4E",X"32",X"AC",X"4E",
		X"32",X"EB",X"4D",X"32",X"40",X"4F",X"3E",X"08",X"32",X"AC",X"4E",X"21",X"A4",X"0F",X"11",X"0A",
		X"4C",X"01",X"04",X"00",X"ED",X"B0",X"CD",X"4B",X"B8",X"C9",X"3A",X"40",X"4F",X"3C",X"47",X"11",
		X"C4",X"0F",X"CD",X"45",X"82",X"C0",X"21",X"40",X"4F",X"34",X"7E",X"FE",X"08",X"30",X"14",X"87",
		X"87",X"21",X"A4",X"0F",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"11",X"0A",X"4C",X"01",X"04",X"00",
		X"ED",X"B0",X"C9",X"36",X"00",X"3E",X"05",X"32",X"B1",X"4D",X"3E",X"1A",X"4F",X"CD",X"B8",X"90",
		X"28",X"04",X"3E",X"C0",X"A9",X"4F",X"69",X"26",X"1C",X"22",X"0A",X"4C",X"C3",X"0E",X"BD",X"3E",
		X"05",X"32",X"B1",X"4D",X"C9",X"3A",X"1A",X"4F",X"D6",X"09",X"0E",X"00",X"38",X"02",X"0E",X"0F",
		X"3A",X"B1",X"4D",X"B1",X"C9",X"2A",X"3B",X"4F",X"22",X"3D",X"4F",X"3E",X"0F",X"32",X"3F",X"4F",
		X"0E",X"04",X"CD",X"E5",X"0A",X"0E",X"05",X"CD",X"E5",X"0A",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
