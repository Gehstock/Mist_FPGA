library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_D7 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(8 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_D7 is
	type rom is array(0 to  511) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"00",X"10",
		X"00",X"60",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"30",X"30",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E1",X"F1",X"F1",X"F0",X"F0",X"60",X"60",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"F1",X"F1",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C1",X"F3",X"F3",X"F1",X"F0",X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C3",X"F7",X"F7",X"F3",X"F1",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F1",X"F7",X"F7",X"F7",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F1",X"F3",X"F7",X"F7",X"C3",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"F1",X"F3",X"F3",X"C1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"F0",X"F0",X"F1",X"F1",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"60",X"F0",X"F0",X"F1",X"F1",X"E1",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"60",
		X"00",X"10",X"00",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",
		X"00",X"30",X"70",X"30",X"30",X"20",X"20",X"30",X"30",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"20",X"60",X"F0",X"30",X"30",X"30",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"81",X"C3",X"F0",X"50",X"60",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"E7",X"F1",X"C0",X"60",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"F7",X"97",X"C5",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F5",X"C7",X"F5",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"C5",X"97",X"F7",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"C0",X"F1",X"E7",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"60",X"50",X"F0",X"C3",X"81",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"30",X"30",X"F0",X"60",X"20",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"30",X"20",X"20",X"30",X"30",X"70",X"30",
		X"00",X"00",X"40",X"80",X"21",X"00",X"12",X"00",X"29",X"00",X"20",X"04",X"40",X"01",X"00",X"20",
		X"20",X"00",X"41",X"10",X"84",X"10",X"44",X"00",X"40",X"24",X"12",X"80",X"01",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
