library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sbagman_program2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sbagman_program2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"82",X"C3",X"C3",X"93",X"C3",X"31",X"F0",X"67",X"3E",X"3F",X"CD",X"A3",X"C3",X"CD",X"B7",
		X"C3",X"3E",X"01",X"32",X"03",X"A0",X"21",X"8C",X"1A",X"11",X"17",X"62",X"01",X"50",X"00",X"ED",
		X"B0",X"21",X"68",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"C3",X"C1",X"EC",X"3A",X"10",
		X"62",X"FE",X"01",X"20",X"3E",X"3A",X"6D",X"62",X"FE",X"20",X"DC",X"47",X"C0",X"FE",X"30",X"DC",
		X"7C",X"C0",X"AF",X"32",X"6D",X"62",X"C9",X"3A",X"6E",X"62",X"FE",X"01",X"28",X"13",X"CD",X"8B",
		X"C0",X"28",X"10",X"11",X"5A",X"57",X"CD",X"67",X"CA",X"CD",X"73",X"C0",X"3E",X"01",X"32",X"6E",
		X"62",X"F1",X"C9",X"11",X"63",X"57",X"CD",X"67",X"CA",X"CD",X"73",X"C0",X"3E",X"01",X"32",X"6E",
		X"62",X"F1",X"C9",X"3E",X"02",X"21",X"40",X"98",X"CD",X"05",X"56",X"C9",X"CD",X"8B",X"C0",X"11",
		X"6C",X"57",X"CD",X"67",X"CA",X"AF",X"32",X"6E",X"62",X"F1",X"C9",X"3A",X"7C",X"61",X"21",X"A0",
		X"93",X"FE",X"01",X"C0",X"21",X"20",X"91",X"C9",X"2B",X"F3",X"CD",X"F3",X"C0",X"23",X"CD",X"F3",
		X"C0",X"0A",X"FB",X"C9",X"C5",X"E5",X"D5",X"AF",X"32",X"0B",X"60",X"11",X"D5",X"35",X"ED",X"52",
		X"20",X"0A",X"CD",X"DF",X"C0",X"28",X"05",X"3E",X"02",X"32",X"0B",X"60",X"D1",X"E1",X"C1",X"C9",
		X"C5",X"E5",X"D5",X"AF",X"32",X"0B",X"60",X"11",X"15",X"36",X"ED",X"52",X"20",X"0A",X"CD",X"DF",
		X"C0",X"28",X"05",X"3E",X"02",X"32",X"0B",X"60",X"D1",X"E1",X"C1",X"C9",X"D1",X"18",X"F9",X"3A",
		X"0D",X"60",X"FE",X"05",X"20",X"F6",X"21",X"F3",X"91",X"7E",X"21",X"DB",X"19",X"01",X"05",X"00",
		X"ED",X"B1",X"C9",X"7E",X"FE",X"51",X"28",X"15",X"FD",X"21",X"12",X"1A",X"11",X"E0",X"19",X"C5",
		X"4F",X"06",X"08",X"1A",X"B9",X"28",X"14",X"13",X"FD",X"23",X"10",X"F7",X"C1",X"03",X"0A",X"3C",
		X"02",X"0B",X"FE",X"03",X"D8",X"AF",X"03",X"02",X"0B",X"02",X"C9",X"C1",X"FD",X"7E",X"00",X"DD",
		X"77",X"03",X"3E",X"01",X"02",X"03",X"AF",X"02",X"0B",X"C9",X"7E",X"FE",X"FF",X"C8",X"CD",X"6D",
		X"C1",X"78",X"32",X"0C",X"60",X"FE",X"00",X"C8",X"FD",X"7E",X"00",X"FE",X"01",X"C8",X"7E",X"FE",
		X"51",X"28",X"0C",X"4F",X"11",X"E8",X"19",X"06",X"30",X"1A",X"B9",X"C8",X"13",X"10",X"FA",X"3A",
		X"0C",X"60",X"FE",X"05",X"30",X"09",X"47",X"DD",X"7E",X"03",X"90",X"DD",X"77",X"03",X"C9",X"2F",
		X"E6",X"07",X"C6",X"01",X"47",X"DD",X"7E",X"03",X"80",X"DD",X"77",X"03",X"C9",X"DD",X"7E",X"03",
		X"CB",X"07",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"06",X"00",X"CB",X"07",X"CB",X"10",
		X"CB",X"07",X"CB",X"10",X"CB",X"07",X"CB",X"10",X"C9",X"CD",X"CD",X"C3",X"3E",X"3F",X"CD",X"A3",
		X"C3",X"3A",X"00",X"B8",X"21",X"00",X"34",X"11",X"00",X"90",X"01",X"00",X"04",X"ED",X"B0",X"21",
		X"82",X"98",X"06",X"06",X"CD",X"61",X"C3",X"CD",X"4D",X"CE",X"CD",X"DD",X"D0",X"CD",X"0E",X"C3",
		X"3A",X"00",X"B8",X"CD",X"DE",X"F8",X"CD",X"7E",X"CA",X"CD",X"F3",X"D0",X"3E",X"63",X"D3",X"58",
		X"C9",X"CD",X"CD",X"C3",X"3E",X"3F",X"CD",X"A3",X"C3",X"3A",X"00",X"B8",X"21",X"00",X"30",X"11",
		X"00",X"90",X"01",X"00",X"04",X"ED",X"B0",X"21",X"02",X"93",X"CD",X"38",X"C3",X"21",X"62",X"98",
		X"06",X"0E",X"CD",X"61",X"C3",X"21",X"1A",X"99",X"06",X"16",X"CD",X"6E",X"C3",X"3E",X"3F",X"32",
		X"57",X"9B",X"CD",X"DD",X"D0",X"21",X"84",X"65",X"3E",X"33",X"77",X"23",X"3E",X"04",X"77",X"23",
		X"3E",X"BF",X"77",X"23",X"3A",X"00",X"B8",X"CD",X"DE",X"F8",X"CD",X"7E",X"CA",X"C9",X"CD",X"CD",
		X"C3",X"3E",X"3F",X"CD",X"A3",X"C3",X"3A",X"00",X"B8",X"21",X"00",X"48",X"11",X"00",X"90",X"01",
		X"00",X"04",X"ED",X"B0",X"21",X"62",X"93",X"CD",X"38",X"C3",X"21",X"42",X"98",X"06",X"0F",X"CD",
		X"61",X"C3",X"21",X"FA",X"98",X"06",X"16",X"CD",X"6E",X"C3",X"21",X"5A",X"98",X"06",X"02",X"CD",
		X"6E",X"C3",X"3E",X"3F",X"32",X"77",X"9A",X"CD",X"DD",X"D0",X"3A",X"00",X"B8",X"3A",X"00",X"B0",
		X"E6",X"20",X"FE",X"20",X"20",X"0F",X"21",X"32",X"92",X"3E",X"34",X"06",X"06",X"77",X"11",X"20",
		X"00",X"19",X"3C",X"10",X"F8",X"CD",X"0E",X"C3",X"CD",X"DE",X"F8",X"CD",X"7E",X"CA",X"CD",X"F3",
		X"D0",X"C9",X"CD",X"CD",X"C3",X"3E",X"3F",X"CD",X"A3",X"C3",X"3A",X"00",X"B8",X"21",X"00",X"44",
		X"11",X"00",X"90",X"01",X"00",X"04",X"ED",X"B0",X"21",X"82",X"91",X"CD",X"38",X"C3",X"21",X"82",
		X"98",X"06",X"07",X"CD",X"61",X"C3",X"21",X"A2",X"9A",X"06",X"09",X"CD",X"61",X"C3",X"3E",X"BE",
		X"32",X"0E",X"93",X"3C",X"32",X"0F",X"93",X"3E",X"24",X"21",X"2C",X"9B",X"11",X"1E",X"00",X"06",
		X"03",X"77",X"23",X"77",X"23",X"77",X"19",X"10",X"F8",X"CD",X"DD",X"D0",X"3A",X"00",X"B8",X"CD",
		X"0E",X"C3",X"CD",X"DE",X"F8",X"CD",X"7E",X"CA",X"C9",X"CD",X"CD",X"C3",X"3E",X"3F",X"CD",X"A3",
		X"C3",X"3A",X"00",X"B8",X"21",X"00",X"40",X"11",X"00",X"90",X"01",X"00",X"04",X"ED",X"B0",X"21",
		X"82",X"91",X"CD",X"38",X"C3",X"21",X"42",X"98",X"06",X"07",X"CD",X"61",X"C3",X"21",X"C2",X"9A",
		X"06",X"07",X"CD",X"61",X"C3",X"CD",X"DD",X"D0",X"3A",X"00",X"B8",X"CD",X"0E",X"C3",X"CD",X"DE",
		X"F8",X"CD",X"7E",X"CA",X"3A",X"10",X"62",X"FE",X"00",X"C8",X"CD",X"F3",X"D0",X"C9",X"21",X"86",
		X"65",X"AF",X"77",X"C9",X"3E",X"01",X"32",X"1A",X"60",X"32",X"1B",X"60",X"3E",X"80",X"32",X"27",
		X"60",X"3E",X"40",X"32",X"67",X"60",X"21",X"1B",X"1A",X"3A",X"00",X"B8",X"11",X"88",X"65",X"01",
		X"14",X"00",X"ED",X"B0",X"CD",X"A3",X"F9",X"C9",X"3E",X"55",X"77",X"23",X"3E",X"51",X"77",X"23",
		X"3E",X"57",X"77",X"11",X"1F",X"00",X"19",X"3E",X"52",X"77",X"2B",X"3E",X"56",X"77",X"7C",X"C6",
		X"08",X"67",X"3E",X"32",X"77",X"23",X"77",X"11",X"E1",X"FF",X"19",X"77",X"2B",X"77",X"2B",X"77",
		X"C9",X"3E",X"38",X"18",X"01",X"C9",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"C9",X"3E",X"2F",
		X"18",X"F4",X"C9",X"C5",X"01",X"E0",X"FF",X"77",X"09",X"C1",X"10",X"F7",X"C9",X"77",X"23",X"10",
		X"FC",X"C9",X"06",X"08",X"21",X"00",X"60",X"AF",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",
		X"C3",X"03",X"C0",X"06",X"08",X"21",X"00",X"60",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",
		X"C3",X"06",X"C0",X"06",X"08",X"21",X"00",X"98",X"0E",X"00",X"77",X"23",X"F5",X"3A",X"00",X"B8",
		X"F1",X"0D",X"20",X"F6",X"10",X"F2",X"C9",X"06",X"04",X"3E",X"E0",X"21",X"00",X"90",X"0E",X"00",
		X"77",X"23",X"F5",X"3A",X"00",X"B8",X"F1",X"0D",X"20",X"F6",X"10",X"F2",X"C9",X"3E",X"E0",X"3E",
		X"E0",X"21",X"E4",X"93",X"06",X"1B",X"E5",X"C5",X"06",X"20",X"CD",X"73",X"C3",X"C1",X"E1",X"23",
		X"10",X"F4",X"C9",X"3E",X"00",X"32",X"03",X"A0",X"06",X"04",X"3E",X"E0",X"21",X"00",X"90",X"CD",
		X"BE",X"C3",X"3E",X"3F",X"CD",X"A3",X"C3",X"3A",X"8C",X"62",X"FE",X"01",X"28",X"09",X"11",X"C3",
		X"56",X"21",X"AF",X"93",X"CD",X"67",X"CA",X"06",X"01",X"21",X"80",X"65",X"3E",X"00",X"CD",X"A8",
		X"C3",X"CD",X"7E",X"CA",X"3E",X"01",X"32",X"03",X"A0",X"C9",X"DD",X"21",X"76",X"61",X"06",X"07",
		X"AF",X"00",X"DD",X"23",X"10",X"FB",X"C9",X"3A",X"63",X"61",X"E6",X"80",X"FE",X"00",X"28",X"09",
		X"3A",X"7C",X"61",X"2F",X"E6",X"01",X"CD",X"E2",X"D8",X"DD",X"21",X"9C",X"60",X"FD",X"21",X"7F",
		X"61",X"06",X"3B",X"CD",X"7E",X"C4",X"DD",X"21",X"C4",X"61",X"FD",X"21",X"FA",X"61",X"06",X"03",
		X"CD",X"7E",X"C4",X"3A",X"56",X"60",X"F5",X"3A",X"7E",X"61",X"32",X"56",X"60",X"F1",X"32",X"7E",
		X"61",X"3A",X"90",X"62",X"F5",X"3A",X"7D",X"62",X"32",X"90",X"62",X"F1",X"32",X"7D",X"62",X"3A",
		X"41",X"63",X"F5",X"3A",X"40",X"63",X"32",X"41",X"63",X"F1",X"32",X"40",X"63",X"C9",X"DD",X"7E",
		X"00",X"F5",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"F1",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",
		X"10",X"EC",X"C9",X"0E",X"0B",X"06",X"07",X"DD",X"7E",X"03",X"C6",X"03",X"91",X"FD",X"BE",X"03",
		X"28",X"06",X"0C",X"10",X"F2",X"3E",X"00",X"C9",X"DD",X"7E",X"02",X"C6",X"08",X"FD",X"BE",X"02",
		X"38",X"F3",X"D6",X"0F",X"FD",X"BE",X"02",X"30",X"EC",X"3E",X"01",X"C9",X"3A",X"98",X"60",X"FE",
		X"05",X"CA",X"B7",X"D9",X"47",X"3A",X"0D",X"60",X"B8",X"C2",X"CB",X"C5",X"E5",X"FD",X"E5",X"FD",
		X"21",X"D1",X"1B",X"FD",X"7E",X"00",X"67",X"FD",X"7E",X"01",X"6F",X"AF",X"ED",X"52",X"28",X"18",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"7E",X"02",X"FE",X"FF",X"20",X"E6",X"2A",X"46",X"61",
		X"AF",X"77",X"FD",X"E1",X"E1",X"C3",X"5A",X"C5",X"3E",X"01",X"2A",X"46",X"61",X"7E",X"FE",X"00",
		X"C2",X"F2",X"C4",X"CD",X"97",X"C5",X"FD",X"E1",X"47",X"FD",X"7E",X"03",X"B8",X"CA",X"8C",X"C5",
		X"2A",X"46",X"61",X"23",X"23",X"23",X"23",X"3E",X"01",X"77",X"E1",X"D5",X"11",X"1C",X"00",X"19",
		X"D1",X"AF",X"77",X"DD",X"7E",X"07",X"3D",X"FD",X"BE",X"03",X"28",X"0C",X"3D",X"FD",X"BE",X"03",
		X"28",X"06",X"2A",X"95",X"60",X"AF",X"77",X"C9",X"3A",X"98",X"60",X"FE",X"05",X"C8",X"2A",X"46",
		X"61",X"23",X"23",X"23",X"23",X"AF",X"77",X"DD",X"7E",X"06",X"2A",X"95",X"60",X"FD",X"BE",X"02",
		X"30",X"04",X"3E",X"40",X"77",X"C9",X"3E",X"80",X"77",X"C9",X"7E",X"FE",X"01",X"28",X"09",X"2A",
		X"46",X"61",X"23",X"23",X"23",X"23",X"77",X"C9",X"2A",X"46",X"61",X"3E",X"01",X"77",X"CD",X"97",
		X"C5",X"47",X"FD",X"7E",X"03",X"B8",X"28",X"15",X"23",X"23",X"23",X"23",X"3E",X"01",X"77",X"3E",
		X"C0",X"FD",X"77",X"02",X"18",X"00",X"2A",X"95",X"60",X"AF",X"77",X"C9",X"E1",X"2A",X"46",X"61",
		X"23",X"23",X"23",X"23",X"AF",X"77",X"C9",X"3A",X"99",X"99",X"3A",X"98",X"60",X"FE",X"04",X"28",
		X"03",X"FE",X"05",X"C8",X"DD",X"7E",X"02",X"FE",X"C0",X"06",X"80",X"30",X"02",X"06",X"40",X"DD",
		X"7E",X"03",X"FE",X"68",X"3E",X"18",X"38",X"0C",X"DD",X"7E",X"03",X"FE",X"C0",X"3E",X"71",X"38",
		X"03",X"3E",X"E1",X"C9",X"E5",X"2A",X"95",X"60",X"70",X"E1",X"C9",X"2A",X"46",X"61",X"23",X"23",
		X"23",X"23",X"AF",X"77",X"C9",X"21",X"00",X"05",X"FB",X"06",X"FF",X"3A",X"00",X"60",X"FE",X"00",
		X"C0",X"3A",X"00",X"B8",X"FB",X"10",X"F4",X"2B",X"7C",X"FE",X"00",X"C8",X"18",X"EB",X"3A",X"ED",
		X"61",X"FE",X"01",X"3E",X"00",X"28",X"22",X"3A",X"78",X"61",X"47",X"3A",X"7C",X"61",X"FE",X"01",
		X"20",X"04",X"3A",X"7B",X"61",X"47",X"3A",X"00",X"B0",X"CB",X"1F",X"CB",X"1F",X"CB",X"1F",X"2F",
		X"E6",X"03",X"80",X"06",X"00",X"CD",X"1D",X"C6",X"78",X"32",X"64",X"61",X"C9",X"FE",X"01",X"D8",
		X"06",X"02",X"FE",X"02",X"D8",X"06",X"04",X"FE",X"03",X"D8",X"06",X"05",X"FE",X"04",X"D8",X"06",
		X"09",X"FE",X"05",X"D8",X"06",X"0A",X"C9",X"DD",X"21",X"94",X"65",X"FD",X"21",X"9C",X"65",X"CD",
		X"93",X"C4",X"FE",X"01",X"20",X"0F",X"3A",X"58",X"61",X"FE",X"01",X"28",X"08",X"3E",X"01",X"32",
		X"37",X"60",X"32",X"08",X"62",X"DD",X"21",X"98",X"65",X"FD",X"21",X"9C",X"65",X"CD",X"93",X"C4",
		X"FE",X"01",X"20",X"0F",X"3A",X"58",X"61",X"FE",X"01",X"28",X"08",X"3E",X"01",X"32",X"77",X"60",
		X"32",X"09",X"62",X"C9",X"3A",X"10",X"62",X"FE",X"01",X"C0",X"FD",X"21",X"76",X"61",X"CD",X"46",
		X"C7",X"78",X"FE",X"05",X"38",X"0B",X"FD",X"21",X"79",X"61",X"CD",X"46",X"C7",X"78",X"FE",X"05",
		X"D0",X"CD",X"98",X"FB",X"CD",X"69",X"C9",X"3A",X"6C",X"62",X"FE",X"01",X"CC",X"27",X"C4",X"CD",
		X"FB",X"C8",X"3E",X"01",X"CD",X"E2",X"D8",X"FD",X"21",X"76",X"61",X"CD",X"46",X"C7",X"78",X"FE",
		X"05",X"D2",X"DF",X"C6",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"D5",X"11",X"F0",X"FF",X"DD",X"19",
		X"D1",X"DD",X"E5",X"23",X"23",X"E5",X"CD",X"72",X"C7",X"3E",X"60",X"32",X"E8",X"61",X"E1",X"CD",
		X"FB",X"C8",X"DD",X"E1",X"3E",X"01",X"32",X"79",X"62",X"CD",X"C6",X"C7",X"CD",X"FB",X"C8",X"3A",
		X"7D",X"61",X"FE",X"01",X"28",X"58",X"3A",X"00",X"B0",X"E6",X"80",X"FE",X"80",X"28",X"05",X"3E",
		X"00",X"CD",X"E2",X"D8",X"3A",X"26",X"60",X"E6",X"80",X"FE",X"80",X"28",X"F7",X"FD",X"21",X"79",
		X"61",X"CD",X"46",X"C7",X"78",X"FE",X"05",X"30",X"35",X"CD",X"FB",X"C8",X"DD",X"23",X"DD",X"23",
		X"DD",X"23",X"D5",X"11",X"F0",X"FF",X"DD",X"19",X"D1",X"DD",X"E5",X"23",X"23",X"E5",X"CD",X"72",
		X"C7",X"3E",X"60",X"32",X"E8",X"61",X"E1",X"CD",X"FB",X"C8",X"DD",X"E1",X"3E",X"00",X"32",X"79",
		X"62",X"CD",X"87",X"C8",X"CD",X"87",X"C8",X"CD",X"87",X"C8",X"CD",X"C6",X"C7",X"C9",X"AF",X"32",
		X"67",X"62",X"32",X"03",X"A0",X"C9",X"DD",X"21",X"17",X"62",X"11",X"10",X"00",X"21",X"0F",X"92",
		X"06",X"05",X"FD",X"7E",X"02",X"DD",X"BE",X"02",X"D8",X"20",X"10",X"FD",X"7E",X"01",X"DD",X"BE",
		X"01",X"D8",X"20",X"07",X"FD",X"7E",X"00",X"DD",X"BE",X"00",X"D8",X"DD",X"19",X"2B",X"2B",X"10",
		X"E1",X"C9",X"C5",X"DD",X"21",X"17",X"62",X"78",X"FE",X"04",X"30",X"11",X"C5",X"06",X"10",X"DD",
		X"7E",X"10",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F6",X"C1",X"04",X"18",X"EA",X"C1",X"DD",X"21",
		X"17",X"62",X"78",X"FE",X"04",X"30",X"05",X"DD",X"19",X"04",X"18",X"F6",X"FD",X"7E",X"00",X"DD",
		X"77",X"00",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"FD",X"7E",X"02",X"DD",X"77",X"02",X"C5",X"06",
		X"0D",X"DD",X"E5",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"3E",X"10",X"DD",X"77",X"00",X"DD",X"23",
		X"10",X"F9",X"DD",X"E1",X"C1",X"C9",X"06",X"11",X"3E",X"00",X"32",X"78",X"62",X"3A",X"79",X"62",
		X"FE",X"01",X"20",X"05",X"CD",X"0A",X"CA",X"18",X"0C",X"3A",X"00",X"B0",X"E6",X"80",X"FE",X"80",
		X"28",X"F2",X"CD",X"26",X"CA",X"3A",X"78",X"62",X"E6",X"10",X"FE",X"10",X"CC",X"20",X"C8",X"3A",
		X"78",X"62",X"E6",X"08",X"FE",X"08",X"CC",X"2F",X"C8",X"3A",X"78",X"62",X"E6",X"40",X"FE",X"40",
		X"CC",X"3E",X"C8",X"3A",X"78",X"62",X"E6",X"20",X"FE",X"20",X"CC",X"5C",X"C8",X"3A",X"78",X"62",
		X"E6",X"80",X"FE",X"80",X"C8",X"3A",X"E8",X"61",X"FE",X"00",X"C8",X"CD",X"78",X"C8",X"18",X"AD",
		X"78",X"FE",X"2A",X"20",X"02",X"06",X"10",X"04",X"CD",X"78",X"C8",X"CD",X"87",X"C8",X"C9",X"78",
		X"FE",X"10",X"20",X"02",X"06",X"2B",X"05",X"CD",X"78",X"C8",X"CD",X"87",X"C8",X"C9",X"7D",X"E6",
		X"F0",X"FE",X"00",X"20",X"04",X"7C",X"FE",X"92",X"C8",X"06",X"10",X"CD",X"78",X"C8",X"11",X"20",
		X"00",X"19",X"DD",X"2B",X"46",X"CD",X"78",X"C8",X"CD",X"87",X"C8",X"C9",X"7D",X"E6",X"F0",X"FE",
		X"C0",X"20",X"04",X"7C",X"FE",X"91",X"C8",X"11",X"20",X"00",X"AF",X"ED",X"52",X"DD",X"23",X"06",
		X"11",X"CD",X"78",X"C8",X"CD",X"87",X"C8",X"C9",X"78",X"DD",X"77",X"00",X"77",X"E5",X"7C",X"C6",
		X"08",X"67",X"3E",X"04",X"77",X"E1",X"C9",X"C5",X"F5",X"E5",X"06",X"70",X"21",X"00",X"03",X"2B",
		X"7C",X"FE",X"00",X"20",X"FA",X"10",X"F5",X"E1",X"F1",X"C1",X"C9",X"21",X"25",X"93",X"11",X"4F",
		X"57",X"CD",X"67",X"CA",X"21",X"05",X"92",X"11",X"55",X"57",X"CD",X"67",X"CA",X"21",X"E3",X"92",
		X"11",X"90",X"56",X"CD",X"67",X"CA",X"21",X"83",X"98",X"3E",X"0E",X"CD",X"05",X"56",X"11",X"00",
		X"4D",X"21",X"82",X"93",X"3E",X"12",X"08",X"CD",X"F0",X"55",X"11",X"1B",X"4D",X"21",X"90",X"93",
		X"3E",X"12",X"08",X"CD",X"F0",X"55",X"06",X"0D",X"3E",X"8B",X"21",X"83",X"93",X"CD",X"EB",X"C8",
		X"3E",X"8E",X"06",X"0D",X"21",X"63",X"90",X"CD",X"EB",X"C8",X"C9",X"77",X"E5",X"F5",X"7C",X"C6",
		X"08",X"67",X"3E",X"10",X"77",X"F1",X"E1",X"23",X"10",X"F1",X"C9",X"DD",X"E5",X"C5",X"E5",X"D5",
		X"CD",X"9B",X"C8",X"11",X"20",X"00",X"21",X"8F",X"92",X"DD",X"21",X"17",X"62",X"06",X"05",X"C5",
		X"E5",X"06",X"03",X"DD",X"7E",X"00",X"E6",X"0F",X"CD",X"7C",X"C8",X"DD",X"7E",X"00",X"0F",X"0F",
		X"0F",X"0F",X"E6",X"0F",X"11",X"20",X"00",X"19",X"CD",X"7C",X"C8",X"DD",X"23",X"19",X"10",X"E3",
		X"E1",X"2B",X"2B",X"C1",X"11",X"0D",X"00",X"DD",X"19",X"10",X"D4",X"11",X"20",X"00",X"DD",X"21",
		X"17",X"62",X"21",X"0F",X"92",X"06",X"05",X"C5",X"E5",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"06",
		X"0D",X"DD",X"7E",X"00",X"CD",X"7C",X"C8",X"DD",X"23",X"ED",X"52",X"10",X"F4",X"E1",X"2B",X"2B",
		X"C1",X"10",X"E4",X"D1",X"E1",X"C1",X"DD",X"E1",X"C9",X"3E",X"01",X"32",X"67",X"62",X"21",X"72",
		X"93",X"11",X"1E",X"57",X"CD",X"67",X"CA",X"21",X"73",X"93",X"11",X"37",X"57",X"CD",X"67",X"CA",
		X"21",X"7D",X"93",X"11",X"75",X"57",X"CD",X"67",X"CA",X"11",X"00",X"4D",X"21",X"91",X"93",X"3E",
		X"12",X"08",X"CD",X"F0",X"55",X"11",X"1B",X"4D",X"21",X"9E",X"93",X"3E",X"12",X"08",X"CD",X"F0",
		X"55",X"06",X"0C",X"21",X"92",X"93",X"3E",X"8B",X"CD",X"EB",X"C8",X"06",X"0C",X"3E",X"8E",X"21",
		X"72",X"90",X"CD",X"EB",X"C8",X"11",X"36",X"4D",X"21",X"75",X"92",X"CD",X"49",X"CA",X"11",X"4A",
		X"4D",X"21",X"B8",X"91",X"CD",X"49",X"CA",X"11",X"5E",X"4D",X"21",X"9B",X"92",X"CD",X"49",X"CA",
		X"11",X"72",X"4D",X"21",X"F8",X"92",X"CD",X"49",X"CA",X"11",X"86",X"4D",X"21",X"58",X"92",X"CD",
		X"42",X"CA",X"11",X"8C",X"4D",X"21",X"16",X"92",X"CD",X"42",X"CA",X"11",X"8E",X"4D",X"21",X"17",
		X"92",X"CD",X"42",X"CA",X"11",X"90",X"4D",X"21",X"19",X"92",X"CD",X"42",X"CA",X"11",X"92",X"4D",
		X"21",X"1A",X"92",X"CD",X"42",X"CA",X"CD",X"9B",X"C8",X"C9",X"AF",X"32",X"07",X"A0",X"3E",X"07",
		X"D3",X"08",X"3E",X"38",X"D3",X"09",X"3E",X"0E",X"D3",X"08",X"DB",X"0C",X"2F",X"32",X"78",X"62",
		X"3E",X"01",X"32",X"07",X"A0",X"C9",X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"38",
		X"D3",X"09",X"3E",X"0F",X"D3",X"08",X"DB",X"0C",X"2F",X"32",X"78",X"62",X"3E",X"01",X"32",X"07",
		X"A0",X"C9",X"3E",X"14",X"08",X"CD",X"F0",X"55",X"C9",X"3E",X"18",X"08",X"CD",X"53",X"CA",X"CD",
		X"F0",X"55",X"C9",X"F5",X"3A",X"00",X"B0",X"E6",X"20",X"FE",X"20",X"20",X"08",X"E5",X"EB",X"11",
		X"0A",X"00",X"19",X"EB",X"E1",X"F1",X"C9",X"F5",X"3A",X"00",X"B0",X"E6",X"20",X"FE",X"20",X"28",
		X"08",X"E5",X"EB",X"11",X"96",X"01",X"19",X"EB",X"E1",X"F1",X"CD",X"D9",X"55",X"C9",X"11",X"5A",
		X"57",X"21",X"A0",X"93",X"CD",X"67",X"CA",X"11",X"63",X"57",X"21",X"20",X"91",X"CD",X"67",X"CA",
		X"C9",X"3A",X"26",X"60",X"FE",X"A5",X"C0",X"11",X"58",X"1A",X"21",X"A2",X"93",X"CD",X"F0",X"55",
		X"11",X"75",X"1A",X"21",X"A3",X"93",X"CD",X"F0",X"55",X"3E",X"00",X"18",X"E4",X"DD",X"21",X"CC",
		X"61",X"AF",X"DD",X"77",X"03",X"32",X"E0",X"61",X"32",X"E1",X"61",X"3E",X"FF",X"32",X"9F",X"65",
		X"C9",X"DD",X"7E",X"00",X"6F",X"DD",X"7E",X"01",X"67",X"3A",X"0D",X"60",X"47",X"DD",X"7E",X"02",
		X"B8",X"C0",X"3A",X"41",X"63",X"FE",X"01",X"28",X"47",X"3E",X"D0",X"77",X"E5",X"CD",X"14",X"CB",
		X"E1",X"23",X"7E",X"FE",X"ED",X"28",X"0C",X"FE",X"EF",X"28",X"08",X"3E",X"D1",X"77",X"E5",X"CD",
		X"14",X"CB",X"E1",X"11",X"20",X"00",X"19",X"7E",X"FE",X"D1",X"C8",X"FE",X"67",X"C8",X"FE",X"27",
		X"C8",X"FE",X"ED",X"C8",X"FE",X"EF",X"C8",X"FE",X"DB",X"C8",X"FE",X"FD",X"C8",X"3E",X"D3",X"77",
		X"CD",X"14",X"CB",X"C9",X"7C",X"FE",X"00",X"C8",X"C6",X"08",X"67",X"3A",X"7A",X"62",X"77",X"C9",
		X"23",X"7E",X"FE",X"ED",X"28",X"0C",X"FE",X"EF",X"28",X"08",X"3E",X"C5",X"77",X"E5",X"CD",X"4D",
		X"CB",X"E1",X"11",X"20",X"00",X"19",X"7E",X"FE",X"D1",X"C8",X"FE",X"67",X"C8",X"FE",X"27",X"C8",
		X"FE",X"ED",X"C8",X"FE",X"EF",X"C8",X"3E",X"C7",X"77",X"CD",X"4D",X"CB",X"C9",X"7C",X"FE",X"00",
		X"C8",X"C6",X"08",X"67",X"3E",X"24",X"77",X"C9",X"DD",X"21",X"94",X"65",X"3A",X"3B",X"60",X"FE",
		X"01",X"C8",X"3A",X"56",X"61",X"FE",X"01",X"C8",X"3A",X"11",X"62",X"FE",X"01",X"C8",X"CD",X"A2",
		X"CB",X"78",X"32",X"99",X"60",X"AF",X"32",X"B5",X"62",X"32",X"B6",X"62",X"C9",X"DD",X"21",X"98",
		X"65",X"3A",X"7B",X"60",X"FE",X"01",X"C8",X"3A",X"57",X"61",X"FE",X"01",X"C8",X"3A",X"12",X"62",
		X"FE",X"01",X"C8",X"CD",X"A2",X"CB",X"78",X"32",X"9A",X"60",X"AF",X"32",X"B9",X"62",X"32",X"BA",
		X"62",X"C9",X"3E",X"80",X"DD",X"77",X"02",X"3E",X"10",X"DD",X"77",X"03",X"06",X"03",X"3A",X"0D",
		X"60",X"FE",X"05",X"C8",X"06",X"02",X"FE",X"04",X"C8",X"06",X"01",X"FE",X"03",X"C8",X"06",X"04",
		X"FE",X"02",X"C8",X"06",X"03",X"C9",X"3A",X"F3",X"61",X"FE",X"00",X"C8",X"3C",X"C5",X"47",X"3A",
		X"75",X"62",X"FE",X"01",X"78",X"C1",X"20",X"06",X"FE",X"30",X"20",X"0B",X"18",X"02",X"FE",X"17",
		X"20",X"05",X"3E",X"00",X"32",X"75",X"62",X"32",X"F3",X"61",X"C9",X"3A",X"82",X"65",X"FE",X"E8",
		X"3E",X"00",X"32",X"85",X"62",X"D4",X"15",X"CC",X"3A",X"82",X"65",X"FE",X"10",X"DC",X"8D",X"CC",
		X"3E",X"00",X"32",X"6F",X"62",X"CD",X"9F",X"D5",X"F3",X"AF",X"32",X"00",X"A0",X"FB",X"3E",X"01",
		X"32",X"00",X"A0",X"00",X"C9",X"CD",X"CC",X"CD",X"3A",X"0D",X"60",X"FE",X"01",X"20",X"16",X"CD",
		X"72",X"C2",X"3E",X"02",X"32",X"0D",X"60",X"3E",X"11",X"32",X"82",X"65",X"CD",X"72",X"FD",X"CD",
		X"1B",X"CE",X"C3",X"1A",X"CD",X"3A",X"0D",X"60",X"FE",X"02",X"20",X"16",X"CD",X"0E",X"C2",X"3E",
		X"03",X"32",X"0D",X"60",X"CD",X"72",X"FD",X"3E",X"11",X"32",X"82",X"65",X"CD",X"1B",X"CE",X"C3",
		X"1A",X"CD",X"3A",X"0D",X"60",X"FE",X"03",X"20",X"16",X"CD",X"C1",X"C1",X"3E",X"04",X"32",X"0D",
		X"60",X"CD",X"72",X"FD",X"3E",X"11",X"32",X"82",X"65",X"CD",X"1B",X"CE",X"C3",X"1A",X"CD",X"3A",
		X"0D",X"60",X"FE",X"04",X"20",X"16",X"CD",X"89",X"C1",X"3E",X"05",X"32",X"0D",X"60",X"CD",X"72",
		X"FD",X"3E",X"11",X"32",X"82",X"65",X"CD",X"1B",X"CE",X"C3",X"1A",X"CD",X"C9",X"3E",X"01",X"32",
		X"85",X"62",X"CD",X"CC",X"CD",X"3A",X"0D",X"60",X"FE",X"01",X"C8",X"FE",X"02",X"20",X"16",X"CD",
		X"C9",X"C2",X"3E",X"01",X"32",X"0D",X"60",X"CD",X"72",X"FD",X"3E",X"E3",X"32",X"82",X"65",X"CD",
		X"1B",X"CE",X"C3",X"1F",X"CD",X"FE",X"03",X"20",X"1E",X"DD",X"21",X"42",X"44",X"DD",X"22",X"81",
		X"62",X"CD",X"72",X"C2",X"3E",X"02",X"32",X"0D",X"60",X"3E",X"E3",X"32",X"82",X"65",X"CD",X"72",
		X"FD",X"CD",X"1B",X"CE",X"C3",X"1F",X"CD",X"FE",X"04",X"20",X"1E",X"DD",X"21",X"42",X"44",X"DD",
		X"22",X"81",X"62",X"CD",X"0E",X"C2",X"3E",X"03",X"32",X"0D",X"60",X"3E",X"E3",X"32",X"82",X"65",
		X"CD",X"72",X"FD",X"CD",X"1B",X"CE",X"C3",X"1F",X"CD",X"FE",X"05",X"C0",X"DD",X"21",X"42",X"44",
		X"DD",X"22",X"81",X"62",X"CD",X"C1",X"C1",X"3E",X"04",X"32",X"0D",X"60",X"3E",X"E3",X"32",X"82",
		X"65",X"CD",X"72",X"FD",X"CD",X"1B",X"CE",X"C3",X"1F",X"CD",X"11",X"28",X"E8",X"18",X"03",X"11",
		X"18",X"C8",X"3A",X"58",X"63",X"FE",X"00",X"C4",X"C9",X"C2",X"3E",X"01",X"32",X"03",X"A0",X"DD",
		X"21",X"94",X"65",X"FD",X"21",X"80",X"65",X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"C2",X"54",X"CD",
		X"DD",X"7E",X"02",X"BA",X"38",X"05",X"CD",X"C5",X"D0",X"18",X"09",X"DD",X"7E",X"02",X"BB",X"30",
		X"03",X"CD",X"C5",X"D0",X"DD",X"21",X"98",X"65",X"FD",X"21",X"80",X"65",X"FD",X"7E",X"03",X"DD",
		X"BE",X"03",X"C2",X"79",X"CD",X"DD",X"7E",X"02",X"BA",X"38",X"05",X"CD",X"D1",X"D0",X"18",X"09",
		X"DD",X"7E",X"02",X"BB",X"30",X"03",X"CD",X"D1",X"D0",X"3A",X"1C",X"60",X"FE",X"01",X"C8",X"3A",
		X"1D",X"60",X"FE",X"01",X"C8",X"3A",X"1E",X"60",X"FE",X"01",X"C8",X"21",X"83",X"65",X"DD",X"21",
		X"8C",X"65",X"7E",X"FE",X"40",X"20",X"05",X"CD",X"C1",X"CD",X"18",X"17",X"DD",X"21",X"88",X"65",
		X"FE",X"E0",X"20",X"05",X"CD",X"C1",X"CD",X"18",X"0A",X"DD",X"21",X"90",X"65",X"FE",X"C8",X"C0",
		X"CD",X"C1",X"CD",X"06",X"30",X"C5",X"CD",X"A6",X"09",X"C1",X"10",X"F9",X"AF",X"32",X"25",X"60",
		X"C9",X"DD",X"7E",X"02",X"FE",X"D8",X"D0",X"FE",X"18",X"D8",X"F1",X"C9",X"AF",X"32",X"03",X"A0",
		X"32",X"8F",X"65",X"32",X"97",X"62",X"32",X"F5",X"62",X"32",X"FA",X"62",X"32",X"23",X"63",X"32",
		X"24",X"63",X"3A",X"C7",X"61",X"FE",X"00",X"CC",X"CC",X"F9",X"3A",X"59",X"61",X"FE",X"00",X"28",
		X"0C",X"3A",X"9F",X"65",X"3C",X"32",X"9F",X"65",X"CD",X"99",X"F1",X"18",X"CF",X"3A",X"3B",X"60",
		X"FE",X"01",X"20",X"08",X"3E",X"01",X"32",X"EB",X"61",X"32",X"3A",X"60",X"3A",X"7B",X"60",X"FE",
		X"01",X"C0",X"3E",X"01",X"32",X"EC",X"61",X"32",X"7A",X"60",X"C9",X"DD",X"21",X"19",X"60",X"21",
		X"82",X"65",X"FD",X"21",X"8A",X"65",X"11",X"04",X"00",X"CD",X"3B",X"CE",X"DD",X"23",X"FD",X"19",
		X"CD",X"3B",X"CE",X"DD",X"23",X"FD",X"19",X"CD",X"3B",X"CE",X"C9",X"DD",X"7E",X"03",X"FE",X"00",
		X"C8",X"7E",X"FD",X"77",X"00",X"3A",X"0D",X"60",X"3D",X"DD",X"77",X"00",X"C9",X"3A",X"7D",X"62",
		X"32",X"F3",X"91",X"FE",X"E0",X"28",X"01",X"3D",X"32",X"F4",X"91",X"3E",X"53",X"E5",X"D5",X"C5",
		X"21",X"B1",X"93",X"11",X"E0",X"FF",X"06",X"06",X"77",X"3D",X"F5",X"E5",X"7C",X"C6",X"08",X"67",
		X"3E",X"1F",X"77",X"E1",X"F1",X"19",X"10",X"F0",X"C1",X"D1",X"E1",X"C9",X"C5",X"47",X"7C",X"FE",
		X"00",X"78",X"C1",X"C8",X"F5",X"7E",X"FE",X"D0",X"28",X"06",X"F1",X"CD",X"A6",X"CE",X"18",X"01",
		X"F1",X"23",X"3C",X"CD",X"A6",X"CE",X"D5",X"11",X"1F",X"00",X"19",X"D1",X"3C",X"CD",X"A6",X"CE",
		X"23",X"3C",X"CD",X"A6",X"CE",X"C9",X"77",X"E5",X"F5",X"7C",X"C6",X"08",X"67",X"08",X"77",X"08",
		X"F1",X"E1",X"C9",X"3A",X"5E",X"61",X"FE",X"01",X"C0",X"DD",X"21",X"94",X"65",X"CD",X"D2",X"CE",
		X"FE",X"01",X"CC",X"F4",X"FC",X"DD",X"21",X"98",X"65",X"CD",X"D2",X"CE",X"FE",X"01",X"CC",X"33",
		X"FD",X"C9",X"FD",X"21",X"9C",X"65",X"FD",X"7E",X"02",X"DD",X"BE",X"02",X"28",X"06",X"3C",X"DD",
		X"BE",X"02",X"20",X"1F",X"FD",X"7E",X"03",X"3C",X"3C",X"DD",X"BE",X"03",X"28",X"18",X"3D",X"DD",
		X"BE",X"03",X"28",X"12",X"3D",X"DD",X"BE",X"03",X"28",X"0C",X"3D",X"DD",X"BE",X"03",X"28",X"06",
		X"3D",X"28",X"03",X"3E",X"00",X"C9",X"3E",X"01",X"C9",X"21",X"04",X"A0",X"FD",X"21",X"E5",X"61",
		X"FD",X"7E",X"00",X"FE",X"00",X"28",X"16",X"FD",X"34",X"01",X"FD",X"7E",X"01",X"FE",X"10",X"38",
		X"0C",X"FE",X"20",X"38",X"0B",X"FD",X"35",X"00",X"AF",X"FD",X"77",X"01",X"C9",X"AF",X"77",X"C9",
		X"3E",X"01",X"77",X"C9",X"3A",X"00",X"A0",X"E6",X"3F",X"47",X"00",X"10",X"FD",X"3A",X"56",X"63",
		X"C9",X"3A",X"00",X"B0",X"E6",X"40",X"FE",X"40",X"3E",X"03",X"28",X"02",X"3E",X"04",X"47",X"3A",
		X"7C",X"61",X"FE",X"01",X"3A",X"78",X"61",X"20",X"03",X"3A",X"7B",X"61",X"B8",X"30",X"05",X"AF",
		X"32",X"86",X"62",X"C9",X"3A",X"86",X"62",X"FE",X"00",X"C0",X"3A",X"56",X"60",X"3C",X"32",X"56",
		X"60",X"3E",X"01",X"32",X"86",X"62",X"C9",X"7E",X"FE",X"E0",X"20",X"23",X"3A",X"0D",X"60",X"B8",
		X"28",X"1D",X"78",X"FE",X"02",X"01",X"65",X"61",X"28",X"05",X"FE",X"03",X"01",X"66",X"61",X"0A",
		X"FE",X"10",X"D8",X"08",X"FE",X"00",X"20",X"03",X"0A",X"3D",X"02",X"1A",X"3D",X"12",X"C9",X"AF",
		X"DD",X"77",X"00",X"FD",X"77",X"00",X"C9",X"21",X"E7",X"61",X"7E",X"D6",X"01",X"27",X"77",X"CB",
		X"19",X"23",X"7E",X"FE",X"00",X"C8",X"CB",X"11",X"DE",X"00",X"27",X"77",X"C9",X"3A",X"D3",X"60",
		X"3C",X"32",X"D3",X"60",X"AF",X"32",X"41",X"63",X"11",X"9C",X"60",X"21",X"15",X"1B",X"FE",X"02",
		X"20",X"03",X"21",X"4E",X"1B",X"01",X"36",X"00",X"ED",X"B0",X"C9",X"11",X"9C",X"60",X"21",X"DC",
		X"1A",X"01",X"36",X"00",X"ED",X"B0",X"C9",X"11",X"7F",X"61",X"21",X"DC",X"1A",X"01",X"36",X"00",
		X"ED",X"B0",X"C9",X"FE",X"E0",X"C8",X"FE",X"4B",X"C8",X"FE",X"4A",X"C8",X"FE",X"49",X"C8",X"FE",
		X"E4",X"C8",X"FE",X"E6",X"C8",X"FE",X"D4",X"C8",X"FE",X"D6",X"C9",X"E5",X"C5",X"01",X"E0",X"FF",
		X"09",X"AF",X"ED",X"52",X"C1",X"E1",X"C9",X"3A",X"7D",X"61",X"FE",X"01",X"C8",X"3E",X"01",X"32",
		X"53",X"60",X"32",X"8C",X"62",X"CD",X"E3",X"C3",X"11",X"5A",X"57",X"21",X"74",X"92",X"CD",X"67",
		X"CA",X"11",X"89",X"56",X"21",X"9F",X"91",X"CD",X"67",X"CA",X"3A",X"7C",X"61",X"3C",X"32",X"94",
		X"91",X"3E",X"08",X"21",X"7F",X"98",X"CD",X"05",X"56",X"3E",X"00",X"32",X"5F",X"98",X"3E",X"05",
		X"21",X"41",X"98",X"CD",X"05",X"56",X"3E",X"02",X"21",X"40",X"98",X"CD",X"05",X"56",X"21",X"93",
		X"92",X"11",X"42",X"1A",X"3E",X"1F",X"08",X"CD",X"F0",X"55",X"21",X"95",X"92",X"11",X"4D",X"1A",
		X"3E",X"1F",X"08",X"CD",X"F0",X"55",X"3E",X"8E",X"32",X"74",X"91",X"3E",X"8B",X"32",X"94",X"92",
		X"3E",X"1F",X"32",X"74",X"99",X"32",X"94",X"9A",X"CD",X"2E",X"16",X"3E",X"00",X"32",X"03",X"98",
		X"32",X"07",X"98",X"32",X"0B",X"98",X"32",X"0F",X"98",X"32",X"13",X"98",X"32",X"17",X"98",X"32",
		X"1B",X"98",X"32",X"1F",X"98",X"21",X"30",X"01",X"06",X"80",X"3A",X"00",X"B8",X"C5",X"E5",X"CD",
		X"2E",X"16",X"E1",X"C1",X"10",X"F4",X"2B",X"7C",X"FE",X"00",X"20",X"EC",X"3E",X"00",X"32",X"53",
		X"60",X"32",X"8C",X"62",X"C9",X"D5",X"06",X"60",X"C5",X"CD",X"C0",X"11",X"C1",X"10",X"F9",X"D1",
		X"C9",X"D5",X"06",X"60",X"C5",X"CD",X"EC",X"11",X"C1",X"10",X"F9",X"D1",X"C9",X"11",X"89",X"56",
		X"21",X"9F",X"91",X"CD",X"67",X"CA",X"3A",X"00",X"B8",X"11",X"05",X"57",X"21",X"40",X"92",X"CD",
		X"67",X"CA",X"C9",X"CD",X"D9",X"D4",X"C0",X"3A",X"53",X"63",X"3C",X"FE",X"03",X"38",X"01",X"AF",
		X"32",X"53",X"63",X"21",X"68",X"3B",X"FE",X"01",X"28",X"0A",X"21",X"00",X"38",X"FE",X"02",X"28",
		X"03",X"21",X"00",X"50",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"C9",X"3A",X"0D",X"60",X"FE",
		X"05",X"C0",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"3A",X"82",X"65",X"FE",X"B3",X"C0",X"C9",X"CD",
		X"69",X"D2",X"79",X"FE",X"00",X"C8",X"3A",X"41",X"63",X"FE",X"01",X"CA",X"D0",X"D1",X"3E",X"00",
		X"32",X"03",X"A0",X"CD",X"B7",X"C3",X"3E",X"04",X"CD",X"A3",X"C3",X"3E",X"01",X"32",X"32",X"63",
		X"32",X"42",X"63",X"DD",X"21",X"13",X"1C",X"3A",X"00",X"B0",X"E6",X"20",X"FE",X"20",X"20",X"04",
		X"DD",X"21",X"6A",X"1C",X"CD",X"2A",X"D8",X"AF",X"32",X"32",X"63",X"32",X"42",X"63",X"F3",X"3E",
		X"01",X"32",X"41",X"63",X"CD",X"51",X"F9",X"CD",X"14",X"C3",X"CD",X"BF",X"DF",X"2A",X"C4",X"61",
		X"E5",X"21",X"00",X"00",X"22",X"C4",X"61",X"E1",X"23",X"3E",X"E0",X"77",X"11",X"20",X"00",X"19",
		X"77",X"DD",X"21",X"B5",X"D1",X"11",X"03",X"00",X"3A",X"00",X"A0",X"E6",X"07",X"3C",X"47",X"DD",
		X"19",X"10",X"FC",X"DD",X"7E",X"00",X"6F",X"DD",X"7E",X"01",X"67",X"DD",X"7E",X"02",X"22",X"9F",
		X"60",X"32",X"A1",X"60",X"C9",X"00",X"00",X"00",X"23",X"91",X"01",X"03",X"92",X"02",X"A3",X"92",
		X"03",X"7C",X"92",X"03",X"03",X"91",X"03",X"F0",X"90",X"03",X"D3",X"92",X"01",X"3C",X"92",X"02",
		X"3A",X"43",X"63",X"FE",X"01",X"28",X"1C",X"AF",X"32",X"88",X"62",X"32",X"54",X"60",X"3E",X"E0",
		X"32",X"0E",X"93",X"32",X"0F",X"93",X"3E",X"01",X"32",X"43",X"63",X"32",X"41",X"63",X"3E",X"E0",
		X"32",X"8E",X"93",X"3E",X"05",X"32",X"99",X"60",X"32",X"9A",X"69",X"3A",X"82",X"65",X"FE",X"10",
		X"C0",X"3A",X"83",X"65",X"FE",X"18",X"C0",X"3E",X"00",X"32",X"43",X"63",X"32",X"53",X"60",X"3E",
		X"01",X"32",X"41",X"63",X"32",X"03",X"A0",X"32",X"32",X"63",X"32",X"42",X"63",X"CD",X"B7",X"C3",
		X"3E",X"04",X"CD",X"A3",X"C3",X"DD",X"21",X"AE",X"1C",X"3A",X"00",X"B0",X"E6",X"20",X"FE",X"20",
		X"20",X"04",X"DD",X"21",X"25",X"1D",X"CD",X"2A",X"D8",X"AF",X"32",X"32",X"63",X"32",X"42",X"63",
		X"32",X"41",X"63",X"3E",X"01",X"32",X"54",X"60",X"3A",X"56",X"60",X"3C",X"32",X"56",X"60",X"F3",
		X"06",X"40",X"21",X"80",X"65",X"3E",X"00",X"77",X"23",X"10",X"FC",X"3E",X"01",X"32",X"54",X"60",
		X"CD",X"BD",X"CF",X"31",X"F0",X"67",X"C3",X"DC",X"EC",X"0E",X"00",X"FD",X"21",X"9C",X"60",X"06",
		X"36",X"FD",X"7E",X"00",X"FE",X"00",X"C0",X"FD",X"23",X"10",X"F6",X"0E",X"01",X"C9",X"21",X"F4",
		X"61",X"7E",X"47",X"3A",X"E8",X"61",X"B8",X"C8",X"FE",X"05",X"D0",X"21",X"94",X"5B",X"22",X"40",
		X"61",X"32",X"F4",X"61",X"AF",X"32",X"42",X"61",X"C9",X"C9",X"3A",X"0D",X"60",X"32",X"98",X"60",
		X"FD",X"21",X"61",X"61",X"DD",X"21",X"84",X"65",X"CD",X"EF",X"EA",X"3A",X"0D",X"60",X"FE",X"04",
		X"28",X"04",X"C9",X"FE",X"05",X"C0",X"DD",X"7E",X"03",X"FE",X"11",X"D8",X"3A",X"0D",X"60",X"FE",
		X"04",X"20",X"11",X"11",X"DE",X"30",X"AF",X"ED",X"5A",X"7C",X"C6",X"2F",X"67",X"11",X"C3",X"90",
		X"06",X"1A",X"18",X"0B",X"11",X"FE",X"34",X"AF",X"ED",X"5A",X"11",X"E4",X"90",X"06",X"1A",X"3E",
		X"FB",X"E5",X"AF",X"ED",X"52",X"E1",X"28",X"09",X"3E",X"FB",X"CD",X"13",X"D3",X"13",X"10",X"EF",
		X"C9",X"DD",X"7E",X"03",X"E6",X"07",X"47",X"3E",X"F3",X"80",X"CD",X"13",X"D3",X"06",X"03",X"13",
		X"C5",X"1A",X"01",X"08",X"00",X"21",X"26",X"D3",X"ED",X"B1",X"3E",X"F3",X"CC",X"13",X"D3",X"C1",
		X"10",X"ED",X"C9",X"12",X"C5",X"47",X"1A",X"B8",X"78",X"C1",X"20",X"F7",X"D5",X"7A",X"C6",X"08",
		X"57",X"3E",X"20",X"12",X"D1",X"C9",X"FB",X"FA",X"F9",X"F8",X"F7",X"F6",X"F5",X"F4",X"2A",X"91",
		X"60",X"22",X"FF",X"61",X"2A",X"93",X"60",X"22",X"01",X"62",X"2A",X"95",X"60",X"22",X"03",X"62",
		X"3A",X"0B",X"60",X"32",X"05",X"62",X"3A",X"98",X"60",X"32",X"F9",X"61",X"C9",X"2A",X"FF",X"61",
		X"22",X"91",X"60",X"2A",X"01",X"62",X"22",X"93",X"60",X"2A",X"03",X"62",X"22",X"95",X"60",X"3A",
		X"05",X"62",X"32",X"0B",X"60",X"3A",X"F9",X"61",X"32",X"98",X"60",X"C9",X"F5",X"D5",X"E5",X"06",
		X"00",X"CD",X"91",X"D3",X"20",X"17",X"23",X"CD",X"91",X"D3",X"20",X"11",X"11",X"1F",X"00",X"19",
		X"CD",X"91",X"D3",X"20",X"08",X"23",X"CD",X"91",X"D3",X"20",X"02",X"06",X"01",X"E1",X"D1",X"F1",
		X"C9",X"7E",X"FE",X"E0",X"C8",X"FE",X"49",X"C8",X"FE",X"4A",X"C8",X"FE",X"4B",X"C8",X"FE",X"51",
		X"C8",X"FE",X"52",X"C8",X"FE",X"57",X"C9",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"E1",X"C9",
		X"DD",X"21",X"CC",X"61",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"03",X"3E",X"FF",
		X"32",X"9F",X"65",X"C9",X"CD",X"BE",X"EA",X"CD",X"81",X"D4",X"28",X"12",X"AF",X"32",X"77",X"60",
		X"3A",X"09",X"62",X"FE",X"01",X"20",X"07",X"CD",X"33",X"FD",X"AF",X"32",X"09",X"62",X"DD",X"21",
		X"8F",X"60",X"FD",X"21",X"57",X"61",X"21",X"E9",X"62",X"D9",X"21",X"98",X"65",X"22",X"15",X"62",
		X"2A",X"78",X"60",X"11",X"7B",X"60",X"3A",X"9A",X"60",X"32",X"98",X"60",X"01",X"12",X"62",X"CD",
		X"41",X"D4",X"CD",X"B1",X"EA",X"CD",X"81",X"D4",X"28",X"12",X"AF",X"32",X"37",X"60",X"3A",X"08",
		X"62",X"FE",X"01",X"20",X"07",X"CD",X"F4",X"FC",X"AF",X"32",X"08",X"62",X"DD",X"21",X"4F",X"60",
		X"FD",X"21",X"56",X"61",X"21",X"ED",X"62",X"D9",X"21",X"94",X"65",X"22",X"15",X"62",X"2A",X"38",
		X"60",X"11",X"3B",X"60",X"3A",X"99",X"60",X"32",X"98",X"60",X"01",X"11",X"62",X"CD",X"41",X"D4",
		X"C9",X"DD",X"7E",X"00",X"FE",X"12",X"38",X"15",X"CD",X"81",X"D4",X"20",X"56",X"1A",X"FE",X"01",
		X"28",X"51",X"D9",X"7E",X"D9",X"FE",X"01",X"28",X"4A",X"3E",X"01",X"02",X"C9",X"0A",X"FE",X"01",
		X"28",X"47",X"AF",X"C9",X"7E",X"E5",X"C5",X"01",X"0A",X"00",X"21",X"77",X"D4",X"ED",X"B1",X"C1",
		X"E1",X"C8",X"AF",X"32",X"08",X"60",X"C9",X"E0",X"FB",X"B3",X"B2",X"B1",X"B0",X"4C",X"4D",X"4E",
		X"4F",X"7E",X"E5",X"C5",X"01",X"14",X"00",X"21",X"8F",X"D4",X"ED",X"B1",X"C1",X"E1",X"C9",X"FF",
		X"FE",X"FD",X"FC",X"FB",X"FA",X"F9",X"E2",X"E1",X"E0",X"DF",X"DE",X"4C",X"4D",X"4E",X"4F",X"B3",
		X"B2",X"B1",X"B0",X"2A",X"15",X"62",X"3E",X"22",X"77",X"AF",X"02",X"DD",X"77",X"00",X"3E",X"01",
		X"FD",X"77",X"00",X"EB",X"11",X"04",X"00",X"AF",X"ED",X"52",X"77",X"21",X"52",X"27",X"22",X"54",
		X"61",X"AF",X"32",X"F5",X"61",X"3A",X"98",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"C0",X"21",X"B1",
		X"D9",X"CD",X"84",X"EC",X"AF",X"32",X"53",X"61",X"C9",X"DD",X"E5",X"DD",X"2A",X"40",X"61",X"DD",
		X"7E",X"03",X"DD",X"E1",X"FE",X"FF",X"C0",X"3A",X"43",X"63",X"FE",X"01",X"C8",X"3A",X"10",X"62",
		X"FE",X"01",X"C8",X"3A",X"00",X"60",X"FE",X"00",X"20",X"0F",X"3A",X"54",X"60",X"FE",X"01",X"28",
		X"08",X"3A",X"00",X"B0",X"E6",X"40",X"FE",X"40",X"C9",X"3E",X"00",X"FE",X"00",X"C9",X"3A",X"54",
		X"60",X"3A",X"00",X"B8",X"DD",X"21",X"80",X"65",X"FD",X"21",X"A8",X"65",X"CD",X"D7",X"D6",X"DD",
		X"21",X"84",X"65",X"FD",X"21",X"A4",X"65",X"CD",X"D7",X"D6",X"DD",X"21",X"88",X"65",X"FD",X"21",
		X"AC",X"65",X"CD",X"D7",X"D6",X"DD",X"21",X"8C",X"65",X"FD",X"21",X"B0",X"65",X"CD",X"D7",X"D6",
		X"DD",X"21",X"90",X"65",X"FD",X"21",X"B4",X"65",X"CD",X"D7",X"D6",X"DD",X"21",X"9C",X"65",X"FD",
		X"21",X"A0",X"65",X"CD",X"D7",X"D6",X"AF",X"32",X"5F",X"98",X"0E",X"01",X"3A",X"FD",X"61",X"FE",
		X"01",X"20",X"02",X"0E",X"FF",X"CD",X"EF",X"D8",X"06",X"08",X"11",X"04",X"00",X"21",X"A3",X"65",
		X"7E",X"FE",X"00",X"28",X"02",X"81",X"77",X"19",X"10",X"F6",X"21",X"AF",X"65",X"06",X"03",X"35",
		X"19",X"10",X"FC",X"79",X"FE",X"FF",X"20",X"16",X"3A",X"0D",X"60",X"FE",X"04",X"20",X"0F",X"3A",
		X"ED",X"61",X"FE",X"01",X"28",X"08",X"3A",X"A6",X"65",X"3C",X"3C",X"32",X"A6",X"65",X"C9",X"3A",
		X"C7",X"61",X"FE",X"00",X"C8",X"3A",X"3A",X"63",X"FE",X"01",X"28",X"14",X"3A",X"82",X"65",X"C6",
		X"0E",X"32",X"9E",X"65",X"3A",X"83",X"65",X"32",X"9F",X"65",X"3E",X"3A",X"32",X"9C",X"65",X"C9",
		X"3A",X"82",X"65",X"C6",X"0D",X"32",X"9E",X"65",X"3A",X"83",X"65",X"C6",X"04",X"32",X"9F",X"65",
		X"3E",X"33",X"32",X"9C",X"65",X"C9",X"3A",X"11",X"63",X"FE",X"00",X"C8",X"3A",X"80",X"65",X"E6",
		X"7F",X"06",X"02",X"FE",X"12",X"28",X"0D",X"06",X"06",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",
		X"20",X"02",X"06",X"F9",X"3A",X"82",X"65",X"80",X"32",X"9E",X"65",X"3A",X"83",X"65",X"32",X"9F",
		X"65",X"3E",X"35",X"32",X"9C",X"65",X"3E",X"24",X"32",X"9D",X"65",X"C9",X"3A",X"43",X"63",X"FE",
		X"00",X"C8",X"3A",X"80",X"65",X"E6",X"7F",X"0E",X"00",X"06",X"00",X"FE",X"12",X"28",X"11",X"0E",
		X"80",X"06",X"06",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",X"20",X"04",X"0E",X"00",X"06",X"F9",
		X"3A",X"82",X"65",X"80",X"32",X"9E",X"65",X"3A",X"83",X"65",X"C6",X"04",X"32",X"9F",X"65",X"3E",
		X"1B",X"B1",X"32",X"9C",X"65",X"3E",X"08",X"32",X"9D",X"65",X"C9",X"3A",X"C7",X"61",X"FE",X"01",
		X"C0",X"CD",X"CE",X"D6",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"06",X"08",X"CD",X"B8",X"D6",X"3A",
		X"C7",X"61",X"FE",X"01",X"C0",X"06",X"10",X"CD",X"C4",X"D6",X"3A",X"C7",X"61",X"FE",X"01",X"C0",
		X"06",X"08",X"CD",X"C4",X"D6",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"06",X"08",X"CD",X"C4",X"D6",
		X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"06",X"08",X"CD",X"C4",X"D6",X"3A",X"C7",X"61",X"FE",X"01",
		X"C0",X"06",X"08",X"CD",X"C4",X"D6",X"06",X"08",X"CD",X"C4",X"D6",X"3A",X"C7",X"61",X"FE",X"01",
		X"C0",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"06",X"40",X"CD",X"B8",X"D6",X"3A",X"C7",X"61",X"FE",
		X"01",X"C0",X"06",X"08",X"CD",X"B8",X"D6",X"C9",X"3A",X"9E",X"65",X"80",X"FE",X"E0",X"D0",X"32",
		X"9E",X"65",X"18",X"0A",X"3A",X"9E",X"65",X"90",X"FE",X"10",X"D8",X"32",X"9E",X"65",X"3E",X"01",
		X"32",X"60",X"61",X"CD",X"BD",X"DA",X"C9",X"06",X"04",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",
		X"23",X"FD",X"23",X"10",X"F4",X"C9",X"3A",X"0D",X"60",X"FE",X"05",X"C0",X"DD",X"7E",X"02",X"FE",
		X"A9",X"D8",X"3A",X"E3",X"62",X"C6",X"08",X"47",X"C6",X"08",X"4F",X"DD",X"7E",X"03",X"B8",X"D8",
		X"B9",X"D0",X"3E",X"01",X"FD",X"77",X"00",X"C9",X"3A",X"0D",X"60",X"FE",X"05",X"20",X"0B",X"DD",
		X"21",X"80",X"65",X"FD",X"21",X"25",X"60",X"CD",X"E6",X"D6",X"3A",X"99",X"60",X"FE",X"05",X"20",
		X"0B",X"DD",X"21",X"94",X"65",X"FD",X"21",X"9F",X"62",X"CD",X"E6",X"D6",X"3A",X"9A",X"60",X"FE",
		X"05",X"C0",X"DD",X"21",X"98",X"65",X"FD",X"21",X"A7",X"62",X"CD",X"E6",X"D6",X"C9",X"3A",X"C7",
		X"61",X"FE",X"01",X"C8",X"3A",X"CF",X"61",X"FE",X"01",X"C8",X"3A",X"11",X"63",X"FE",X"01",X"C8",
		X"3A",X"58",X"61",X"FE",X"01",X"C9",X"AF",X"32",X"97",X"60",X"32",X"88",X"62",X"32",X"08",X"60",
		X"32",X"13",X"60",X"32",X"29",X"60",X"32",X"2A",X"60",X"32",X"4E",X"60",X"32",X"77",X"60",X"32",
		X"28",X"60",X"32",X"E0",X"61",X"32",X"E1",X"61",X"32",X"14",X"60",X"32",X"13",X"60",X"32",X"B5",
		X"62",X"32",X"B6",X"62",X"32",X"B9",X"62",X"32",X"BA",X"62",X"32",X"AF",X"62",X"32",X"B0",X"62",
		X"32",X"D2",X"62",X"32",X"D6",X"62",X"32",X"DA",X"62",X"32",X"D3",X"62",X"32",X"BD",X"62",X"32",
		X"F6",X"61",X"32",X"F7",X"61",X"32",X"11",X"63",X"C9",X"3A",X"D3",X"60",X"FE",X"02",X"D8",X"3E",
		X"06",X"32",X"94",X"62",X"32",X"9C",X"62",X"32",X"A4",X"62",X"3E",X"01",X"32",X"93",X"62",X"32",
		X"9B",X"62",X"32",X"A3",X"62",X"32",X"99",X"62",X"C9",X"AF",X"32",X"C7",X"61",X"32",X"CF",X"61",
		X"32",X"14",X"60",X"32",X"1C",X"60",X"32",X"58",X"61",X"32",X"40",X"63",X"32",X"41",X"63",X"3E",
		X"01",X"32",X"D3",X"60",X"32",X"B6",X"61",X"C9",X"DD",X"E5",X"F5",X"D5",X"C5",X"DD",X"21",X"01",
		X"90",X"FD",X"21",X"00",X"90",X"11",X"20",X"00",X"06",X"20",X"DD",X"E5",X"FD",X"E5",X"C5",X"06",
		X"1F",X"DD",X"7E",X"00",X"4F",X"DD",X"7E",X"00",X"B9",X"20",X"F6",X"FD",X"77",X"00",X"DD",X"23",
		X"FD",X"23",X"10",X"ED",X"3E",X"0A",X"FD",X"77",X"00",X"C1",X"FD",X"E1",X"DD",X"E1",X"DD",X"19",
		X"FD",X"19",X"10",X"D6",X"C1",X"D1",X"F1",X"DD",X"E1",X"C9",X"AF",X"06",X"20",X"21",X"00",X"98",
		X"77",X"23",X"10",X"FC",X"32",X"5F",X"98",X"3E",X"01",X"32",X"03",X"A0",X"CD",X"E2",X"D8",X"21",
		X"B0",X"93",X"22",X"2F",X"63",X"ED",X"56",X"FB",X"3E",X"01",X"32",X"00",X"A0",X"DD",X"7E",X"00",
		X"FE",X"FF",X"28",X"1F",X"CD",X"A2",X"D8",X"CD",X"D4",X"D8",X"DD",X"23",X"DD",X"7E",X"00",X"FE",
		X"FE",X"CC",X"86",X"D8",X"3A",X"42",X"63",X"FE",X"01",X"28",X"E2",X"3A",X"00",X"60",X"FE",X"00",
		X"C0",X"18",X"DA",X"CD",X"D4",X"D8",X"CD",X"D4",X"D8",X"CD",X"D4",X"D8",X"CD",X"D4",X"D8",X"CD",
		X"D4",X"D8",X"CD",X"D4",X"D8",X"C9",X"2A",X"2F",X"63",X"F5",X"7D",X"FE",X"BF",X"20",X"05",X"CD",
		X"E8",X"D7",X"18",X"01",X"23",X"22",X"2F",X"63",X"F1",X"DD",X"23",X"CD",X"E8",X"D7",X"CD",X"CD",
		X"D8",X"C9",X"DD",X"7E",X"00",X"D6",X"30",X"FE",X"0A",X"CC",X"D4",X"D8",X"77",X"FE",X"0A",X"C4",
		X"C0",X"D8",X"E5",X"11",X"00",X"08",X"19",X"3E",X"04",X"77",X"E1",X"11",X"E0",X"FF",X"19",X"C9",
		X"E5",X"C5",X"D5",X"21",X"7B",X"D9",X"CD",X"84",X"EC",X"D1",X"C1",X"E1",X"C9",X"E5",X"F5",X"21",
		X"00",X"60",X"18",X"05",X"E5",X"F5",X"21",X"00",X"30",X"2B",X"7C",X"FE",X"00",X"20",X"FA",X"F1",
		X"E1",X"C9",X"F5",X"00",X"00",X"00",X"00",X"32",X"01",X"A0",X"32",X"02",X"A0",X"F1",X"C9",X"C9",
		X"79",X"2F",X"3C",X"4F",X"C9",X"00",X"00",X"B2",X"05",X"61",X"05",X"14",X"05",X"CC",X"04",X"86",
		X"04",X"45",X"04",X"08",X"04",X"CE",X"03",X"97",X"03",X"63",X"03",X"34",X"03",X"05",X"03",X"D9",
		X"02",X"B0",X"02",X"8A",X"02",X"66",X"02",X"43",X"02",X"22",X"02",X"04",X"02",X"E7",X"01",X"CB",
		X"01",X"B2",X"01",X"99",X"01",X"82",X"01",X"6D",X"01",X"58",X"01",X"45",X"01",X"33",X"01",X"22",
		X"01",X"11",X"01",X"02",X"01",X"F4",X"00",X"E6",X"00",X"D9",X"00",X"CD",X"00",X"C1",X"00",X"B6",
		X"00",X"AC",X"00",X"A2",X"00",X"9A",X"00",X"91",X"00",X"89",X"00",X"81",X"00",X"7A",X"00",X"73",
		X"00",X"6C",X"00",X"66",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"00",X"00",X"01",
		X"00",X"01",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"2A",X"3D",X"63",X"7E",X"FE",X"01",X"20",X"0D",X"7E",
		X"23",X"77",X"2A",X"46",X"61",X"23",X"23",X"23",X"23",X"AF",X"77",X"C9",X"FD",X"E5",X"FD",X"21",
		X"A8",X"23",X"FD",X"7E",X"00",X"67",X"FD",X"7E",X"01",X"6F",X"AF",X"ED",X"52",X"28",X"14",X"FD",
		X"23",X"FD",X"23",X"FD",X"7E",X"01",X"FE",X"FF",X"20",X"E8",X"2A",X"3D",X"63",X"7E",X"23",X"77",
		X"FD",X"E1",X"C9",X"FD",X"E1",X"2A",X"3D",X"63",X"23",X"7E",X"2A",X"46",X"61",X"FE",X"01",X"20",
		X"21",X"2A",X"95",X"60",X"3E",X"40",X"77",X"C9",X"06",X"80",X"FD",X"7E",X"03",X"FE",X"98",X"28",
		X"02",X"06",X"40",X"2A",X"95",X"60",X"78",X"77",X"2A",X"46",X"61",X"23",X"23",X"23",X"23",X"AF",
		X"77",X"C9",X"3A",X"0D",X"60",X"FE",X"05",X"20",X"DF",X"FD",X"7E",X"03",X"23",X"23",X"23",X"23",
		X"47",X"3A",X"E3",X"62",X"B8",X"28",X"15",X"3D",X"B8",X"28",X"11",X"3E",X"01",X"77",X"7D",X"21",
		X"57",X"60",X"FE",X"48",X"28",X"03",X"21",X"97",X"60",X"AF",X"77",X"C9",X"AF",X"77",X"2A",X"95",
		X"60",X"3E",X"80",X"77",X"C9",X"3A",X"34",X"63",X"FE",X"01",X"C8",X"2A",X"26",X"63",X"7E",X"FE",
		X"D4",X"28",X"07",X"3E",X"D4",X"08",X"3E",X"24",X"18",X"05",X"3E",X"D0",X"08",X"3E",X"2C",X"08",
		X"77",X"E5",X"F5",X"7C",X"C6",X"08",X"67",X"F1",X"08",X"77",X"E1",X"11",X"20",X"00",X"19",X"08",
		X"3C",X"3C",X"77",X"7C",X"C6",X"08",X"67",X"08",X"77",X"C9",X"3A",X"CF",X"61",X"FE",X"00",X"C8",
		X"2A",X"E0",X"61",X"7D",X"FE",X"00",X"20",X"06",X"7C",X"FE",X"00",X"20",X"01",X"C9",X"23",X"22",
		X"E0",X"61",X"11",X"FF",X"01",X"ED",X"52",X"C0",X"21",X"00",X"00",X"22",X"E0",X"61",X"3E",X"00",
		X"DD",X"21",X"CC",X"61",X"DD",X"77",X"03",X"3E",X"FF",X"32",X"9F",X"65",X"C9",X"3A",X"60",X"61",
		X"FE",X"01",X"C0",X"3A",X"34",X"63",X"FE",X"01",X"C8",X"3A",X"CF",X"61",X"FE",X"01",X"28",X"28",
		X"3A",X"58",X"61",X"FE",X"01",X"28",X"21",X"3A",X"11",X"63",X"FE",X"01",X"CA",X"65",X"DB",X"01",
		X"C7",X"61",X"FD",X"21",X"C4",X"61",X"3E",X"3A",X"FD",X"77",X"04",X"3E",X"28",X"FD",X"77",X"05",
		X"3E",X"EC",X"32",X"CA",X"61",X"CD",X"CC",X"FB",X"06",X"04",X"FD",X"21",X"D0",X"61",X"3A",X"C7",
		X"61",X"FE",X"01",X"CA",X"4F",X"DB",X"C5",X"FD",X"E5",X"01",X"CF",X"61",X"FD",X"21",X"CC",X"61",
		X"3E",X"37",X"FD",X"77",X"04",X"3E",X"20",X"FD",X"77",X"05",X"3A",X"00",X"B8",X"3E",X"E4",X"32",
		X"D2",X"61",X"CD",X"CC",X"FB",X"FD",X"E1",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"CD",X"C2",X"DB",
		X"C1",X"10",X"D3",X"01",X"CF",X"61",X"FD",X"21",X"CC",X"61",X"3E",X"37",X"FD",X"77",X"04",X"3E",
		X"20",X"FD",X"77",X"05",X"3A",X"00",X"B8",X"3E",X"E4",X"32",X"D2",X"61",X"CD",X"CC",X"FB",X"3A",
		X"60",X"61",X"FE",X"01",X"C0",X"3A",X"C7",X"61",X"FE",X"01",X"CA",X"B4",X"DB",X"3A",X"CF",X"61",
		X"FE",X"01",X"CA",X"B4",X"DB",X"06",X"04",X"FD",X"21",X"12",X"63",X"C5",X"FD",X"E5",X"01",X"11",
		X"63",X"FD",X"21",X"0E",X"63",X"3E",X"35",X"FD",X"77",X"04",X"3E",X"24",X"FD",X"77",X"05",X"3A",
		X"00",X"B8",X"3E",X"D4",X"32",X"14",X"63",X"CD",X"CC",X"FB",X"FD",X"E1",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"CD",X"B5",X"DB",X"C1",X"10",X"D3",X"01",X"11",X"63",X"FD",X"21",X"0E",X"63",X"3E",
		X"32",X"FD",X"77",X"04",X"3E",X"24",X"FD",X"77",X"05",X"3A",X"00",X"B8",X"3E",X"D4",X"32",X"14",
		X"63",X"CD",X"CC",X"FB",X"C9",X"C5",X"FD",X"E5",X"DD",X"E5",X"06",X"03",X"DD",X"21",X"0E",X"63",
		X"18",X"0B",X"C5",X"FD",X"E5",X"DD",X"E5",X"06",X"03",X"DD",X"21",X"CC",X"61",X"DD",X"7E",X"00",
		X"08",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"08",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"10",
		X"EC",X"DD",X"E1",X"FD",X"E1",X"C1",X"C9",X"3A",X"F5",X"62",X"FE",X"01",X"C0",X"AF",X"32",X"51",
		X"63",X"2A",X"26",X"63",X"22",X"F6",X"61",X"CD",X"F3",X"F3",X"2A",X"26",X"63",X"11",X"40",X"00",
		X"19",X"22",X"F8",X"62",X"21",X"B6",X"DE",X"22",X"F6",X"62",X"FD",X"2A",X"F8",X"62",X"DD",X"21",
		X"FC",X"62",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"FD",X"7E",
		X"E0",X"DD",X"77",X"02",X"FD",X"7E",X"E1",X"DD",X"77",X"03",X"FD",X"7E",X"C0",X"DD",X"77",X"04",
		X"FD",X"7E",X"C1",X"DD",X"77",X"05",X"FD",X"7E",X"A0",X"DD",X"77",X"06",X"FD",X"7E",X"A1",X"DD",
		X"77",X"07",X"E5",X"C5",X"FD",X"E5",X"06",X"08",X"FD",X"21",X"FC",X"62",X"16",X"0B",X"FD",X"7E",
		X"00",X"BA",X"DC",X"F3",X"DC",X"FD",X"23",X"10",X"F5",X"18",X"00",X"FD",X"E1",X"C1",X"E1",X"FD",
		X"2A",X"F8",X"62",X"11",X"00",X"08",X"FD",X"19",X"DD",X"21",X"04",X"63",X"FD",X"7E",X"00",X"DD",
		X"77",X"00",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"FD",X"7E",X"E0",X"DD",X"77",X"02",X"FD",X"7E",
		X"E1",X"DD",X"77",X"03",X"FD",X"7E",X"C0",X"DD",X"77",X"04",X"FD",X"7E",X"C1",X"DD",X"77",X"05",
		X"FD",X"7E",X"A0",X"DD",X"77",X"06",X"FD",X"7E",X"A1",X"DD",X"77",X"07",X"CD",X"3B",X"DE",X"06",
		X"08",X"DD",X"21",X"FC",X"62",X"FD",X"21",X"04",X"63",X"CD",X"DD",X"DC",X"DD",X"23",X"FD",X"23",
		X"10",X"F7",X"3E",X"01",X"32",X"F5",X"62",X"3A",X"54",X"60",X"FE",X"00",X"C8",X"3E",X"1F",X"32",
		X"4C",X"63",X"3E",X"07",X"32",X"4D",X"63",X"3A",X"48",X"63",X"FE",X"01",X"C8",X"21",X"DC",X"3F",
		X"22",X"4E",X"63",X"AF",X"32",X"42",X"61",X"3E",X"03",X"32",X"48",X"63",X"C9",X"DD",X"7E",X"00",
		X"FE",X"49",X"28",X"09",X"FE",X"4A",X"28",X"05",X"FE",X"4B",X"28",X"01",X"C9",X"3E",X"1F",X"FD",
		X"77",X"00",X"C9",X"3E",X"E0",X"FD",X"77",X"00",X"3E",X"3F",X"FD",X"77",X"08",X"3A",X"0D",X"60",
		X"FE",X"05",X"C0",X"CD",X"77",X"EA",X"CD",X"77",X"EA",X"CD",X"77",X"EA",X"CD",X"77",X"EA",X"CD",
		X"77",X"EA",X"C9",X"3A",X"F5",X"62",X"FE",X"01",X"C0",X"3A",X"34",X"63",X"FE",X"01",X"C8",X"3A",
		X"FA",X"62",X"FE",X"00",X"28",X"05",X"3D",X"32",X"FA",X"62",X"C9",X"FD",X"2A",X"F6",X"62",X"2A",
		X"F8",X"62",X"FD",X"7E",X"00",X"77",X"CD",X"AC",X"DE",X"11",X"E0",X"FF",X"19",X"FD",X"23",X"FD",
		X"7E",X"00",X"77",X"CD",X"AC",X"DE",X"19",X"FD",X"23",X"FD",X"7E",X"00",X"77",X"CD",X"AC",X"DE",
		X"19",X"FD",X"23",X"FD",X"7E",X"00",X"77",X"CD",X"AC",X"DE",X"FD",X"23",X"11",X"61",X"00",X"19",
		X"FD",X"7E",X"00",X"77",X"CD",X"AC",X"DE",X"FD",X"23",X"11",X"E0",X"FF",X"19",X"FD",X"7E",X"00",
		X"77",X"CD",X"AC",X"DE",X"FD",X"23",X"19",X"FD",X"7E",X"00",X"77",X"CD",X"AC",X"DE",X"FD",X"23",
		X"FD",X"7E",X"00",X"19",X"77",X"CD",X"AC",X"DE",X"FD",X"23",X"FD",X"22",X"F6",X"62",X"3E",X"03",
		X"32",X"FA",X"62",X"FD",X"7E",X"00",X"FE",X"FF",X"C0",X"AF",X"32",X"F5",X"62",X"FD",X"2A",X"F8",
		X"62",X"DD",X"21",X"FC",X"62",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"FD",X"77",
		X"01",X"DD",X"7E",X"02",X"FD",X"77",X"E0",X"DD",X"7E",X"03",X"FD",X"77",X"E1",X"DD",X"7E",X"04",
		X"FD",X"77",X"C0",X"DD",X"7E",X"05",X"FD",X"77",X"C1",X"DD",X"7E",X"06",X"FD",X"77",X"A0",X"DD",
		X"7E",X"07",X"FD",X"77",X"A1",X"FD",X"2A",X"F8",X"62",X"11",X"00",X"08",X"FD",X"19",X"DD",X"21",
		X"04",X"63",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"DD",X"7E",
		X"02",X"FD",X"77",X"E0",X"DD",X"7E",X"03",X"FD",X"77",X"E1",X"DD",X"7E",X"04",X"FD",X"77",X"C0",
		X"DD",X"7E",X"05",X"FD",X"77",X"C1",X"DD",X"7E",X"06",X"FD",X"77",X"A0",X"DD",X"7E",X"07",X"FD",
		X"77",X"A1",X"3A",X"36",X"63",X"FE",X"01",X"20",X"03",X"32",X"25",X"60",X"3A",X"37",X"63",X"FE",
		X"01",X"20",X"03",X"32",X"9F",X"62",X"3A",X"38",X"63",X"FE",X"01",X"20",X"03",X"32",X"A7",X"62",
		X"AF",X"32",X"36",X"63",X"32",X"37",X"63",X"32",X"38",X"63",X"C9",X"2A",X"F8",X"62",X"CD",X"64",
		X"EB",X"FD",X"21",X"36",X"63",X"DD",X"21",X"80",X"65",X"CD",X"4E",X"EB",X"FD",X"7E",X"00",X"FE",
		X"01",X"20",X"08",X"3E",X"01",X"32",X"60",X"61",X"CD",X"99",X"E3",X"FD",X"21",X"37",X"63",X"DD",
		X"21",X"94",X"65",X"CD",X"4E",X"EB",X"FD",X"7E",X"00",X"FE",X"01",X"CC",X"21",X"E3",X"FD",X"21",
		X"38",X"63",X"DD",X"21",X"98",X"65",X"CD",X"4E",X"EB",X"FD",X"7E",X"00",X"FE",X"01",X"CC",X"7D",
		X"E3",X"C9",X"3A",X"0D",X"60",X"D5",X"47",X"11",X"A6",X"DE",X"13",X"10",X"FD",X"1A",X"47",X"7C",
		X"90",X"67",X"D1",X"C9",X"3A",X"0D",X"60",X"D5",X"47",X"11",X"A6",X"DE",X"13",X"10",X"FD",X"1A",
		X"47",X"7C",X"80",X"67",X"D1",X"C9",X"00",X"50",X"4C",X"48",X"60",X"5C",X"E5",X"7C",X"C6",X"08",
		X"67",X"3E",X"38",X"77",X"E1",X"C9",X"E0",X"7D",X"7C",X"7B",X"E0",X"79",X"78",X"77",X"76",X"75",
		X"74",X"73",X"72",X"71",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"69",X"68",X"67",X"6E",X"6D",
		X"6C",X"6B",X"6A",X"69",X"68",X"67",X"76",X"75",X"74",X"73",X"72",X"71",X"70",X"6F",X"76",X"75",
		X"74",X"73",X"72",X"71",X"70",X"6F",X"E0",X"7D",X"7C",X"7B",X"E0",X"79",X"78",X"77",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"3A",X"43",X"63",X"FE",X"01",X"C8",X"3A",X"F0",X"62",
		X"3C",X"32",X"F0",X"62",X"FE",X"0C",X"C0",X"AF",X"32",X"F0",X"62",X"3A",X"0D",X"60",X"FE",X"02",
		X"C0",X"2A",X"F1",X"62",X"23",X"22",X"F1",X"62",X"7E",X"FE",X"FF",X"20",X"07",X"21",X"2D",X"DF",
		X"22",X"F1",X"62",X"7E",X"32",X"8E",X"93",X"3E",X"08",X"32",X"8E",X"9B",X"C9",X"78",X"7C",X"74",
		X"72",X"6E",X"6A",X"76",X"7E",X"7A",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"FF",X"DD",X"21",X"80",X"65",X"FD",X"21",X"E5",X"62",X"3A",X"0D",X"60",X"CD",X"6D",X"DF",
		X"DD",X"21",X"94",X"65",X"FD",X"21",X"E9",X"62",X"3A",X"99",X"60",X"CD",X"6D",X"DF",X"DD",X"21",
		X"98",X"65",X"FD",X"21",X"ED",X"62",X"3A",X"9A",X"60",X"CD",X"6D",X"DF",X"C9",X"47",X"DD",X"7E",
		X"02",X"FE",X"A9",X"38",X"13",X"78",X"FE",X"05",X"20",X"0E",X"3A",X"E3",X"62",X"DD",X"BE",X"03",
		X"20",X"06",X"3E",X"01",X"FD",X"77",X"00",X"C9",X"AF",X"FD",X"77",X"00",X"C9",X"21",X"C7",X"90",
		X"22",X"DD",X"62",X"21",X"04",X"E0",X"22",X"DB",X"62",X"3E",X"BB",X"32",X"E0",X"62",X"3E",X"FF",
		X"32",X"DF",X"62",X"3E",X"28",X"32",X"E3",X"62",X"3A",X"0D",X"60",X"FE",X"05",X"C0",X"3E",X"B2",
		X"32",X"C6",X"90",X"32",X"06",X"91",X"3E",X"B3",X"32",X"E6",X"90",X"32",X"26",X"91",X"C9",X"CD",
		X"8D",X"DF",X"21",X"2D",X"DF",X"22",X"F1",X"62",X"21",X"63",X"92",X"22",X"0E",X"63",X"3E",X"01",
		X"32",X"10",X"63",X"21",X"3C",X"91",X"22",X"15",X"63",X"3E",X"02",X"32",X"17",X"63",X"21",X"54",
		X"92",X"22",X"18",X"63",X"3E",X"03",X"32",X"1A",X"63",X"21",X"2E",X"91",X"22",X"1B",X"63",X"3E",
		X"04",X"32",X"1D",X"63",X"21",X"7C",X"92",X"22",X"1E",X"63",X"3E",X"05",X"32",X"20",X"63",X"CD",
		X"8C",X"E5",X"C9",X"FE",X"AC",X"A8",X"A4",X"A0",X"9C",X"98",X"94",X"90",X"AE",X"AA",X"A6",X"A2",
		X"9E",X"9A",X"96",X"92",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"8D",X"DF",X"2A",X"DD",X"62",X"7D",
		X"FE",X"C7",X"38",X"F5",X"FE",X"DE",X"30",X"F1",X"3A",X"E1",X"62",X"FE",X"00",X"28",X"05",X"3D",
		X"32",X"E1",X"62",X"C9",X"3A",X"DF",X"62",X"FE",X"00",X"C8",X"47",X"3A",X"E3",X"62",X"90",X"32",
		X"E3",X"62",X"47",X"3A",X"E5",X"62",X"FE",X"00",X"28",X"04",X"78",X"32",X"83",X"65",X"3A",X"E9",
		X"62",X"FE",X"00",X"28",X"04",X"78",X"32",X"97",X"65",X"3A",X"ED",X"62",X"FE",X"00",X"28",X"04",
		X"78",X"32",X"9B",X"65",X"3A",X"DF",X"62",X"47",X"2A",X"DD",X"62",X"CD",X"88",X"E1",X"DD",X"2A",
		X"DB",X"62",X"3A",X"DF",X"62",X"FE",X"FF",X"DD",X"7E",X"12",X"28",X"03",X"DD",X"7E",X"24",X"FE",
		X"01",X"CC",X"C7",X"E0",X"DD",X"2A",X"DB",X"62",X"2A",X"DD",X"62",X"DD",X"7E",X"00",X"CD",X"F7",
		X"E0",X"CD",X"72",X"E1",X"2A",X"DB",X"62",X"CD",X"EC",X"E0",X"22",X"DB",X"62",X"2A",X"DD",X"62",
		X"CD",X"37",X"E1",X"CD",X"51",X"E1",X"C9",X"DD",X"7E",X"00",X"FE",X"FF",X"CC",X"DE",X"E0",X"FE",
		X"FE",X"CC",X"E5",X"E0",X"2A",X"DD",X"62",X"CD",X"EC",X"E0",X"22",X"DD",X"62",X"C9",X"21",X"04",
		X"E0",X"22",X"DB",X"62",X"C9",X"21",X"13",X"E0",X"22",X"DB",X"62",X"C9",X"3A",X"DF",X"62",X"FE",
		X"FF",X"28",X"02",X"2B",X"C9",X"23",X"C9",X"F5",X"FE",X"AE",X"28",X"0E",X"FE",X"AC",X"28",X"0A",
		X"FE",X"90",X"28",X"27",X"FE",X"92",X"28",X"23",X"18",X"2B",X"7D",X"1E",X"49",X"FE",X"CB",X"CC",
		X"AA",X"E1",X"1E",X"71",X"FE",X"D0",X"CC",X"AA",X"E1",X"1E",X"99",X"FE",X"D5",X"CC",X"AA",X"E1",
		X"1E",X"29",X"FE",X"C7",X"20",X"0F",X"CD",X"AA",X"E1",X"18",X"0A",X"7D",X"1E",X"E0",X"FE",X"DD",
		X"20",X"03",X"CD",X"AA",X"E1",X"F1",X"C9",X"3A",X"DF",X"62",X"FE",X"01",X"C0",X"7D",X"FE",X"C7",
		X"C0",X"DD",X"7E",X"00",X"FE",X"AC",X"C0",X"2A",X"DB",X"62",X"23",X"23",X"22",X"DB",X"62",X"18",
		X"18",X"3A",X"DF",X"62",X"FE",X"FF",X"C0",X"7D",X"FE",X"DD",X"C0",X"DD",X"7E",X"00",X"FE",X"90",
		X"C0",X"2A",X"DB",X"62",X"2B",X"2B",X"22",X"DB",X"62",X"3A",X"DF",X"62",X"2F",X"3C",X"32",X"DF",
		X"62",X"C9",X"08",X"3A",X"0D",X"60",X"FE",X"05",X"C0",X"08",X"77",X"11",X"20",X"00",X"19",X"3C",
		X"77",X"19",X"3D",X"77",X"19",X"3C",X"77",X"C9",X"3A",X"0D",X"60",X"FE",X"05",X"C0",X"CD",X"A1",
		X"E1",X"11",X"20",X"00",X"19",X"CD",X"A1",X"E1",X"19",X"CD",X"A1",X"E1",X"19",X"CD",X"A1",X"E1",
		X"C9",X"E5",X"C1",X"78",X"D6",X"5C",X"47",X"0A",X"77",X"C9",X"3E",X"50",X"32",X"E1",X"62",X"7B",
		X"32",X"E3",X"62",X"C9",X"DD",X"21",X"80",X"65",X"FD",X"21",X"D2",X"62",X"CD",X"D8",X"E1",X"C9",
		X"DD",X"21",X"94",X"65",X"FD",X"21",X"D6",X"62",X"CD",X"D8",X"E1",X"C9",X"DD",X"21",X"98",X"65",
		X"FD",X"21",X"DA",X"62",X"CD",X"D8",X"E1",X"C9",X"FD",X"7E",X"00",X"FE",X"01",X"C0",X"DD",X"7E",
		X"02",X"3C",X"DD",X"77",X"02",X"DD",X"7E",X"03",X"3C",X"DD",X"77",X"03",X"C9",X"DD",X"21",X"80",
		X"65",X"FD",X"21",X"D2",X"62",X"11",X"0D",X"60",X"06",X"1C",X"3A",X"08",X"60",X"FE",X"01",X"28",
		X"08",X"3A",X"BD",X"62",X"FE",X"01",X"C4",X"64",X"E2",X"CD",X"43",X"E2",X"C9",X"DD",X"21",X"94",
		X"65",X"FD",X"21",X"D6",X"62",X"11",X"99",X"60",X"3A",X"37",X"60",X"FE",X"01",X"28",X"05",X"06",
		X"3F",X"CD",X"64",X"E2",X"CD",X"43",X"E2",X"C9",X"DD",X"21",X"98",X"65",X"FD",X"21",X"DA",X"62",
		X"11",X"9A",X"60",X"06",X"3F",X"3A",X"77",X"60",X"FE",X"01",X"28",X"03",X"CD",X"64",X"E2",X"CD",
		X"43",X"E2",X"C9",X"FD",X"7E",X"00",X"FE",X"01",X"C0",X"1A",X"FE",X"03",X"28",X"0B",X"DD",X"7E",
		X"02",X"FE",X"81",X"D8",X"AF",X"FD",X"77",X"00",X"C9",X"DD",X"7E",X"02",X"FE",X"73",X"D8",X"AF",
		X"FD",X"77",X"00",X"C9",X"FD",X"7E",X"00",X"FE",X"01",X"C8",X"DD",X"7E",X"03",X"FE",X"38",X"20",
		X"24",X"1A",X"FE",X"02",X"C0",X"DD",X"7E",X"02",X"FE",X"50",X"D8",X"DD",X"7E",X"02",X"FE",X"55",
		X"D0",X"3E",X"01",X"FD",X"77",X"00",X"DD",X"7E",X"00",X"E6",X"80",X"B0",X"DD",X"77",X"00",X"3E",
		X"20",X"FD",X"77",X"01",X"C9",X"FE",X"50",X"20",X"0F",X"1A",X"FE",X"03",X"C0",X"DD",X"7E",X"02",
		X"FE",X"41",X"D8",X"FE",X"50",X"D0",X"18",X"D9",X"FE",X"53",X"D8",X"FE",X"70",X"D0",X"1A",X"FE",
		X"03",X"C0",X"DD",X"7E",X"02",X"FE",X"4B",X"D8",X"FE",X"60",X"D0",X"DD",X"7E",X"02",X"C6",X"10",
		X"DD",X"77",X"03",X"18",X"BC",X"11",X"99",X"60",X"DD",X"21",X"94",X"65",X"21",X"27",X"60",X"CD",
		X"EC",X"E2",X"78",X"FE",X"01",X"CC",X"21",X"E3",X"11",X"9A",X"60",X"DD",X"21",X"98",X"65",X"21",
		X"67",X"60",X"CD",X"EC",X"E2",X"78",X"FE",X"01",X"CC",X"7D",X"E3",X"C9",X"FD",X"21",X"2D",X"E3",
		X"06",X"00",X"1A",X"FD",X"BE",X"02",X"20",X"19",X"DD",X"7E",X"02",X"FD",X"BE",X"00",X"20",X"11",
		X"DD",X"7E",X"03",X"FD",X"BE",X"01",X"20",X"09",X"7E",X"FD",X"BE",X"03",X"20",X"03",X"06",X"01",
		X"C9",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"7E",X"00",X"FE",X"FF",X"C8",X"18",
		X"D1",X"DD",X"21",X"94",X"65",X"FD",X"21",X"C4",X"62",X"CD",X"87",X"E4",X"C9",X"92",X"C0",X"02",
		X"40",X"81",X"C0",X"02",X"80",X"5A",X"C0",X"02",X"40",X"49",X"C0",X"02",X"80",X"A2",X"68",X"02",
		X"40",X"90",X"68",X"02",X"80",X"92",X"80",X"03",X"40",X"7A",X"80",X"03",X"80",X"32",X"50",X"04",
		X"40",X"20",X"50",X"04",X"80",X"38",X"70",X"04",X"80",X"B8",X"18",X"04",X"80",X"B8",X"70",X"04",
		X"80",X"C2",X"18",X"04",X"40",X"C2",X"70",X"04",X"40",X"FF",X"FF",X"FF",X"FF",X"DD",X"21",X"94",
		X"65",X"FD",X"21",X"C4",X"62",X"ED",X"5B",X"38",X"60",X"CD",X"F0",X"E3",X"C9",X"DD",X"21",X"98",
		X"65",X"FD",X"21",X"CB",X"62",X"CD",X"87",X"E4",X"C9",X"DD",X"21",X"98",X"65",X"FD",X"21",X"CB",
		X"62",X"ED",X"5B",X"78",X"60",X"CD",X"F0",X"E3",X"C9",X"DD",X"21",X"80",X"65",X"FD",X"21",X"BD",
		X"62",X"3A",X"08",X"60",X"FE",X"00",X"C0",X"3A",X"1C",X"60",X"FE",X"01",X"C8",X"3A",X"2A",X"60",
		X"FE",X"01",X"C8",X"3A",X"60",X"61",X"FE",X"01",X"C0",X"3A",X"AF",X"62",X"FE",X"01",X"C8",X"3A",
		X"B0",X"62",X"FE",X"01",X"C8",X"CD",X"63",X"E4",X"C9",X"3A",X"BC",X"62",X"FE",X"01",X"20",X"08",
		X"AF",X"32",X"BC",X"62",X"CD",X"63",X"E4",X"C9",X"3A",X"BC",X"62",X"3C",X"32",X"BC",X"62",X"C9",
		X"DD",X"21",X"80",X"65",X"FD",X"21",X"BD",X"62",X"ED",X"5B",X"09",X"60",X"CD",X"F0",X"E3",X"C9",
		X"FD",X"7E",X"00",X"FE",X"00",X"C8",X"FD",X"66",X"01",X"FD",X"6E",X"02",X"7E",X"FE",X"FF",X"28",
		X"5D",X"DD",X"E5",X"FD",X"E5",X"E5",X"EB",X"FD",X"7E",X"03",X"FE",X"80",X"20",X"05",X"CD",X"CC",
		X"0D",X"18",X"03",X"CD",X"71",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"E1",X"FD",X"E1",X"DD",X"E1",
		X"20",X"3C",X"7E",X"47",X"FD",X"7E",X"03",X"B0",X"DD",X"77",X"00",X"23",X"7E",X"47",X"FD",X"7E",
		X"04",X"FE",X"00",X"28",X"05",X"3D",X"FD",X"77",X"04",X"04",X"FD",X"7E",X"03",X"FE",X"80",X"20",
		X"04",X"78",X"2F",X"3C",X"47",X"DD",X"7E",X"02",X"80",X"DD",X"77",X"02",X"23",X"7E",X"47",X"DD",
		X"7E",X"03",X"80",X"DD",X"77",X"03",X"23",X"FD",X"74",X"01",X"FD",X"75",X"02",X"C9",X"AF",X"FD",
		X"77",X"00",X"C9",X"CD",X"E3",X"F4",X"78",X"FE",X"01",X"C0",X"FD",X"7E",X"00",X"FE",X"00",X"C0",
		X"3E",X"01",X"FD",X"77",X"00",X"21",X"A4",X"E4",X"FD",X"74",X"01",X"FD",X"75",X"02",X"DD",X"7E",
		X"00",X"E6",X"80",X"FD",X"77",X"03",X"C9",X"FD",X"7E",X"00",X"FE",X"00",X"C0",X"3E",X"01",X"FD",
		X"77",X"00",X"21",X"01",X"E5",X"FD",X"74",X"01",X"FD",X"75",X"02",X"DD",X"7E",X"00",X"E6",X"80",
		X"FD",X"77",X"03",X"C9",X"1F",X"01",X"00",X"1F",X"00",X"00",X"1F",X"01",X"00",X"1F",X"00",X"00",
		X"1F",X"01",X"00",X"1F",X"00",X"00",X"1F",X"01",X"00",X"1D",X"00",X"00",X"1D",X"01",X"00",X"1D",
		X"00",X"00",X"1D",X"01",X"00",X"1D",X"00",X"00",X"1D",X"01",X"00",X"1D",X"00",X"00",X"1D",X"01",
		X"00",X"1E",X"00",X"00",X"1E",X"01",X"00",X"1E",X"01",X"00",X"1E",X"00",X"00",X"1E",X"01",X"00",
		X"1E",X"01",X"00",X"1E",X"01",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",
		X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"FF",X"FF",
		X"FF",X"2E",X"01",X"00",X"2E",X"01",X"00",X"2E",X"01",X"00",X"2E",X"01",X"00",X"2E",X"01",X"00",
		X"2E",X"01",X"00",X"2E",X"01",X"00",X"2F",X"01",X"00",X"2F",X"01",X"00",X"2F",X"01",X"00",X"2F",
		X"01",X"00",X"2F",X"01",X"00",X"2F",X"01",X"00",X"2F",X"01",X"00",X"2F",X"01",X"00",X"2F",X"00",
		X"00",X"2F",X"01",X"00",X"2F",X"01",X"00",X"2F",X"00",X"00",X"2F",X"01",X"00",X"30",X"01",X"00",
		X"30",X"01",X"00",X"30",X"00",X"00",X"31",X"00",X"00",X"31",X"00",X"00",X"31",X"00",X"00",X"31",
		X"00",X"00",X"31",X"00",X"00",X"31",X"00",X"00",X"31",X"00",X"00",X"FF",X"FF",X"FF",X"FE",X"01",
		X"20",X"04",X"7C",X"C6",X"50",X"C9",X"FE",X"02",X"20",X"04",X"7C",X"C6",X"4C",X"C9",X"FE",X"03",
		X"20",X"04",X"7C",X"C6",X"48",X"C9",X"FE",X"04",X"20",X"04",X"7C",X"C6",X"60",X"C9",X"FE",X"05",
		X"C0",X"7C",X"C6",X"5C",X"C9",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F9",X"AF",X"DD",X"21",X"93",
		X"62",X"06",X"24",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F9",X"AF",X"32",X"F5",X"62",X"32",X"F6",
		X"62",X"32",X"F7",X"62",X"32",X"F8",X"62",X"32",X"F9",X"62",X"32",X"FA",X"62",X"32",X"FB",X"62",
		X"32",X"23",X"63",X"32",X"24",X"63",X"32",X"26",X"63",X"32",X"27",X"63",X"32",X"E5",X"62",X"32",
		X"E9",X"62",X"32",X"EA",X"62",X"32",X"ED",X"62",X"32",X"EE",X"62",X"32",X"D2",X"62",X"CD",X"CC",
		X"F9",X"C9",X"06",X"00",X"3A",X"54",X"60",X"FE",X"00",X"28",X"30",X"3A",X"FD",X"61",X"FE",X"01",
		X"28",X"16",X"3A",X"50",X"60",X"E6",X"04",X"FE",X"04",X"28",X"0C",X"3A",X"26",X"60",X"E6",X"04",
		X"FE",X"04",X"20",X"03",X"06",X"01",X"C9",X"C9",X"3A",X"52",X"60",X"E6",X"04",X"FE",X"04",X"C8",
		X"3A",X"51",X"60",X"E6",X"04",X"FE",X"04",X"C0",X"06",X"01",X"C9",X"3A",X"50",X"60",X"E6",X"04",
		X"FE",X"04",X"C0",X"06",X"01",X"C9",X"11",X"95",X"62",X"CD",X"29",X"E6",X"11",X"9D",X"62",X"CD",
		X"29",X"E6",X"11",X"A5",X"62",X"CD",X"29",X"E6",X"C9",X"1A",X"FE",X"00",X"C8",X"3D",X"12",X"C9",
		X"3A",X"0D",X"60",X"FE",X"03",X"C0",X"DD",X"21",X"80",X"65",X"DD",X"7E",X"03",X"FE",X"A0",X"20",
		X"26",X"DD",X"7E",X"02",X"FE",X"58",X"38",X"1F",X"FE",X"60",X"30",X"1B",X"3E",X"01",X"32",X"93",
		X"62",X"3E",X"06",X"32",X"94",X"62",X"32",X"9C",X"62",X"32",X"A4",X"62",X"3E",X"E0",X"32",X"95",
		X"92",X"3E",X"3F",X"32",X"95",X"9A",X"C9",X"3A",X"94",X"62",X"FE",X"00",X"C0",X"3E",X"BD",X"32",
		X"95",X"92",X"3E",X"36",X"32",X"95",X"9A",X"C9",X"AF",X"32",X"46",X"63",X"C9",X"DD",X"21",X"98",
		X"65",X"FD",X"21",X"A3",X"62",X"3A",X"99",X"62",X"FE",X"01",X"C0",X"3A",X"97",X"62",X"FE",X"01",
		X"C8",X"3A",X"A4",X"62",X"FE",X"00",X"C8",X"CD",X"53",X"E8",X"78",X"FE",X"01",X"C8",X"3A",X"7C",
		X"60",X"FE",X"80",X"20",X"0A",X"DD",X"7E",X"00",X"E6",X"80",X"FE",X"00",X"C0",X"18",X"08",X"DD",
		X"7E",X"00",X"E6",X"80",X"FE",X"00",X"C8",X"3A",X"9A",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"C0",
		X"3A",X"57",X"61",X"FE",X"00",X"20",X"B1",X"3A",X"46",X"63",X"FE",X"0F",X"38",X"10",X"0E",X"28",
		X"DD",X"7E",X"00",X"E6",X"80",X"B1",X"DD",X"77",X"00",X"3E",X"20",X"FD",X"77",X"02",X"CD",X"2C",
		X"E8",X"3A",X"46",X"63",X"3C",X"32",X"46",X"63",X"B8",X"D8",X"AF",X"32",X"46",X"63",X"3E",X"28",
		X"4F",X"C3",X"B4",X"E7",X"AF",X"32",X"45",X"63",X"C9",X"DD",X"21",X"94",X"65",X"FD",X"21",X"9B",
		X"62",X"3A",X"99",X"62",X"FE",X"01",X"C0",X"3A",X"97",X"62",X"FE",X"01",X"C8",X"3A",X"9C",X"62",
		X"FE",X"00",X"C8",X"CD",X"53",X"E8",X"78",X"FE",X"01",X"C8",X"3A",X"3C",X"60",X"FE",X"80",X"20",
		X"0A",X"DD",X"7E",X"00",X"E6",X"80",X"FE",X"00",X"C0",X"18",X"08",X"DD",X"7E",X"00",X"E6",X"80",
		X"FE",X"00",X"C8",X"3A",X"99",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"C0",X"3A",X"56",X"61",X"FE",
		X"00",X"20",X"B1",X"3A",X"45",X"63",X"FE",X"0F",X"38",X"10",X"0E",X"28",X"DD",X"7E",X"00",X"E6",
		X"80",X"B1",X"DD",X"77",X"00",X"3E",X"20",X"FD",X"77",X"02",X"CD",X"2C",X"E8",X"3A",X"45",X"63",
		X"3C",X"32",X"45",X"63",X"B8",X"D8",X"AF",X"32",X"45",X"63",X"3E",X"28",X"4F",X"18",X"45",X"3A",
		X"93",X"62",X"FE",X"01",X"C0",X"3E",X"BD",X"32",X"1F",X"92",X"3E",X"35",X"32",X"1F",X"9A",X"3A",
		X"94",X"62",X"FE",X"00",X"20",X"05",X"3E",X"E0",X"32",X"1F",X"92",X"3A",X"52",X"63",X"C6",X"04",
		X"32",X"52",X"63",X"FE",X"80",X"38",X"05",X"3E",X"E0",X"32",X"1F",X"92",X"3A",X"97",X"62",X"FE",
		X"00",X"C0",X"CD",X"D2",X"E5",X"78",X"FE",X"00",X"C8",X"3E",X"11",X"4F",X"DD",X"21",X"80",X"65",
		X"FD",X"21",X"93",X"62",X"FD",X"7E",X"01",X"FE",X"00",X"C8",X"FD",X"7E",X"01",X"3D",X"FD",X"77",
		X"01",X"3E",X"01",X"32",X"97",X"62",X"06",X"01",X"DD",X"7E",X"00",X"E6",X"80",X"FE",X"80",X"20",
		X"02",X"06",X"FF",X"78",X"32",X"98",X"62",X"DD",X"7E",X"00",X"E6",X"80",X"B1",X"DD",X"77",X"00",
		X"DD",X"7E",X"02",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"32",X"8E",
		X"65",X"DD",X"7E",X"03",X"32",X"8F",X"65",X"3E",X"10",X"32",X"8C",X"65",X"3E",X"0F",X"32",X"8D",
		X"65",X"3E",X"30",X"FD",X"77",X"02",X"3A",X"48",X"63",X"FE",X"01",X"C8",X"3A",X"54",X"60",X"FE",
		X"00",X"C8",X"21",X"28",X"54",X"22",X"4E",X"63",X"AF",X"32",X"42",X"61",X"3E",X"02",X"32",X"48",
		X"63",X"3E",X"0F",X"32",X"4C",X"63",X"3E",X"01",X"32",X"4D",X"63",X"C9",X"3A",X"64",X"61",X"06",
		X"18",X"C9",X"06",X"38",X"FE",X"00",X"C8",X"06",X"30",X"FE",X"01",X"C8",X"06",X"28",X"FE",X"02",
		X"C8",X"06",X"20",X"FE",X"03",X"C8",X"06",X"18",X"FE",X"04",X"C8",X"06",X"10",X"FE",X"05",X"C8",
		X"06",X"08",X"C9",X"DD",X"7E",X"02",X"06",X"01",X"FE",X"D8",X"D0",X"FE",X"18",X"D8",X"06",X"00",
		X"C9",X"3A",X"97",X"62",X"FE",X"01",X"C0",X"18",X"1F",X"3A",X"97",X"62",X"FE",X"01",X"C0",X"3A",
		X"ED",X"61",X"FE",X"01",X"C8",X"CD",X"CB",X"EA",X"11",X"1F",X"00",X"19",X"7E",X"CD",X"05",X"0E",
		X"3A",X"0B",X"60",X"FE",X"02",X"C2",X"14",X"E9",X"3A",X"8E",X"65",X"FE",X"10",X"DA",X"14",X"E9",
		X"FE",X"F0",X"D2",X"14",X"E9",X"DD",X"E5",X"3A",X"0D",X"60",X"32",X"98",X"60",X"DD",X"21",X"80",
		X"65",X"21",X"25",X"60",X"11",X"25",X"60",X"CD",X"DE",X"E8",X"3A",X"99",X"60",X"32",X"98",X"60",
		X"DD",X"21",X"94",X"65",X"21",X"9F",X"62",X"11",X"56",X"61",X"CD",X"DE",X"E8",X"3A",X"9A",X"60",
		X"32",X"98",X"60",X"DD",X"21",X"98",X"65",X"21",X"A7",X"62",X"11",X"57",X"61",X"CD",X"DE",X"E8",
		X"DD",X"E1",X"3A",X"98",X"62",X"47",X"3A",X"8E",X"65",X"80",X"32",X"8E",X"65",X"C9",X"3A",X"98",
		X"60",X"47",X"3A",X"0D",X"60",X"B8",X"C0",X"1A",X"FE",X"01",X"C8",X"DD",X"7E",X"02",X"D6",X"08",
		X"47",X"C6",X"10",X"4F",X"3A",X"8E",X"65",X"B8",X"D8",X"B9",X"D0",X"3A",X"8F",X"65",X"C6",X"07",
		X"47",X"D6",X"0E",X"4F",X"DD",X"7E",X"03",X"B8",X"D0",X"B9",X"D8",X"3E",X"01",X"77",X"32",X"99",
		X"62",X"18",X"01",X"C9",X"AF",X"32",X"97",X"62",X"32",X"8F",X"65",X"C9",X"DD",X"21",X"80",X"65",
		X"FD",X"21",X"AF",X"62",X"3A",X"0D",X"60",X"CD",X"4F",X"E9",X"DD",X"21",X"94",X"65",X"FD",X"21",
		X"B5",X"62",X"3A",X"99",X"60",X"CD",X"4F",X"E9",X"DD",X"21",X"98",X"65",X"FD",X"21",X"B9",X"62",
		X"3A",X"9A",X"60",X"CD",X"4F",X"E9",X"C9",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"C9",X"FE",
		X"01",X"20",X"F4",X"CD",X"7C",X"E9",X"CD",X"BF",X"E9",X"CD",X"9E",X"E9",X"FD",X"7E",X"00",X"FE",
		X"00",X"C8",X"FD",X"7E",X"01",X"FE",X"01",X"28",X"0B",X"F3",X"DD",X"7E",X"03",X"FE",X"39",X"38",
		X"03",X"DD",X"35",X"03",X"DD",X"34",X"02",X"DD",X"34",X"02",X"FB",X"C9",X"DD",X"7E",X"02",X"FE",
		X"48",X"D8",X"FE",X"50",X"D0",X"DD",X"7E",X"03",X"FE",X"70",X"C0",X"3A",X"AD",X"62",X"FE",X"00",
		X"C0",X"3E",X"01",X"FD",X"77",X"00",X"DD",X"7E",X"03",X"3C",X"DD",X"77",X"03",X"C9",X"DD",X"7E",
		X"02",X"FE",X"B8",X"D8",X"FE",X"C0",X"D0",X"DD",X"7E",X"03",X"FE",X"38",X"28",X"08",X"FE",X"37",
		X"C0",X"3E",X"38",X"DD",X"77",X"03",X"3E",X"01",X"FD",X"77",X"00",X"FD",X"77",X"01",X"C9",X"FD",
		X"7E",X"00",X"FE",X"01",X"C0",X"DD",X"7E",X"03",X"FE",X"39",X"D0",X"AF",X"FD",X"77",X"00",X"FD",
		X"77",X"01",X"C9",X"3A",X"AC",X"62",X"FE",X"03",X"D8",X"AF",X"32",X"AC",X"62",X"3A",X"0D",X"60",
		X"FE",X"01",X"C0",X"3A",X"ED",X"61",X"FE",X"01",X"C8",X"DD",X"21",X"87",X"1B",X"ED",X"5B",X"AD",
		X"62",X"DD",X"19",X"21",X"D0",X"92",X"CD",X"3C",X"EA",X"DD",X"21",X"87",X"1B",X"DD",X"19",X"21",
		X"8F",X"92",X"CD",X"3C",X"EA",X"21",X"4E",X"92",X"CD",X"3C",X"EA",X"21",X"0D",X"92",X"CD",X"3C",
		X"EA",X"21",X"CC",X"91",X"CD",X"3C",X"EA",X"21",X"8B",X"91",X"CD",X"3C",X"EA",X"21",X"4A",X"91",
		X"CD",X"3C",X"EA",X"D5",X"CD",X"1C",X"E9",X"D1",X"13",X"13",X"13",X"13",X"ED",X"53",X"AD",X"62",
		X"7B",X"FE",X"20",X"D8",X"11",X"00",X"00",X"ED",X"53",X"AD",X"62",X"C9",X"DD",X"7E",X"00",X"77",
		X"2B",X"DD",X"7E",X"02",X"77",X"D5",X"11",X"E0",X"FF",X"19",X"D1",X"DD",X"7E",X"03",X"77",X"23",
		X"DD",X"7E",X"01",X"77",X"C9",X"3A",X"0D",X"60",X"FE",X"05",X"C0",X"3A",X"83",X"65",X"FE",X"98",
		X"C0",X"3A",X"82",X"65",X"FE",X"88",X"C0",X"3A",X"CF",X"61",X"FE",X"00",X"C8",X"3A",X"9C",X"65",
		X"FE",X"B8",X"28",X"03",X"FE",X"B7",X"C0",X"3A",X"F3",X"91",X"FE",X"E0",X"C8",X"FE",X"E6",X"C8",
		X"FE",X"E4",X"C8",X"FE",X"D0",X"C8",X"3A",X"F3",X"91",X"FE",X"02",X"28",X"0B",X"3D",X"3D",X"32",
		X"F3",X"91",X"3D",X"32",X"F4",X"91",X"18",X"08",X"3E",X"E0",X"32",X"F3",X"91",X"32",X"F4",X"91",
		X"3A",X"F3",X"91",X"32",X"7D",X"62",X"C9",X"DD",X"21",X"80",X"65",X"FD",X"21",X"09",X"60",X"18",
		X"34",X"DD",X"21",X"94",X"65",X"FD",X"21",X"38",X"60",X"3A",X"99",X"60",X"18",X"2A",X"DD",X"21",
		X"98",X"65",X"FD",X"21",X"78",X"60",X"3A",X"9A",X"60",X"18",X"1D",X"DD",X"21",X"8C",X"65",X"FD",
		X"21",X"B2",X"62",X"3A",X"0D",X"60",X"18",X"10",X"DD",X"21",X"9C",X"65",X"FD",X"21",X"5A",X"61",
		X"3A",X"0D",X"60",X"18",X"03",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",X"EF",X"EA",X"C9",X"CD",
		X"0E",X"EB",X"CD",X"FC",X"EA",X"FD",X"75",X"00",X"FD",X"74",X"01",X"C9",X"DD",X"7E",X"03",X"C6",
		X"10",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"C9",X"DD",X"7E",
		X"02",X"C6",X"07",X"2F",X"E6",X"F8",X"26",X"00",X"6F",X"CB",X"25",X"CB",X"14",X"CB",X"25",X"CB",
		X"14",X"7C",X"F6",X"40",X"67",X"3A",X"98",X"60",X"FE",X"01",X"C8",X"FE",X"02",X"20",X"05",X"7C",
		X"C6",X"04",X"67",X"C9",X"FE",X"03",X"20",X"05",X"7C",X"C6",X"08",X"67",X"C9",X"FE",X"04",X"20",
		X"05",X"7C",X"D6",X"10",X"67",X"C9",X"FE",X"05",X"C0",X"7C",X"D6",X"0C",X"67",X"C9",X"DD",X"7E",
		X"02",X"B8",X"D8",X"B9",X"D0",X"D9",X"DD",X"7E",X"03",X"B8",X"D8",X"B9",X"D0",X"D9",X"3E",X"01",
		X"FD",X"77",X"00",X"C9",X"7D",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"D6",X"08",X"47",X"C6",X"10",
		X"4F",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"7D",X"D9",X"E6",X"F8",X"C6",X"07",X"2F",
		X"D6",X"08",X"47",X"C6",X"25",X"4F",X"C9",X"06",X"50",X"FE",X"01",X"C8",X"06",X"4C",X"FE",X"02",
		X"C8",X"06",X"48",X"FE",X"03",X"C8",X"06",X"60",X"FE",X"04",X"C8",X"06",X"5C",X"C9",X"3A",X"C7",
		X"61",X"FE",X"01",X"C0",X"CD",X"E9",X"EB",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"3A",X"9E",X"65",
		X"D6",X"20",X"32",X"9E",X"65",X"CD",X"E9",X"EB",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"3A",X"9E",
		X"65",X"D6",X"08",X"32",X"9E",X"65",X"CD",X"E9",X"EB",X"3A",X"C7",X"61",X"FE",X"01",X"C0",X"3A",
		X"9E",X"65",X"D6",X"08",X"32",X"9E",X"65",X"CD",X"E9",X"EB",X"3A",X"C7",X"61",X"FE",X"01",X"C0",
		X"3A",X"9E",X"65",X"C6",X"30",X"32",X"9E",X"65",X"C9",X"C5",X"FD",X"E5",X"01",X"C7",X"61",X"D9",
		X"FD",X"21",X"C4",X"61",X"3E",X"28",X"FD",X"77",X"05",X"3E",X"EC",X"FD",X"77",X"06",X"CD",X"55",
		X"FC",X"FD",X"E1",X"C1",X"C9",X"3A",X"41",X"63",X"FE",X"01",X"28",X"14",X"23",X"7E",X"FE",X"ED",
		X"C8",X"FE",X"EF",X"C8",X"7D",X"C6",X"20",X"6F",X"7C",X"CE",X"00",X"67",X"7E",X"FE",X"ED",X"C9",
		X"23",X"7E",X"FE",X"BF",X"C8",X"D5",X"11",X"20",X"00",X"19",X"7E",X"FE",X"BF",X"28",X"06",X"19",
		X"7E",X"FE",X"BF",X"28",X"00",X"D1",X"C9",X"3A",X"83",X"65",X"D6",X"02",X"32",X"9F",X"65",X"3A",
		X"80",X"65",X"E6",X"7F",X"FE",X"12",X"C8",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",X"28",X"0E",
		X"3A",X"82",X"65",X"C6",X"08",X"32",X"9E",X"65",X"3E",X"31",X"32",X"9C",X"65",X"C9",X"3A",X"82",
		X"65",X"D6",X"08",X"32",X"9E",X"65",X"3E",X"B1",X"32",X"9C",X"65",X"C9",X"21",X"6E",X"92",X"11",
		X"A1",X"56",X"CD",X"67",X"CA",X"C9",X"06",X"18",X"21",X"00",X"30",X"2B",X"7C",X"FE",X"00",X"20",
		X"FA",X"10",X"F5",X"C9",X"3A",X"10",X"62",X"FE",X"01",X"28",X"0F",X"3A",X"54",X"60",X"FE",X"01",
		X"28",X"08",X"3A",X"00",X"B0",X"E6",X"40",X"FE",X"40",X"C0",X"11",X"BD",X"61",X"01",X"06",X"00",
		X"ED",X"B0",X"3E",X"01",X"32",X"F3",X"61",X"C9",X"AF",X"32",X"00",X"A0",X"F3",X"3C",X"C3",X"00",
		X"C0",X"21",X"00",X"05",X"CD",X"D9",X"C5",X"3E",X"01",X"CD",X"E2",X"D8",X"3E",X"40",X"32",X"E8",
		X"61",X"CD",X"18",X"12",X"CD",X"DB",X"CF",X"CD",X"E7",X"CF",X"21",X"3C",X"51",X"22",X"40",X"61",
		X"22",X"4E",X"63",X"3E",X"38",X"32",X"4D",X"63",X"AF",X"32",X"48",X"63",X"F3",X"3A",X"00",X"B8",
		X"CD",X"51",X"F9",X"CD",X"14",X"C3",X"AF",X"32",X"25",X"60",X"3C",X"32",X"9A",X"60",X"3E",X"03",
		X"32",X"99",X"60",X"CD",X"BF",X"DF",X"CD",X"A9",X"D7",X"3E",X"01",X"ED",X"56",X"32",X"00",X"A0",
		X"FB",X"3A",X"00",X"A8",X"CD",X"34",X"CF",X"CD",X"2E",X"C0",X"DD",X"21",X"80",X"65",X"FD",X"21",
		X"94",X"65",X"11",X"04",X"00",X"3A",X"0D",X"60",X"47",X"3A",X"99",X"60",X"B8",X"20",X"13",X"CD",
		X"37",X"55",X"FE",X"00",X"28",X"0C",X"3A",X"56",X"61",X"FE",X"00",X"20",X"05",X"3E",X"01",X"32",
		X"25",X"60",X"DD",X"21",X"80",X"65",X"FD",X"21",X"98",X"65",X"11",X"04",X"00",X"3A",X"0D",X"60",
		X"47",X"3A",X"9A",X"60",X"B8",X"20",X"13",X"CD",X"37",X"55",X"FE",X"00",X"28",X"0C",X"3A",X"57",
		X"61",X"FE",X"00",X"20",X"05",X"3E",X"01",X"32",X"25",X"60",X"3A",X"54",X"60",X"FE",X"01",X"28",
		X"64",X"3E",X"01",X"CD",X"E2",X"D8",X"3A",X"53",X"60",X"FE",X"01",X"20",X"58",X"3A",X"10",X"62",
		X"FE",X"01",X"28",X"51",X"F3",X"3A",X"55",X"60",X"FE",X"01",X"28",X"23",X"3A",X"00",X"B8",X"CD",
		X"E3",X"C3",X"CD",X"A4",X"F8",X"CD",X"2E",X"16",X"21",X"68",X"5B",X"22",X"40",X"61",X"AF",X"32",
		X"42",X"61",X"3E",X"01",X"32",X"55",X"60",X"3A",X"54",X"60",X"FE",X"01",X"CA",X"F9",X"EC",X"3A",
		X"10",X"62",X"FE",X"01",X"28",X"1F",X"3A",X"00",X"60",X"FE",X"01",X"20",X"0C",X"11",X"DF",X"56",
		X"21",X"11",X"93",X"CD",X"67",X"CA",X"C3",X"F9",X"EC",X"11",X"F2",X"56",X"21",X"11",X"93",X"CD",
		X"67",X"CA",X"C3",X"F9",X"EC",X"CD",X"F7",X"F8",X"FE",X"01",X"CA",X"DC",X"EC",X"3A",X"E8",X"61",
		X"FE",X"00",X"20",X"08",X"CD",X"2D",X"F9",X"FE",X"01",X"CA",X"DC",X"EC",X"CD",X"37",X"F9",X"32",
		X"00",X"B8",X"CD",X"F2",X"F6",X"3A",X"A3",X"58",X"32",X"73",X"62",X"3A",X"00",X"B8",X"3A",X"0D",
		X"60",X"47",X"3A",X"99",X"60",X"B8",X"CC",X"6D",X"F6",X"FB",X"CD",X"8B",X"F7",X"3A",X"0F",X"57",
		X"32",X"70",X"62",X"3A",X"00",X"B8",X"3A",X"00",X"B8",X"3A",X"0D",X"60",X"47",X"3A",X"9A",X"60",
		X"B8",X"CC",X"56",X"F7",X"FB",X"32",X"00",X"B0",X"3A",X"99",X"60",X"32",X"98",X"60",X"FD",X"21",
		X"94",X"65",X"FD",X"22",X"93",X"60",X"DD",X"21",X"27",X"60",X"DD",X"22",X"95",X"60",X"DD",X"21",
		X"35",X"60",X"FD",X"21",X"94",X"65",X"ED",X"5B",X"38",X"60",X"ED",X"53",X"91",X"60",X"3A",X"00",
		X"B8",X"CD",X"0B",X"F5",X"DD",X"21",X"3B",X"60",X"21",X"57",X"60",X"11",X"48",X"61",X"CD",X"2E",
		X"F4",X"3A",X"48",X"61",X"FE",X"00",X"20",X"2D",X"3A",X"57",X"60",X"FE",X"F0",X"D4",X"58",X"CB",
		X"FE",X"10",X"FD",X"21",X"94",X"65",X"FD",X"22",X"93",X"60",X"DD",X"21",X"27",X"60",X"DD",X"22",
		X"95",X"60",X"FD",X"21",X"94",X"65",X"ED",X"5B",X"38",X"60",X"ED",X"53",X"91",X"60",X"DD",X"21",
		X"35",X"60",X"D4",X"B8",X"FB",X"3A",X"9A",X"60",X"32",X"98",X"60",X"FD",X"21",X"98",X"65",X"FD",
		X"22",X"93",X"60",X"DD",X"21",X"67",X"60",X"DD",X"22",X"95",X"60",X"DD",X"21",X"75",X"60",X"FD",
		X"21",X"98",X"65",X"ED",X"5B",X"78",X"60",X"ED",X"53",X"91",X"60",X"3A",X"00",X"B8",X"3A",X"0C",
		X"57",X"32",X"71",X"62",X"CD",X"0B",X"F5",X"DD",X"21",X"7B",X"60",X"21",X"97",X"60",X"11",X"49",
		X"61",X"CD",X"2E",X"F4",X"3A",X"49",X"61",X"FE",X"00",X"20",X"2D",X"3A",X"97",X"60",X"FE",X"F0",
		X"D4",X"7D",X"CB",X"FE",X"10",X"FD",X"21",X"98",X"65",X"FD",X"22",X"93",X"60",X"DD",X"21",X"67",
		X"60",X"DD",X"22",X"95",X"60",X"FD",X"21",X"98",X"65",X"ED",X"5B",X"78",X"60",X"ED",X"53",X"91",
		X"60",X"DD",X"21",X"75",X"60",X"D4",X"B8",X"FB",X"FB",X"3A",X"ED",X"62",X"FE",X"01",X"28",X"10",
		X"2A",X"78",X"60",X"CD",X"8E",X"F1",X"CA",X"0B",X"EF",X"18",X"05",X"3E",X"01",X"32",X"77",X"60",
		X"2A",X"38",X"60",X"3A",X"E9",X"62",X"FE",X"01",X"28",X"0C",X"CD",X"8E",X"F1",X"28",X"02",X"18",
		X"05",X"3E",X"01",X"32",X"37",X"60",X"2A",X"38",X"60",X"FD",X"21",X"37",X"60",X"DD",X"21",X"94",
		X"65",X"CD",X"2A",X"C1",X"01",X"E0",X"FF",X"2A",X"38",X"60",X"DD",X"21",X"94",X"65",X"CD",X"98",
		X"C0",X"2A",X"78",X"60",X"FD",X"21",X"77",X"60",X"DD",X"21",X"98",X"65",X"CD",X"2A",X"C1",X"01",
		X"E0",X"FF",X"2A",X"78",X"60",X"DD",X"21",X"98",X"65",X"CD",X"98",X"C0",X"3A",X"00",X"B8",X"2A",
		X"09",X"60",X"FB",X"CD",X"8E",X"F1",X"28",X"0E",X"3A",X"4E",X"60",X"FE",X"01",X"28",X"0C",X"3E",
		X"00",X"32",X"08",X"60",X"18",X"05",X"3E",X"01",X"32",X"08",X"60",X"2A",X"09",X"60",X"FD",X"21",
		X"08",X"60",X"DD",X"21",X"80",X"65",X"CD",X"2A",X"C1",X"2A",X"09",X"60",X"DD",X"21",X"80",X"65",
		X"01",X"3A",X"63",X"CD",X"98",X"C0",X"3E",X"01",X"32",X"6F",X"62",X"3A",X"00",X"B8",X"CD",X"EB",
		X"CB",X"3E",X"00",X"32",X"6F",X"62",X"CD",X"2D",X"F8",X"FE",X"01",X"CA",X"DC",X"EC",X"DD",X"21",
		X"3C",X"60",X"06",X"04",X"DD",X"7E",X"00",X"FE",X"00",X"20",X"30",X"DD",X"23",X"10",X"F5",X"21",
		X"E9",X"62",X"22",X"3D",X"63",X"21",X"27",X"60",X"22",X"95",X"60",X"21",X"44",X"61",X"22",X"46",
		X"61",X"3A",X"99",X"60",X"32",X"98",X"60",X"DD",X"21",X"80",X"65",X"FD",X"21",X"94",X"65",X"ED",
		X"5B",X"38",X"60",X"21",X"3B",X"60",X"CD",X"BC",X"C4",X"18",X"04",X"AF",X"32",X"48",X"61",X"DD",
		X"21",X"7C",X"60",X"06",X"04",X"DD",X"7E",X"00",X"FE",X"00",X"20",X"30",X"DD",X"23",X"10",X"F5",
		X"21",X"ED",X"62",X"22",X"3D",X"63",X"21",X"67",X"60",X"22",X"95",X"60",X"21",X"45",X"61",X"22",
		X"46",X"61",X"3A",X"9A",X"60",X"32",X"98",X"60",X"DD",X"21",X"80",X"65",X"FD",X"21",X"98",X"65",
		X"ED",X"5B",X"78",X"60",X"21",X"7B",X"60",X"CD",X"BC",X"C4",X"18",X"04",X"AF",X"32",X"49",X"61",
		X"3A",X"60",X"61",X"32",X"2A",X"63",X"2A",X"09",X"60",X"CD",X"CB",X"F2",X"F3",X"CD",X"BD",X"DA",
		X"CD",X"3E",X"D7",X"28",X"03",X"CD",X"99",X"E3",X"FB",X"3A",X"CF",X"61",X"FE",X"00",X"28",X"27",
		X"3A",X"99",X"60",X"47",X"3A",X"70",X"62",X"B8",X"3A",X"0D",X"60",X"B8",X"20",X"19",X"DD",X"21",
		X"94",X"65",X"FD",X"21",X"9C",X"65",X"0E",X"00",X"06",X"06",X"CD",X"97",X"C4",X"FE",X"01",X"20",
		X"06",X"CD",X"F4",X"FC",X"CD",X"AD",X"CA",X"3A",X"9F",X"62",X"FE",X"01",X"CC",X"F4",X"FC",X"AF",
		X"32",X"9F",X"62",X"3A",X"CF",X"61",X"FE",X"00",X"28",X"23",X"DD",X"21",X"98",X"65",X"FD",X"21",
		X"9C",X"65",X"3A",X"9A",X"60",X"47",X"3A",X"0D",X"60",X"B8",X"20",X"11",X"0E",X"00",X"06",X"06",
		X"CD",X"97",X"C4",X"FE",X"01",X"20",X"06",X"CD",X"33",X"FD",X"CD",X"AD",X"CA",X"3A",X"A7",X"62",
		X"FE",X"01",X"CC",X"33",X"FD",X"AF",X"32",X"A7",X"62",X"DD",X"21",X"80",X"65",X"FD",X"21",X"84",
		X"65",X"CD",X"93",X"C4",X"FE",X"01",X"20",X"11",X"3E",X"01",X"32",X"25",X"60",X"AF",X"32",X"29",
		X"60",X"CD",X"2D",X"F8",X"FE",X"01",X"CA",X"DC",X"EC",X"FB",X"CD",X"EE",X"C5",X"CD",X"7E",X"D2",
		X"3A",X"ED",X"61",X"FE",X"00",X"CC",X"72",X"FD",X"3A",X"7C",X"60",X"47",X"3A",X"7D",X"60",X"B0",
		X"FE",X"00",X"C4",X"7D",X"E6",X"3A",X"3C",X"60",X"47",X"3A",X"3D",X"60",X"B0",X"FE",X"00",X"C4",
		X"F9",X"E6",X"CD",X"C5",X"E2",X"CD",X"ED",X"E1",X"CD",X"0D",X"E2",X"CD",X"28",X"E2",X"CD",X"F7",
		X"DE",X"CD",X"08",X"D7",X"3A",X"43",X"63",X"FE",X"01",X"CC",X"2F",X"D1",X"3A",X"11",X"63",X"FE",
		X"01",X"28",X"2F",X"3A",X"23",X"63",X"FE",X"01",X"20",X"32",X"3A",X"34",X"63",X"FE",X"01",X"28",
		X"2B",X"3A",X"24",X"63",X"3D",X"32",X"24",X"63",X"FE",X"00",X"20",X"11",X"3E",X"01",X"32",X"F5",
		X"62",X"3E",X"01",X"32",X"51",X"63",X"AF",X"32",X"23",X"63",X"C3",X"5C",X"F1",X"CD",X"55",X"DA",
		X"18",X"0A",X"3E",X"01",X"32",X"23",X"63",X"3E",X"20",X"32",X"24",X"63",X"3A",X"B6",X"62",X"FE",
		X"01",X"20",X"05",X"3E",X"80",X"32",X"27",X"60",X"3A",X"BA",X"62",X"FE",X"01",X"20",X"05",X"3E",
		X"80",X"32",X"67",X"60",X"3A",X"56",X"61",X"FE",X"00",X"28",X"04",X"AF",X"32",X"57",X"60",X"3A",
		X"57",X"61",X"FE",X"00",X"28",X"04",X"AF",X"32",X"97",X"60",X"00",X"C3",X"F9",X"EC",X"7E",X"21",
		X"9E",X"23",X"23",X"01",X"09",X"00",X"ED",X"B1",X"C9",X"3A",X"5E",X"61",X"FE",X"00",X"20",X"06",
		X"3A",X"59",X"61",X"FE",X"00",X"C8",X"DD",X"21",X"9C",X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",
		X"60",X"32",X"98",X"60",X"DD",X"35",X"03",X"CD",X"EF",X"EA",X"DD",X"21",X"9C",X"65",X"DD",X"34",
		X"03",X"7E",X"E5",X"21",X"24",X"5B",X"01",X"07",X"00",X"ED",X"B9",X"E1",X"C2",X"D9",X"F1",X"3E",
		X"01",X"32",X"5E",X"61",X"AF",X"32",X"59",X"61",X"C9",X"AF",X"32",X"5E",X"61",X"3C",X"32",X"59",
		X"61",X"DD",X"21",X"9C",X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",
		X"EF",X"EA",X"7E",X"E5",X"21",X"E3",X"21",X"01",X"17",X"00",X"ED",X"B9",X"E1",X"C8",X"AF",X"32",
		X"5E",X"61",X"32",X"59",X"61",X"FD",X"2A",X"5C",X"61",X"3A",X"0D",X"60",X"FD",X"77",X"02",X"CD",
		X"B2",X"F2",X"7E",X"EB",X"21",X"E3",X"21",X"01",X"17",X"00",X"ED",X"B9",X"EB",X"28",X"06",X"11",
		X"20",X"00",X"19",X"18",X"21",X"11",X"20",X"00",X"E5",X"19",X"7E",X"E1",X"FE",X"EC",X"28",X"16",
		X"FE",X"EE",X"28",X"12",X"EB",X"21",X"E3",X"21",X"01",X"17",X"00",X"ED",X"B9",X"EB",X"28",X"06",
		X"11",X"20",X"00",X"AF",X"ED",X"52",X"F3",X"FD",X"75",X"00",X"7D",X"FE",X"C0",X"20",X"02",X"3E",
		X"68",X"FD",X"74",X"01",X"3A",X"0D",X"60",X"FD",X"77",X"02",X"FB",X"CD",X"05",X"EC",X"28",X"02",
		X"18",X"42",X"DD",X"E5",X"CD",X"C2",X"F2",X"3A",X"9D",X"65",X"FE",X"24",X"20",X"0B",X"3E",X"20",
		X"32",X"9D",X"65",X"CD",X"C2",X"F2",X"CD",X"C2",X"F2",X"21",X"81",X"D9",X"CD",X"84",X"EC",X"CD",
		X"D9",X"D4",X"20",X"0A",X"21",X"78",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"DD",X"E1",
		X"F3",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FB",X"3E",X"40",X"32",X"E8",
		X"61",X"CD",X"2F",X"D1",X"AF",X"DD",X"21",X"9C",X"65",X"DD",X"77",X"02",X"3E",X"FF",X"DD",X"77",
		X"03",X"C9",X"CD",X"87",X"EB",X"7C",X"80",X"67",X"AF",X"7D",X"D6",X"22",X"6F",X"7C",X"DE",X"00",
		X"67",X"C9",X"2A",X"E7",X"61",X"2E",X"00",X"CD",X"90",X"5C",X"C9",X"3A",X"D2",X"62",X"FE",X"01",
		X"C8",X"3A",X"3A",X"63",X"FE",X"01",X"C8",X"3A",X"58",X"61",X"FE",X"00",X"C2",X"A7",X"F4",X"3A",
		X"CF",X"61",X"FE",X"01",X"C8",X"3A",X"C7",X"61",X"FE",X"01",X"C8",X"3A",X"59",X"61",X"FE",X"01",
		X"C8",X"3A",X"11",X"63",X"FE",X"01",X"C8",X"3A",X"5E",X"61",X"FE",X"01",X"C8",X"3A",X"34",X"63",
		X"FE",X"01",X"C8",X"FD",X"21",X"9C",X"60",X"06",X"12",X"2A",X"09",X"60",X"3E",X"24",X"32",X"7B",
		X"62",X"FD",X"7E",X"02",X"C5",X"47",X"3A",X"0D",X"60",X"B8",X"C1",X"C2",X"35",X"F3",X"FD",X"56",
		X"01",X"FD",X"5E",X"00",X"13",X"13",X"CD",X"7B",X"F4",X"AF",X"E5",X"ED",X"52",X"E1",X"28",X"13",
		X"CD",X"0B",X"D0",X"28",X"0E",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"3E",X"20",X"32",X"7B",X"62",
		X"10",X"CF",X"C9",X"CD",X"E3",X"F4",X"78",X"FE",X"00",X"C8",X"3A",X"CF",X"61",X"FE",X"00",X"28",
		X"1F",X"FD",X"E5",X"E5",X"01",X"CF",X"61",X"FD",X"21",X"CC",X"61",X"3E",X"38",X"FD",X"77",X"04",
		X"3E",X"28",X"FD",X"77",X"05",X"3E",X"E4",X"32",X"D2",X"61",X"CD",X"55",X"FC",X"E1",X"FD",X"E1",
		X"DD",X"21",X"80",X"65",X"3A",X"41",X"63",X"FE",X"01",X"20",X"1A",X"3E",X"31",X"DD",X"77",X"1C",
		X"3E",X"24",X"DD",X"77",X"1D",X"DD",X"7E",X"03",X"DD",X"77",X"1F",X"DD",X"7E",X"02",X"D6",X"08",
		X"DD",X"77",X"1E",X"18",X"19",X"3E",X"3F",X"DD",X"77",X"1C",X"3A",X"7B",X"62",X"DD",X"77",X"1D",
		X"DD",X"7E",X"03",X"DD",X"77",X"1F",X"DD",X"7E",X"02",X"D6",X"08",X"DD",X"77",X"1E",X"CD",X"D9",
		X"D4",X"20",X"0A",X"21",X"A8",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"3E",X"01",X"32",
		X"58",X"61",X"FD",X"22",X"5C",X"61",X"FD",X"66",X"01",X"FD",X"6E",X"00",X"22",X"F6",X"61",X"AF",
		X"32",X"7E",X"62",X"F3",X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FB",X"3A",X"7B",
		X"62",X"FE",X"24",X"3E",X"00",X"20",X"02",X"3E",X"01",X"32",X"7C",X"62",X"C9",X"3A",X"7E",X"62",
		X"FE",X"07",X"D0",X"2A",X"F6",X"61",X"7C",X"FE",X"00",X"C8",X"7D",X"E6",X"1F",X"FE",X"00",X"C8",
		X"CD",X"65",X"F4",X"CD",X"3B",X"F4",X"23",X"CD",X"65",X"F4",X"CD",X"3B",X"F4",X"11",X"20",X"00",
		X"19",X"CD",X"65",X"F4",X"CD",X"3B",X"F4",X"2B",X"CD",X"65",X"F4",X"CD",X"3B",X"F4",X"3A",X"7E",
		X"62",X"3C",X"32",X"7E",X"62",X"3A",X"0D",X"60",X"FE",X"05",X"CC",X"4D",X"CE",X"C9",X"DD",X"7E",
		X"00",X"FE",X"01",X"C8",X"7E",X"FE",X"F0",X"D8",X"AF",X"12",X"C9",X"06",X"1F",X"7E",X"FE",X"49",
		X"28",X"16",X"FE",X"4A",X"28",X"12",X"FE",X"4B",X"28",X"0E",X"FE",X"51",X"28",X"13",X"FE",X"52",
		X"28",X"0F",X"FE",X"57",X"28",X"0B",X"06",X"3F",X"E5",X"7C",X"C6",X"08",X"67",X"78",X"77",X"E1",
		X"C9",X"06",X"32",X"18",X"F3",X"7C",X"57",X"7D",X"5F",X"CD",X"7B",X"F4",X"1A",X"77",X"1A",X"BE",
		X"20",X"FA",X"E5",X"7C",X"C6",X"08",X"67",X"AF",X"77",X"E1",X"C9",X"3A",X"0D",X"60",X"FE",X"01",
		X"20",X"05",X"7A",X"D6",X"50",X"57",X"C9",X"FE",X"02",X"20",X"05",X"7A",X"D6",X"4C",X"57",X"C9",
		X"FE",X"03",X"20",X"05",X"7A",X"D6",X"48",X"57",X"C9",X"FE",X"04",X"20",X"05",X"7A",X"D6",X"60",
		X"57",X"C9",X"7A",X"D6",X"5C",X"57",X"C9",X"3A",X"59",X"61",X"FE",X"01",X"C8",X"3A",X"9E",X"65",
		X"FE",X"E0",X"D0",X"FE",X"18",X"D8",X"CD",X"E3",X"F4",X"78",X"FE",X"00",X"C8",X"DD",X"21",X"9C",
		X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",X"EF",X"EA",X"FB",X"2B",
		X"7E",X"E5",X"CD",X"F2",X"F4",X"E1",X"C0",X"AF",X"32",X"58",X"61",X"32",X"7C",X"62",X"3C",X"32",
		X"59",X"61",X"C9",X"06",X"00",X"3A",X"60",X"61",X"FE",X"00",X"C8",X"AF",X"32",X"60",X"61",X"06",
		X"01",X"C9",X"21",X"84",X"23",X"01",X"13",X"00",X"F5",X"3A",X"41",X"63",X"FE",X"01",X"CB",X"1B",
		X"F1",X"CB",X"13",X"38",X"03",X"01",X"15",X"00",X"ED",X"B9",X"C9",X"FD",X"E5",X"CD",X"18",X"19",
		X"FD",X"7E",X"00",X"67",X"FD",X"7E",X"01",X"6F",X"AF",X"ED",X"52",X"28",X"17",X"FD",X"23",X"FD",
		X"23",X"FD",X"23",X"3A",X"00",X"B8",X"FD",X"7E",X"02",X"FE",X"FF",X"20",X"E3",X"AF",X"DD",X"77",
		X"11",X"FD",X"E1",X"C9",X"DD",X"E5",X"FD",X"22",X"4B",X"60",X"3A",X"98",X"60",X"47",X"3A",X"0D",
		X"60",X"B8",X"28",X"03",X"CD",X"3A",X"19",X"06",X"08",X"DD",X"7E",X"11",X"FE",X"01",X"CA",X"44",
		X"F6",X"DD",X"7E",X"07",X"FE",X"00",X"C2",X"44",X"F6",X"DD",X"23",X"10",X"F4",X"DD",X"E1",X"AF",
		X"DD",X"77",X"15",X"3A",X"47",X"60",X"FE",X"00",X"CA",X"95",X"F5",X"3A",X"82",X"65",X"47",X"FD",
		X"E1",X"FD",X"7E",X"02",X"FD",X"E5",X"B8",X"F5",X"D4",X"49",X"F6",X"F1",X"DC",X"52",X"F6",X"3A",
		X"83",X"65",X"47",X"FD",X"E1",X"FD",X"7E",X"03",X"FD",X"E5",X"B8",X"F5",X"DC",X"64",X"F6",X"F1",
		X"D4",X"5B",X"F6",X"18",X"58",X"3A",X"00",X"A0",X"E5",X"21",X"85",X"23",X"E6",X"03",X"85",X"6F",
		X"7C",X"CE",X"00",X"67",X"3A",X"00",X"B8",X"7E",X"C5",X"DD",X"E5",X"DD",X"2A",X"95",X"60",X"47",
		X"DD",X"7E",X"00",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"E6",X"0F",X"FE",X"01",X"20",
		X"04",X"3E",X"02",X"18",X"16",X"FE",X"02",X"20",X"04",X"3E",X"01",X"18",X"0E",X"FE",X"04",X"20",
		X"04",X"3E",X"08",X"18",X"06",X"FE",X"08",X"20",X"02",X"3E",X"04",X"B8",X"20",X"07",X"DD",X"E1",
		X"C1",X"E1",X"C3",X"95",X"F5",X"DD",X"E1",X"78",X"C1",X"E1",X"DD",X"77",X"15",X"AF",X"FD",X"2A",
		X"4B",X"60",X"FD",X"7E",X"02",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"47",X"DD",X"7E",
		X"15",X"A0",X"CB",X"0F",X"2A",X"91",X"60",X"32",X"44",X"60",X"FD",X"21",X"94",X"65",X"FD",X"22",
		X"93",X"60",X"2A",X"95",X"60",X"30",X"05",X"CD",X"E8",X"F6",X"18",X"20",X"CB",X"0F",X"30",X"05",
		X"CD",X"DE",X"F6",X"18",X"17",X"CB",X"0F",X"30",X"05",X"CD",X"C0",X"F6",X"18",X"07",X"CB",X"0F",
		X"30",X"0A",X"CD",X"A2",X"F6",X"3A",X"0B",X"60",X"FE",X"02",X"20",X"05",X"3E",X"01",X"DD",X"77",
		X"11",X"FD",X"E1",X"C9",X"DD",X"E1",X"FD",X"E1",X"C9",X"DD",X"7E",X"15",X"F6",X"04",X"DD",X"77",
		X"15",X"C9",X"DD",X"7E",X"15",X"F6",X"08",X"DD",X"77",X"15",X"C9",X"DD",X"7E",X"15",X"F6",X"01",
		X"DD",X"77",X"15",X"C9",X"DD",X"7E",X"15",X"F6",X"02",X"DD",X"77",X"15",X"C9",X"2A",X"38",X"60",
		X"22",X"91",X"60",X"FD",X"21",X"94",X"65",X"FD",X"22",X"93",X"60",X"21",X"27",X"60",X"22",X"95",
		X"60",X"3A",X"3C",X"60",X"FE",X"00",X"C4",X"A2",X"F6",X"3A",X"3D",X"60",X"FE",X"00",X"C4",X"C0",
		X"F6",X"3A",X"3E",X"60",X"FE",X"00",X"C4",X"E8",X"F6",X"3A",X"3F",X"60",X"FE",X"00",X"C4",X"DE",
		X"F6",X"C9",X"2A",X"91",X"60",X"DD",X"E5",X"DD",X"2A",X"93",X"60",X"CD",X"71",X"0D",X"DD",X"E1",
		X"3A",X"0B",X"60",X"FE",X"02",X"C0",X"E5",X"2A",X"95",X"60",X"AF",X"CB",X"FF",X"77",X"E1",X"C9",
		X"2A",X"91",X"60",X"DD",X"E5",X"DD",X"2A",X"93",X"60",X"CD",X"CC",X"0D",X"DD",X"E1",X"3A",X"0B",
		X"60",X"FE",X"02",X"C0",X"E5",X"2A",X"95",X"60",X"AF",X"CB",X"F7",X"77",X"E1",X"C9",X"AF",X"E5",
		X"2A",X"95",X"60",X"CB",X"EF",X"77",X"E1",X"C9",X"AF",X"E5",X"2A",X"95",X"60",X"CB",X"E7",X"77",
		X"E1",X"C9",X"3A",X"0D",X"60",X"47",X"3A",X"99",X"60",X"B8",X"C0",X"DD",X"21",X"3D",X"60",X"2A",
		X"38",X"60",X"01",X"E0",X"FF",X"3A",X"CF",X"61",X"FE",X"00",X"3E",X"40",X"20",X"06",X"DD",X"21",
		X"3C",X"60",X"3E",X"80",X"08",X"CD",X"F5",X"F7",X"2A",X"38",X"60",X"DD",X"21",X"3C",X"60",X"01",
		X"20",X"00",X"3A",X"CF",X"61",X"FE",X"00",X"3E",X"80",X"20",X"06",X"DD",X"21",X"3D",X"60",X"3E",
		X"40",X"08",X"CD",X"F5",X"F7",X"2A",X"38",X"60",X"01",X"FF",X"FF",X"3E",X"10",X"08",X"DD",X"21",
		X"3E",X"60",X"CD",X"F5",X"F7",X"2A",X"38",X"60",X"DD",X"21",X"3F",X"60",X"01",X"01",X"00",X"3E",
		X"20",X"08",X"CD",X"F5",X"F7",X"C9",X"2A",X"78",X"60",X"22",X"91",X"60",X"FD",X"21",X"98",X"65",
		X"FD",X"22",X"93",X"60",X"21",X"67",X"60",X"22",X"95",X"60",X"3A",X"7C",X"60",X"FE",X"00",X"C4",
		X"A2",X"F6",X"3A",X"7D",X"60",X"FE",X"00",X"C4",X"C0",X"F6",X"3A",X"7E",X"60",X"FE",X"00",X"C4",
		X"E8",X"F6",X"3A",X"7F",X"60",X"FE",X"00",X"C4",X"DE",X"F6",X"C9",X"3A",X"0D",X"60",X"47",X"3A",
		X"9A",X"60",X"B8",X"C0",X"DD",X"21",X"7D",X"60",X"2A",X"78",X"60",X"01",X"E0",X"FF",X"3A",X"CF",
		X"61",X"FE",X"00",X"3E",X"40",X"20",X"06",X"DD",X"21",X"7C",X"60",X"3E",X"80",X"08",X"CD",X"F5",
		X"F7",X"2A",X"78",X"60",X"01",X"20",X"00",X"DD",X"21",X"7C",X"60",X"3A",X"CF",X"61",X"FE",X"00",
		X"3A",X"B2",X"91",X"32",X"72",X"62",X"3E",X"80",X"20",X"06",X"DD",X"21",X"7D",X"60",X"3E",X"40",
		X"08",X"CD",X"F5",X"F7",X"2A",X"78",X"60",X"01",X"FF",X"FF",X"3E",X"10",X"08",X"DD",X"21",X"7E",
		X"60",X"CD",X"F5",X"F7",X"2A",X"78",X"60",X"DD",X"21",X"7F",X"60",X"01",X"01",X"00",X"3E",X"20",
		X"08",X"CD",X"F5",X"F7",X"C9",X"2B",X"2B",X"AF",X"DD",X"77",X"00",X"ED",X"4A",X"7E",X"C5",X"06",
		X"15",X"FD",X"21",X"89",X"23",X"FD",X"BE",X"00",X"28",X"06",X"FD",X"23",X"10",X"F7",X"C1",X"C9",
		X"C1",X"E5",X"ED",X"5B",X"09",X"60",X"1B",X"1B",X"AF",X"ED",X"52",X"E1",X"28",X"0A",X"E5",X"13",
		X"AF",X"ED",X"52",X"E1",X"28",X"02",X"18",X"CF",X"08",X"DD",X"77",X"00",X"C9",X"3A",X"29",X"60",
		X"FE",X"01",X"28",X"08",X"3A",X"25",X"60",X"FE",X"01",X"CA",X"E1",X"F9",X"AF",X"C9",X"3A",X"25",
		X"60",X"FE",X"01",X"C8",X"3A",X"29",X"60",X"FE",X"01",X"C8",X"DD",X"21",X"82",X"65",X"FD",X"21",
		X"8A",X"65",X"21",X"22",X"60",X"11",X"04",X"00",X"3A",X"2A",X"60",X"FE",X"01",X"C8",X"CD",X"62",
		X"F8",X"C9",X"FD",X"7E",X"01",X"D6",X"04",X"DD",X"BE",X"01",X"D0",X"FD",X"7E",X"01",X"C6",X"0E",
		X"DD",X"BE",X"01",X"D8",X"FD",X"7E",X"00",X"D6",X"0D",X"47",X"C6",X"04",X"4F",X"CD",X"96",X"F8",
		X"32",X"25",X"60",X"FE",X"01",X"C8",X"FD",X"7E",X"00",X"C6",X"0A",X"47",X"C6",X"04",X"4F",X"CD",
		X"96",X"F8",X"32",X"25",X"60",X"C9",X"DD",X"7E",X"00",X"B8",X"38",X"06",X"B9",X"30",X"03",X"3E",
		X"01",X"C9",X"AF",X"C9",X"11",X"80",X"56",X"21",X"A0",X"93",X"CD",X"67",X"CA",X"11",X"80",X"56",
		X"21",X"20",X"91",X"CD",X"67",X"CA",X"11",X"05",X"57",X"21",X"40",X"92",X"CD",X"67",X"CA",X"3E",
		X"02",X"21",X"40",X"90",X"77",X"11",X"89",X"56",X"21",X"9F",X"91",X"CD",X"67",X"CA",X"3A",X"04",
		X"60",X"32",X"9F",X"90",X"3A",X"05",X"60",X"32",X"BF",X"90",X"CD",X"DE",X"F8",X"C9",X"3E",X"02",
		X"21",X"40",X"98",X"CD",X"05",X"56",X"3E",X"08",X"21",X"5F",X"98",X"CD",X"05",X"56",X"3E",X"05",
		X"21",X"41",X"98",X"CD",X"05",X"56",X"C9",X"3A",X"4D",X"60",X"FE",X"12",X"38",X"25",X"3E",X"01",
		X"32",X"4E",X"60",X"2A",X"09",X"60",X"7E",X"FE",X"F8",X"E5",X"21",X"A7",X"23",X"01",X"0A",X"00",
		X"ED",X"B9",X"E1",X"20",X"10",X"3A",X"14",X"60",X"FE",X"01",X"28",X"11",X"3A",X"E5",X"62",X"FE",
		X"01",X"28",X"0A",X"AF",X"C9",X"3A",X"83",X"65",X"D6",X"02",X"32",X"83",X"65",X"AF",X"32",X"08",
		X"60",X"CD",X"E1",X"F9",X"3E",X"01",X"C9",X"3A",X"54",X"60",X"FE",X"01",X"28",X"0C",X"3A",X"00",
		X"60",X"FE",X"00",X"28",X"06",X"3E",X"01",X"32",X"53",X"60",X"C9",X"3E",X"00",X"32",X"53",X"60",
		X"C9",X"21",X"60",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"CD",X"E7",X"D4",X"20",X"0D",
		X"21",X"68",X"3B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"32",X"48",X"63",X"AF",X"32",X"03",
		X"A0",X"CD",X"C9",X"C2",X"3E",X"01",X"32",X"16",X"60",X"CD",X"A4",X"F8",X"3E",X"01",X"32",X"0D",
		X"60",X"32",X"03",X"A0",X"3E",X"20",X"21",X"80",X"65",X"77",X"23",X"3E",X"08",X"77",X"23",X"3E",
		X"29",X"77",X"23",X"3E",X"D8",X"77",X"32",X"29",X"60",X"3E",X"40",X"32",X"65",X"61",X"3E",X"C8",
		X"32",X"66",X"61",X"11",X"C7",X"61",X"21",X"FB",X"1B",X"01",X"18",X"00",X"ED",X"B0",X"3E",X"40",
		X"32",X"E8",X"61",X"3E",X"01",X"32",X"86",X"62",X"32",X"19",X"60",X"3E",X"B0",X"32",X"9A",X"65",
		X"CD",X"BF",X"DF",X"3E",X"38",X"32",X"4D",X"63",X"CD",X"56",X"D7",X"C9",X"3A",X"C5",X"61",X"FE",
		X"00",X"28",X"01",X"C9",X"3A",X"41",X"63",X"FE",X"01",X"C8",X"21",X"C3",X"92",X"22",X"C4",X"61",
		X"C9",X"CD",X"4B",X"D6",X"3E",X"01",X"32",X"F1",X"61",X"CD",X"69",X"D2",X"79",X"FE",X"01",X"CC",
		X"BD",X"CF",X"3A",X"7C",X"61",X"32",X"6C",X"62",X"2A",X"09",X"60",X"FD",X"21",X"08",X"60",X"DD",
		X"21",X"80",X"65",X"CD",X"2A",X"C1",X"3E",X"01",X"32",X"51",X"61",X"32",X"00",X"A0",X"21",X"79",
		X"27",X"22",X"54",X"61",X"21",X"5D",X"D9",X"AF",X"32",X"52",X"61",X"FB",X"CD",X"84",X"EC",X"3A",
		X"56",X"60",X"FE",X"00",X"28",X"0F",X"21",X"38",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",
		X"32",X"48",X"63",X"18",X"16",X"CD",X"E7",X"D4",X"20",X"11",X"F3",X"21",X"60",X"3F",X"22",X"40",
		X"61",X"AF",X"32",X"42",X"61",X"3E",X"01",X"32",X"48",X"63",X"FB",X"3A",X"52",X"61",X"FE",X"01",
		X"20",X"F9",X"21",X"00",X"E0",X"2B",X"7C",X"FE",X"00",X"20",X"FA",X"3A",X"56",X"60",X"FE",X"00",
		X"20",X"06",X"CD",X"6C",X"EC",X"CD",X"76",X"EC",X"CD",X"EA",X"FA",X"DD",X"21",X"9C",X"65",X"DD",
		X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"3E",X"FF",X"DD",X"77",X"03",X"AF",X"32",X"58",
		X"61",X"32",X"C7",X"61",X"32",X"11",X"63",X"CD",X"BF",X"DF",X"3A",X"7D",X"61",X"FE",X"01",X"28",
		X"14",X"3A",X"7C",X"61",X"C6",X"01",X"E6",X"01",X"32",X"7C",X"61",X"3A",X"7D",X"61",X"47",X"FE",
		X"02",X"78",X"CC",X"27",X"C4",X"3A",X"56",X"60",X"FE",X"00",X"20",X"1B",X"3A",X"7C",X"61",X"C6",
		X"01",X"E6",X"01",X"32",X"7C",X"61",X"3A",X"7D",X"61",X"47",X"FE",X"02",X"78",X"CC",X"27",X"C4",
		X"3A",X"56",X"60",X"FE",X"00",X"28",X"51",X"3D",X"32",X"56",X"60",X"CD",X"17",X"D0",X"AF",X"32",
		X"08",X"60",X"32",X"4E",X"60",X"32",X"4D",X"60",X"32",X"8F",X"60",X"32",X"77",X"60",X"32",X"37",
		X"60",X"32",X"4F",X"60",X"CD",X"14",X"C3",X"3E",X"01",X"C9",X"DD",X"21",X"44",X"61",X"3E",X"00",
		X"06",X"06",X"CD",X"85",X"E5",X"AF",X"32",X"52",X"61",X"32",X"51",X"61",X"32",X"25",X"60",X"32",
		X"28",X"60",X"32",X"4E",X"60",X"32",X"29",X"60",X"32",X"13",X"60",X"32",X"4D",X"60",X"32",X"59",
		X"61",X"32",X"5E",X"61",X"32",X"C7",X"61",X"C9",X"CD",X"6C",X"EC",X"AF",X"32",X"54",X"60",X"06",
		X"16",X"21",X"00",X"30",X"2B",X"FB",X"3E",X"01",X"32",X"53",X"60",X"32",X"F1",X"61",X"7C",X"FE",
		X"00",X"20",X"F1",X"10",X"EC",X"CD",X"74",X"C6",X"AF",X"32",X"10",X"62",X"32",X"7C",X"61",X"3A",
		X"00",X"60",X"FE",X"00",X"20",X"35",X"CD",X"98",X"FB",X"11",X"AC",X"56",X"21",X"5A",X"93",X"CD",
		X"67",X"CA",X"11",X"53",X"23",X"21",X"B5",X"93",X"CD",X"D9",X"55",X"3E",X"0E",X"21",X"9A",X"98",
		X"CD",X"05",X"56",X"3E",X"03",X"21",X"55",X"98",X"CD",X"05",X"56",X"3E",X"11",X"32",X"B5",X"9B",
		X"CD",X"FB",X"C8",X"3E",X"01",X"32",X"00",X"A0",X"CD",X"D5",X"C5",X"F3",X"CD",X"DB",X"CF",X"CD",
		X"E7",X"CF",X"CD",X"1A",X"C4",X"AF",X"32",X"53",X"60",X"32",X"F1",X"61",X"3A",X"00",X"60",X"FE",
		X"00",X"CC",X"18",X"12",X"FB",X"3E",X"01",X"C9",X"3E",X"00",X"32",X"03",X"A0",X"CD",X"B7",X"C3",
		X"3E",X"30",X"CD",X"A3",X"C3",X"06",X"01",X"21",X"80",X"65",X"3E",X"00",X"CD",X"A8",X"C3",X"CD",
		X"A4",X"F8",X"3E",X"01",X"32",X"03",X"A0",X"C9",X"3A",X"00",X"A0",X"21",X"70",X"59",X"E6",X"03",
		X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",X"2A",X"95",X"60",X"77",X"C9",X"3A",X"59",X"61",X"FE",
		X"01",X"C8",X"3A",X"5E",X"61",X"FE",X"01",X"C8",X"0A",X"D9",X"FE",X"00",X"C2",X"3C",X"FC",X"2A",
		X"09",X"60",X"3A",X"0D",X"60",X"FD",X"BE",X"02",X"C0",X"FD",X"56",X"01",X"FD",X"5E",X"00",X"D5",
		X"13",X"13",X"CD",X"7B",X"F4",X"E5",X"AF",X"ED",X"52",X"E1",X"28",X"07",X"CD",X"0B",X"D0",X"28",
		X"02",X"D1",X"C9",X"D1",X"CD",X"E3",X"F4",X"78",X"FE",X"00",X"C8",X"62",X"6B",X"22",X"F6",X"61",
		X"AF",X"32",X"7E",X"62",X"DD",X"21",X"80",X"65",X"FD",X"7E",X"04",X"DD",X"77",X"1C",X"FD",X"7E",
		X"05",X"DD",X"77",X"1D",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",X"7E",X"04",X"FE",X"37",
		X"20",X"05",X"3E",X"01",X"FD",X"77",X"14",X"3E",X"01",X"D9",X"02",X"C9",X"FD",X"7E",X"00",X"FE",
		X"00",X"C0",X"3A",X"82",X"65",X"FE",X"D0",X"D0",X"3A",X"3A",X"63",X"FE",X"01",X"C8",X"CD",X"E3",
		X"F4",X"78",X"FE",X"00",X"C8",X"DD",X"21",X"9C",X"65",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",
		X"EF",X"EA",X"3A",X"11",X"63",X"FE",X"01",X"CA",X"E7",X"FC",X"E5",X"3A",X"0D",X"60",X"FD",X"77",
		X"02",X"CD",X"5E",X"E5",X"67",X"AF",X"7D",X"D6",X"22",X"6F",X"7C",X"DE",X"00",X"67",X"FD",X"75",
		X"00",X"FD",X"74",X"01",X"3A",X"0D",X"60",X"FD",X"77",X"02",X"C5",X"CD",X"6C",X"D3",X"78",X"C1",
		X"FE",X"00",X"CA",X"A7",X"D3",X"E1",X"7E",X"FE",X"E0",X"E5",X"CA",X"A7",X"D3",X"E1",X"E5",X"AF",
		X"7D",X"D6",X"20",X"7C",X"DE",X"00",X"67",X"E1",X"7E",X"FE",X"E0",X"C8",X"D9",X"3A",X"C7",X"61",
		X"FE",X"01",X"20",X"05",X"3E",X"28",X"08",X"18",X"1A",X"3E",X"20",X"08",X"3A",X"CF",X"61",X"FE",
		X"01",X"28",X"10",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"AF",X"D9",X"02",X"3E",X"01",X"32",
		X"34",X"63",X"C9",X"AF",X"02",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"FD",X"7E",X"06",X"CD",X"7C",
		X"CE",X"3E",X"FF",X"32",X"9F",X"65",X"C9",X"2B",X"C5",X"7E",X"E5",X"CD",X"F2",X"F4",X"E1",X"C1",
		X"C0",X"C3",X"C3",X"FC",X"FD",X"21",X"56",X"61",X"FD",X"7E",X"00",X"FE",X"01",X"C8",X"3A",X"99",
		X"60",X"32",X"98",X"60",X"DD",X"E5",X"21",X"00",X"05",X"CD",X"90",X"5C",X"21",X"6F",X"D9",X"CD",
		X"84",X"EC",X"DD",X"E1",X"DD",X"21",X"4F",X"60",X"CD",X"A9",X"D4",X"AF",X"32",X"57",X"60",X"3E",
		X"21",X"32",X"94",X"65",X"2A",X"38",X"60",X"FD",X"21",X"37",X"60",X"DD",X"21",X"94",X"65",X"CD",
		X"2A",X"C1",X"C9",X"FD",X"21",X"57",X"61",X"FD",X"7E",X"00",X"FE",X"01",X"C8",X"3A",X"9A",X"60",
		X"32",X"98",X"60",X"DD",X"E5",X"21",X"00",X"05",X"CD",X"90",X"5C",X"21",X"6F",X"D9",X"CD",X"84",
		X"EC",X"DD",X"E1",X"DD",X"21",X"8F",X"60",X"CD",X"A9",X"D4",X"AF",X"32",X"97",X"60",X"3E",X"21",
		X"32",X"98",X"65",X"2A",X"78",X"60",X"FD",X"21",X"77",X"60",X"DD",X"21",X"98",X"65",X"CD",X"2A",
		X"C1",X"C9",X"DD",X"21",X"9C",X"60",X"3E",X"04",X"32",X"7A",X"62",X"06",X"13",X"DD",X"E5",X"C5",
		X"CD",X"C1",X"CA",X"C1",X"DD",X"E1",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"3E",X"01",X"32",X"7A",
		X"62",X"10",X"EA",X"3A",X"C7",X"61",X"FE",X"01",X"28",X"1C",X"3A",X"0D",X"60",X"47",X"FD",X"21",
		X"C4",X"61",X"FD",X"7E",X"02",X"B8",X"20",X"0E",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"3E",X"28",
		X"08",X"3E",X"EC",X"CD",X"7C",X"CE",X"3A",X"0D",X"60",X"47",X"FD",X"21",X"CC",X"61",X"FD",X"7E",
		X"02",X"B8",X"20",X"22",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"7E",X"CD",X"F3",X"CF",X"20",X"16",
		X"E5",X"D5",X"11",X"20",X"00",X"19",X"7E",X"CD",X"F3",X"CF",X"D1",X"E1",X"20",X"08",X"3E",X"20",
		X"08",X"3E",X"E4",X"CD",X"7C",X"CE",X"06",X"04",X"FD",X"21",X"D3",X"61",X"11",X"CC",X"61",X"C5",
		X"FD",X"E5",X"D5",X"CD",X"C2",X"DB",X"1A",X"6F",X"13",X"1A",X"67",X"1B",X"3A",X"0D",X"60",X"FD",
		X"E1",X"FD",X"BE",X"02",X"FD",X"E5",X"20",X"1C",X"7E",X"CD",X"F3",X"CF",X"20",X"16",X"E5",X"D5",
		X"11",X"20",X"00",X"19",X"7E",X"CD",X"F3",X"CF",X"D1",X"E1",X"20",X"08",X"3E",X"20",X"08",X"3E",
		X"E4",X"CD",X"7C",X"CE",X"D1",X"FD",X"E1",X"C1",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"BF",
		X"3A",X"FF",X"FF",X"3A",X"0D",X"60",X"47",X"FD",X"21",X"0E",X"63",X"FD",X"7E",X"02",X"B8",X"20",
		X"22",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"7E",X"CD",X"F3",X"CF",X"20",X"16",X"E5",X"D5",X"11",
		X"20",X"00",X"19",X"7E",X"CD",X"F3",X"CF",X"D1",X"E1",X"20",X"08",X"3E",X"24",X"08",X"3E",X"D4",
		X"CD",X"7C",X"CE",X"06",X"04",X"FD",X"21",X"15",X"63",X"11",X"0E",X"63",X"C5",X"FD",X"E5",X"D5",
		X"CD",X"B5",X"DB",X"1A",X"6F",X"13",X"1A",X"67",X"1B",X"3A",X"0D",X"60",X"FD",X"E1",X"FD",X"BE",
		X"02",X"FD",X"E5",X"20",X"1C",X"7E",X"CD",X"F3",X"CF",X"20",X"16",X"E5",X"D5",X"11",X"20",X"00",
		X"19",X"7E",X"CD",X"F3",X"CF",X"D1",X"E1",X"20",X"08",X"3E",X"24",X"08",X"3E",X"D4",X"CD",X"7C",
		X"CE",X"D1",X"FD",X"E1",X"C1",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"BF",X"C9",X"3A",X"34",
		X"63",X"FE",X"00",X"C8",X"DD",X"21",X"9C",X"65",X"FD",X"21",X"5A",X"61",X"3A",X"0D",X"60",X"32",
		X"98",X"60",X"CD",X"EF",X"EA",X"7E",X"E5",X"21",X"E3",X"21",X"01",X"17",X"00",X"ED",X"B9",X"E1",
		X"C8",X"3A",X"0D",X"60",X"CD",X"B2",X"F2",X"22",X"26",X"63",X"3E",X"24",X"08",X"3E",X"D4",X"CD",
		X"7C",X"CE",X"3E",X"00",X"32",X"34",X"63",X"3E",X"FF",X"32",X"9F",X"65",X"C9",X"05",X"08",X"4E",
		X"20",X"48",X"03",X"41",X"30",X"08",X"01",X"DC",X"08",X"0C",X"30",X"45",X"10",X"46",X"31",X"4D",
		X"00",X"44",X"02",X"4F",X"20",X"41",X"A3",X"CA",X"00",X"14",X"08",X"47",X"00",X"03",X"01",X"D9",
		X"10",X"43",X"14",X"7F",X"80",X"4D",X"05",X"CD",X"91",X"4C",X"A4",X"E6",X"00",X"41",X"90",X"6F",
		X"68",X"04",X"3E",X"55",X"18",X"4E",X"79",X"84",X"00",X"C1",X"30",X"5B",X"61",X"CD",X"7C",X"4B",
		X"21",X"47",X"21",X"8F",X"09",X"DC",X"B7",X"4F",X"B0",X"46",X"23",X"CE",X"20",X"4C",X"B4",X"0E",
		X"02",X"0F",X"08",X"47",X"08",X"9D",X"AA",X"4B",X"00",X"E3",X"AA",X"CF",X"00",X"0E",X"C0",X"4F",
		X"19",X"46",X"24",X"CF",X"04",X"1D",X"A0",X"CB",X"09",X"46",X"21",X"07",X"00",X"42",X"E4",X"E4",
		X"20",X"13",X"0E",X"46",X"00",X"C8",X"12",X"DC",X"01",X"55",X"9B",X"63",X"30",X"88",X"29",X"4F",
		X"10",X"45",X"04",X"4C",X"03",X"67",X"02",X"4E",X"88",X"4F",X"38",X"56",X"80",X"49",X"05",X"47",
		X"08",X"48",X"0B",X"EC",X"29",X"48",X"11",X"6E",X"20",X"50",X"A3",X"6A",X"21",X"65",X"20",X"0C",
		X"80",X"48",X"0A",X"6B",X"64",X"48",X"6B",X"4E",X"20",X"4B",X"22",X"49",X"09",X"A4",X"2F",X"17",
		X"A6",X"CE",X"09",X"4F",X"0B",X"E9",X"01",X"C7",X"3D",X"5D",X"26",X"DD",X"68",X"EF",X"A5",X"45",
		X"25",X"07",X"3F",X"85",X"14",X"44",X"B0",X"CC",X"80",X"59",X"31",X"51",X"77",X"B4",X"FB",X"F7",
		X"21",X"09",X"69",X"2D",X"20",X"18",X"1A",X"4A",X"10",X"41",X"72",X"49",X"04",X"41",X"20",X"12",
		X"00",X"4F",X"00",X"17",X"00",X"EE",X"74",X"2A",X"01",X"53",X"00",X"5F",X"F7",X"3B",X"F7",X"BB",
		X"00",X"01",X"2D",X"6E",X"A1",X"0C",X"22",X"43",X"11",X"6D",X"16",X"06",X"20",X"CE",X"B8",X"D5",
		X"00",X"43",X"02",X"82",X"20",X"4B",X"12",X"5E",X"00",X"0D",X"15",X"84",X"FF",X"8C",X"EF",X"3E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
