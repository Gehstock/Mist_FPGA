library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity g1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of g1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",
		X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",
		X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",
		X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",X"1F",X"24",
		X"1F",X"24",X"3F",X"24",X"5F",X"24",X"7F",X"24",X"9F",X"24",X"BF",X"24",X"DF",X"24",X"FF",X"24",
		X"1F",X"25",X"3F",X"25",X"5F",X"25",X"7F",X"25",X"9F",X"25",X"BF",X"25",X"DF",X"25",X"FF",X"25",
		X"1F",X"26",X"3F",X"26",X"5F",X"26",X"7F",X"26",X"9F",X"26",X"BF",X"26",X"DF",X"26",X"FF",X"26",
		X"1F",X"27",X"3F",X"27",X"5F",X"27",X"7F",X"27",X"9F",X"27",X"BF",X"27",X"DF",X"27",X"FF",X"27",
		X"1F",X"28",X"3F",X"28",X"5F",X"28",X"7F",X"28",X"9F",X"28",X"BF",X"28",X"DF",X"28",X"FF",X"28",
		X"1F",X"29",X"3F",X"29",X"5F",X"29",X"7F",X"29",X"9F",X"29",X"BF",X"29",X"DF",X"29",X"FF",X"29",
		X"1F",X"2A",X"3F",X"2A",X"5F",X"2A",X"7F",X"2A",X"9F",X"2A",X"BF",X"2A",X"DF",X"2A",X"FF",X"2A",
		X"1F",X"2B",X"3F",X"2B",X"5F",X"2B",X"7F",X"2B",X"9F",X"2B",X"BF",X"2B",X"DF",X"2B",X"FF",X"2B",
		X"1F",X"2C",X"3F",X"2C",X"5F",X"2C",X"7F",X"2C",X"9F",X"2C",X"BF",X"2C",X"DF",X"2C",X"FF",X"2C",
		X"1F",X"2D",X"3F",X"2D",X"5F",X"2D",X"7F",X"2D",X"9F",X"2D",X"BF",X"2D",X"DF",X"2D",X"FF",X"2D",
		X"1F",X"2E",X"3F",X"2E",X"5F",X"2E",X"7F",X"2E",X"9F",X"2E",X"BF",X"2E",X"DF",X"2E",X"FF",X"2E",
		X"1F",X"2F",X"3F",X"2F",X"5F",X"2F",X"7F",X"2F",X"9F",X"2F",X"BF",X"2F",X"DF",X"2F",X"FF",X"2F",
		X"1F",X"30",X"3F",X"30",X"5F",X"30",X"7F",X"30",X"9F",X"30",X"BF",X"30",X"DF",X"30",X"FF",X"30",
		X"1F",X"31",X"3F",X"31",X"5F",X"31",X"7F",X"31",X"9F",X"31",X"BF",X"31",X"DF",X"31",X"FF",X"31",
		X"1F",X"32",X"3F",X"32",X"5F",X"32",X"7F",X"32",X"9F",X"32",X"BF",X"32",X"DF",X"32",X"FF",X"32",
		X"1F",X"33",X"3F",X"33",X"5F",X"33",X"7F",X"33",X"9F",X"33",X"BF",X"33",X"DF",X"33",X"FF",X"33",
		X"1F",X"34",X"3F",X"34",X"5F",X"34",X"7F",X"34",X"9F",X"34",X"BF",X"34",X"DF",X"34",X"FF",X"34",
		X"1F",X"35",X"3F",X"35",X"5F",X"35",X"7F",X"35",X"9F",X"35",X"BF",X"35",X"DF",X"35",X"FF",X"35",
		X"1F",X"36",X"3F",X"36",X"5F",X"36",X"7F",X"36",X"9F",X"36",X"BF",X"36",X"DF",X"36",X"FF",X"36",
		X"1F",X"37",X"3F",X"37",X"5F",X"37",X"7F",X"37",X"9F",X"37",X"BF",X"37",X"DF",X"37",X"FF",X"37",
		X"1F",X"38",X"3F",X"38",X"5F",X"38",X"7F",X"38",X"9F",X"38",X"BF",X"38",X"DF",X"38",X"FF",X"38",
		X"1F",X"39",X"3F",X"39",X"5F",X"39",X"7F",X"39",X"9F",X"39",X"BF",X"39",X"DF",X"39",X"FF",X"39",
		X"1F",X"3A",X"3F",X"3A",X"5F",X"3A",X"7F",X"3A",X"9F",X"3A",X"BF",X"3A",X"DF",X"3A",X"FF",X"3A",
		X"1F",X"3B",X"3F",X"3B",X"5F",X"3B",X"7F",X"3B",X"9F",X"3B",X"BF",X"3B",X"DF",X"3B",X"FF",X"3B",
		X"1F",X"3C",X"3F",X"3C",X"5F",X"3C",X"7F",X"3C",X"9F",X"3C",X"BF",X"3C",X"DF",X"3C",X"FF",X"3C",
		X"1F",X"3D",X"3F",X"3D",X"5F",X"3D",X"7F",X"3D",X"9F",X"3D",X"BF",X"3D",X"DF",X"3D",X"FF",X"3D",
		X"1F",X"3E",X"3F",X"3E",X"5F",X"3E",X"7F",X"3E",X"9F",X"3E",X"BF",X"3E",X"DF",X"3E",X"FF",X"3E",
		X"1F",X"3F",X"3F",X"3F",X"5F",X"3F",X"7F",X"3F",X"9F",X"3F",X"9F",X"3F",X"9F",X"3F",X"9F",X"3F",
		X"9F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"04",
		X"00",X"04",X"00",X"0A",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"1F",X"0A",X"1F",
		X"0A",X"0A",X"00",X"04",X"1E",X"05",X"0E",X"14",X"0F",X"04",X"00",X"03",X"13",X"08",X"04",X"02",
		X"19",X"18",X"00",X"02",X"05",X"05",X"02",X"15",X"09",X"16",X"00",X"04",X"04",X"04",X"00",X"00",
		X"00",X"00",X"00",X"04",X"02",X"01",X"01",X"01",X"02",X"04",X"00",X"04",X"08",X"10",X"10",X"10",
		X"08",X"04",X"00",X"04",X"15",X"0E",X"04",X"0E",X"15",X"04",X"00",X"00",X"04",X"04",X"1F",X"04",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"11",X"11",X"11",X"11",X"11",X"0E",X"00",X"04",X"06",X"04",X"04",X"04",
		X"04",X"0E",X"00",X"0E",X"11",X"10",X"0C",X"02",X"01",X"1F",X"00",X"1F",X"10",X"08",X"0C",X"10",
		X"11",X"0E",X"00",X"08",X"0C",X"0A",X"09",X"1F",X"08",X"08",X"00",X"1F",X"01",X"0F",X"10",X"10",
		X"11",X"0E",X"00",X"1C",X"02",X"01",X"0F",X"11",X"11",X"0E",X"00",X"1F",X"10",X"08",X"04",X"02",
		X"02",X"02",X"00",X"0E",X"11",X"11",X"0E",X"11",X"11",X"0E",X"00",X"0E",X"11",X"11",X"1E",X"10",
		X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",
		X"04",X"02",X"00",X"08",X"04",X"02",X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"1F",X"00",X"1F",
		X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"08",X"04",X"02",X"00",X"0E",X"11",X"08",X"04",X"04",
		X"00",X"04",X"00",X"0E",X"11",X"15",X"1D",X"0D",X"01",X"1E",X"00",X"04",X"0A",X"11",X"11",X"1F",
		X"11",X"11",X"00",X"0F",X"11",X"11",X"0F",X"11",X"11",X"0F",X"00",X"0E",X"11",X"01",X"01",X"01",
		X"11",X"0E",X"00",X"0F",X"11",X"11",X"11",X"11",X"11",X"0F",X"00",X"1F",X"01",X"01",X"0F",X"01",
		X"01",X"1F",X"00",X"1F",X"01",X"01",X"0F",X"01",X"01",X"01",X"00",X"1E",X"01",X"01",X"01",X"19",
		X"11",X"1E",X"00",X"11",X"11",X"11",X"1F",X"11",X"11",X"11",X"00",X"0E",X"04",X"04",X"04",X"04",
		X"04",X"0E",X"00",X"10",X"10",X"10",X"10",X"10",X"11",X"0E",X"00",X"11",X"09",X"05",X"03",X"05",
		X"09",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"1F",X"00",X"11",X"1B",X"15",X"15",X"11",
		X"11",X"11",X"00",X"11",X"11",X"13",X"15",X"19",X"11",X"11",X"00",X"0E",X"11",X"11",X"11",X"11",
		X"11",X"0E",X"00",X"0F",X"11",X"11",X"0F",X"01",X"01",X"01",X"00",X"0E",X"11",X"11",X"11",X"15",
		X"09",X"16",X"00",X"0F",X"11",X"11",X"0F",X"05",X"09",X"11",X"00",X"0E",X"11",X"01",X"0E",X"10",
		X"11",X"0E",X"00",X"1F",X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"11",X"11",X"11",X"11",X"11",
		X"11",X"0E",X"00",X"11",X"11",X"11",X"11",X"11",X"0A",X"04",X"00",X"11",X"11",X"11",X"15",X"15",
		X"1B",X"11",X"00",X"11",X"11",X"0A",X"04",X"0A",X"11",X"11",X"00",X"11",X"11",X"0A",X"04",X"04",
		X"04",X"04",X"00",X"1F",X"10",X"08",X"04",X"02",X"01",X"1F",X"00",X"1F",X"03",X"03",X"03",X"03",
		X"03",X"1F",X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"00",X"00",X"1F",X"18",X"18",X"18",X"18",
		X"18",X"1F",X"00",X"00",X"00",X"04",X"0A",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"26",X"9E",X"26",X"D3",X"27",X"C6",X"27",X"5A",X"28",X"AD",X"27",X"DD",X"28",X"C1",X"28",
		X"85",X"2B",X"9B",X"29",X"42",X"2A",X"B4",X"2A",X"D8",X"2A",X"08",X"2B",X"D0",X"2A",X"0C",X"2B",
		X"43",X"2B",X"95",X"2B",X"D9",X"2B",X"06",X"2C",X"54",X"2C",X"8A",X"2C",X"DD",X"2C",X"16",X"2D",
		X"44",X"2D",X"87",X"2D",X"C9",X"2D",X"18",X"2E",X"57",X"2E",X"99",X"2E",X"D8",X"2E",X"16",X"2F",
		X"46",X"2F",X"8A",X"2F",X"D5",X"2F",X"11",X"30",X"5C",X"30",X"87",X"30",X"C4",X"30",X"05",X"31",
		X"4B",X"31",X"8E",X"31",X"D3",X"31",X"17",X"32",X"9B",X"32",X"CD",X"32",X"02",X"33",X"43",X"33",
		X"87",X"33",X"D0",X"33",X"0B",X"34",X"55",X"34",X"99",X"34",X"D0",X"34",X"17",X"35",X"4E",X"35",
		X"85",X"35",X"C8",X"35",X"11",X"36",X"56",X"36",X"98",X"36",X"CE",X"36",X"04",X"37",X"47",X"37",
		X"8D",X"37",X"D6",X"37",X"1D",X"38",X"59",X"38",X"94",X"38",X"D0",X"38",X"05",X"39",X"4F",X"39",
		X"96",X"39",X"CC",X"39",X"09",X"3A",X"5C",X"3A",X"98",X"3A",X"D4",X"3A",X"10",X"3B",X"4C",X"3B",
		X"84",X"3B",X"C6",X"3B",X"08",X"3C",X"4A",X"3C",X"96",X"3C",X"DC",X"3C",X"19",X"3D",X"4A",X"3D",
		X"90",X"3D",X"C6",X"3D",X"0C",X"3E",X"54",X"3E",X"9A",X"3E",X"CF",X"3E",X"09",X"3E",X"44",X"3F",
		X"8C",X"3F",X"D0",X"3F",X"CD",X"CE",X"0C",X"CD",X"CB",X"0F",X"CD",X"5A",X"0D",X"C9",X"21",X"97",
		X"21",X"DF",X"C2",X"F0",X"0C",X"36",X"02",X"06",X"02",X"21",X"99",X"21",X"11",X"0A",X"20",X"7E",
		X"80",X"80",X"77",X"1A",X"D6",X"1A",X"BE",X"D2",X"EC",X"0C",X"36",X"00",X"7E",X"CD",X"27",X"0D",
		X"11",X"0A",X"20",X"3A",X"D7",X"20",X"B7",X"CA",X"05",X"0D",X"1A",X"06",X"06",X"90",X"90",X"D6",
		X"1A",X"CD",X"27",X"0D",X"C9",X"1A",X"06",X"02",X"D6",X"1A",X"F3",X"21",X"00",X"00",X"39",X"22",
		X"95",X"21",X"26",X"0C",X"E6",X"FE",X"6F",X"F9",X"E1",X"7E",X"E6",X"FE",X"77",X"05",X"C2",X"18",
		X"0D",X"2A",X"95",X"21",X"F9",X"FB",X"C9",X"21",X"00",X"00",X"F3",X"39",X"22",X"95",X"21",X"26",
		X"0C",X"E6",X"FE",X"6F",X"F9",X"E1",X"7E",X"F6",X"01",X"77",X"05",X"C2",X"35",X"0D",X"2A",X"95",
		X"21",X"F9",X"FB",X"C9",X"21",X"11",X"2D",X"7E",X"F6",X"01",X"77",X"21",X"CD",X"2D",X"7E",X"F6",
		X"01",X"77",X"21",X"92",X"2C",X"7E",X"F6",X"01",X"77",X"C9",X"21",X"9B",X"21",X"DF",X"C0",X"3A",
		X"12",X"20",X"E6",X"0F",X"C6",X"0F",X"77",X"3A",X"99",X"21",X"E6",X"FE",X"26",X"0C",X"6F",X"5E",
		X"23",X"56",X"1A",X"E6",X"FE",X"12",X"C9",X"2A",X"80",X"21",X"7D",X"B4",X"C8",X"7E",X"23",X"22",
		X"80",X"21",X"FE",X"FF",X"C2",X"92",X"0D",X"21",X"00",X"00",X"22",X"80",X"21",X"AF",X"32",X"84",
		X"21",X"C9",X"FE",X"C0",X"C2",X"9D",X"0D",X"3E",X"FF",X"32",X"84",X"21",X"C9",X"07",X"0F",X"D2",
		X"CD",X"0D",X"2A",X"82",X"21",X"47",X"CD",X"C2",X"0D",X"78",X"E6",X"1F",X"47",X"7D",X"E6",X"1F",
		X"80",X"47",X"CD",X"C2",X"0D",X"78",X"E6",X"1F",X"47",X"7D",X"E6",X"E0",X"B0",X"6F",X"22",X"82",
		X"21",X"C9",X"E6",X"60",X"EB",X"26",X"00",X"6F",X"29",X"29",X"29",X"19",X"C9",X"D6",X"20",X"26",
		X"00",X"6F",X"29",X"29",X"29",X"11",X"02",X"0A",X"19",X"EB",X"2A",X"82",X"21",X"06",X"08",X"3A",
		X"84",X"21",X"B7",X"C2",X"F7",X"0D",X"CD",X"0A",X"0E",X"11",X"00",X"FF",X"19",X"3E",X"01",X"00",
		X"CD",X"A5",X"0D",X"22",X"82",X"21",X"C9",X"1A",X"2F",X"77",X"13",X"7D",X"C6",X"20",X"D2",X"02",
		X"0E",X"24",X"6F",X"05",X"C2",X"F7",X"0D",X"C3",X"E9",X"0D",X"1A",X"77",X"13",X"7D",X"C6",X"20",
		X"D2",X"14",X"0E",X"24",X"6F",X"05",X"C2",X"0A",X"0E",X"C9",X"CD",X"06",X"0F",X"CD",X"44",X"0E",
		X"3A",X"12",X"20",X"07",X"E6",X"0E",X"21",X"34",X"0E",X"85",X"D2",X"2E",X"0E",X"24",X"6F",X"5E",
		X"23",X"56",X"EB",X"E9",X"7E",X"0E",X"89",X"0E",X"96",X"0E",X"A1",X"0E",X"AE",X"0E",X"B9",X"0E",
		X"C6",X"0E",X"D7",X"0E",X"3A",X"12",X"20",X"E6",X"0F",X"C0",X"3A",X"12",X"20",X"E6",X"10",X"CA",
		X"65",X"0E",X"3A",X"2A",X"20",X"B7",X"C2",X"5B",X"0E",X"3E",X"0A",X"07",X"07",X"07",X"11",X"C3",
		X"25",X"CD",X"47",X"0F",X"C9",X"3A",X"50",X"23",X"B7",X"C0",X"3A",X"30",X"20",X"B7",X"C2",X"73",
		X"0E",X"3E",X"0A",X"07",X"07",X"07",X"2A",X"37",X"20",X"2B",X"CD",X"31",X"0F",X"C9",X"3A",X"29",
		X"20",X"0F",X"11",X"C4",X"25",X"CD",X"47",X"0F",X"C9",X"3A",X"29",X"20",X"07",X"07",X"07",X"11",
		X"C5",X"25",X"CD",X"47",X"0F",X"C9",X"3A",X"28",X"20",X"0F",X"11",X"C6",X"25",X"CD",X"47",X"0F",
		X"C9",X"3A",X"28",X"20",X"07",X"07",X"07",X"11",X"C7",X"25",X"CD",X"47",X"0F",X"C9",X"3A",X"39",
		X"20",X"0F",X"11",X"D9",X"25",X"CD",X"47",X"0F",X"C9",X"3A",X"39",X"20",X"07",X"07",X"07",X"11",
		X"DA",X"25",X"CD",X"47",X"0F",X"C9",X"3A",X"51",X"23",X"FE",X"01",X"D0",X"3A",X"2F",X"20",X"0F",
		X"2A",X"37",X"20",X"CD",X"31",X"0F",X"C9",X"3A",X"51",X"23",X"FE",X"02",X"D0",X"3A",X"2F",X"20",
		X"07",X"07",X"07",X"2A",X"37",X"20",X"23",X"CD",X"31",X"0F",X"C9",X"3A",X"50",X"23",X"B7",X"C8",
		X"3A",X"51",X"23",X"FE",X"05",X"D0",X"3E",X"0A",X"07",X"07",X"07",X"2A",X"37",X"20",X"23",X"23",
		X"23",X"23",X"CD",X"31",X"0F",X"C9",X"CD",X"EB",X"0E",X"3A",X"51",X"23",X"FE",X"04",X"D0",X"3A",
		X"2E",X"20",X"07",X"07",X"07",X"2A",X"37",X"20",X"23",X"23",X"23",X"CD",X"31",X"0F",X"2A",X"37",
		X"20",X"23",X"23",X"3A",X"51",X"23",X"FE",X"03",X"D0",X"3A",X"2E",X"20",X"0F",X"CD",X"31",X"0F",
		X"C9",X"E6",X"78",X"C6",X"80",X"EB",X"21",X"02",X"0A",X"85",X"D2",X"3E",X"0F",X"24",X"6F",X"23",
		X"EB",X"06",X"07",X"CD",X"0A",X"0E",X"C9",X"E6",X"78",X"47",X"0F",X"0F",X"80",X"21",X"5D",X"0F",
		X"85",X"D2",X"55",X"0F",X"24",X"6F",X"EB",X"06",X"0A",X"CD",X"0A",X"0E",X"C9",X"1C",X"36",X"63",
		X"63",X"63",X"63",X"63",X"63",X"36",X"1C",X"10",X"18",X"1C",X"10",X"10",X"10",X"10",X"10",X"10",
		X"7E",X"1C",X"36",X"63",X"60",X"30",X"18",X"0C",X"06",X"03",X"7F",X"7E",X"40",X"20",X"10",X"18",
		X"30",X"60",X"63",X"36",X"1C",X"30",X"28",X"24",X"22",X"21",X"7F",X"20",X"20",X"20",X"20",X"7F",
		X"01",X"01",X"01",X"1F",X"30",X"60",X"63",X"36",X"1C",X"30",X"18",X"0C",X"06",X"1F",X"37",X"63",
		X"63",X"36",X"1C",X"7F",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"1C",X"36",X"63",
		X"36",X"1C",X"36",X"63",X"63",X"36",X"1C",X"1C",X"36",X"63",X"63",X"76",X"7C",X"30",X"18",X"0C",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"E3",X"21",X"FE",X"03",
		X"D0",X"C3",X"44",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
