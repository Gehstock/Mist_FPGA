library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity skyskip_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of skyskip_sp_bits_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7E",X"9C",X"80",X"40",X"E0",X"C0",X"00",X"00",X"0C",X"1C",X"1C",X"94",
		X"74",X"F4",X"C4",X"8C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"07",X"03",X"03",X"E0",X"F0",
		X"F1",X"F3",X"E3",X"07",X"07",X"07",X"03",X"01",X"00",X"01",X"01",X"03",X"03",X"07",X"03",X"00",
		X"01",X"01",X"01",X"01",X"01",X"81",X"42",X"E3",X"E3",X"00",X"00",X"00",X"1B",X"30",X"E0",X"00",
		X"00",X"C0",X"E0",X"70",X"38",X"1D",X"0F",X"07",X"07",X"0D",X"1C",X"18",X"38",X"33",X"E7",X"6E",
		X"FD",X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"FC",X"23",X"DF",X"EF",X"FF",X"FF",X"DF",X"EF",X"F3",
		X"E3",X"E7",X"E7",X"E3",X"F3",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"8F",X"DF",X"7F",X"FE",
		X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"01",X"01",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"04",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"03",X"07",X"00",X"0F",
		X"1F",X"1F",X"BC",X"73",X"07",X"0F",X"1F",X"1B",X"1B",X"17",X"07",X"07",X"0F",X"17",X"1B",X"1B",
		X"13",X"1F",X"0E",X"0E",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7C",X"78",X"01",X"03",X"03",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"9C",X"FF",X"FF",X"FF",X"FF",X"FE",X"C8",X"F0",X"88",X"8B",X"8B",X"77",X"07",X"8F",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"FD",X"F0",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EF",X"F6",X"F9",X"F9",X"F6",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"90",X"00",
		X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",
		X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"01",X"0F",X"3F",X"38",
		X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"79",X"08",X"10",X"21",X"41",X"78",X"00",X"02",X"00",X"00",X"02",
		X"01",X"03",X"07",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"0F",X"0F",
		X"40",X"C0",X"E0",X"70",X"38",X"1C",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"E0",X"70",X"38",X"1C",X"0F",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"73",X"00",X"00",X"00",X"00",X"00",
		X"60",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"20",X"20",X"2C",X"2C",X"28",X"F8",X"FB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FB",X"3F",X"07",X"07",X"03",X"03",
		X"3C",X"FC",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"C0",X"C0",
		X"60",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"60",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FB",X"3F",X"87",X"87",X"83",X"83",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"87",X"0F",X"1F",X"3F",X"3F",X"3C",X"3C",X"3C",X"1C",X"1C",X"18",X"00",X"00",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"18",X"3F",X"3F",X"3F",X"3F",
		X"0F",X"0F",X"07",X"07",X"83",X"81",X"C4",X"E2",X"F9",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"3F",X"0F",X"07",X"07",X"83",X"81",X"C0",X"EC",X"FE",X"FE",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",
		X"3F",X"0F",X"07",X"07",X"83",X"81",X"C4",X"E2",X"F9",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EF",X"EF",X"2D",X"0D",X"05",X"01",X"01",X"01",X"05",X"1D",X"3B",X"F3",X"F1",X"F0",X"FA",
		X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"F6",X"F8",X"88",X"8C",X"8C",X"9F",X"FF",X"FF",X"9F",X"07",X"07",X"0F",X"0E",X"06",X"03",X"01",
		X"FF",X"FF",X"87",X"87",X"8F",X"9F",X"FF",X"FF",X"FF",X"97",X"07",X"0F",X"0E",X"06",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"7F",X"7F",X"BF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DE",X"CC",X"00",X"20",X"40",X"80",X"80",X"40",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"CF",X"07",X"23",X"43",X"83",X"81",X"41",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"23",X"23",X"23",X"23",X"23",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F6",X"F9",X"F9",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"63",X"03",X"03",X"07",X"0F",X"1F",X"12",X"12",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"0F",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"38",X"00",X"00",X"00",
		X"30",X"3F",X"1F",X"FF",X"FF",X"7F",X"1F",X"FF",X"FF",X"FF",X"67",X"0E",X"1E",X"1E",X"1C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",X"03",X"07",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"1F",X"3B",X"3B",X"37",X"07",X"0E",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"0A",X"0B",X"09",X"0E",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"1E",X"3C",X"3C",X"00",X"30",X"00",X"18",X"1C",X"0C",
		X"0D",X"0D",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"0D",X"0D",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"77",X"FC",X"E0",X"00",X"04",X"04",X"08",X"00",X"00",X"00",X"00",X"01",X"07",X"07",
		X"00",X"00",X"C0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"3F",X"FF",X"FF",
		X"0F",X"0F",X"2F",X"2F",X"3F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"3E",X"3E",X"BE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F0",X"E0",X"F0",X"00",X"00",X"00",X"E0",X"F8",X"FF",X"FF",X"FF",X"F8",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F0",X"F0",X"F0",
		X"F9",X"FF",X"BF",X"1F",X"0F",X"1F",X"3F",X"17",X"07",X"06",X"02",X"02",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"BF",X"1F",X"07",X"07",X"1F",X"1F",X"37",X"2D",X"09",X"00",X"00",X"00",X"00",X"00",
		X"79",X"7F",X"3F",X"3F",X"0F",X"1F",X"3F",X"7F",X"9F",X"38",X"20",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"02",X"03",X"70",X"78",X"3C",X"1E",X"0F",X"0F",
		X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"BF",X"FF",X"FF",X"FF",
		X"07",X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F4",X"F4",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"3F",X"FF",X"FF",X"7F",X"9F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7B",X"F8",X"F0",X"70",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"FB",X"F1",X"E0",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"C3",X"80",X"00",X"00",
		X"0F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"01",
		X"00",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"E0",X"E0",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"07",X"07",X"E7",X"E7",X"07",X"07",X"E7",X"E7",X"07",X"07",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"7C",X"7C",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"3C",X"1C",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"1B",X"1B",X"07",X"07",X"0F",X"1F",X"1F",X"3F",X"9F",X"DF",X"7F",X"3F",
		X"1F",X"3F",X"3F",X"01",X"3D",X"1A",X"07",X"07",X"47",X"47",X"42",X"62",X"62",X"36",X"18",X"08",
		X"00",X"FC",X"FF",X"67",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"9F",X"DF",X"FF",X"7F",X"1F",
		X"1F",X"3F",X"3F",X"01",X"3D",X"1A",X"07",X"07",X"07",X"07",X"06",X"42",X"C2",X"E2",X"7E",X"1C",
		X"F8",X"3C",X"38",X"3F",X"3E",X"70",X"61",X"60",X"43",X"47",X"47",X"47",X"43",X"40",X"41",X"79",
		X"70",X"7C",X"7E",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"5F",X"5F",X"CF",X"E9",X"EB",X"AB",X"06",
		X"FC",X"7C",X"3C",X"3F",X"7E",X"70",X"61",X"40",X"7B",X"7F",X"FF",X"D7",X"C3",X"C0",X"C1",X"79",
		X"70",X"7C",X"7E",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0B",X"0B",X"09",X"06",
		X"00",X"00",X"00",X"00",X"01",X"47",X"EF",X"6F",X"7F",X"DF",X"BF",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"3E",X"3C",X"3E",X"1C",X"1D",X"0F",X"03",X"03",X"03",X"07",X"05",X"01",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3E",X"3C",X"1E",X"1C",X"0F",X"03",X"03",X"03",X"07",X"05",X"01",
		X"01",X"00",X"00",X"00",X"7F",X"1F",X"1D",X"18",X"18",X"1A",X"1A",X"1D",X"1F",X"1F",X"0F",X"07",
		X"7E",X"7E",X"3E",X"0C",X"00",X"00",X"03",X"01",X"00",X"47",X"EF",X"EF",X"CF",X"EF",X"67",X"23",
		X"01",X"7F",X"1F",X"1D",X"18",X"18",X"1A",X"1A",X"1D",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",
		X"38",X"78",X"F8",X"F8",X"DC",X"00",X"00",X"03",X"01",X"00",X"07",X"0F",X"2F",X"6F",X"EF",X"CF",
		X"C3",X"E1",X"C0",X"00",X"7F",X"1F",X"1D",X"18",X"18",X"1A",X"1A",X"1D",X"1F",X"1F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0C",X"1D",X"06",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"37",X"7F",X"3F",X"7F",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"09",X"05",X"02",X"06",X"37",X"7F",X"3F",X"7F",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3F",X"3F",X"19",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"07",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"1B",X"19",X"1F",X"1C",X"18",X"0C",X"0F",X"07",X"03",X"01",X"00",
		X"03",X"07",X"07",X"07",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"04",X"05",X"01",X"02",X"02",X"06",X"07",X"03",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"1F",X"3F",X"03",X"01",X"01",X"08",X"1C",X"1E",X"0F",X"07",X"03",X"01",X"00",
		X"07",X"0F",X"10",X"00",X"00",X"01",X"01",X"00",X"04",X"0E",X"0E",X"07",X"03",X"01",X"00",X"00",
		X"01",X"03",X"01",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",
		X"41",X"C3",X"67",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"1B",X"1F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"3F",X"78",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"78",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"78",X"F0",
		X"19",X"3B",X"33",X"32",X"1B",X"1B",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F8",X"F8",X"FC",X"FC",X"7F",X"7E",X"7C",X"7C",X"3E",X"3E",X"1F",X"0F",X"03",X"00",
		X"00",X"80",X"80",X"E0",X"7C",X"1E",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"1F",X"0F",X"07",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"01",X"80",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F8",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"1C",X"1C",X"0E",X"0E",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"78",X"78",X"3C",X"3C",X"1C",X"1E",X"0E",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"19",X"09",X"19",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"19",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"39",X"39",X"19",X"00",X"00",X"00",X"00",
		X"FF",X"C6",X"C6",X"C7",X"C7",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"CE",X"CE",X"CE",
		X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",
		X"C6",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"FF",
		X"FF",X"CF",X"D6",X"C6",X"C6",X"C7",X"C7",X"C6",X"C6",X"CE",X"CE",X"C7",X"C7",X"C7",X"C6",X"C6",
		X"FF",X"C6",X"C7",X"DF",X"FF",X"C7",X"C7",X"CD",X"CC",X"DC",X"DE",X"DF",X"DF",X"DB",X"D9",X"D8",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"FF",
		X"D9",X"DB",X"D9",X"CF",X"CD",X"CF",X"CC",X"CC",X"CC",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"07",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"1F",X"3F",X"5F",X"6F",X"F7",X"F7",X"F7",X"F7",X"6F",X"5F",X"3F",X"1F",X"0F",X"03",
		X"03",X"0F",X"17",X"3B",X"7C",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7C",X"3B",X"17",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"20",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"1F",X"3E",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"3E",X"18",
		X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"07",X"07",X"03",
		X"C0",X"60",X"60",X"1C",X"1C",X"1E",X"02",X"C1",X"71",X"38",X"0C",X"F0",X"F8",X"FC",X"0C",X"0E",
		X"40",X"80",X"20",X"0C",X"1C",X"1E",X"00",X"C1",X"70",X"38",X"0C",X"F0",X"F8",X"FC",X"0C",X"0E",
		X"06",X"07",X"83",X"E3",X"E9",X"ED",X"DC",X"58",X"80",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"08",X"0C",X"06",X"C3",X"F1",X"3C",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"08",X"0C",X"06",X"C3",X"F1",X"3C",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"C0",X"E0",X"B0",X"98",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"0F",X"1F",X"3F",X"3F",X"3F",X"1F",X"17",X"17",X"1B",X"0B",X"0F",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",
		X"00",X"02",X"07",X"00",X"00",X"00",X"C0",X"E1",X"FF",X"BF",X"DF",X"DF",X"EF",X"F7",X"F7",X"FB",
		X"00",X"02",X"07",X"00",X"00",X"00",X"C0",X"E1",X"FF",X"BF",X"DF",X"DF",X"EF",X"F7",X"F7",X"FB",
		X"7B",X"01",X"01",X"00",X"00",X"00",X"00",X"FC",X"07",X"00",X"01",X"01",X"03",X"03",X"06",X"06",
		X"7B",X"01",X"01",X"00",X"00",X"00",X"00",X"FC",X"07",X"00",X"01",X"01",X"03",X"03",X"06",X"06",
		X"1F",X"1F",X"3F",X"3F",X"1F",X"1B",X"1B",X"1D",X"0D",X"0D",X"0F",X"0E",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",
		X"1F",X"2F",X"30",X"3D",X"3D",X"3D",X"3D",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"1F",X"2F",X"30",X"3D",X"3D",X"3D",X"3D",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"02",X"03",
		X"D8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"F8",X"78",X"70",X"70",X"F0",X"FC",X"FF",X"FF",
		X"07",X"06",X"06",X"00",X"01",X"00",X"20",X"32",X"18",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"06",X"06",X"00",X"01",X"00",X"00",X"02",X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"DE",X"E1",X"F7",X"F7",X"F7",X"77",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"08",X"00",X"02",X"00",X"00",
		X"03",X"07",X"07",X"03",X"1F",X"6F",X"DF",X"DF",X"BF",X"7F",X"FF",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"F0",X"AC",X"8E",X"B7",X"B7",X"DF",X"DF",X"DF",X"7F",X"3E",X"1C",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"20",X"00",X"0C",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"0C",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"00",X"00",X"00",X"C0",X"C0",X"80",X"81",X"47",X"47",X"47",X"27",X"23",X"13",X"33",
		X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"C7",X"47",X"87",X"47",X"23",X"13",X"33",
		X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"59",
		X"85",X"0C",X"0A",X"0A",X"FE",X"FC",X"B8",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"80",X"00",
		X"33",X"31",X"01",X"11",X"11",X"18",X"10",X"08",X"08",X"08",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"33",X"31",X"01",X"11",X"09",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"11",X"01",X"11",X"01",X"11",X"19",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"11",X"21",X"11",X"21",X"01",X"19",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"07",X"F3",X"3D",X"1C",X"00",X"04",X"0E",X"0A",X"7A",X"7E",X"7E",X"3C",X"80",X"00",X"00",X"00",
		X"11",X"01",X"11",X"01",X"11",X"10",X"10",X"18",X"18",X"10",X"30",X"30",X"03",X"00",X"00",X"00",
		X"01",X"09",X"11",X"21",X"11",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
