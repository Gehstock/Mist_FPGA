`define BUILD_DATE "190417"
`define BUILD_TIME "161535"
