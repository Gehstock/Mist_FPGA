library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MoonWar_program2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MoonWar_program2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"2A",X"AE",X"F8",X"7C",X"B5",X"C0",X"EB",X"22",X"AE",X"F8",X"C9",X"D5",X"CD",X"7C",X"2E",X"D1",
		X"07",X"07",X"EE",X"09",X"E6",X"0F",X"90",X"FA",X"1C",X"C0",X"18",X"FA",X"80",X"28",X"0C",X"47",
		X"7E",X"CB",X"7F",X"20",X"03",X"23",X"18",X"F8",X"23",X"10",X"F5",X"7E",X"47",X"E6",X"7F",X"12",
		X"13",X"CB",X"78",X"23",X"28",X"F5",X"C9",X"2A",X"AE",X"F8",X"7C",X"B5",X"C0",X"21",X"B1",X"F8",
		X"35",X"C0",X"CD",X"7C",X"2E",X"07",X"07",X"07",X"07",X"E6",X"0F",X"C6",X"01",X"77",X"21",X"2E",
		X"F9",X"CD",X"7C",X"2E",X"E6",X"07",X"F6",X"78",X"77",X"23",X"36",X"21",X"EB",X"21",X"72",X"C0",
		X"06",X"0B",X"CD",X"0B",X"C0",X"EB",X"36",X"47",X"23",X"36",X"FF",X"21",X"2E",X"F9",X"22",X"AE",
		X"F8",X"C9",X"01",X"02",X"0B",X"8C",X"00",X"21",X"01",X"0F",X"98",X"03",X"84",X"15",X"22",X"03",
		X"84",X"05",X"A3",X"05",X"02",X"08",X"87",X"0D",X"0E",X"0F",X"90",X"01",X"02",X"86",X"05",X"02",
		X"86",X"00",X"00",X"1A",X"92",X"0E",X"02",X"89",X"45",X"FF",X"7C",X"11",X"12",X"13",X"14",X"45",
		X"FF",X"7C",X"01",X"02",X"06",X"45",X"FF",X"7C",X"05",X"02",X"06",X"45",X"FF",X"7C",X"03",X"02",
		X"09",X"45",X"FF",X"7C",X"03",X"02",X"0A",X"45",X"FF",X"7C",X"08",X"07",X"17",X"21",X"15",X"45",
		X"FF",X"7C",X"07",X"04",X"21",X"00",X"24",X"24",X"24",X"45",X"FF",X"7C",X"1A",X"1B",X"1C",X"20",
		X"45",X"FF",X"7C",X"1A",X"1B",X"1D",X"20",X"45",X"FF",X"7C",X"1A",X"1B",X"1E",X"20",X"45",X"FF",
		X"7C",X"1A",X"1B",X"1F",X"20",X"45",X"FF",X"7C",X"00",X"00",X"21",X"03",X"02",X"19",X"45",X"FF",
		X"7C",X"15",X"22",X"0F",X"08",X"07",X"16",X"17",X"45",X"FF",X"7C",X"15",X"22",X"0F",X"06",X"16",
		X"04",X"45",X"FF",X"3A",X"E1",X"43",X"B7",X"C0",X"3A",X"EC",X"43",X"B7",X"28",X"04",X"DB",X"4A",
		X"18",X"02",X"DB",X"48",X"08",X"DB",X"60",X"0E",X"1F",X"CB",X"5F",X"28",X"02",X"CB",X"A1",X"CB",
		X"5F",X"3E",X"0F",X"28",X"02",X"A9",X"4F",X"08",X"A9",X"47",X"E6",X"0F",X"21",X"EF",X"43",X"4E",
		X"77",X"91",X"F2",X"38",X"C1",X"2F",X"C6",X"01",X"FE",X"08",X"DA",X"42",X"C1",X"F6",X"F0",X"2F",
		X"C6",X"01",X"21",X"EE",X"43",X"4F",X"CB",X"29",X"81",X"CB",X"60",X"20",X"04",X"86",X"77",X"18",
		X"04",X"47",X"7E",X"90",X"77",X"C9",X"7B",X"BD",X"38",X"01",X"EB",X"42",X"4B",X"E5",X"2E",X"00",
		X"60",X"E3",X"FD",X"E1",X"E5",X"2E",X"00",X"61",X"E3",X"7C",X"90",X"16",X"00",X"30",X"01",X"15",
		X"5F",X"7D",X"91",X"06",X"00",X"30",X"01",X"05",X"4F",X"E1",X"7B",X"B1",X"3E",X"01",X"28",X"21",
		X"3E",X"FF",X"08",X"7B",X"AA",X"17",X"38",X"0F",X"79",X"A8",X"17",X"38",X"0A",X"CB",X"23",X"CB",
		X"21",X"08",X"CB",X"3F",X"C3",X"82",X"C1",X"08",X"3C",X"C5",X"01",X"80",X"00",X"09",X"FD",X"09",
		X"C1",X"08",X"7C",X"FD",X"E5",X"D9",X"E1",X"6F",X"06",X"10",X"CD",X"68",X"2F",X"36",X"80",X"D9",
		X"08",X"09",X"FD",X"19",X"3D",X"C2",X"A1",X"C1",X"C9",X"EC",X"2A",X"AE",X"F8",X"7C",X"B5",X"C0",
		X"EB",X"22",X"AE",X"F8",X"C9",X"01",X"D8",X"01",X"F8",X"DE",X"F8",X"DE",X"D8",X"01",X"D8",X"FE",
		X"02",X"DB",X"44",X"DB",X"FE",X"02",X"DC",X"44",X"DC",X"FE",X"02",X"DD",X"44",X"DD",X"FE",X"02",
		X"DE",X"44",X"DE",X"FE",X"02",X"DF",X"44",X"DF",X"FE",X"02",X"E0",X"44",X"E0",X"FE",X"02",X"E3",
		X"44",X"E3",X"FE",X"02",X"E4",X"44",X"E4",X"FE",X"02",X"E5",X"44",X"E5",X"FE",X"02",X"E6",X"44",
		X"E6",X"FE",X"02",X"E7",X"44",X"E7",X"FE",X"02",X"E8",X"44",X"E8",X"FE",X"03",X"F8",X"03",X"EE",
		X"44",X"EE",X"44",X"F8",X"FF",X"01",X"23",X"1C",X"12",X"1E",X"10",X"10",X"10",X"00",X"0C",X"12",
		X"12",X"12",X"12",X"0C",X"00",X"11",X"11",X"11",X"15",X"15",X"0E",X"00",X"1E",X"10",X"18",X"10",
		X"10",X"1E",X"00",X"1C",X"12",X"1E",X"18",X"14",X"12",X"00",X"01",X"23",X"0E",X"09",X"0E",X"0E",
		X"09",X"0E",X"00",X"06",X"09",X"09",X"09",X"09",X"06",X"00",X"09",X"0D",X"0D",X"0B",X"0B",X"09",
		X"00",X"09",X"09",X"09",X"09",X"09",X"06",X"00",X"07",X"08",X"06",X"01",X"01",X"0E",X"00",X"01",
		X"23",X"06",X"09",X"0F",X"09",X"09",X"09",X"00",X"09",X"0D",X"0D",X"0B",X"0B",X"09",X"00",X"07",
		X"08",X"08",X"0B",X"09",X"06",X"00",X"08",X"08",X"08",X"08",X"08",X"0F",X"00",X"0F",X"08",X"0C",
		X"08",X"08",X"0F",X"00",X"02",X"05",X"08",X"BA",X"0D",X"93",X"0A",X"92",X"08",X"92",X"08",X"BA",
		X"02",X"05",X"5C",X"60",X"50",X"80",X"DC",X"40",X"50",X"20",X"5C",X"C0",X"02",X"04",X"0F",X"1E",
		X"0F",X"1E",X"0F",X"1E",X"0F",X"1E",X"02",X"04",X"3C",X"78",X"3C",X"78",X"3C",X"78",X"3C",X"78",
		X"02",X"05",X"0E",X"7A",X"09",X"4A",X"0E",X"4A",X"09",X"4A",X"0E",X"7B",X"02",X"05",X"3E",X"60",
		X"08",X"80",X"08",X"40",X"08",X"20",X"C8",X"C0",X"02",X"05",X"07",X"0C",X"04",X"92",X"07",X"1E",
		X"05",X"12",X"04",X"92",X"02",X"05",X"32",X"40",X"42",X"80",X"43",X"00",X"42",X"80",X"32",X"40",
		X"02",X"05",X"04",X"1E",X"04",X"10",X"04",X"18",X"04",X"10",X"07",X"9E",X"02",X"05",X"79",X"C0",
		X"40",X"80",X"60",X"80",X"40",X"80",X"40",X"80",X"02",X"05",X"1C",X"E6",X"21",X"09",X"19",X"09",
		X"05",X"09",X"38",X"E6",X"02",X"05",X"73",X"9C",X"4A",X"20",X"73",X"18",X"52",X"04",X"4B",X"B8",
		X"01",X"3B",X"00",X"16",X"F0",X"3E",X"AA",X"E6",X"0F",X"5F",X"3E",X"08",X"CD",X"B9",X"CC",X"01",
		X"3B",X"01",X"16",X"F0",X"3E",X"BB",X"E6",X"0F",X"5F",X"3E",X"06",X"CD",X"B9",X"CC",X"01",X"FB",
		X"01",X"16",X"F0",X"3E",X"99",X"E6",X"0F",X"5F",X"3E",X"02",X"CD",X"B9",X"CC",X"01",X"3C",X"00",
		X"16",X"F0",X"3E",X"AA",X"E6",X"0F",X"5F",X"3E",X"0C",X"CD",X"B9",X"CC",X"01",X"BC",X"01",X"16",
		X"F0",X"3E",X"BB",X"E6",X"0F",X"5F",X"3E",X"03",X"CD",X"B9",X"CC",X"01",X"1C",X"02",X"16",X"F0",
		X"3E",X"99",X"E6",X"0F",X"5F",X"3E",X"01",X"CD",X"B9",X"CC",X"01",X"3E",X"00",X"16",X"F0",X"3E",
		X"99",X"E6",X"0F",X"5F",X"3E",X"10",X"CD",X"B9",X"CC",X"01",X"3E",X"00",X"16",X"0F",X"3E",X"99",
		X"E6",X"F0",X"5F",X"3E",X"10",X"CD",X"B9",X"CC",X"01",X"C5",X"C1",X"CD",X"4F",X"C6",X"21",X"D9",
		X"48",X"11",X"15",X"C2",X"CD",X"E0",X"C6",X"01",X"5B",X"02",X"16",X"F0",X"3E",X"22",X"E6",X"0F",
		X"5F",X"3E",X"09",X"CD",X"B9",X"CC",X"01",X"5C",X"02",X"16",X"0F",X"3E",X"22",X"E6",X"F0",X"5F",
		X"3E",X"09",X"CD",X"B9",X"CC",X"21",X"E0",X"48",X"11",X"3A",X"C2",X"CD",X"E0",X"C6",X"01",X"5C",
		X"02",X"16",X"F0",X"3E",X"BB",X"E6",X"0F",X"5F",X"3E",X"09",X"CD",X"B9",X"CC",X"21",X"EC",X"48",
		X"11",X"5F",X"C2",X"CD",X"E0",X"C6",X"01",X"5E",X"02",X"16",X"0F",X"3E",X"EE",X"E6",X"F0",X"5F",
		X"3E",X"09",X"CD",X"B9",X"CC",X"21",X"D9",X"6F",X"11",X"84",X"C2",X"CD",X"E0",X"C6",X"21",X"E9",
		X"6F",X"11",X"90",X"C2",X"CD",X"E0",X"C6",X"01",X"DB",X"03",X"16",X"AA",X"1E",X"00",X"3E",X"07",
		X"CD",X"EF",X"CC",X"21",X"D8",X"78",X"11",X"9C",X"C2",X"CD",X"E0",X"C6",X"21",X"E8",X"78",X"11",
		X"A6",X"C2",X"CD",X"E0",X"C6",X"21",X"D9",X"80",X"11",X"B0",X"C2",X"CD",X"E0",X"C6",X"21",X"E9",
		X"80",X"11",X"BC",X"C2",X"CD",X"E0",X"C6",X"01",X"5B",X"04",X"16",X"AA",X"1E",X"00",X"3E",X"07",
		X"CD",X"EF",X"CC",X"21",X"D8",X"88",X"11",X"9C",X"C2",X"CD",X"E0",X"C6",X"21",X"E8",X"88",X"11",
		X"A6",X"C2",X"CD",X"E0",X"C6",X"01",X"9B",X"04",X"16",X"55",X"1E",X"00",X"3E",X"06",X"CD",X"EF",
		X"CC",X"01",X"BB",X"04",X"16",X"55",X"1E",X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"21",X"D9",X"90",
		X"11",X"C8",X"C2",X"CD",X"E0",X"C6",X"21",X"E9",X"90",X"11",X"D4",X"C2",X"CD",X"E0",X"C6",X"21",
		X"BE",X"43",X"11",X"E2",X"98",X"06",X"02",X"CD",X"B5",X"30",X"01",X"DB",X"04",X"16",X"33",X"1E",
		X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"01",X"FB",X"04",X"16",X"33",X"1E",X"00",X"3E",X"06",X"CD",
		X"EF",X"CC",X"01",X"1B",X"05",X"16",X"55",X"1E",X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"01",X"3B",
		X"05",X"16",X"55",X"1E",X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"21",X"D9",X"A2",X"11",X"E0",X"C2",
		X"CD",X"E0",X"C6",X"21",X"E9",X"A2",X"11",X"EC",X"C2",X"CD",X"E0",X"C6",X"21",X"BF",X"43",X"11",
		X"E2",X"AA",X"06",X"02",X"CD",X"B5",X"30",X"01",X"5B",X"05",X"16",X"33",X"1E",X"00",X"3E",X"06",
		X"CD",X"EF",X"CC",X"01",X"7B",X"05",X"16",X"33",X"1E",X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"21",
		X"D9",X"B5",X"11",X"F8",X"C2",X"CD",X"E0",X"C6",X"21",X"E9",X"B5",X"11",X"04",X"C3",X"CD",X"E0",
		X"C6",X"01",X"FB",X"05",X"16",X"DD",X"1E",X"00",X"3E",X"07",X"CD",X"EF",X"CC",X"01",X"1B",X"06",
		X"16",X"DD",X"1E",X"00",X"3E",X"07",X"CD",X"EF",X"CC",X"01",X"5B",X"06",X"16",X"EE",X"1E",X"00",
		X"3E",X"07",X"CD",X"EF",X"CC",X"01",X"7B",X"06",X"16",X"EE",X"1E",X"00",X"3E",X"07",X"CD",X"EF",
		X"CC",X"21",X"73",X"43",X"11",X"D6",X"D5",X"06",X"06",X"CD",X"B5",X"30",X"01",X"1F",X"00",X"16",
		X"F0",X"3E",X"00",X"E6",X"0F",X"5F",X"3E",X"37",X"CD",X"B9",X"CC",X"3E",X"FF",X"32",X"E0",X"43",
		X"C9",X"01",X"1B",X"05",X"16",X"55",X"1E",X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"01",X"3B",X"05",
		X"16",X"55",X"1E",X"00",X"3E",X"06",X"CD",X"EF",X"CC",X"01",X"5B",X"05",X"16",X"11",X"1E",X"00",
		X"3E",X"06",X"CD",X"EF",X"CC",X"01",X"7B",X"05",X"16",X"11",X"1E",X"00",X"3E",X"06",X"CD",X"EF",
		X"CC",X"C9",X"3A",X"E0",X"43",X"B7",X"28",X"18",X"CD",X"72",X"C6",X"21",X"E2",X"AA",X"06",X"03",
		X"0E",X"08",X"CD",X"AF",X"C6",X"21",X"BF",X"43",X"11",X"E2",X"AA",X"06",X"02",X"CD",X"B5",X"30",
		X"CD",X"06",X"C7",X"CD",X"0D",X"C6",X"CD",X"1D",X"C6",X"C9",X"0E",X"99",X"18",X"02",X"0E",X"22",
		X"C5",X"47",X"79",X"21",X"5A",X"85",X"CD",X"2A",X"C7",X"28",X"03",X"21",X"A5",X"83",X"CB",X"78",
		X"CB",X"B8",X"28",X"0B",X"21",X"DA",X"84",X"CD",X"2A",X"C7",X"28",X"03",X"21",X"25",X"84",X"48",
		X"06",X"00",X"CD",X"2A",X"C7",X"28",X"0C",X"B7",X"ED",X"42",X"0D",X"20",X"0E",X"E6",X"F0",X"F6",
		X"07",X"18",X"08",X"09",X"0D",X"20",X"04",X"E6",X"0F",X"F6",X"70",X"77",X"C1",X"C9",X"C5",X"F5",
		X"3A",X"F6",X"43",X"6F",X"0E",X"00",X"CD",X"F5",X"C5",X"F1",X"32",X"F6",X"43",X"6F",X"0E",X"FF",
		X"CD",X"F5",X"C5",X"C1",X"C9",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"11",X"9E",X"44",X"CD",
		X"2A",X"C7",X"28",X"06",X"11",X"61",X"5F",X"CD",X"8F",X"21",X"19",X"71",X"C9",X"21",X"9B",X"44",
		X"CD",X"2A",X"C7",X"28",X"03",X"21",X"64",X"5F",X"3A",X"C1",X"43",X"18",X"0E",X"21",X"9C",X"44",
		X"CD",X"2A",X"C7",X"28",X"03",X"21",X"63",X"5F",X"3A",X"C0",X"43",X"0E",X"0F",X"06",X"40",X"11",
		X"20",X"00",X"CD",X"2A",X"C7",X"28",X"05",X"11",X"E0",X"FF",X"0E",X"F0",X"B8",X"38",X"06",X"08",
		X"7E",X"B1",X"77",X"18",X"05",X"08",X"7E",X"B1",X"A9",X"77",X"08",X"19",X"10",X"EE",X"C9",X"0A",
		X"03",X"57",X"0A",X"03",X"5F",X"0A",X"03",X"67",X"0A",X"03",X"6F",X"E5",X"C5",X"CD",X"56",X"C1",
		X"C1",X"D1",X"0A",X"FE",X"FD",X"DA",X"55",X"C6",X"03",X"3C",X"C8",X"3C",X"CA",X"4F",X"C6",X"C3",
		X"55",X"C6",X"CD",X"96",X"C6",X"AF",X"32",X"E0",X"43",X"11",X"D6",X"BE",X"21",X"AF",X"43",X"06",
		X"06",X"CD",X"B5",X"30",X"3A",X"E9",X"43",X"FE",X"02",X"C0",X"11",X"D6",X"C8",X"21",X"B2",X"43",
		X"06",X"06",X"CD",X"B5",X"30",X"C9",X"26",X"BE",X"2E",X"D8",X"0E",X"10",X"06",X"04",X"CD",X"AF",
		X"C6",X"FD",X"E5",X"11",X"D8",X"BD",X"21",X"D8",X"CF",X"CD",X"56",X"C1",X"FD",X"E1",X"C9",X"C5",
		X"CD",X"2A",X"C7",X"28",X"08",X"3E",X"E0",X"80",X"5F",X"16",X"FF",X"18",X"06",X"3E",X"20",X"90",
		X"5F",X"16",X"00",X"06",X"00",X"CD",X"68",X"2F",X"C1",X"78",X"08",X"08",X"47",X"08",X"36",X"00",
		X"CD",X"2A",X"C7",X"20",X"03",X"23",X"18",X"01",X"2B",X"10",X"F3",X"19",X"0D",X"20",X"EC",X"C9",
		X"CD",X"66",X"2F",X"EB",X"CD",X"07",X"2D",X"C9",X"21",X"C0",X"43",X"7E",X"FE",X"40",X"D0",X"34",
		X"C9",X"21",X"C0",X"43",X"7E",X"FE",X"1F",X"20",X"08",X"D9",X"11",X"AD",X"C0",X"CD",X"BA",X"C1",
		X"D9",X"7E",X"B7",X"C8",X"35",X"C9",X"21",X"C1",X"43",X"7E",X"FE",X"20",X"20",X"DD",X"D9",X"11",
		X"B9",X"C0",X"CD",X"BA",X"C1",X"D9",X"18",X"D3",X"21",X"C1",X"43",X"7E",X"FE",X"1F",X"20",X"E1",
		X"D9",X"11",X"B3",X"C0",X"CD",X"BA",X"C1",X"D9",X"18",X"D7",X"E5",X"21",X"EC",X"43",X"CB",X"46",
		X"E1",X"C9",X"D9",X"C1",X"D1",X"E1",X"19",X"E5",X"C5",X"D9",X"C9",X"D9",X"C1",X"D1",X"E1",X"B7",
		X"ED",X"52",X"E5",X"C5",X"D9",X"C9",X"D9",X"C1",X"D1",X"7A",X"16",X"00",X"21",X"00",X"00",X"C5",
		X"06",X"08",X"29",X"CB",X"17",X"30",X"01",X"19",X"10",X"F8",X"C1",X"E5",X"C5",X"D9",X"C9",X"21",
		X"5D",X"F9",X"06",X"04",X"34",X"23",X"10",X"FC",X"3A",X"E4",X"43",X"FE",X"FF",X"20",X"04",X"AF",
		X"32",X"E4",X"43",X"47",X"3A",X"BF",X"43",X"90",X"38",X"1D",X"28",X"1B",X"3A",X"E4",X"43",X"B7",
		X"28",X"0D",X"FE",X"05",X"30",X"11",X"3A",X"5D",X"F9",X"21",X"BA",X"43",X"BE",X"38",X"08",X"AF",
		X"32",X"5D",X"F9",X"CD",X"CB",X"27",X"C9",X"B7",X"C9",X"3A",X"E1",X"43",X"B7",X"C0",X"21",X"C7",
		X"C7",X"3A",X"BE",X"43",X"4F",X"DB",X"62",X"06",X"06",X"CB",X"3F",X"10",X"FC",X"3D",X"81",X"BE",
		X"28",X"0B",X"3E",X"FF",X"BE",X"C8",X"11",X"07",X"00",X"19",X"C3",X"A1",X"C7",X"23",X"01",X"06",
		X"00",X"11",X"B7",X"43",X"ED",X"B0",X"C9",X"02",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"10",
		X"00",X"01",X"10",X"20",X"24",X"04",X"20",X"00",X"02",X"0F",X"18",X"20",X"05",X"30",X"01",X"02",
		X"13",X"10",X"1C",X"06",X"40",X"01",X"02",X"12",X"10",X"18",X"07",X"50",X"01",X"02",X"10",X"10",
		X"14",X"08",X"60",X"01",X"02",X"10",X"0F",X"10",X"09",X"80",X"01",X"02",X"10",X"0E",X"10",X"10",
		X"FF",X"01",X"02",X"0F",X"0D",X"10",X"11",X"FF",X"01",X"02",X"0F",X"0C",X"10",X"15",X"FF",X"02",
		X"02",X"0F",X"0A",X"10",X"FF",X"3A",X"B9",X"43",X"47",X"3A",X"F0",X"43",X"B8",X"D0",X"3A",X"BB",
		X"43",X"21",X"5E",X"F9",X"BE",X"D0",X"AF",X"32",X"5E",X"F9",X"21",X"BC",X"43",X"FD",X"21",X"77",
		X"40",X"FD",X"7E",X"0B",X"DD",X"96",X"0B",X"C6",X"07",X"F2",X"3E",X"C8",X"ED",X"44",X"BE",X"DA",
		X"97",X"C7",X"FD",X"7E",X"11",X"DD",X"96",X"11",X"C6",X"07",X"F2",X"4F",X"C8",X"ED",X"44",X"BE",
		X"DA",X"97",X"C7",X"CD",X"CB",X"27",X"C9",X"CD",X"6A",X"29",X"DD",X"CB",X"00",X"DE",X"CD",X"EF",
		X"CB",X"21",X"20",X"0A",X"06",X"15",X"0E",X"3C",X"CD",X"AF",X"C6",X"CD",X"05",X"1F",X"2D",X"C9",
		X"54",X"C9",X"7F",X"C9",X"A7",X"C9",X"CD",X"92",X"C8",X"CD",X"B9",X"C8",X"CD",X"72",X"C6",X"21",
		X"BE",X"43",X"7E",X"C6",X"01",X"27",X"77",X"3E",X"8C",X"CD",X"40",X"28",X"21",X"B6",X"43",X"7E",
		X"B7",X"C9",X"21",X"20",X"AA",X"06",X"16",X"0E",X"18",X"CD",X"AF",X"C6",X"21",X"60",X"B0",X"11",
		X"86",X"08",X"CD",X"E0",X"C6",X"CD",X"40",X"2F",X"00",X"70",X"B4",X"20",X"2D",X"20",X"00",X"08",
		X"06",X"02",X"21",X"B6",X"43",X"CD",X"AA",X"2F",X"C9",X"CD",X"40",X"2F",X"00",X"20",X"28",X"42",
		X"6F",X"6E",X"75",X"73",X"20",X"2D",X"20",X"20",X"20",X"20",X"20",X"30",X"00",X"21",X"40",X"40",
		X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"2B",X"2B",X"DD",X"21",X"C0",X"43",X"DD",X"7E",
		X"00",X"B7",X"C8",X"CD",X"BE",X"3D",X"DD",X"E5",X"3A",X"BE",X"43",X"F5",X"21",X"42",X"40",X"06",
		X"04",X"0E",X"05",X"CD",X"21",X"C9",X"01",X"05",X"00",X"CD",X"C3",X"2E",X"F1",X"3D",X"20",X"EB",
		X"21",X"40",X"40",X"06",X"06",X"11",X"58",X"28",X"CD",X"A0",X"2F",X"CD",X"D4",X"3D",X"DD",X"E1",
		X"DD",X"35",X"00",X"F5",X"CD",X"1D",X"C6",X"F1",X"28",X"04",X"DD",X"E5",X"18",X"CA",X"C3",X"51",
		X"3A",X"79",X"86",X"27",X"77",X"D0",X"2B",X"05",X"C8",X"0E",X"01",X"18",X"F4",X"CD",X"40",X"2F",
		X"00",X"20",X"14",X"52",X"61",X"63",X"6B",X"20",X"00",X"06",X"02",X"21",X"BE",X"43",X"CD",X"AA",
		X"2F",X"CD",X"40",X"2F",X"00",X"60",X"14",X"20",X"63",X"6F",X"6D",X"70",X"6C",X"65",X"74",X"65",
		X"64",X"2E",X"00",X"C9",X"CD",X"40",X"2F",X"00",X"00",X"14",X"20",X"00",X"06",X"02",X"21",X"BE",
		X"43",X"CD",X"AA",X"2F",X"CD",X"40",X"2F",X"00",X"28",X"14",X"52",X"75",X"6E",X"64",X"65",X"20",
		X"61",X"62",X"67",X"65",X"73",X"63",X"68",X"6C",X"6F",X"73",X"73",X"65",X"6E",X"00",X"C9",X"CD",
		X"40",X"2F",X"00",X"20",X"14",X"4D",X"61",X"6E",X"63",X"68",X"65",X"20",X"00",X"06",X"02",X"21",
		X"BE",X"43",X"CD",X"AA",X"2F",X"CD",X"40",X"2F",X"00",X"70",X"14",X"20",X"74",X"65",X"72",X"6D",
		X"69",X"6E",X"65",X"65",X"2E",X"00",X"C9",X"CD",X"40",X"2F",X"00",X"08",X"14",X"50",X"61",X"72",
		X"74",X"69",X"64",X"61",X"20",X"6E",X"6F",X"2E",X"20",X"00",X"06",X"02",X"21",X"BE",X"43",X"CD",
		X"AA",X"2F",X"CD",X"40",X"2F",X"00",X"80",X"14",X"20",X"74",X"65",X"72",X"6D",X"69",X"6E",X"61",
		X"64",X"61",X"00",X"C9",X"21",X"00",X"00",X"39",X"31",X"86",X"F8",X"E5",X"3A",X"BD",X"43",X"3C",
		X"32",X"BD",X"43",X"E1",X"F9",X"C3",X"1B",X"25",X"C5",X"D5",X"CD",X"E4",X"05",X"7E",X"B7",X"28",
		X"08",X"D1",X"7A",X"C6",X"0E",X"57",X"C1",X"18",X"EF",X"D1",X"C1",X"C9",X"CD",X"B0",X"28",X"CD",
		X"0B",X"28",X"CD",X"8D",X"CA",X"E5",X"CD",X"21",X"3C",X"E1",X"CD",X"0A",X"CB",X"21",X"F0",X"43",
		X"34",X"21",X"B7",X"43",X"CD",X"7C",X"2E",X"BE",X"30",X"17",X"DD",X"CB",X"14",X"C6",X"21",X"AC",
		X"19",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"CB",X"14",X"EE",X"DD",X"36",X"15",X"05",X"18",
		X"0D",X"21",X"9E",X"19",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"36",X"15",X"4B",X"DD",X"CB",
		X"00",X"CE",X"DD",X"E5",X"E1",X"FD",X"E5",X"CD",X"D1",X"2B",X"FD",X"E1",X"DD",X"CB",X"00",X"D6",
		X"DD",X"E5",X"CD",X"4B",X"28",X"DD",X"E1",X"DD",X"CB",X"00",X"7E",X"20",X"1D",X"DD",X"CB",X"14",
		X"7E",X"20",X"1E",X"CD",X"AA",X"20",X"DD",X"CB",X"14",X"46",X"20",X"05",X"DD",X"35",X"15",X"28",
		X"09",X"DD",X"E5",X"3E",X"01",X"CD",X"40",X"28",X"18",X"DB",X"21",X"F0",X"43",X"35",X"C3",X"4F",
		X"17",X"21",X"F0",X"43",X"35",X"CD",X"BD",X"28",X"CD",X"4B",X"28",X"18",X"FB",X"FD",X"21",X"77",
		X"40",X"DD",X"E5",X"DD",X"2A",X"F1",X"43",X"26",X"00",X"FD",X"6E",X"0B",X"16",X"00",X"1E",X"08",
		X"19",X"DD",X"5E",X"0B",X"ED",X"52",X"EB",X"26",X"00",X"FD",X"6E",X"11",X"06",X"00",X"0E",X"05",
		X"09",X"DD",X"4E",X"11",X"ED",X"42",X"7D",X"F6",X"01",X"6F",X"7B",X"AA",X"E6",X"80",X"20",X"0D",
		X"7D",X"AC",X"E6",X"80",X"20",X"07",X"CB",X"23",X"CB",X"25",X"C3",X"BA",X"CA",X"FD",X"E1",X"FD",
		X"72",X"09",X"FD",X"73",X"08",X"DD",X"36",X"07",X"00",X"DD",X"36",X"06",X"00",X"CD",X"02",X"CB",
		X"DD",X"72",X"09",X"DD",X"73",X"08",X"FD",X"74",X"0F",X"FD",X"75",X"0E",X"DD",X"36",X"0D",X"00",
		X"DD",X"36",X"0C",X"00",X"CD",X"02",X"CB",X"DD",X"72",X"0F",X"DD",X"73",X"0E",X"FD",X"E5",X"DD",
		X"E1",X"C9",X"7A",X"2F",X"57",X"7B",X"2F",X"5F",X"13",X"C9",X"16",X"08",X"1E",X"08",X"DD",X"7E",
		X"09",X"B7",X"F2",X"19",X"CB",X"7A",X"ED",X"44",X"57",X"DD",X"7E",X"0F",X"B7",X"F2",X"24",X"CB",
		X"7B",X"ED",X"44",X"5F",X"FD",X"2A",X"F1",X"43",X"FD",X"7E",X"0B",X"82",X"C6",X"04",X"DD",X"77",
		X"0B",X"FD",X"7E",X"11",X"83",X"C6",X"04",X"DD",X"77",X"11",X"C9",X"CD",X"39",X"CD",X"CD",X"71",
		X"CC",X"1B",X"00",X"38",X"05",X"77",X"C9",X"CD",X"71",X"CC",X"00",X"00",X"04",X"20",X"AA",X"CD",
		X"71",X"CC",X"80",X"00",X"01",X"20",X"FF",X"CD",X"71",X"CC",X"A0",X"00",X"29",X"20",X"11",X"CD",
		X"71",X"CC",X"A0",X"00",X"29",X"09",X"99",X"CD",X"71",X"CC",X"A9",X"00",X"29",X"08",X"BB",X"CD",
		X"71",X"CC",X"B0",X"00",X"29",X"10",X"55",X"CD",X"71",X"CC",X"C0",X"05",X"0A",X"20",X"77",X"CD",
		X"71",X"CC",X"80",X"06",X"04",X"0A",X"DD",X"CD",X"71",X"CC",X"96",X"06",X"04",X"0A",X"EE",X"C9",
		X"CD",X"71",X"CC",X"00",X"00",X"38",X"20",X"AA",X"C9",X"CD",X"71",X"CC",X"00",X"00",X"38",X"20",
		X"FF",X"C9",X"CD",X"71",X"CC",X"E0",X"05",X"04",X"20",X"33",X"C9",X"CD",X"71",X"CC",X"E0",X"05",
		X"04",X"20",X"99",X"C9",X"CD",X"71",X"CC",X"E0",X"05",X"04",X"20",X"66",X"C9",X"CD",X"71",X"CC",
		X"00",X"00",X"08",X"20",X"BB",X"CD",X"71",X"CC",X"00",X"01",X"10",X"20",X"66",X"CD",X"71",X"CC",
		X"00",X"03",X"04",X"20",X"FF",X"CD",X"71",X"CC",X"80",X"03",X"1C",X"20",X"AA",X"C9",X"CD",X"71",
		X"CC",X"00",X"00",X"2F",X"20",X"CC",X"CD",X"71",X"CC",X"E0",X"05",X"09",X"20",X"AA",X"C9",X"DD",
		X"E5",X"E1",X"CB",X"5E",X"CA",X"15",X"CC",X"CB",X"9E",X"E5",X"2A",X"61",X"F9",X"11",X"63",X"F9",
		X"3E",X"05",X"08",X"06",X"03",X"1A",X"13",X"77",X"23",X"10",X"FA",X"01",X"1D",X"00",X"09",X"08",
		X"3D",X"C2",X"02",X"CC",X"E1",X"CB",X"66",X"C8",X"CB",X"A6",X"E5",X"11",X"0B",X"00",X"19",X"5E",
		X"23",X"23",X"23",X"23",X"23",X"23",X"3A",X"EC",X"43",X"B7",X"7E",X"28",X"0A",X"ED",X"44",X"C6",
		X"D0",X"08",X"3E",X"F1",X"93",X"5F",X"08",X"CB",X"3F",X"CB",X"3F",X"67",X"6B",X"CB",X"3C",X"CB",
		X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"01",X"00",X"81",X"09",X"22",X"61",X"F9",
		X"3A",X"EB",X"43",X"11",X"1D",X"00",X"FD",X"21",X"63",X"F9",X"0E",X"05",X"06",X"03",X"08",X"7E",
		X"FD",X"77",X"00",X"FD",X"23",X"08",X"77",X"23",X"10",X"F4",X"19",X"0D",X"C2",X"5C",X"CC",X"E1",
		X"C9",X"E1",X"5E",X"23",X"56",X"23",X"E5",X"3A",X"EC",X"43",X"B7",X"20",X"06",X"21",X"00",X"81",
		X"19",X"18",X"05",X"21",X"FF",X"87",X"ED",X"52",X"EB",X"E1",X"4E",X"23",X"08",X"7E",X"23",X"08",
		X"B7",X"7E",X"23",X"E5",X"EB",X"20",X"11",X"11",X"20",X"00",X"08",X"47",X"08",X"E5",X"77",X"23",
		X"10",X"FC",X"E1",X"19",X"0D",X"20",X"F3",X"C9",X"11",X"E0",X"FF",X"08",X"47",X"08",X"E5",X"77",
		X"2B",X"10",X"FC",X"E1",X"19",X"0D",X"20",X"F3",X"C9",X"08",X"3A",X"EC",X"43",X"B7",X"28",X"1C",
		X"08",X"B7",X"21",X"FF",X"87",X"ED",X"42",X"01",X"E0",X"FF",X"CB",X"0A",X"CB",X"0A",X"CB",X"0A",
		X"CB",X"0A",X"CB",X"0B",X"CB",X"0B",X"CB",X"0B",X"CB",X"0B",X"18",X"08",X"08",X"21",X"00",X"81",
		X"09",X"01",X"20",X"00",X"08",X"7E",X"A2",X"B3",X"77",X"09",X"08",X"3D",X"20",X"F6",X"C9",X"CD",
		X"2A",X"C7",X"28",X"0D",X"B7",X"21",X"FF",X"87",X"ED",X"42",X"08",X"7B",X"2F",X"5F",X"08",X"18",
		X"04",X"21",X"00",X"81",X"09",X"47",X"4B",X"CB",X"41",X"C5",X"28",X"14",X"7E",X"1E",X"0F",X"A3",
		X"08",X"3E",X"F0",X"A2",X"5F",X"08",X"B3",X"77",X"CD",X"2A",X"C7",X"28",X"15",X"2B",X"18",X"12",
		X"7E",X"1E",X"F0",X"A3",X"08",X"3E",X"0F",X"A2",X"5F",X"08",X"B3",X"77",X"CD",X"2A",X"C7",X"20",
		X"01",X"23",X"C1",X"79",X"2F",X"4F",X"10",X"CF",X"C9",X"21",X"6E",X"CD",X"16",X"00",X"3A",X"BE",
		X"43",X"47",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"80",X"27",X"E6",X"07",X"5F",X"19",
		X"56",X"7A",X"32",X"EA",X"43",X"06",X"38",X"21",X"00",X"00",X"C5",X"E5",X"C1",X"C5",X"3E",X"40",
		X"1E",X"FF",X"CD",X"EF",X"CC",X"E1",X"01",X"20",X"00",X"09",X"C1",X"10",X"ED",X"C9",X"FF",X"AA",
		X"BB",X"DD",X"CC",X"77",X"EE",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
