library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_vec_rom3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_vec_rom3 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3B",X"44",X"23",X"43",X"35",X"43",X"07",X"59",X"00",X"C0",X"1C",X"49",X"3E",X"55",X"24",X"43",
		X"22",X"59",X"24",X"41",X"3E",X"46",X"24",X"41",X"36",X"47",X"04",X"57",X"00",X"C0",X"00",X"4A",
		X"3C",X"54",X"3C",X"54",X"28",X"44",X"28",X"5C",X"3C",X"4C",X"3C",X"4C",X"00",X"56",X"00",X"C0",
		X"04",X"49",X"38",X"57",X"37",X"56",X"29",X"41",X"26",X"59",X"21",X"4D",X"21",X"4C",X"1C",X"57",
		X"00",X"C0",X"07",X"47",X"35",X"5A",X"34",X"5B",X"29",X"5D",X"23",X"57",X"25",X"4C",X"26",X"4B",
		X"19",X"59",X"00",X"C0",X"09",X"44",X"34",X"5F",X"33",X"5F",X"27",X"5A",X"3F",X"57",X"2A",X"49",
		X"29",X"48",X"17",X"5C",X"00",X"C0",X"0A",X"40",X"34",X"44",X"34",X"44",X"24",X"58",X"3C",X"58",
		X"2C",X"44",X"2C",X"44",X"16",X"40",X"00",X"C0",X"09",X"5C",X"37",X"48",X"36",X"49",X"21",X"57",
		X"39",X"5A",X"2D",X"5F",X"2C",X"5F",X"17",X"44",X"00",X"C0",X"07",X"59",X"3A",X"4B",X"3B",X"4C",
		X"3D",X"57",X"37",X"5D",X"2C",X"5B",X"2B",X"5A",X"19",X"47",X"00",X"C0",X"04",X"57",X"3F",X"4C",
		X"3F",X"4D",X"3A",X"59",X"37",X"41",X"29",X"56",X"28",X"57",X"1C",X"49",X"00",X"C0",X"00",X"56",
		X"24",X"4C",X"24",X"4C",X"38",X"5C",X"38",X"44",X"24",X"54",X"24",X"54",X"00",X"4A",X"00",X"C0",
		X"1C",X"57",X"28",X"49",X"29",X"4A",X"37",X"5F",X"3A",X"47",X"3F",X"53",X"3F",X"54",X"04",X"49",
		X"00",X"C0",X"19",X"59",X"2B",X"46",X"2C",X"45",X"37",X"43",X"3D",X"49",X"3B",X"54",X"3A",X"55",
		X"07",X"47",X"00",X"C0",X"17",X"5C",X"2C",X"41",X"2D",X"41",X"39",X"46",X"21",X"49",X"36",X"57",
		X"37",X"58",X"09",X"44",X"00",X"C0",X"16",X"40",X"2C",X"5C",X"2C",X"5C",X"3C",X"48",X"24",X"48",
		X"34",X"5C",X"34",X"5C",X"0A",X"40",X"00",X"C0",X"17",X"44",X"29",X"58",X"2A",X"57",X"3F",X"49",
		X"27",X"46",X"33",X"41",X"34",X"41",X"09",X"5C",X"00",X"C0",X"19",X"47",X"26",X"55",X"25",X"54",
		X"23",X"49",X"29",X"43",X"34",X"45",X"35",X"46",X"07",X"59",X"00",X"C0",X"1C",X"49",X"21",X"54",
		X"21",X"53",X"26",X"47",X"29",X"5F",X"37",X"4A",X"38",X"49",X"04",X"57",X"00",X"C0",X"1E",X"43",
		X"3E",X"5D",X"21",X"5D",X"20",X"5E",X"3E",X"5E",X"20",X"5A",X"25",X"43",X"25",X"5D",X"20",X"46",
		X"3E",X"42",X"20",X"42",X"21",X"43",X"3E",X"43",X"3F",X"41",X"3E",X"40",X"3F",X"5F",X"02",X"5D",
		X"00",X"C0",X"1F",X"44",X"3D",X"5E",X"20",X"5C",X"3F",X"5F",X"3E",X"5E",X"3D",X"5B",X"26",X"41",
		X"24",X"5B",X"22",X"46",X"3D",X"42",X"23",X"42",X"22",X"42",X"3F",X"44",X"3F",X"41",X"3D",X"41",
		X"20",X"40",X"01",X"5C",X"00",X"C0",X"1F",X"44",X"3E",X"5F",X"3F",X"5D",X"3E",X"5F",X"3E",X"40",
		X"3B",X"5B",X"26",X"5F",X"21",X"5A",X"25",X"45",X"20",X"42",X"21",X"42",X"23",X"41",X"21",X"44",
		X"20",X"41",X"3E",X"42",X"3D",X"40",X"01",X"5C",X"00",X"C0",X"02",X"43",X"3C",X"41",X"3E",X"5E",
		X"3E",X"5F",X"3E",X"41",X"3A",X"5E",X"25",X"5C",X"3F",X"5A",X"25",X"43",X"22",X"42",X"21",X"41",
		X"24",X"40",X"22",X"45",X"20",X"40",X"3F",X"41",X"3F",X"41",X"1E",X"5D",X"00",X"C0",X"03",X"42",
		X"3D",X"42",X"3D",X"5F",X"3E",X"40",X"3E",X"42",X"3A",X"40",X"23",X"5B",X"3D",X"5B",X"26",X"40",
		X"22",X"42",X"22",X"40",X"23",X"5F",X"23",X"42",X"21",X"43",X"20",X"40",X"3F",X"41",X"1D",X"5E",
		X"00",X"C0",X"04",X"41",X"3E",X"43",X"3C",X"40",X"3F",X"41",X"3E",X"42",X"3B",X"43",X"21",X"5A",
		X"3B",X"5C",X"26",X"5E",X"22",X"43",X"22",X"5D",X"22",X"5E",X"24",X"41",X"21",X"41",X"21",X"43",
		X"20",X"40",X"1C",X"5F",X"00",X"C0",X"04",X"41",X"3F",X"42",X"3D",X"41",X"3F",X"42",X"20",X"42",
		X"3B",X"45",X"3F",X"5A",X"3A",X"5F",X"25",X"5B",X"22",X"40",X"22",X"5F",X"21",X"5D",X"22",X"5F",
		X"23",X"40",X"22",X"42",X"20",X"43",X"1C",X"5F",X"00",X"C0",X"03",X"5E",X"21",X"44",X"3E",X"42",
		X"3D",X"42",X"23",X"42",X"3E",X"46",X"3C",X"5B",X"3A",X"41",X"23",X"5B",X"22",X"5E",X"21",X"5F",
		X"20",X"5C",X"23",X"5E",X"20",X"40",X"23",X"41",X"21",X"41",X"1D",X"42",X"00",X"C0",X"02",X"5D",
		X"22",X"43",X"3F",X"43",X"20",X"42",X"22",X"42",X"20",X"46",X"3B",X"5D",X"3B",X"43",X"20",X"5A",
		X"22",X"5E",X"20",X"5E",X"3F",X"5D",X"22",X"5D",X"21",X"5F",X"22",X"40",X"21",X"41",X"1E",X"43",
		X"00",X"C0",X"1F",X"5C",X"25",X"42",X"20",X"44",X"21",X"41",X"22",X"42",X"23",X"45",X"3A",X"5F",
		X"3C",X"45",X"3E",X"5A",X"21",X"5E",X"3F",X"5E",X"3E",X"5E",X"21",X"5C",X"21",X"5F",X"21",X"5F",
		X"20",X"40",X"01",X"44",X"00",X"C0",X"1F",X"5C",X"24",X"41",X"21",X"43",X"22",X"41",X"22",X"40",
		X"25",X"45",X"3A",X"41",X"3F",X"46",X"3B",X"5B",X"20",X"5E",X"3F",X"5E",X"3D",X"5F",X"3F",X"5E",
		X"20",X"5D",X"22",X"5E",X"21",X"40",X"01",X"44",X"00",X"C0",X"1E",X"5D",X"24",X"5F",X"22",X"42",
		X"22",X"43",X"22",X"5D",X"26",X"42",X"3B",X"44",X"21",X"46",X"3B",X"5D",X"3E",X"5E",X"3F",X"5F",
		X"3C",X"40",X"3E",X"5D",X"20",X"40",X"21",X"5D",X"21",X"5F",X"02",X"43",X"00",X"C0",X"1D",X"5E",
		X"23",X"5E",X"23",X"41",X"22",X"40",X"22",X"5E",X"26",X"40",X"3D",X"45",X"23",X"45",X"3A",X"40",
		X"3E",X"5E",X"3E",X"40",X"3D",X"41",X"3D",X"5E",X"3F",X"5F",X"20",X"40",X"21",X"5D",X"03",X"42",
		X"00",X"C0",X"1C",X"41",X"22",X"5B",X"24",X"40",X"21",X"5F",X"22",X"5E",X"25",X"5D",X"3F",X"46",
		X"25",X"44",X"3A",X"42",X"3E",X"5F",X"3E",X"41",X"3E",X"42",X"3C",X"5F",X"3F",X"5F",X"3F",X"5F",
		X"20",X"40",X"04",X"5F",X"00",X"C0",X"1C",X"41",X"21",X"5C",X"23",X"5F",X"21",X"5E",X"20",X"5E",
		X"25",X"5B",X"21",X"46",X"26",X"41",X"3B",X"45",X"3E",X"40",X"3E",X"41",X"3F",X"43",X"3C",X"41",
		X"3F",X"40",X"3E",X"5E",X"20",X"5F",X"04",X"5F",X"00",X"C0",X"1D",X"42",X"3F",X"5C",X"22",X"5E",
		X"21",X"5E",X"3F",X"5E",X"22",X"5A",X"24",X"45",X"26",X"5F",X"3D",X"45",X"3E",X"42",X"3F",X"41",
		X"20",X"44",X"3B",X"42",X"20",X"40",X"3F",X"5F",X"3F",X"5F",X"03",X"5E",X"00",X"C0",X"1E",X"43",
		X"3A",X"5A",X"20",X"5A",X"26",X"5A",X"24",X"40",X"26",X"46",X"20",X"46",X"3A",X"46",X"1E",X"5D",
		X"00",X"C0",X"1F",X"44",X"38",X"5C",X"3E",X"5B",X"23",X"58",X"24",X"5E",X"28",X"44",X"22",X"45",
		X"3D",X"48",X"1D",X"5E",X"00",X"C0",X"1F",X"44",X"39",X"40",X"3C",X"5D",X"20",X"56",X"23",X"5D",
		X"28",X"40",X"25",X"44",X"20",X"49",X"1C",X"5F",X"00",X"C0",X"02",X"43",X"38",X"43",X"3B",X"5E",
		X"3C",X"58",X"22",X"5C",X"28",X"5D",X"25",X"42",X"24",X"4A",X"1C",X"5F",X"00",X"C0",X"03",X"42",
		X"3A",X"46",X"3A",X"40",X"3A",X"5A",X"20",X"5C",X"26",X"5A",X"26",X"40",X"26",X"46",X"1D",X"42",
		X"00",X"C0",X"04",X"41",X"3C",X"48",X"3B",X"42",X"38",X"5D",X"3E",X"5C",X"24",X"58",X"25",X"5E",
		X"28",X"43",X"1E",X"43",X"00",X"C0",X"04",X"41",X"20",X"47",X"3B",X"44",X"38",X"40",X"3D",X"5D",
		X"20",X"58",X"24",X"5B",X"27",X"40",X"01",X"44",X"00",X"C0",X"03",X"5E",X"23",X"48",X"3E",X"45",
		X"38",X"44",X"3C",X"5E",X"3D",X"58",X"22",X"5B",X"28",X"5C",X"01",X"44",X"00",X"C0",X"02",X"5D",
		X"26",X"46",X"20",X"46",X"3A",X"46",X"3C",X"40",X"3A",X"5A",X"20",X"5A",X"26",X"5A",X"02",X"43",
		X"00",X"C0",X"1F",X"5C",X"2A",X"44",X"22",X"45",X"3D",X"48",X"3C",X"42",X"38",X"5C",X"3E",X"5B",
		X"23",X"58",X"03",X"42",X"00",X"C0",X"1F",X"5C",X"29",X"40",X"24",X"45",X"20",X"48",X"3D",X"43",
		X"36",X"40",X"3D",X"5C",X"20",X"59",X"04",X"5F",X"00",X"C0",X"1E",X"5D",X"28",X"5D",X"25",X"42",
		X"24",X"48",X"3E",X"44",X"38",X"43",X"3B",X"5E",X"3C",X"58",X"04",X"5F",X"00",X"C0",X"1D",X"5E",
		X"26",X"5A",X"26",X"40",X"26",X"46",X"20",X"44",X"3A",X"46",X"3A",X"40",X"3A",X"5A",X"03",X"5E",
		X"00",X"C0",X"1C",X"41",X"24",X"56",X"25",X"5E",X"28",X"43",X"22",X"44",X"3C",X"48",X"3B",X"42",
		X"38",X"5D",X"02",X"5D",X"00",X"C0",X"1C",X"41",X"20",X"57",X"23",X"5C",X"2A",X"40",X"23",X"43",
		X"20",X"4A",X"3C",X"43",X"37",X"40",X"01",X"5C",X"00",X"C0",X"1D",X"42",X"3D",X"58",X"22",X"5B",
		X"28",X"5C",X"24",X"42",X"23",X"48",X"3E",X"45",X"36",X"44",X"01",X"5C",X"00",X"C0",X"02",X"43",
		X"22",X"43",X"3F",X"43",X"3E",X"41",X"21",X"5E",X"20",X"5E",X"3E",X"5E",X"3E",X"42",X"20",X"42",
		X"21",X"42",X"3E",X"5F",X"3F",X"5D",X"22",X"5D",X"02",X"5D",X"00",X"C0",X"03",X"42",X"23",X"42",
		X"20",X"43",X"3F",X"42",X"20",X"5E",X"3F",X"5E",X"3E",X"5F",X"3E",X"42",X"21",X"42",X"22",X"42",
		X"3C",X"5F",X"20",X"5E",X"20",X"5D",X"01",X"5C",X"00",X"C0",X"04",X"41",X"23",X"40",X"21",X"43",
		X"20",X"42",X"3F",X"5E",X"3F",X"5F",X"3D",X"40",X"20",X"43",X"21",X"41",X"22",X"41",X"3E",X"40",
		X"3D",X"5F",X"3E",X"5D",X"01",X"5C",X"00",X"C0",X"04",X"41",X"23",X"5E",X"22",X"42",X"21",X"42",
		X"3E",X"5E",X"3E",X"5F",X"3E",X"42",X"21",X"42",X"22",X"41",X"22",X"40",X"3E",X"41",X"3D",X"40",
		X"3E",X"5D",X"1E",X"5D",X"00",X"C0",X"4E",X"00",X"03",X"5E",X"23",X"5E",X"23",X"41",X"21",X"44",
		X"3E",X"5D",X"3E",X"40",X"3E",X"42",X"22",X"42",X"22",X"40",X"22",X"5F",X"3F",X"42",X"3D",X"41",
		X"3D",X"5E",X"1D",X"5E",X"00",X"C0",X"02",X"5D",X"22",X"5D",X"23",X"40",X"22",X"41",X"3E",X"40",
		X"3E",X"41",X"3F",X"42",X"22",X"42",X"22",X"5F",X"22",X"5E",X"3F",X"44",X"3E",X"40",X"3D",X"40",
		X"1C",X"5F",X"00",X"C0",X"1F",X"5C",X"22",X"5D",X"23",X"5F",X"22",X"40",X"3E",X"41",X"3F",X"41",
		X"20",X"43",X"23",X"40",X"21",X"5F",X"21",X"5E",X"20",X"42",X"3F",X"43",X"3D",X"42",X"1C",X"5F",
		X"00",X"C0",X"1F",X"5C",X"20",X"5D",X"20",X"5E",X"24",X"5F",X"3E",X"42",X"3F",X"42",X"22",X"42",
		X"22",X"5F",X"21",X"5E",X"20",X"5E",X"21",X"42",X"20",X"43",X"3D",X"42",X"1D",X"42",X"00",X"C0",
		X"1E",X"5D",X"3E",X"5D",X"21",X"5D",X"22",X"5F",X"3F",X"42",X"20",X"42",X"22",X"42",X"22",X"5E",
		X"20",X"5E",X"3F",X"5E",X"22",X"41",X"21",X"43",X"3E",X"43",X"1E",X"43",X"00",X"C0",X"1D",X"5E",
		X"3D",X"5E",X"20",X"5D",X"21",X"5E",X"20",X"42",X"21",X"42",X"22",X"41",X"22",X"5E",X"3F",X"5E",
		X"3E",X"5E",X"22",X"41",X"22",X"42",X"3E",X"43",X"01",X"44",X"00",X"C0",X"1C",X"41",X"3D",X"5E",
		X"3F",X"5D",X"20",X"5E",X"21",X"42",X"21",X"41",X"23",X"40",X"20",X"5D",X"3F",X"5F",X"3E",X"5F",
		X"22",X"40",X"23",X"41",X"20",X"43",X"01",X"44",X"00",X"C0",X"1C",X"41",X"3D",X"40",X"3E",X"40",
		X"3F",X"5C",X"22",X"42",X"22",X"41",X"22",X"5E",X"3F",X"5E",X"3E",X"5F",X"3E",X"40",X"22",X"5F",
		X"23",X"40",X"22",X"43",X"02",X"43",X"00",X"C0",X"1D",X"42",X"3D",X"42",X"3D",X"5F",X"3F",X"5E",
		X"22",X"41",X"22",X"40",X"22",X"5E",X"3E",X"5E",X"3E",X"40",X"3E",X"43",X"21",X"5C",X"23",X"5F",
		X"23",X"42",X"03",X"42",X"00",X"C0",X"1E",X"43",X"3E",X"43",X"3D",X"40",X"3E",X"5F",X"22",X"40",
		X"22",X"5F",X"21",X"5E",X"3E",X"5E",X"3E",X"41",X"3E",X"42",X"21",X"5E",X"22",X"5E",X"23",X"42",
		X"04",X"5F",X"00",X"C0",X"1F",X"44",X"20",X"43",X"3D",X"41",X"3E",X"40",X"22",X"5F",X"21",X"5F",
		X"20",X"5D",X"3D",X"40",X"3F",X"41",X"3F",X"42",X"20",X"5E",X"21",X"5D",X"23",X"40",X"04",X"5F",
		X"00",X"C0",X"1F",X"44",X"22",X"43",X"3E",X"42",X"3E",X"41",X"22",X"5E",X"21",X"5E",X"3E",X"5E",
		X"3E",X"41",X"3F",X"42",X"20",X"42",X"3F",X"5E",X"20",X"5D",X"23",X"5E",X"03",X"5E",X"00",X"C0",
		X"02",X"43",X"23",X"43",X"3F",X"43",X"3E",X"41",X"21",X"5E",X"20",X"5E",X"3D",X"5E",X"3D",X"42",
		X"20",X"42",X"21",X"42",X"3E",X"5F",X"3F",X"5D",X"23",X"5D",X"02",X"5D",X"00",X"C0",X"03",X"42",
		X"24",X"42",X"20",X"43",X"3F",X"41",X"20",X"5E",X"3F",X"5E",X"3D",X"40",X"3E",X"43",X"20",X"42",
		X"22",X"41",X"3E",X"40",X"3E",X"5D",X"21",X"5D",X"01",X"5C",X"00",X"C0",X"04",X"41",X"24",X"40",
		X"21",X"43",X"3F",X"42",X"20",X"5E",X"3E",X"5E",X"3D",X"41",X"3F",X"43",X"22",X"42",X"22",X"40",
		X"3E",X"41",X"3B",X"5F",X"20",X"5C",X"01",X"5C",X"00",X"C0",X"04",X"41",X"23",X"5D",X"23",X"42",
		X"20",X"42",X"3F",X"5E",X"3E",X"40",X"3D",X"42",X"20",X"43",X"22",X"41",X"22",X"40",X"3F",X"41",
		X"3D",X"40",X"3E",X"5C",X"1E",X"5D",X"00",X"C0",X"03",X"5E",X"23",X"5D",X"23",X"41",X"21",X"42",
		X"3E",X"5F",X"3E",X"40",X"3E",X"43",X"22",X"43",X"22",X"40",X"22",X"5F",X"3F",X"42",X"3D",X"41",
		X"3D",X"5D",X"1D",X"5E",X"00",X"C0",X"02",X"5D",X"22",X"5C",X"23",X"40",X"21",X"41",X"3E",X"40",
		X"3E",X"41",X"20",X"43",X"23",X"42",X"22",X"40",X"21",X"5E",X"20",X"42",X"3D",X"42",X"3D",X"5F",
		X"1C",X"5F",X"00",X"C0",X"1F",X"5C",X"20",X"5C",X"25",X"5F",X"22",X"41",X"3E",X"40",X"3E",X"42",
		X"21",X"43",X"23",X"41",X"22",X"5E",X"20",X"5E",X"21",X"42",X"3F",X"45",X"3C",X"40",X"1C",X"5F",
		X"00",X"C0",X"1F",X"5C",X"3F",X"5D",X"22",X"5D",X"22",X"40",X"3E",X"41",X"20",X"42",X"22",X"43",
		X"23",X"40",X"21",X"5E",X"20",X"5E",X"21",X"41",X"20",X"43",X"3C",X"42",X"1D",X"42",X"00",X"C0",
		X"1E",X"5D",X"3D",X"5D",X"21",X"5D",X"22",X"5F",X"3F",X"42",X"20",X"42",X"23",X"42",X"23",X"5E",
		X"20",X"5E",X"3F",X"5E",X"22",X"41",X"21",X"43",X"3D",X"43",X"1E",X"43",X"00",X"C0",X"1D",X"5E",
		X"3C",X"5E",X"20",X"5D",X"21",X"5F",X"20",X"42",X"21",X"42",X"23",X"40",X"22",X"5D",X"20",X"5E",
		X"3E",X"5F",X"22",X"40",X"22",X"43",X"3D",X"43",X"01",X"44",X"00",X"C0",X"1C",X"41",X"3C",X"40",
		X"3F",X"5B",X"21",X"5E",X"20",X"42",X"22",X"42",X"23",X"5F",X"21",X"5D",X"3E",X"5E",X"3E",X"40",
		X"22",X"5F",X"23",X"41",X"20",X"44",X"01",X"44",X"00",X"C0",X"1C",X"41",X"3D",X"41",X"3D",X"5E",
		X"20",X"5E",X"21",X"42",X"22",X"40",X"23",X"5E",X"20",X"5D",X"3E",X"5F",X"3E",X"40",X"21",X"5F",
		X"23",X"40",X"22",X"44",X"02",X"43",X"00",X"C0",X"1D",X"42",X"3D",X"43",X"3D",X"5F",X"3F",X"5E",
		X"22",X"41",X"22",X"40",X"22",X"5D",X"3E",X"5D",X"3E",X"40",X"3E",X"41",X"21",X"5E",X"23",X"5F",
		X"23",X"43",X"03",X"42",X"00",X"C0",X"1E",X"43",X"3E",X"44",X"3D",X"40",X"3F",X"5F",X"22",X"40",
		X"22",X"5F",X"20",X"5D",X"3D",X"5E",X"3E",X"40",X"3F",X"42",X"20",X"5E",X"23",X"5E",X"23",X"43",
		X"04",X"5F",X"00",X"C0",X"1F",X"44",X"20",X"44",X"3D",X"41",X"3E",X"5F",X"22",X"40",X"22",X"5E",
		X"3F",X"5D",X"3D",X"5F",X"3E",X"42",X"20",X"42",X"3F",X"5E",X"21",X"5D",X"24",X"40",X"04",X"5F",
		X"00",X"C0",X"1F",X"44",X"23",X"43",X"3E",X"43",X"3E",X"40",X"22",X"5F",X"20",X"5E",X"3E",X"5D",
		X"3D",X"40",X"3F",X"42",X"20",X"42",X"3F",X"5F",X"20",X"5D",X"24",X"5E",X"03",X"5E",X"00",X"C0",
		X"02",X"43",X"23",X"43",X"20",X"43",X"3E",X"41",X"21",X"5E",X"3F",X"5E",X"3D",X"5E",X"3D",X"42",
		X"3F",X"42",X"21",X"42",X"3E",X"5F",X"20",X"5D",X"23",X"5D",X"02",X"5D",X"00",X"C0",X"03",X"42",
		X"24",X"42",X"21",X"42",X"3F",X"42",X"20",X"5E",X"3E",X"5E",X"3D",X"40",X"3E",X"43",X"3F",X"42",
		X"22",X"41",X"3E",X"40",X"3F",X"5D",X"21",X"5D",X"01",X"5C",X"00",X"C0",X"04",X"41",X"24",X"40",
		X"22",X"42",X"3F",X"42",X"3F",X"5E",X"3E",X"5F",X"3D",X"41",X"3F",X"43",X"21",X"42",X"22",X"41",
		X"3E",X"41",X"3C",X"5E",X"20",X"5C",X"01",X"5C",X"00",X"C0",X"04",X"41",X"23",X"5D",X"23",X"41",
		X"20",X"42",X"3F",X"40",X"3E",X"5F",X"3D",X"42",X"20",X"43",X"22",X"42",X"22",X"40",X"3E",X"41",
		X"3E",X"5F",X"3E",X"5C",X"1E",X"5D",X"00",X"C0",X"03",X"5E",X"23",X"5D",X"23",X"40",X"21",X"42",
		X"3E",X"5F",X"3E",X"41",X"3E",X"43",X"22",X"43",X"22",X"41",X"22",X"5F",X"3F",X"42",X"3D",X"40",
		X"3D",X"5D",X"1D",X"5E",X"00",X"C0",X"02",X"5D",X"22",X"5C",X"22",X"5F",X"22",X"41",X"3E",X"40",
		X"3E",X"42",X"20",X"43",X"23",X"42",X"22",X"41",X"21",X"5E",X"20",X"42",X"3D",X"41",X"3D",X"5F",
		X"1C",X"5F",X"00",X"C0",X"1F",X"5C",X"20",X"5C",X"24",X"5E",X"22",X"41",X"3E",X"41",X"3F",X"42",
		X"21",X"43",X"23",X"41",X"22",X"5F",X"21",X"5E",X"21",X"42",X"3E",X"44",X"3C",X"40",X"1C",X"5F",
		X"00",X"C0",X"1F",X"5C",X"3F",X"5D",X"21",X"5D",X"22",X"40",X"3E",X"41",X"21",X"42",X"22",X"43",
		X"23",X"40",X"22",X"5E",X"20",X"5E",X"21",X"42",X"3F",X"42",X"3C",X"42",X"1D",X"42",X"00",X"C0",
		X"1E",X"5D",X"3D",X"5D",X"20",X"5D",X"22",X"5F",X"3F",X"42",X"21",X"42",X"23",X"42",X"23",X"5E",
		X"21",X"5E",X"3F",X"5E",X"22",X"41",X"20",X"43",X"3D",X"43",X"1E",X"43",X"00",X"C0",X"1D",X"5E",
		X"3C",X"5E",X"3F",X"5E",X"21",X"5E",X"20",X"42",X"22",X"42",X"23",X"40",X"22",X"5D",X"3F",X"5E",
		X"20",X"5F",X"22",X"40",X"21",X"43",X"3D",X"43",X"01",X"44",X"00",X"C0",X"1C",X"41",X"3C",X"40",
		X"3E",X"5C",X"21",X"5E",X"21",X"42",X"22",X"41",X"23",X"5F",X"21",X"5D",X"3F",X"5E",X"3E",X"5F",
		X"22",X"5F",X"22",X"42",X"20",X"44",X"01",X"44",X"00",X"C0",X"1C",X"41",X"3D",X"41",X"3D",X"5F",
		X"20",X"5E",X"21",X"42",X"22",X"5F",X"23",X"5E",X"20",X"5D",X"3E",X"5E",X"3E",X"40",X"22",X"5F",
		X"22",X"41",X"22",X"44",X"02",X"43",X"00",X"C0",X"1D",X"42",X"3D",X"43",X"3D",X"40",X"3F",X"5E",
		X"22",X"41",X"22",X"5F",X"22",X"5D",X"3E",X"5D",X"3E",X"5F",X"3E",X"41",X"21",X"5E",X"23",X"40",
		X"23",X"43",X"03",X"42",X"00",X"C0",X"1E",X"43",X"3E",X"44",X"3E",X"41",X"3E",X"5F",X"22",X"40",
		X"22",X"5E",X"20",X"5D",X"3D",X"5E",X"3E",X"41",X"3F",X"40",X"20",X"5E",X"23",X"5F",X"23",X"43",
		X"04",X"5F",X"00",X"C0",X"1F",X"44",X"20",X"44",X"3E",X"42",X"3E",X"5F",X"22",X"5F",X"21",X"5E",
		X"3F",X"5D",X"3D",X"5F",X"3E",X"41",X"3F",X"42",X"3F",X"5E",X"22",X"5E",X"24",X"40",X"04",X"5F",
		X"00",X"C0",X"1F",X"44",X"23",X"43",X"3F",X"43",X"3E",X"40",X"20",X"5F",X"21",X"5E",X"3E",X"5D",
		X"3D",X"40",X"3E",X"42",X"20",X"42",X"3F",X"5E",X"21",X"5E",X"24",X"5E",X"03",X"5E",X"00",X"C0",
		X"1E",X"43",X"3D",X"45",X"3F",X"44",X"02",X"54",X"3C",X"43",X"3C",X"5E",X"09",X"5C",X"3A",X"41",
		X"3D",X"5C",X"0C",X"40",X"0C",X"40",X"3D",X"44",X"3A",X"5F",X"01",X"43",X"24",X"43",X"24",X"5E",
		X"16",X"42",X"23",X"45",X"21",X"44",X"1A",X"54",X"00",X"C0",X"1F",X"44",X"3F",X"45",X"21",X"44",
		X"1D",X"55",X"3E",X"44",X"3B",X"40",X"07",X"58",X"3B",X"44",X"3C",X"5F",X"0B",X"59",X"0B",X"5C",
		X"3F",X"45",X"3A",X"41",X"02",X"42",X"25",X"42",X"22",X"5C",X"18",X"46",X"25",X"43",X"22",X"44",
		X"16",X"57",X"00",X"C0",X"1F",X"44",X"23",X"45",X"22",X"44",X"19",X"56",X"3F",X"45",X"3C",X"41",
		X"04",X"57",X"3C",X"45",X"3B",X"5F",X"09",X"58",X"08",X"57",X"21",X"45",X"3B",X"44",X"03",X"41",
		X"25",X"5F",X"21",X"5C",X"1B",X"49",X"25",X"41",X"24",X"42",X"13",X"5C",X"00",X"C0",X"02",X"43",
		X"23",X"45",X"24",X"42",X"15",X"5A",X"22",X"45",X"3C",X"42",X"00",X"57",X"3F",X"46",X"3B",X"41",
		X"04",X"55",X"05",X"55",X"23",X"44",X"3C",X"45",X"04",X"40",X"24",X"5E",X"20",X"5B",X"1E",X"4C",
		X"25",X"5D",X"24",X"43",X"13",X"5F",X"00",X"C0",X"03",X"42",X"25",X"43",X"24",X"41",X"14",X"5E",
		X"23",X"44",X"3C",X"44",X"1E",X"57",X"21",X"46",X"3C",X"43",X"00",X"54",X"00",X"54",X"24",X"43",
		X"3F",X"46",X"03",X"5F",X"23",X"5C",X"3E",X"5C",X"02",X"4A",X"25",X"5D",X"24",X"5F",X"14",X"46",
		X"00",X"C0",X"04",X"41",X"25",X"41",X"24",X"5F",X"15",X"43",X"24",X"42",X"20",X"45",X"18",X"59",
		X"24",X"45",X"3D",X"44",X"1B",X"55",X"1C",X"55",X"25",X"41",X"21",X"46",X"02",X"5E",X"22",X"5B",
		X"3C",X"5E",X"06",X"48",X"23",X"5B",X"24",X"5E",X"17",X"4A",X"00",X"C0",X"04",X"41",X"25",X"5D",
		X"24",X"5E",X"16",X"47",X"25",X"41",X"21",X"44",X"17",X"5C",X"25",X"44",X"3F",X"45",X"18",X"57",
		X"17",X"58",X"25",X"5F",X"24",X"45",X"01",X"5D",X"3F",X"5B",X"3C",X"5F",X"07",X"45",X"23",X"5B",
		X"22",X"5C",X"1C",X"4D",X"00",X"C0",X"03",X"5E",X"25",X"5D",X"22",X"5C",X"1A",X"4B",X"25",X"5E",
		X"22",X"44",X"17",X"40",X"26",X"41",X"21",X"45",X"15",X"5C",X"15",X"5B",X"24",X"5D",X"25",X"44",
		X"00",X"5C",X"3E",X"5C",X"3B",X"40",X"0A",X"42",X"3F",X"5B",X"21",X"5C",X"01",X"4D",X"00",X"C0",
		X"02",X"5D",X"23",X"5B",X"21",X"5C",X"1E",X"4C",X"24",X"5D",X"24",X"44",X"17",X"42",X"26",X"5F",
		X"23",X"44",X"14",X"40",X"14",X"40",X"23",X"5C",X"26",X"41",X"1F",X"5D",X"3C",X"5D",X"3C",X"42",
		X"0A",X"5E",X"3D",X"5B",X"3F",X"5C",X"06",X"4C",X"00",X"C0",X"1F",X"5C",X"23",X"5B",X"3D",X"5C",
		X"05",X"4B",X"22",X"5C",X"25",X"40",X"19",X"48",X"25",X"5C",X"24",X"43",X"15",X"45",X"15",X"44",
		X"21",X"5B",X"26",X"5F",X"1E",X"5E",X"3B",X"5E",X"3E",X"44",X"08",X"5A",X"3B",X"5D",X"3E",X"5C",
		X"0A",X"49",X"00",X"C0",X"1F",X"5C",X"3F",X"5B",X"3E",X"5C",X"07",X"4A",X"21",X"5B",X"24",X"5F",
		X"1C",X"49",X"24",X"5B",X"25",X"41",X"17",X"48",X"18",X"49",X"3F",X"5B",X"25",X"5C",X"1D",X"5F",
		X"3B",X"41",X"3F",X"44",X"05",X"59",X"3B",X"5D",X"3C",X"5E",X"0D",X"44",X"00",X"C0",X"1E",X"5D",
		X"3D",X"5B",X"3C",X"5E",X"0B",X"46",X"3E",X"5B",X"24",X"5E",X"00",X"49",X"21",X"5A",X"25",X"5F",
		X"1C",X"4B",X"19",X"4B",X"3F",X"5C",X"24",X"5B",X"1C",X"40",X"3C",X"42",X"20",X"45",X"02",X"56",
		X"3B",X"41",X"3C",X"5F",X"0D",X"5F",X"00",X"C0",X"1D",X"5E",X"3B",X"5D",X"3C",X"5F",X"0C",X"42",
		X"3D",X"5C",X"22",X"5C",X"04",X"49",X"3F",X"5A",X"24",X"5D",X"00",X"4C",X"00",X"4C",X"3C",X"5D",
		X"21",X"5A",X"1D",X"41",X"3D",X"44",X"22",X"44",X"1E",X"56",X"3B",X"43",X"3C",X"41",X"0C",X"5A",
		X"00",X"C0",X"1C",X"41",X"3B",X"5D",X"3C",X"43",X"0B",X"5B",X"3C",X"5E",X"20",X"5B",X"08",X"47",
		X"3C",X"5B",X"21",X"5C",X"07",X"4B",X"04",X"4B",X"3B",X"5F",X"3F",X"5A",X"1E",X"42",X"3E",X"45",
		X"24",X"42",X"1A",X"58",X"3D",X"45",X"3C",X"42",X"09",X"56",X"00",X"C0",X"1C",X"41",X"3B",X"41",
		X"3C",X"42",X"0A",X"59",X"3B",X"5F",X"3F",X"5C",X"09",X"44",X"3B",X"5C",X"21",X"5B",X"08",X"49",
		X"09",X"48",X"3B",X"41",X"3C",X"5B",X"1F",X"43",X"21",X"45",X"24",X"41",X"17",X"5B",X"3F",X"45",
		X"3E",X"44",X"04",X"53",X"00",X"C0",X"1D",X"42",X"3B",X"43",X"3E",X"44",X"06",X"55",X"3B",X"42",
		X"3E",X"5C",X"09",X"40",X"3A",X"5F",X"3F",X"5B",X"0B",X"44",X"0B",X"47",X"3C",X"41",X"3B",X"5C",
		X"00",X"44",X"22",X"44",X"25",X"40",X"14",X"5E",X"23",X"45",X"3D",X"44",X"01",X"53",X"00",X"C0",
		X"1E",X"43",X"3B",X"43",X"3E",X"44",X"05",X"56",X"3B",X"5F",X"3E",X"5C",X"08",X"42",X"3B",X"5D",
		X"3E",X"5B",X"0A",X"40",X"0A",X"40",X"3E",X"45",X"3B",X"43",X"08",X"5E",X"3E",X"44",X"3B",X"41",
		X"1E",X"43",X"25",X"43",X"22",X"44",X"17",X"56",X"00",X"C0",X"1F",X"44",X"3D",X"44",X"20",X"45",
		X"00",X"55",X"3B",X"41",X"3D",X"5D",X"08",X"5E",X"3A",X"40",X"3D",X"5C",X"09",X"5C",X"09",X"5C",
		X"20",X"45",X"3D",X"45",X"06",X"5B",X"20",X"45",X"3C",X"42",X"1F",X"44",X"26",X"41",X"23",X"43",
		X"14",X"5A",X"00",X"C0",X"1F",X"44",X"20",X"45",X"20",X"44",X"1E",X"56",X"3C",X"43",X"3C",X"5E",
		X"07",X"5C",X"3A",X"41",X"3B",X"40",X"07",X"57",X"07",X"59",X"22",X"45",X"3F",X"46",X"04",X"59",
		X"22",X"44",X"3D",X"44",X"01",X"44",X"25",X"40",X"24",X"40",X"13",X"5F",X"00",X"C0",X"02",X"43",
		X"21",X"46",X"23",X"43",X"18",X"58",X"3E",X"44",X"3B",X"40",X"05",X"5A",X"3B",X"43",X"3B",X"40",
		X"04",X"57",X"04",X"57",X"24",X"43",X"20",X"46",X"02",X"58",X"23",X"43",X"3F",X"45",X"02",X"45",
		X"24",X"5B",X"25",X"40",X"13",X"44",X"00",X"C0",X"03",X"42",X"23",X"45",X"24",X"42",X"16",X"5B",
		X"3F",X"45",X"3C",X"42",X"02",X"58",X"3D",X"45",X"3B",X"42",X"00",X"56",X"00",X"56",X"25",X"42",
		X"23",X"45",X"1E",X"58",X"24",X"42",X"21",X"45",X"03",X"42",X"23",X"5B",X"24",X"5E",X"16",X"49",
		X"00",X"C0",X"04",X"41",X"24",X"43",X"25",X"40",X"15",X"40",X"21",X"45",X"3D",X"43",X"1E",X"58",
		X"20",X"46",X"3C",X"43",X"1C",X"57",X"1C",X"57",X"25",X"40",X"25",X"43",X"1B",X"5A",X"25",X"40",
		X"22",X"44",X"04",X"41",X"21",X"5A",X"23",X"5D",X"1A",X"4C",X"00",X"C0",X"04",X"41",X"25",X"40",
		X"24",X"40",X"16",X"42",X"23",X"44",X"3E",X"44",X"1C",X"59",X"21",X"46",X"3E",X"45",X"19",X"59",
		X"19",X"59",X"25",X"5E",X"26",X"41",X"19",X"5C",X"24",X"5E",X"24",X"43",X"02",X"5F",X"20",X"5B",
		X"20",X"5C",X"01",X"4D",X"00",X"C0",X"03",X"5E",X"26",X"5F",X"23",X"5D",X"18",X"48",X"24",X"42",
		X"20",X"45",X"1A",X"5B",X"23",X"45",X"20",X"45",X"17",X"5C",X"17",X"5C",X"23",X"5C",X"26",X"40",
		X"18",X"5E",X"23",X"5D",X"25",X"41",X"03",X"5E",X"3D",X"5C",X"20",X"5B",X"04",X"4D",X"00",X"C0",
		X"02",X"5D",X"25",X"5D",X"22",X"5C",X"1B",X"4A",X"25",X"41",X"22",X"44",X"18",X"5E",X"25",X"43",
		X"22",X"45",X"16",X"40",X"16",X"40",X"22",X"5B",X"25",X"5D",X"18",X"42",X"22",X"5C",X"25",X"5F",
		X"02",X"5D",X"3B",X"5D",X"3E",X"5C",X"09",X"4A",X"00",X"C0",X"1F",X"5C",X"25",X"5C",X"20",X"5B",
		X"00",X"4B",X"25",X"5F",X"23",X"43",X"18",X"42",X"26",X"40",X"23",X"44",X"17",X"44",X"17",X"44",
		X"20",X"5B",X"23",X"5B",X"1A",X"45",X"20",X"5B",X"24",X"5E",X"01",X"5C",X"3A",X"5F",X"3D",X"5D",
		X"0C",X"46",X"00",X"C0",X"1F",X"5C",X"20",X"5B",X"20",X"5C",X"04",X"4A",X"24",X"5D",X"24",X"42",
		X"19",X"44",X"26",X"5F",X"25",X"42",X"19",X"47",X"17",X"47",X"20",X"5B",X"21",X"5A",X"1C",X"47",
		X"3E",X"5C",X"23",X"5C",X"1F",X"5E",X"3B",X"40",X"3C",X"40",X"0D",X"5F",X"00",X"C0",X"1E",X"5D",
		X"3F",X"5A",X"3D",X"5D",X"08",X"48",X"22",X"5C",X"25",X"40",X"1B",X"46",X"25",X"5D",X"25",X"40",
		X"1C",X"49",X"1C",X"49",X"3C",X"5D",X"20",X"5A",X"1E",X"48",X"3D",X"5D",X"21",X"5B",X"1E",X"5D",
		X"3C",X"43",X"3B",X"40",X"0D",X"5C",X"00",X"C0",X"1D",X"5E",X"3D",X"5B",X"3C",X"5E",X"0A",X"45",
		X"3F",X"5B",X"26",X"5E",X"1E",X"48",X"23",X"5B",X"25",X"5E",X"00",X"4A",X"00",X"4A",X"3B",X"5E",
		X"3D",X"5B",X"02",X"48",X"3C",X"5E",X"3F",X"5B",X"1D",X"5E",X"3D",X"45",X"3C",X"42",X"0A",X"57",
		X"00",X"C0",X"1C",X"41",X"3C",X"5B",X"3B",X"40",X"0B",X"40",X"3F",X"5B",X"23",X"5D",X"02",X"48",
		X"20",X"5A",X"24",X"5D",X"04",X"49",X"04",X"49",X"3B",X"40",X"3B",X"5D",X"05",X"46",X"3B",X"40",
		X"3E",X"5C",X"1C",X"5F",X"3F",X"46",X"3D",X"43",X"06",X"54",X"00",X"C0",X"1C",X"41",X"3B",X"40",
		X"3C",X"40",X"0A",X"5C",X"3D",X"5C",X"22",X"5C",X"04",X"47",X"3F",X"5A",X"20",X"5B",X"09",X"47",
		X"07",X"49",X"3B",X"40",X"3A",X"5F",X"07",X"44",X"3C",X"42",X"3C",X"5D",X"1C",X"41",X"20",X"45",
		X"20",X"44",X"01",X"53",X"00",X"C0",X"1D",X"42",X"3A",X"41",X"3D",X"43",X"08",X"58",X"3C",X"5E",
		X"20",X"5B",X"06",X"45",X"3D",X"5B",X"20",X"5B",X"09",X"44",X"09",X"44",X"3D",X"44",X"3A",X"40",
		X"08",X"42",X"3D",X"43",X"3B",X"5F",X"1B",X"42",X"25",X"44",X"20",X"45",X"1C",X"53",X"00",X"C0",
		X"1E",X"43",X"3A",X"41",X"3E",X"44",X"06",X"58",X"3C",X"5D",X"3E",X"5C",X"07",X"44",X"3C",X"5C",
		X"3F",X"5B",X"08",X"40",X"08",X"40",X"3F",X"45",X"3C",X"44",X"07",X"5C",X"3E",X"44",X"3C",X"43",
		X"1E",X"43",X"26",X"41",X"22",X"44",X"16",X"58",X"00",X"C0",X"1F",X"44",X"3B",X"43",X"20",X"44",
		X"02",X"57",X"3B",X"5E",X"3D",X"5D",X"08",X"41",X"3B",X"5E",X"3D",X"5C",X"07",X"5D",X"08",X"5D",
		X"21",X"45",X"3E",X"45",X"05",X"5A",X"3F",X"44",X"3E",X"44",X"1F",X"44",X"26",X"5F",X"23",X"43",
		X"14",X"5C",X"00",X"C0",X"1F",X"44",X"3E",X"44",X"22",X"45",X"1E",X"56",X"3B",X"41",X"3C",X"5E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
