library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"32",X"01",X"70",X"C3",X"82",X"01",X"84",X"AF",X"21",X"06",X"70",X"77",X"23",X"77",X"C9",
		X"F5",X"C5",X"D5",X"E5",X"5E",X"23",X"56",X"23",X"E5",X"C1",X"EB",X"11",X"20",X"00",X"0A",X"FE",
		X"FF",X"28",X"07",X"D6",X"30",X"77",X"03",X"19",X"18",X"F4",X"E1",X"D1",X"C1",X"F1",X"C9",X"67",
		X"21",X"07",X"42",X"06",X"1B",X"71",X"23",X"23",X"10",X"FB",X"3A",X"00",X"78",X"21",X"00",X"42",
		X"11",X"40",X"42",X"06",X"20",X"AF",X"77",X"12",X"13",X"23",X"23",X"10",X"F9",X"06",X"20",X"12",
		X"13",X"10",X"FC",X"C9",X"DB",X"28",X"0C",X"D9",X"CD",X"12",X"DA",X"D9",X"28",X"0A",X"CD",X"3A",
		X"84",X"18",X"DF",X"CD",X"35",X"84",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"01",X"70",X"3A",X"00",X"78",X"21",X"00",X"42",X"01",X"60",X"00",X"11",X"00",X"58",X"ED",X"B0",
		X"21",X"BB",X"42",X"34",X"21",X"84",X"42",X"CD",X"E2",X"00",X"CD",X"2F",X"31",X"21",X"60",X"42",
		X"01",X"20",X"00",X"11",X"60",X"58",X"ED",X"B0",X"CD",X"1F",X"34",X"3A",X"CE",X"42",X"B7",X"C4",
		X"F4",X"00",X"CD",X"0B",X"01",X"CD",X"67",X"01",X"CD",X"8A",X"36",X"21",X"02",X"70",X"3E",X"FF",
		X"77",X"00",X"00",X"C3",X"97",X"20",X"AF",X"21",X"02",X"70",X"77",X"7A",X"B7",X"28",X"0E",X"31",
		X"00",X"48",X"21",X"22",X"04",X"E5",X"3E",X"01",X"32",X"01",X"70",X"ED",X"45",X"FD",X"E1",X"DD",
		X"E1",X"E1",X"D1",X"C1",X"3E",X"01",X"32",X"01",X"70",X"F1",X"ED",X"45",X"3A",X"00",X"60",X"CB",
		X"47",X"C9",X"34",X"7E",X"FE",X"3C",X"C0",X"36",X"00",X"23",X"34",X"C9",X"3A",X"86",X"42",X"E6",
		X"03",X"FE",X"03",X"C9",X"3A",X"BB",X"42",X"CB",X"5F",X"20",X"08",X"FD",X"66",X"0B",X"FD",X"6E",
		X"0A",X"D7",X"C9",X"FD",X"66",X"0D",X"FD",X"6E",X"0C",X"D7",X"C9",X"3A",X"84",X"42",X"B7",X"C0",
		X"3A",X"BD",X"42",X"CB",X"47",X"28",X"0D",X"21",X"BC",X"42",X"35",X"20",X"07",X"21",X"8F",X"42",
		X"CB",X"9E",X"CB",X"87",X"CB",X"4F",X"28",X"08",X"21",X"A5",X"42",X"35",X"20",X"02",X"CB",X"8F",
		X"CB",X"57",X"28",X"08",X"21",X"A4",X"42",X"35",X"20",X"02",X"CB",X"97",X"CB",X"5F",X"28",X"23",
		X"21",X"A6",X"42",X"35",X"20",X"1D",X"4F",X"21",X"9E",X"42",X"CB",X"3E",X"7E",X"CB",X"3E",X"86",
		X"77",X"21",X"9F",X"42",X"CB",X"3E",X"7E",X"CB",X"3E",X"86",X"77",X"21",X"CA",X"42",X"CB",X"D6",
		X"79",X"CB",X"9F",X"32",X"BD",X"42",X"C9",X"3A",X"8B",X"42",X"B7",X"C8",X"21",X"CA",X"42",X"CB",
		X"46",X"C0",X"21",X"CC",X"42",X"CB",X"46",X"C0",X"21",X"CA",X"42",X"CB",X"C6",X"21",X"8B",X"42",
		X"35",X"C9",X"31",X"00",X"48",X"CD",X"97",X"37",X"21",X"00",X"40",X"36",X"00",X"3A",X"00",X"78",
		X"23",X"7C",X"FE",X"71",X"20",X"F5",X"32",X"00",X"78",X"32",X"1F",X"49",X"3A",X"AB",X"C0",X"FE",
		X"CF",X"00",X"00",X"00",X"21",X"00",X"50",X"06",X"10",X"0E",X"54",X"CD",X"FD",X"04",X"21",X"03",
		X"42",X"3E",X"07",X"77",X"23",X"23",X"77",X"21",X"07",X"05",X"D7",X"21",X"21",X"05",X"D7",X"21",
		X"3D",X"42",X"3E",X"05",X"77",X"23",X"23",X"77",X"21",X"52",X"05",X"D7",X"3A",X"00",X"78",X"21",
		X"D2",X"05",X"01",X"07",X"00",X"11",X"87",X"40",X"ED",X"B0",X"21",X"DA",X"05",X"01",X"07",X"00",
		X"11",X"87",X"41",X"ED",X"B0",X"3A",X"00",X"78",X"21",X"35",X"38",X"01",X"E0",X"00",X"11",X"D2",
		X"42",X"ED",X"B0",X"CD",X"DF",X"0C",X"3A",X"00",X"70",X"47",X"3A",X"00",X"68",X"17",X"CB",X"10",
		X"17",X"CB",X"10",X"78",X"32",X"86",X"42",X"21",X"86",X"42",X"ED",X"6F",X"47",X"ED",X"67",X"78",
		X"E6",X"03",X"3C",X"32",X"87",X"42",X"3A",X"86",X"42",X"CB",X"5F",X"28",X"05",X"21",X"87",X"41",
		X"36",X"00",X"3E",X"EA",X"32",X"A7",X"42",X"3E",X"01",X"32",X"01",X"70",X"CD",X"EC",X"00",X"CA",
		X"22",X"04",X"31",X"00",X"48",X"CF",X"0E",X"1B",X"CD",X"DC",X"04",X"0E",X"01",X"F7",X"CD",X"D7",
		X"0B",X"21",X"88",X"0B",X"D7",X"21",X"C4",X"05",X"D7",X"06",X"05",X"CD",X"C8",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"20",X"00",X"21",
		X"46",X"50",X"06",X"1C",X"C5",X"E5",X"06",X"08",X"36",X"50",X"23",X"10",X"FB",X"E1",X"19",X"C1",
		X"10",X"F2",X"21",X"68",X"53",X"11",X"C2",X"03",X"06",X"18",X"C5",X"E5",X"06",X"04",X"1A",X"77",
		X"23",X"13",X"10",X"FA",X"E1",X"01",X"20",X"00",X"A7",X"ED",X"42",X"C1",X"10",X"EC",X"06",X"03",
		X"CD",X"C8",X"0C",X"21",X"E4",X"53",X"22",X"91",X"42",X"21",X"8E",X"42",X"36",X"00",X"21",X"5C",
		X"42",X"36",X"00",X"23",X"36",X"3A",X"23",X"36",X"05",X"23",X"36",X"20",X"3E",X"11",X"CD",X"97",
		X"03",X"CD",X"F3",X"22",X"CD",X"A9",X"07",X"06",X"28",X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",
		X"47",X"20",X"EE",X"3E",X"43",X"CD",X"97",X"03",X"CD",X"A8",X"22",X"CD",X"A9",X"07",X"06",X"28",
		X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",X"47",X"20",X"EE",X"3A",X"5F",X"42",X"FE",X"60",X"20",
		X"E2",X"3E",X"13",X"CD",X"97",X"03",X"CD",X"F3",X"22",X"CD",X"A9",X"07",X"06",X"28",X"CD",X"C0",
		X"0C",X"3A",X"8F",X"42",X"CB",X"47",X"20",X"EE",X"3A",X"5C",X"42",X"DD",X"21",X"08",X"53",X"FE",
		X"40",X"CC",X"A1",X"03",X"DD",X"21",X"88",X"52",X"FE",X"60",X"CC",X"A1",X"03",X"DD",X"21",X"08",
		X"52",X"FE",X"80",X"CC",X"A1",X"03",X"DD",X"21",X"88",X"51",X"FE",X"A0",X"CC",X"A1",X"03",X"DD",
		X"21",X"08",X"51",X"FE",X"C0",X"CC",X"A1",X"03",X"DD",X"21",X"88",X"50",X"FE",X"E0",X"CC",X"A1",
		X"03",X"FE",X"E0",X"20",X"AC",X"3E",X"83",X"CD",X"97",X"03",X"CD",X"5D",X"22",X"CD",X"A9",X"07",
		X"06",X"28",X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",X"47",X"20",X"EE",X"3A",X"5F",X"42",X"FE",
		X"30",X"20",X"E2",X"3E",X"87",X"CD",X"97",X"03",X"CD",X"5D",X"22",X"CD",X"A9",X"07",X"06",X"28",
		X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",X"47",X"20",X"EE",X"3E",X"11",X"CD",X"97",X"03",X"CD",
		X"F3",X"22",X"CD",X"A9",X"07",X"06",X"28",X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",X"47",X"20",
		X"EE",X"06",X"08",X"CD",X"C8",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C3",X"32",X"02",X"21",X"8F",X"42",X"77",X"3E",X"08",X"32",X"9B",X"42",
		X"C9",X"F5",X"06",X"06",X"DD",X"7E",X"03",X"DD",X"77",X"05",X"DD",X"7E",X"23",X"DD",X"77",X"25",
		X"DD",X"7E",X"43",X"DD",X"77",X"45",X"DD",X"7E",X"63",X"DD",X"77",X"65",X"DD",X"2B",X"10",X"E4",
		X"F1",X"C9",X"F2",X"F7",X"F7",X"F3",X"F4",X"E6",X"E7",X"F5",X"F4",X"E4",X"E5",X"F5",X"F0",X"F6",
		X"F6",X"F1",X"F2",X"F7",X"F7",X"F3",X"F4",X"E2",X"E3",X"F5",X"F4",X"E0",X"E1",X"F5",X"F0",X"F6",
		X"F6",X"F1",X"F2",X"F7",X"F7",X"F3",X"F4",X"EA",X"EB",X"F5",X"F4",X"E8",X"E9",X"F5",X"F0",X"F6",
		X"F6",X"F1",X"F2",X"F7",X"F7",X"F3",X"F4",X"E6",X"E7",X"F5",X"F4",X"E4",X"E5",X"F5",X"F0",X"F6",
		X"F6",X"F1",X"F2",X"F7",X"F7",X"F3",X"F4",X"EE",X"EF",X"F5",X"F4",X"EC",X"ED",X"F5",X"F0",X"F6",
		X"F6",X"F1",X"F2",X"F7",X"F7",X"F3",X"F4",X"EA",X"EB",X"F5",X"F4",X"E8",X"E9",X"F5",X"F0",X"F6",
		X"F6",X"F1",X"31",X"00",X"48",X"CF",X"0E",X"1B",X"CD",X"DC",X"04",X"0E",X"02",X"F7",X"21",X"5A",
		X"05",X"D7",X"21",X"90",X"05",X"D7",X"21",X"AA",X"05",X"D7",X"21",X"C4",X"05",X"D7",X"21",X"95",
		X"51",X"3A",X"87",X"42",X"77",X"CD",X"EC",X"00",X"28",X"3C",X"21",X"3A",X"05",X"D7",X"3A",X"88",
		X"42",X"FE",X"02",X"38",X"05",X"21",X"7F",X"05",X"18",X"03",X"21",X"6E",X"05",X"D7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"88",X"42",X"47",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"BE",X"52",X"78",X"E6",X"0F",X"32",X"9E",
		X"52",X"CD",X"93",X"04",X"18",X"C8",X"21",X"46",X"05",X"D7",X"21",X"7F",X"05",X"D7",X"CD",X"93",
		X"04",X"18",X"FB",X"21",X"00",X"68",X"CB",X"46",X"20",X"1F",X"CB",X"4E",X"20",X"01",X"C9",X"CD",
		X"EC",X"00",X"28",X"06",X"3A",X"88",X"42",X"FE",X"02",X"D8",X"21",X"E8",X"05",X"D7",X"21",X"03",
		X"06",X"D7",X"3E",X"02",X"32",X"8D",X"42",X"18",X"0D",X"21",X"F4",X"05",X"D7",X"21",X"15",X"06",
		X"D7",X"3E",X"01",X"32",X"8D",X"42",X"21",X"FA",X"05",X"D7",X"47",X"CD",X"EC",X"00",X"CA",X"A5",
		X"08",X"3A",X"88",X"42",X"90",X"27",X"32",X"88",X"42",X"C3",X"A5",X"08",X"E5",X"C5",X"21",X"00",
		X"50",X"23",X"23",X"23",X"41",X"3E",X"10",X"77",X"23",X"10",X"FC",X"3A",X"00",X"78",X"79",X"FE",
		X"1D",X"28",X"02",X"23",X"23",X"7C",X"FE",X"54",X"20",X"E7",X"C1",X"E1",X"C9",X"70",X"3A",X"00",
		X"78",X"23",X"7C",X"B9",X"20",X"F7",X"C9",X"81",X"50",X"50",X"55",X"32",X"40",X"40",X"40",X"40",
		X"45",X"52",X"4F",X"43",X"53",X"40",X"48",X"47",X"49",X"48",X"40",X"40",X"40",X"50",X"55",X"31",
		X"FF",X"62",X"50",X"30",X"30",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"30",X"30",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"30",X"30",X"FF",X"9E",X"52",X"40",X"40",X"40",X"54",
		X"49",X"44",X"45",X"52",X"43",X"FF",X"9E",X"52",X"59",X"41",X"4C",X"50",X"40",X"45",X"45",X"52",
		X"46",X"FF",X"DE",X"50",X"44",X"4E",X"55",X"4F",X"52",X"FF",X"0E",X"51",X"4E",X"4F",X"54",X"54",
		X"55",X"42",X"40",X"54",X"52",X"41",X"54",X"53",X"40",X"48",X"53",X"55",X"50",X"FF",X"31",X"51",
		X"40",X"59",X"4C",X"4E",X"4F",X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",X"31",X"FF",X"31",
		X"51",X"53",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",X"32",X"40",X"52",X"4F",X"40",X"31",X"FF",
		X"95",X"50",X"53",X"54",X"50",X"40",X"30",X"30",X"30",X"30",X"40",X"40",X"52",X"4F",X"46",X"40",
		X"53",X"55",X"4E",X"4F",X"42",X"40",X"54",X"53",X"31",X"FF",X"97",X"50",X"53",X"54",X"50",X"40",
		X"30",X"30",X"30",X"30",X"36",X"40",X"52",X"4F",X"46",X"40",X"53",X"55",X"4E",X"4F",X"42",X"40",
		X"44",X"4E",X"32",X"FF",X"1B",X"51",X"32",X"38",X"39",X"31",X"40",X"40",X"58",X"41",X"4C",X"40",
		X"B0",X"FF",X"00",X"82",X"53",X"E2",X"05",X"EE",X"05",X"00",X"01",X"02",X"51",X"E8",X"05",X"F4",
		X"05",X"00",X"01",X"53",X"50",X"55",X"31",X"FF",X"81",X"50",X"50",X"55",X"32",X"FF",X"01",X"53",
		X"40",X"40",X"40",X"FF",X"81",X"50",X"40",X"40",X"40",X"FF",X"E2",X"52",X"30",X"30",X"40",X"40",
		X"40",X"40",X"FF",X"62",X"50",X"30",X"30",X"40",X"40",X"40",X"40",X"FF",X"E2",X"52",X"40",X"40",
		X"40",X"40",X"40",X"40",X"FF",X"62",X"50",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"FD",X"7E",
		X"03",X"F5",X"0E",X"00",X"11",X"20",X"00",X"21",X"9E",X"50",X"CD",X"89",X"07",X"F1",X"11",X"40",
		X"00",X"4F",X"A7",X"28",X"3B",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"47",X"79",X"E6",X"0F",X"FE",
		X"05",X"F5",X"38",X"02",X"D6",X"05",X"4F",X"DD",X"21",X"44",X"50",X"78",X"A7",X"28",X"09",X"3E",
		X"BC",X"CD",X"AF",X"06",X"DD",X"19",X"10",X"F7",X"F1",X"38",X"07",X"3E",X"B8",X"CD",X"AF",X"06",
		X"DD",X"19",X"79",X"41",X"A7",X"28",X"09",X"3E",X"B4",X"CD",X"AF",X"06",X"DD",X"19",X"10",X"F7",
		X"DD",X"E5",X"E1",X"7C",X"FE",X"54",X"D0",X"3E",X"10",X"CD",X"BF",X"06",X"DD",X"19",X"18",X"F0",
		X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"7E",X"05",X"11",X"C0",X"FF",X"DD",X"21",X"9E",X"53",X"0E",
		X"09",X"47",X"A7",X"28",X"0A",X"3E",X"F8",X"CD",X"AF",X"06",X"DD",X"19",X"0D",X"10",X"F6",X"3E",
		X"10",X"CD",X"BF",X"06",X"DD",X"19",X"0D",X"20",X"F6",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"DD",
		X"77",X"00",X"3C",X"DD",X"77",X"01",X"3C",X"DD",X"77",X"20",X"3C",X"DD",X"77",X"21",X"C9",X"DD",
		X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"20",X"DD",X"77",X"21",X"C9",X"F5",X"C5",X"D5",X"E5",
		X"DD",X"E5",X"FD",X"E5",X"E1",X"7A",X"86",X"27",X"77",X"79",X"23",X"8E",X"27",X"77",X"78",X"23",
		X"8E",X"27",X"77",X"47",X"FD",X"7E",X"04",X"E6",X"03",X"FE",X"03",X"28",X"3C",X"4F",X"78",X"FE",
		X"06",X"38",X"1C",X"FD",X"CB",X"04",X"CE",X"FD",X"34",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"21",X"CA",X"42",X"CB",X"CE",X"E1",X"CB",
		X"41",X"20",X"16",X"3A",X"87",X"42",X"4F",X"78",X"B9",X"38",X"0E",X"FD",X"CB",X"04",X"C6",X"FD",
		X"34",X"05",X"E5",X"21",X"CA",X"42",X"CB",X"CE",X"E1",X"CD",X"80",X"06",X"DD",X"21",X"80",X"42",
		X"11",X"82",X"42",X"EB",X"CD",X"3F",X"07",X"CD",X"3F",X"07",X"CD",X"3F",X"07",X"18",X"1B",X"46",
		X"1A",X"B8",X"1B",X"2B",X"C8",X"C1",X"38",X"12",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"FD",X"7E",
		X"01",X"DD",X"77",X"01",X"FD",X"7E",X"02",X"DD",X"77",X"02",X"21",X"42",X"52",X"CD",X"74",X"07",
		X"FD",X"E5",X"DD",X"E1",X"FD",X"66",X"09",X"FD",X"6E",X"08",X"CD",X"74",X"07",X"DD",X"E1",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"C5",X"D5",X"11",X"20",X"00",X"01",X"00",X"03",X"DD",X"7E",X"02",X"CD",
		X"89",X"07",X"DD",X"2B",X"10",X"F6",X"D1",X"C1",X"C9",X"F5",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CD",X"98",X"07",X"F1",X"E6",X"0F",X"20",X"08",X"CB",X"41",X"20",X"04",X"3E",X"10",
		X"18",X"02",X"CB",X"C1",X"77",X"A7",X"ED",X"52",X"C9",X"21",X"8E",X"42",X"7E",X"E6",X"C3",X"20",
		X"2F",X"3A",X"9B",X"42",X"E6",X"01",X"47",X"CD",X"DE",X"33",X"4F",X"28",X"11",X"3E",X"36",X"CB",
		X"59",X"20",X"02",X"3E",X"3A",X"80",X"CB",X"61",X"20",X"13",X"CB",X"FF",X"18",X"0F",X"3E",X"34",
		X"CB",X"59",X"20",X"02",X"3E",X"38",X"80",X"CB",X"79",X"20",X"02",X"F6",X"C0",X"32",X"5D",X"42",
		X"CD",X"10",X"2B",X"CD",X"1F",X"2B",X"D8",X"79",X"E6",X"0B",X"20",X"F7",X"CB",X"51",X"20",X"3A",
		X"CB",X"58",X"28",X"0F",X"CB",X"48",X"28",X"04",X"3E",X"19",X"18",X"02",X"3E",X"19",X"CD",X"44",
		X"08",X"18",X"24",X"CB",X"48",X"28",X"04",X"3E",X"15",X"18",X"02",X"3E",X"17",X"CD",X"44",X"08",
		X"57",X"78",X"E6",X"30",X"28",X"09",X"7A",X"CB",X"60",X"20",X"0C",X"CB",X"FF",X"18",X"08",X"23",
		X"7E",X"E6",X"C0",X"B2",X"77",X"18",X"BC",X"23",X"18",X"FA",X"DD",X"7E",X"08",X"E5",X"CB",X"48",
		X"28",X"05",X"21",X"4B",X"08",X"18",X"03",X"21",X"50",X"08",X"3D",X"28",X"03",X"23",X"18",X"FA",
		X"7E",X"E1",X"18",X"CC",X"DD",X"CB",X"03",X"56",X"C8",X"3C",X"C9",X"15",X"0D",X"0E",X"0F",X"10",
		X"17",X"11",X"12",X"13",X"14",X"3A",X"8E",X"42",X"CB",X"47",X"C0",X"CB",X"77",X"C8",X"3A",X"AB",
		X"42",X"B7",X"C0",X"21",X"9D",X"42",X"7E",X"B7",X"CC",X"93",X"08",X"35",X"C0",X"36",X"C0",X"21",
		X"9B",X"42",X"35",X"46",X"20",X"0B",X"21",X"8E",X"42",X"CB",X"C6",X"3E",X"00",X"32",X"5D",X"42",
		X"C9",X"21",X"8F",X"08",X"05",X"28",X"03",X"23",X"18",X"FA",X"7E",X"32",X"5D",X"42",X"C9",X"3F",
		X"3E",X"3D",X"3C",X"E5",X"21",X"40",X"42",X"06",X"18",X"AF",X"77",X"23",X"10",X"FC",X"21",X"CB",
		X"42",X"CB",X"DE",X"E1",X"C9",X"31",X"00",X"48",X"08",X"3E",X"60",X"08",X"0E",X"1B",X"CD",X"DC",
		X"04",X"0E",X"07",X"F7",X"CD",X"D7",X"0B",X"FD",X"21",X"80",X"40",X"CD",X"0B",X"0C",X"3A",X"8D",
		X"42",X"FE",X"01",X"28",X"07",X"FD",X"21",X"80",X"41",X"CD",X"0B",X"0C",X"FD",X"21",X"80",X"40",
		X"31",X"00",X"48",X"FD",X"7E",X"07",X"CD",X"09",X"00",X"CD",X"DF",X"0C",X"CD",X"97",X"0B",X"CD",
		X"1E",X"06",X"CD",X"80",X"06",X"CD",X"81",X"0D",X"CD",X"F0",X"0C",X"FD",X"CB",X"04",X"76",X"C2",
		X"8F",X"09",X"FD",X"CB",X"04",X"F6",X"06",X"03",X"CD",X"C8",X"0C",X"FD",X"35",X"05",X"CD",X"80",
		X"06",X"21",X"CB",X"42",X"CB",X"F6",X"21",X"E4",X"53",X"22",X"91",X"42",X"21",X"8E",X"42",X"36",
		X"00",X"21",X"5C",X"42",X"36",X"00",X"23",X"36",X"3A",X"23",X"36",X"05",X"23",X"36",X"20",X"21",
		X"8F",X"42",X"36",X"11",X"3E",X"01",X"32",X"9D",X"42",X"3E",X"08",X"32",X"9B",X"42",X"CD",X"F3",
		X"22",X"CD",X"A9",X"07",X"06",X"1C",X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",X"47",X"20",X"EE",
		X"3A",X"5C",X"42",X"FE",X"70",X"20",X"D8",X"21",X"8F",X"42",X"36",X"43",X"3E",X"08",X"32",X"9B",
		X"42",X"CD",X"A8",X"22",X"CD",X"A9",X"07",X"06",X"1C",X"CD",X"C0",X"0C",X"3A",X"8F",X"42",X"CB",
		X"47",X"20",X"EE",X"3A",X"5F",X"42",X"FE",X"80",X"20",X"DD",X"21",X"8F",X"42",X"36",X"47",X"3E",
		X"08",X"32",X"9B",X"42",X"CD",X"A8",X"22",X"CD",X"A9",X"07",X"06",X"1C",X"CD",X"C0",X"0C",X"3A",
		X"8F",X"42",X"CB",X"47",X"20",X"EE",X"3A",X"CD",X"42",X"CB",X"77",X"20",X"F9",X"18",X"0B",X"06",
		X"02",X"CD",X"C8",X"0C",X"FD",X"35",X"05",X"CD",X"80",X"06",X"CD",X"2B",X"0C",X"CD",X"DF",X"0C",
		X"21",X"5C",X"42",X"36",X"70",X"23",X"36",X"3A",X"23",X"36",X"05",X"23",X"36",X"90",X"06",X"01",
		X"CD",X"C8",X"0C",X"21",X"00",X"19",X"22",X"7C",X"43",X"3E",X"46",X"32",X"7F",X"43",X"3E",X"03",
		X"32",X"B7",X"42",X"3E",X"08",X"32",X"B9",X"42",X"08",X"32",X"BA",X"42",X"08",X"3E",X"02",X"32",
		X"B8",X"42",X"32",X"CE",X"42",X"32",X"BE",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"32",X"AB",X"42",X"32",X"BF",X"42",
		X"3E",X"0E",X"32",X"BD",X"42",X"21",X"CB",X"42",X"CB",X"EE",X"CB",X"E6",X"CD",X"97",X"20",X"CD",
		X"A9",X"07",X"CD",X"97",X"25",X"CD",X"DD",X"28",X"CD",X"B3",X"31",X"CD",X"97",X"35",X"CD",X"44",
		X"0C",X"06",X"40",X"10",X"FE",X"3A",X"AB",X"42",X"A7",X"20",X"E1",X"3A",X"8E",X"42",X"CB",X"77",
		X"20",X"4D",X"FD",X"7E",X"06",X"A7",X"20",X"D4",X"AF",X"32",X"BD",X"42",X"32",X"BE",X"42",X"CD",
		X"64",X"0A",X"FD",X"CB",X"04",X"BE",X"FD",X"34",X"05",X"CD",X"D5",X"0C",X"CD",X"DF",X"0C",X"06",
		X"01",X"CD",X"C8",X"0C",X"21",X"CB",X"42",X"CB",X"CE",X"CB",X"4E",X"20",X"FC",X"21",X"CD",X"42",
		X"CB",X"4E",X"20",X"FC",X"06",X"02",X"CD",X"C8",X"0C",X"06",X"04",X"21",X"5F",X"42",X"CD",X"69",
		X"0A",X"C3",X"D0",X"08",X"06",X"18",X"21",X"77",X"42",X"AF",X"77",X"2B",X"10",X"FC",X"C9",X"AF",
		X"32",X"BE",X"42",X"32",X"BD",X"42",X"06",X"0C",X"CD",X"66",X"0A",X"CD",X"FD",X"20",X"06",X"01",
		X"CD",X"C8",X"0C",X"CD",X"64",X"0A",X"CD",X"DF",X"0C",X"06",X"03",X"CD",X"C8",X"0C",X"CD",X"55",
		X"08",X"06",X"01",X"CD",X"C0",X"0C",X"3A",X"8E",X"42",X"CB",X"47",X"28",X"F1",X"CD",X"10",X"2B",
		X"CD",X"1F",X"2B",X"38",X"0D",X"CB",X"59",X"28",X"F7",X"DD",X"CB",X"00",X"C6",X"FD",X"35",X"06",
		X"18",X"EE",X"AF",X"32",X"CE",X"42",X"FD",X"66",X"0B",X"FD",X"6E",X"0A",X"D7",X"CD",X"DF",X"0C",
		X"06",X"06",X"CD",X"C8",X"0C",X"FD",X"7E",X"06",X"B7",X"CC",X"D5",X"0C",X"FD",X"7E",X"05",X"B7",
		X"20",X"3D",X"21",X"CB",X"42",X"CB",X"FE",X"CB",X"7E",X"20",X"FC",X"21",X"CD",X"42",X"CB",X"7E",
		X"20",X"FC",X"21",X"88",X"0B",X"D7",X"06",X"05",X"CD",X"C8",X"0C",X"3A",X"8D",X"42",X"FE",X"01",
		X"28",X"09",X"CD",X"A6",X"0C",X"FD",X"7E",X"05",X"B7",X"20",X"3D",X"AF",X"32",X"8D",X"42",X"CD",
		X"EC",X"00",X"CA",X"22",X"04",X"3A",X"88",X"42",X"B7",X"C2",X"22",X"04",X"C3",X"32",X"02",X"3A",
		X"8D",X"42",X"FE",X"01",X"20",X"14",X"FD",X"7E",X"06",X"B7",X"20",X"07",X"FD",X"CB",X"04",X"BE",
		X"C3",X"D0",X"08",X"FD",X"CB",X"04",X"FE",X"C3",X"D0",X"08",X"CD",X"A6",X"0C",X"FD",X"7E",X"05",
		X"B7",X"20",X"05",X"CD",X"A6",X"0C",X"18",X"DE",X"CD",X"A6",X"0C",X"FD",X"7E",X"06",X"B7",X"20",
		X"08",X"FD",X"CB",X"04",X"BE",X"0E",X"00",X"18",X"06",X"FD",X"CB",X"04",X"FE",X"0E",X"01",X"CD",
		X"A6",X"0C",X"FD",X"7E",X"04",X"FD",X"CB",X"04",X"7E",X"28",X"02",X"CB",X"C9",X"06",X"1C",X"21",
		X"46",X"50",X"DD",X"21",X"B2",X"43",X"C5",X"06",X"18",X"56",X"DD",X"5E",X"00",X"CB",X"41",X"28",
		X"03",X"DD",X"72",X"00",X"CB",X"49",X"28",X"01",X"73",X"23",X"DD",X"23",X"10",X"EB",X"11",X"08",
		X"00",X"19",X"C1",X"10",X"E1",X"C3",X"D0",X"08",X"51",X"51",X"40",X"52",X"45",X"56",X"4F",X"40",
		X"40",X"45",X"4D",X"41",X"47",X"40",X"FF",X"FD",X"CB",X"04",X"7E",X"C0",X"21",X"3E",X"50",X"11",
		X"08",X"00",X"06",X"1C",X"19",X"C5",X"06",X"18",X"36",X"50",X"23",X"10",X"FB",X"C1",X"10",X"F4",
		X"DD",X"21",X"32",X"52",X"CD",X"3B",X"0E",X"FD",X"CB",X"04",X"76",X"C8",X"DD",X"21",X"06",X"52",
		X"06",X"0C",X"DD",X"36",X"00",X"4B",X"DD",X"36",X"20",X"4A",X"DD",X"23",X"10",X"F4",X"DD",X"36",
		X"00",X"10",X"DD",X"36",X"20",X"10",X"C9",X"21",X"07",X"42",X"01",X"02",X"03",X"CD",X"F5",X"0B",
		X"01",X"00",X"08",X"CD",X"F5",X"0B",X"06",X"06",X"0C",X"CD",X"F5",X"0B",X"06",X"06",X"0C",X"CD",
		X"F5",X"0B",X"06",X"04",X"0C",X"71",X"23",X"23",X"10",X"FB",X"C9",X"77",X"F5",X"23",X"3C",X"77",
		X"11",X"1F",X"00",X"19",X"3C",X"77",X"23",X"3C",X"77",X"F1",X"C9",X"AF",X"FD",X"77",X"00",X"FD",
		X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",X"04",X"3C",X"FD",X"77",X"03",X"3A",X"86",X"42",X"CB",
		X"3F",X"CB",X"3F",X"E6",X"01",X"C6",X"03",X"FD",X"77",X"05",X"C9",X"21",X"8F",X"42",X"36",X"10",
		X"3E",X"01",X"32",X"9B",X"42",X"32",X"9D",X"42",X"21",X"32",X"52",X"22",X"91",X"42",X"21",X"8E",
		X"42",X"36",X"00",X"C9",X"21",X"8E",X"42",X"CB",X"46",X"C0",X"CB",X"4E",X"C0",X"CB",X"76",X"C0",
		X"21",X"B9",X"42",X"35",X"C0",X"36",X"08",X"DD",X"21",X"5C",X"42",X"DD",X"56",X"00",X"DD",X"5E",
		X"03",X"CD",X"10",X"2B",X"CD",X"1F",X"2B",X"D8",X"CB",X"41",X"20",X"F8",X"CB",X"59",X"20",X"F4",
		X"CB",X"51",X"20",X"F0",X"CD",X"B3",X"2B",X"7A",X"CD",X"9C",X"0C",X"30",X"E7",X"7B",X"41",X"CD",
		X"9C",X"0C",X"30",X"E0",X"CD",X"5B",X"33",X"CD",X"8A",X"2B",X"3A",X"8E",X"42",X"CB",X"F7",X"32",
		X"8E",X"42",X"3E",X"05",X"32",X"9B",X"42",X"AF",X"32",X"9D",X"42",X"C9",X"B8",X"30",X"03",X"67",
		X"78",X"44",X"90",X"FE",X"05",X"C9",X"C5",X"FD",X"E5",X"C1",X"78",X"2F",X"C6",X"82",X"47",X"C5",
		X"FD",X"E1",X"3A",X"86",X"42",X"CB",X"5F",X"20",X"05",X"08",X"2F",X"C6",X"C9",X"08",X"C1",X"C9",
		X"0E",X"00",X"0D",X"20",X"FD",X"10",X"F9",X"C9",X"16",X"00",X"1E",X"00",X"1D",X"20",X"FD",X"15",
		X"20",X"F8",X"10",X"F4",X"C9",X"FD",X"7E",X"03",X"C6",X"01",X"27",X"FD",X"77",X"03",X"C9",X"21",
		X"CA",X"42",X"7E",X"E6",X"01",X"77",X"23",X"36",X"00",X"21",X"00",X"00",X"22",X"CC",X"42",X"C9",
		X"FD",X"E5",X"E1",X"01",X"80",X"00",X"A7",X"ED",X"42",X"22",X"A9",X"42",X"E5",X"DD",X"E1",X"21",
		X"1D",X"39",X"FD",X"CB",X"03",X"46",X"20",X"03",X"21",X"2F",X"39",X"06",X"03",X"FD",X"4E",X"04",
		X"CB",X"79",X"28",X"19",X"DD",X"CB",X"00",X"46",X"28",X"13",X"E5",X"5E",X"23",X"56",X"AF",X"12",
		X"13",X"12",X"13",X"12",X"13",X"12",X"E1",X"11",X"06",X"00",X"19",X"18",X"1B",X"DD",X"36",X"00",
		X"00",X"5E",X"DD",X"73",X"01",X"23",X"56",X"DD",X"72",X"02",X"23",X"CD",X"66",X"0D",X"7E",X"DD",
		X"77",X"05",X"23",X"7E",X"DD",X"77",X"06",X"23",X"11",X"07",X"00",X"DD",X"19",X"10",X"C1",X"FD",
		X"CB",X"04",X"7E",X"C0",X"01",X"15",X"39",X"FD",X"CB",X"03",X"46",X"20",X"04",X"03",X"03",X"03",
		X"03",X"CD",X"76",X"0D",X"18",X"10",X"7E",X"23",X"12",X"13",X"3E",X"2C",X"12",X"13",X"3E",X"04",
		X"12",X"13",X"7E",X"23",X"12",X"C9",X"0A",X"6F",X"03",X"0A",X"67",X"03",X"3E",X"4C",X"C3",X"FB",
		X"0B",X"FD",X"E5",X"E1",X"01",X"50",X"00",X"A7",X"ED",X"42",X"22",X"A0",X"42",X"22",X"A2",X"42",
		X"E5",X"DD",X"E1",X"11",X"40",X"00",X"21",X"41",X"39",X"FD",X"7E",X"03",X"FE",X"09",X"38",X"0A",
		X"CB",X"47",X"20",X"04",X"3E",X"08",X"18",X"02",X"3E",X"07",X"3D",X"28",X"03",X"19",X"18",X"FA",
		X"7E",X"32",X"9E",X"42",X"23",X"7E",X"32",X"9F",X"42",X"23",X"7E",X"32",X"A4",X"42",X"23",X"7E",
		X"32",X"A5",X"42",X"23",X"7E",X"32",X"A6",X"42",X"23",X"7E",X"FD",X"CB",X"04",X"7E",X"20",X"03",
		X"FD",X"77",X"06",X"23",X"47",X"5E",X"DD",X"73",X"04",X"23",X"56",X"DD",X"72",X"05",X"23",X"FD",
		X"CB",X"04",X"7E",X"20",X"0B",X"4E",X"DD",X"E5",X"D5",X"DD",X"E1",X"CD",X"37",X"0E",X"DD",X"E1",
		X"23",X"5E",X"DD",X"73",X"06",X"23",X"56",X"DD",X"72",X"07",X"23",X"FD",X"CB",X"04",X"7E",X"28",
		X"0B",X"DD",X"CB",X"00",X"46",X"28",X"05",X"23",X"23",X"23",X"18",X"1F",X"DD",X"E5",X"D5",X"DD",
		X"E1",X"56",X"23",X"5E",X"23",X"7E",X"23",X"CD",X"95",X"0E",X"DD",X"E1",X"DD",X"77",X"00",X"DD",
		X"36",X"01",X"00",X"DD",X"36",X"02",X"01",X"DD",X"36",X"08",X"00",X"11",X"0A",X"00",X"DD",X"19",
		X"10",X"A3",X"DD",X"36",X"00",X"00",X"C9",X"CB",X"41",X"20",X"2D",X"DD",X"36",X"A0",X"46",X"DD",
		X"36",X"A1",X"47",X"DD",X"36",X"40",X"44",X"DD",X"36",X"41",X"45",X"0E",X"48",X"DD",X"71",X"C0",
		X"DD",X"71",X"E0",X"DD",X"71",X"00",X"DD",X"71",X"20",X"0E",X"49",X"DD",X"71",X"C1",X"DD",X"71",
		X"E1",X"DD",X"71",X"01",X"DD",X"71",X"21",X"C9",X"DD",X"36",X"DE",X"46",X"DD",X"36",X"E3",X"47",
		X"DD",X"36",X"FE",X"44",X"DD",X"36",X"03",X"45",X"0E",X"4B",X"DD",X"71",X"DF",X"DD",X"71",X"E0",
		X"DD",X"71",X"E1",X"DD",X"71",X"E2",X"0E",X"4A",X"DD",X"71",X"FF",X"DD",X"71",X"00",X"DD",X"71",
		X"01",X"DD",X"71",X"02",X"C9",X"DD",X"72",X"00",X"DD",X"73",X"03",X"16",X"17",X"1E",X"07",X"CB",
		X"4F",X"28",X"04",X"16",X"15",X"1E",X"06",X"DD",X"72",X"01",X"DD",X"73",X"02",X"C9",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"00",X"18",X"09",X"04",X"10",X"10",X"10",X"05",X"08",X"F8",X"02",X"32",X"87",X"00",X"0D",
		X"01",X"1B",X"02",X"7F",X"00",X"FE",X"00",X"FC",X"01",X"6B",X"00",X"D6",X"00",X"AC",X"01",X"55",
		X"00",X"AA",X"00",X"53",X"01",X"47",X"00",X"8F",X"00",X"1D",X"01",X"55",X"00",X"AA",X"00",X"53",
		X"01",X"6B",X"00",X"D6",X"00",X"AC",X"01",X"7F",X"00",X"FE",X"00",X"FC",X"01",X"00",X"00",X"AF",
		X"CD",X"14",X"95",X"DD",X"7E",X"00",X"CD",X"14",X"95",X"82",X"57",X"23",X"DD",X"23",X"0B",X"1D",
		X"20",X"F1",X"AF",X"92",X"CD",X"14",X"95",X"18",X"C2",X"3E",X"3A",X"CD",X"31",X"95",X"AF",X"1E",
		X"03",X"CD",X"14",X"95",X"1D",X"20",X"FA",X"3C",X"CD",X"14",X"95",X"CD",X"4E",X"95",X"3E",X"FF",
		X"CD",X"14",X"95",X"CD",X"4E",X"95",X"3E",X"0D",X"CD",X"14",X"95",X"CD",X"4E",X"95",X"3E",X"0A",
		X"03",X"00",X"18",X"09",X"04",X"10",X"10",X"10",X"05",X"08",X"F8",X"02",X"42",X"87",X"00",X"0D",
		X"01",X"1B",X"02",X"7F",X"00",X"FE",X"00",X"FC",X"01",X"6B",X"00",X"D6",X"00",X"AC",X"01",X"55",
		X"00",X"AA",X"00",X"53",X"01",X"47",X"00",X"8F",X"00",X"1D",X"01",X"00",X"00",X"00",X"00",X"28",
		X"FA",X"DB",X"20",X"C9",X"FE",X"0A",X"30",X"03",X"F6",X"30",X"C9",X"C6",X"37",X"C9",X"21",X"00",
		X"80",X"2B",X"7C",X"B5",X"20",X"FB",X"C9",X"DD",X"21",X"00",X"A0",X"01",X"00",X"10",X"3A",X"F5",
		X"8F",X"FE",X"04",X"28",X"03",X"01",X"00",X"08",X"C9",X"3A",X"07",X"42",X"FE",X"00",X"28",X"25",
		X"FE",X"01",X"C2",X"CB",X"26",X"21",X"08",X"42",X"7E",X"B7",X"28",X"04",X"36",X"00",X"18",X"15",
		X"3E",X"01",X"77",X"32",X"05",X"42",X"3E",X"03",X"32",X"06",X"42",X"C3",X"87",X"00",X"21",X"49",
		X"03",X"00",X"18",X"09",X"04",X"01",X"10",X"10",X"05",X"00",X"FC",X"02",X"44",X"6B",X"00",X"D6",
		X"00",X"AC",X"01",X"04",X"01",X"01",X"01",X"47",X"00",X"8F",X"00",X"1D",X"01",X"04",X"10",X"10",
		X"10",X"47",X"00",X"8F",X"00",X"1D",X"01",X"6B",X"00",X"D6",X"00",X"AC",X"01",X"47",X"00",X"8F",
		X"00",X"1D",X"01",X"71",X"00",X"E2",X"00",X"C5",X"01",X"04",X"01",X"01",X"01",X"39",X"00",X"71",
		X"00",X"E2",X"00",X"04",X"10",X"10",X"10",X"39",X"00",X"71",X"00",X"E2",X"00",X"02",X"02",X"B4",
		X"00",X"68",X"01",X"CF",X"02",X"6B",X"00",X"D6",X"00",X"AC",X"01",X"02",X"06",X"32",X"00",X"39",
		X"00",X"71",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"8F",X"00",X"1D",X"01",X"20",X"32",X"01",
		X"01",X"01",X"01",X"02",X"06",X"6B",X"00",X"D6",X"00",X"32",X"3A",X"00",X"00",X"6B",X"61",X"76",
		X"03",X"00",X"18",X"09",X"04",X"10",X"10",X"10",X"05",X"08",X"F8",X"02",X"11",X"AA",X"00",X"97",
		X"00",X"8F",X"00",X"B4",X"00",X"A0",X"00",X"97",X"00",X"BE",X"00",X"AA",X"00",X"A0",X"00",X"CA",
		X"00",X"B4",X"00",X"AA",X"00",X"D6",X"00",X"BE",X"00",X"B4",X"00",X"E2",X"00",X"CA",X"00",X"BE",
		X"00",X"F0",X"00",X"D6",X"00",X"CA",X"00",X"FE",X"00",X"E2",X"00",X"D6",X"00",X"0D",X"01",X"F0",
		X"00",X"E2",X"00",X"1D",X"01",X"FE",X"00",X"F0",X"00",X"2E",X"01",X"0D",X"01",X"FE",X"00",X"00",
		X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"45",X"4E",
		X"44",X"0D",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"03",X"00",X"0A",X"09",X"04",X"10",X"10",X"10",X"05",X"00",X"F0",X"02",X"45",X"AC",X"01",X"7D",
		X"01",X"53",X"01",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"B4",X"00",X"B4",X"00",X"D6",
		X"00",X"D6",X"00",X"D6",X"00",X"00",X"00",X"20",X"20",X"4E",X"4D",X"49",X"52",X"45",X"54",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"3B",X"4A",X"6D",X"70",X"20",X"74",X"6F",
		X"20",X"4D",X"61",X"69",X"6E",X"20",X"4E",X"6D",X"69",X"20",X"50",X"47",X"2E",X"00",X"6F",X"72",
		X"6B",X"20",X"41",X"64",X"64",X"72",X"65",X"73",X"00",X"41",X"64",X"64",X"72",X"65",X"73",X"00",
		X"45",X"52",X"00",X"00",X"DE",X"20",X"B5",X"DD",X"CC",X"DF",X"29",X"0D",X"09",X"44",X"42",X"20",
		X"20",X"20",X"20",X"20",X"20",X"34",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"3B",X"4E",X"6F",
		X"69",X"73",X"65",X"20",X"34",X"0D",X"09",X"44",X"42",X"20",X"20",X"20",X"20",X"20",X"20",X"30",
		X"42",X"38",X"48",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"3B",X"4D",X"69",X"78",X"65",X"72",X"20",X"33",X"63",
		X"68",X"20",X"54",X"75",X"6E",X"65",X"20",X"49",X"2F",X"4F",X"20",X"3D",X"20",X"41",X"28",X"49",
		X"4E",X"29",X"00",X"00",X"27",X"02",X"81",X"80",X"62",X"D0",X"00",X"00",X"62",X"01",X"C5",X"00",
		X"01",X"01",X"62",X"CF",X"10",X"12",X"66",X"E7",X"01",X"01",X"00",X"00",X"27",X"02",X"00",X"00",
		X"27",X"02",X"81",X"80",X"BC",X"D1",X"00",X"00",X"62",X"01",X"C5",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"30",X"08",X"04",X"10",X"10",X"10",X"05",X"00",X"F0",X"02",X"43",X"1D",X"01",X"53",
		X"01",X"AC",X"01",X"00",X"00",X"AC",X"01",X"D6",X"00",X"50",X"00",X"A0",X"01",X"A0",X"00",X"71",
		X"00",X"C5",X"01",X"E2",X"00",X"47",X"00",X"1D",X"01",X"8F",X"00",X"6B",X"00",X"AC",X"01",X"D6",
		X"00",X"00",X"00",X"41",X"4D",X"45",X"4E",X"44",X"FF",X"43",X"00",X"00",X"49",X"4E",X"41",X"43",
		X"54",X"56",X"00",X"48",X"00",X"00",X"54",X"56",X"44",X"20",X"20",X"20",X"00",X"50",X"00",X"00",
		X"50",X"4F",X"52",X"54",X"31",X"20",X"00",X"60",X"00",X"00",X"50",X"4F",X"52",X"54",X"32",X"20",
		X"00",X"68",X"00",X"00",X"50",X"4F",X"52",X"54",X"33",X"20",X"00",X"70",X"00",X"00",X"43",X"55",
		X"50",X"20",X"20",X"20",X"80",X"40",X"00",X"00",X"43",X"44",X"57",X"20",X"20",X"20",X"C0",X"40",
		X"00",X"00",X"4D",X"49",X"53",X"53",X"20",X"20",X"60",X"68",X"00",X"00",X"4E",X"4D",X"49",X"20",
		X"20",X"20",X"01",X"70",X"00",X"00",X"4C",X"4F",X"43",X"41",X"54",X"45",X"06",X"70",X"00",X"00",
		X"52",X"45",X"53",X"45",X"54",X"20",X"00",X"78",X"00",X"00",X"50",X"53",X"55",X"44",X"20",X"20",
		X"06",X"00",X"00",X"00",X"50",X"53",X"55",X"44",X"32",X"20",X"03",X"00",X"00",X"00",X"50",X"53",
		X"4C",X"46",X"20",X"20",X"06",X"00",X"00",X"00",X"50",X"53",X"4C",X"46",X"32",X"20",X"03",X"00",
		X"00",X"00",X"49",X"53",X"55",X"44",X"20",X"20",X"02",X"00",X"00",X"00",X"4F",X"53",X"55",X"44",
		X"20",X"20",X"06",X"00",X"00",X"00",X"49",X"53",X"42",X"4B",X"20",X"20",X"08",X"00",X"00",X"00",
		X"46",X"43",X"45",X"58",X"20",X"20",X"14",X"00",X"00",X"00",X"43",X"53",X"44",X"4C",X"59",X"20",
		X"03",X"00",X"0A",X"09",X"04",X"10",X"10",X"10",X"05",X"00",X"F8",X"02",X"21",X"D6",X"00",X"AC",
		X"01",X"57",X"03",X"04",X"01",X"01",X"01",X"53",X"01",X"00",X"00",X"4C",X"55",X"04",X"10",X"10",
		X"10",X"D6",X"00",X"AC",X"01",X"57",X"03",X"8F",X"00",X"1D",X"01",X"3B",X"02",X"00",X"00",X"49",
		X"4D",X"45",X"0A",X"00",X"00",X"00",X"50",X"4C",X"41",X"59",X"31",X"20",X"00",X"40",X"00",X"00",
		X"50",X"4C",X"41",X"59",X"32",X"20",X"00",X"41",X"00",X"00",X"53",X"43",X"52",X"45",X"45",X"4E",
		X"03",X"00",X"00",X"00",X"53",X"52",X"56",X"46",X"4C",X"47",X"04",X"00",X"00",X"00",X"50",X"41",
		X"43",X"4B",X"4D",X"4E",X"05",X"00",X"00",X"00",X"54",X"45",X"4E",X"53",X"4F",X"20",X"06",X"00",
		X"00",X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",X"07",X"00",X"00",X"00",X"42",X"4E",X"53",X"50",
		X"4F",X"54",X"09",X"00",X"00",X"00",X"54",X"56",X"20",X"20",X"20",X"20",X"77",X"00",X"00",X"00",
		X"50",X"41",X"43",X"50",X"4F",X"54",X"78",X"00",X"00",X"00",X"54",X"45",X"4E",X"44",X"54",X"20",
		X"7A",X"00",X"00",X"00",X"55",X"50",X"41",X"44",X"52",X"20",X"7C",X"00",X"00",X"00",X"53",X"43",
		X"52",X"41",X"44",X"52",X"7E",X"00",X"00",X"00",X"53",X"50",X"45",X"45",X"44",X"20",X"80",X"41",
		X"00",X"00",X"4F",X"49",X"4B",X"41",X"4B",X"45",X"98",X"41",X"00",X"00",X"42",X"4E",X"53",X"41",
		X"44",X"44",X"DA",X"41",X"00",X"00",X"48",X"49",X"53",X"43",X"4F",X"52",X"00",X"42",X"00",X"00",
		X"50",X"4C",X"59",X"4E",X"55",X"4D",X"03",X"42",X"00",X"00",X"43",X"52",X"45",X"44",X"49",X"54",
		X"04",X"42",X"00",X"00",X"43",X"4F",X"49",X"4E",X"54",X"4D",X"05",X"42",X"00",X"00",X"43",X"43",
		X"03",X"00",X"0A",X"09",X"04",X"10",X"10",X"10",X"05",X"00",X"F8",X"02",X"11",X"AC",X"01",X"C5",
		X"01",X"FC",X"01",X"94",X"01",X"AC",X"01",X"E0",X"01",X"7D",X"01",X"94",X"01",X"C5",X"01",X"68",
		X"01",X"7D",X"01",X"AC",X"01",X"53",X"01",X"68",X"01",X"94",X"01",X"40",X"01",X"53",X"01",X"7D",
		X"01",X"2E",X"01",X"40",X"01",X"68",X"01",X"1D",X"01",X"2E",X"01",X"53",X"01",X"0D",X"01",X"1D",
		X"01",X"40",X"01",X"FE",X"00",X"0D",X"01",X"2E",X"01",X"F0",X"00",X"FE",X"00",X"1D",X"01",X"E2",
		X"00",X"F0",X"00",X"0D",X"01",X"D6",X"00",X"E2",X"00",X"FE",X"00",X"CA",X"00",X"D6",X"00",X"F0",
		X"00",X"BE",X"00",X"CA",X"00",X"E2",X"00",X"B4",X"00",X"BE",X"00",X"D6",X"00",X"AA",X"00",X"B4",
		X"00",X"CA",X"00",X"A0",X"00",X"AA",X"00",X"BE",X"00",X"97",X"00",X"A0",X"00",X"B4",X"00",X"8F",
		X"00",X"97",X"00",X"AA",X"00",X"00",X"00",X"00",X"02",X"FE",X"00",X"FC",X"01",X"FC",X"01",X"0D",
		X"01",X"1B",X"02",X"1B",X"02",X"FE",X"00",X"FC",X"01",X"FC",X"01",X"F0",X"00",X"E0",X"01",X"E0",
		X"01",X"E2",X"00",X"C5",X"01",X"C5",X"01",X"F0",X"00",X"E0",X"01",X"E0",X"01",X"E2",X"00",X"C5",
		X"01",X"C5",X"01",X"02",X"08",X"D6",X"00",X"AC",X"01",X"AC",X"01",X"00",X"00",X"50",X"41",X"43",
		X"4B",X"20",X"1A",X"42",X"00",X"00",X"50",X"4F",X"57",X"45",X"52",X"31",X"1B",X"42",X"00",X"00",
		X"50",X"4F",X"57",X"45",X"52",X"32",X"1C",X"42",X"00",X"00",X"50",X"4F",X"57",X"45",X"52",X"33",
		X"1D",X"42",X"00",X"00",X"54",X"49",X"4D",X"45",X"52",X"33",X"1E",X"42",X"00",X"00",X"54",X"49",
		X"4D",X"45",X"52",X"34",X"1F",X"42",X"00",X"00",X"4F",X"49",X"4B",X"41",X"54",X"4D",X"21",X"42",
		X"03",X"00",X"0A",X"09",X"04",X"10",X"10",X"01",X"05",X"00",X"F8",X"02",X"12",X"1B",X"02",X"35",
		X"04",X"3B",X"02",X"FC",X"01",X"F9",X"03",X"5D",X"02",X"FC",X"01",X"F9",X"03",X"3B",X"02",X"E0",
		X"01",X"C0",X"03",X"1B",X"02",X"E0",X"01",X"C0",X"03",X"FC",X"01",X"C5",X"01",X"8A",X"03",X"1B",
		X"02",X"C5",X"01",X"8A",X"03",X"FC",X"01",X"02",X"04",X"AC",X"01",X"57",X"03",X"02",X"04",X"00",
		X"00",X"C5",X"01",X"C5",X"01",X"02",X"02",X"F0",X"00",X"E0",X"01",X"E0",X"01",X"FE",X"00",X"FC",
		X"01",X"FC",X"01",X"02",X"06",X"FE",X"00",X"FC",X"01",X"FC",X"01",X"02",X"02",X"FE",X"00",X"FC",
		X"01",X"FC",X"01",X"0D",X"01",X"1B",X"02",X"1B",X"02",X"FE",X"00",X"FC",X"01",X"FC",X"01",X"F0",
		X"00",X"E0",X"01",X"E0",X"01",X"E2",X"00",X"C5",X"01",X"C5",X"01",X"F0",X"00",X"01",X"E0",X"01",
		X"03",X"00",X"18",X"09",X"04",X"10",X"10",X"01",X"05",X"00",X"F8",X"02",X"51",X"AA",X"00",X"53",
		X"01",X"AA",X"00",X"A0",X"00",X"40",X"01",X"AA",X"00",X"97",X"00",X"2E",X"01",X"AA",X"00",X"02",
		X"02",X"04",X"10",X"10",X"10",X"8F",X"00",X"1D",X"01",X"EB",X"08",X"04",X"10",X"10",X"01",X"AA",
		X"00",X"53",X"01",X"AA",X"00",X"04",X"10",X"10",X"10",X"A0",X"00",X"40",X"01",X"6B",X"08",X"04",
		X"10",X"10",X"01",X"BE",X"00",X"7D",X"01",X"AA",X"00",X"04",X"10",X"10",X"10",X"AA",X"00",X"53",
		X"01",X"F2",X"07",X"04",X"10",X"10",X"01",X"D6",X"00",X"AC",X"01",X"AA",X"00",X"04",X"10",X"10",
		X"10",X"BE",X"00",X"7D",X"01",X"14",X"07",X"04",X"10",X"10",X"01",X"E2",X"00",X"C5",X"01",X"AA",
		X"00",X"04",X"10",X"10",X"10",X"04",X"10",X"10",X"10",X"D6",X"00",X"AC",X"01",X"AE",X"00",X"04",
		X"01",X"01",X"01",X"AA",X"00",X"AA",X"01",X"AA",X"02",X"04",X"10",X"10",X"01",X"6B",X"00",X"D6",
		X"00",X"AA",X"00",X"04",X"10",X"10",X"10",X"D6",X"00",X"AC",X"01",X"AE",X"06",X"00",X"00",X"02",
		X"02",X"04",X"10",X"10",X"10",X"8F",X"00",X"1D",X"01",X"EB",X"08",X"04",X"10",X"10",X"01",X"AA",
		X"00",X"53",X"01",X"AA",X"00",X"04",X"10",X"10",X"10",X"A0",X"00",X"40",X"01",X"6B",X"08",X"04",
		X"10",X"10",X"01",X"BE",X"00",X"7D",X"01",X"AA",X"00",X"04",X"10",X"10",X"10",X"AA",X"00",X"53",
		X"01",X"F2",X"07",X"04",X"10",X"10",X"01",X"D6",X"00",X"AC",X"01",X"AA",X"00",X"04",X"10",X"10",
		X"10",X"BE",X"00",X"7D",X"01",X"14",X"07",X"04",X"10",X"10",X"01",X"E2",X"00",X"C5",X"01",X"AA",
		X"00",X"04",X"10",X"10",X"10",X"04",X"10",X"10",X"10",X"D6",X"00",X"AC",X"01",X"AE",X"00",X"04",
		X"01",X"01",X"01",X"AA",X"00",X"AA",X"01",X"AA",X"02",X"04",X"10",X"10",X"01",X"6B",X"00",X"D6",
		X"00",X"AA",X"00",X"04",X"10",X"10",X"10",X"D6",X"00",X"AC",X"01",X"AE",X"06",X"00",X"FF",X"53",
		X"01",X"02",X"06",X"D6",X"00",X"1D",X"01",X"53",X"01",X"AA",X"00",X"D6",X"00",X"1D",X"01",X"02",
		X"04",X"AA",X"00",X"D6",X"00",X"1D",X"01",X"AA",X"00",X"D6",X"00",X"1D",X"01",X"02",X"06",X"AA",
		X"00",X"D6",X"00",X"1D",X"01",X"8F",X"00",X"AA",X"00",X"D6",X"00",X"8F",X"00",X"AA",X"00",X"D6",
		X"00",X"8F",X"00",X"AA",X"00",X"D6",X"00",X"02",X"08",X"6B",X"00",X"8F",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"4C",X"43",X"54",X"20",X"20",X"20",X"09",X"00",X"00",X"00",X"4F",X"55",X"54",X"53",
		X"54",X"52",X"10",X"00",X"00",X"00",X"4F",X"55",X"54",X"53",X"54",X"31",X"17",X"00",X"00",X"00",
		X"03",X"00",X"20",X"09",X"04",X"10",X"10",X"10",X"05",X"00",X"F8",X"02",X"42",X"4C",X"00",X"5A",
		X"00",X"7F",X"00",X"50",X"00",X"5F",X"00",X"87",X"00",X"55",X"00",X"65",X"00",X"8F",X"00",X"5A",
		X"00",X"6B",X"00",X"97",X"00",X"5F",X"00",X"71",X"00",X"A0",X"00",X"65",X"00",X"78",X"00",X"AA",
		X"00",X"6B",X"00",X"7F",X"00",X"B4",X"00",X"02",X"06",X"40",X"00",X"5A",X"00",X"6B",X"00",X"00",
		X"00",X"20",X"5E",X"00",X"00",X"00",X"4E",X"4D",X"49",X"30",X"31",X"20",X"78",X"00",X"00",X"00",
		X"4E",X"4D",X"49",X"52",X"45",X"54",X"87",X"00",X"00",X"00",X"4E",X"4D",X"49",X"30",X"32",X"20",
		X"9D",X"00",X"00",X"00",X"4D",X"41",X"49",X"4E",X"20",X"20",X"AF",X"00",X"00",X"00",X"4D",X"41",
		X"49",X"4E",X"31",X"20",X"C7",X"00",X"00",X"00",X"4D",X"41",X"49",X"4E",X"32",X"20",X"D2",X"00",
		X"02",X"24",X"03",X"00",X"05",X"04",X"04",X"0F",X"0F",X"0F",X"05",X"04",X"B8",X"00",X"00",X"4E",
		X"35",X"20",X"FE",X"00",X"00",X"00",X"4D",X"41",X"49",X"4E",X"35",X"31",X"06",X"01",X"00",X"00",
		X"4D",X"41",X"49",X"4E",X"36",X"20",X"11",X"01",X"00",X"00",X"4D",X"41",X"49",X"4E",X"37",X"20",
		X"02",X"24",X"03",X"00",X"05",X"04",X"04",X"0F",X"0F",X"0F",X"05",X"04",X"B8",X"00",X"00",X"45",
		X"41",X"44",X"32",X"20",X"98",X"01",X"00",X"00",X"44",X"45",X"41",X"44",X"33",X"20",X"9E",X"01",
		X"00",X"00",X"44",X"45",X"41",X"44",X"33",X"30",X"AE",X"01",X"00",X"00",X"44",X"45",X"41",X"44",
		X"02",X"24",X"03",X"00",X"05",X"04",X"04",X"0F",X"0F",X"0F",X"05",X"04",X"B8",X"00",X"00",X"00",
		X"44",X"45",X"4D",X"4F",X"20",X"20",X"F8",X"01",X"00",X"00",X"4D",X"49",X"53",X"43",X"4C",X"52",
		X"03",X"00",X"09",X"09",X"04",X"10",X"10",X"10",X"05",X"08",X"F8",X"02",X"02",X"97",X"00",X"2E",
		X"01",X"AE",X"06",X"8F",X"00",X"1D",X"01",X"75",X"04",X"8F",X"00",X"1D",X"01",X"AE",X"06",X"8F",
		X"00",X"1D",X"01",X"75",X"04",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"14",X"07",X"04",
		X"10",X"10",X"10",X"8F",X"00",X"1D",X"01",X"75",X"04",X"8F",X"00",X"1D",X"01",X"14",X"07",X"8F",
		X"00",X"1D",X"01",X"75",X"04",X"8F",X"00",X"1D",X"01",X"80",X"07",X"8F",X"00",X"1D",X"01",X"75",
		X"04",X"8F",X"00",X"1D",X"01",X"80",X"07",X"8F",X"00",X"1D",X"01",X"75",X"04",X"04",X"01",X"01",
		X"10",X"AA",X"00",X"AA",X"01",X"F2",X"07",X"04",X"10",X"10",X"10",X"8F",X"00",X"1D",X"01",X"75",
		X"04",X"8F",X"00",X"1D",X"01",X"F2",X"07",X"8F",X"00",X"1D",X"01",X"75",X"04",X"AA",X"00",X"53",
		X"01",X"6B",X"08",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"06",X"05",X"04",X"10",X"10",
		X"10",X"BE",X"00",X"7D",X"01",X"6B",X"08",X"AA",X"00",X"53",X"01",X"06",X"05",X"04",X"01",X"01",
		X"10",X"AA",X"00",X"AA",X"01",X"6B",X"08",X"04",X"10",X"10",X"10",X"BE",X"00",X"7D",X"01",X"06",
		X"05",X"AA",X"00",X"53",X"01",X"6B",X"08",X"BE",X"00",X"7D",X"01",X"06",X"05",X"AA",X"00",X"53",
		X"01",X"EB",X"08",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"06",X"05",X"AA",X"00",X"AA",
		X"01",X"EB",X"08",X"AA",X"00",X"AA",X"01",X"06",X"05",X"04",X"10",X"10",X"10",X"BE",X"00",X"7D",
		X"01",X"F2",X"07",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"06",X"05",X"AA",X"00",X"AA",
		X"01",X"F2",X"07",X"AA",X"00",X"AA",X"01",X"06",X"05",X"04",X"10",X"10",X"10",X"B4",X"00",X"68",
		X"01",X"AE",X"06",X"AA",X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"AE",X"06",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"14",X"07",X"04",
		X"10",X"10",X"10",X"AA",X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"14",X"07",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"80",X"07",X"AA",X"00",X"53",X"01",X"75",
		X"04",X"AA",X"00",X"53",X"01",X"80",X"07",X"AA",X"00",X"53",X"01",X"75",X"04",X"04",X"01",X"01",
		X"10",X"AA",X"00",X"AA",X"01",X"F2",X"07",X"04",X"10",X"10",X"10",X"AA",X"00",X"53",X"01",X"75",
		X"04",X"AA",X"00",X"53",X"01",X"F2",X"07",X"AA",X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",
		X"01",X"6B",X"08",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"06",X"05",X"04",X"10",X"10",
		X"10",X"BE",X"00",X"7D",X"01",X"6B",X"08",X"AA",X"00",X"53",X"01",X"06",X"05",X"04",X"01",X"01",
		X"10",X"AA",X"00",X"AA",X"01",X"6B",X"08",X"04",X"10",X"10",X"10",X"BE",X"00",X"7D",X"01",X"06",
		X"05",X"AA",X"00",X"53",X"01",X"6B",X"08",X"BE",X"00",X"7D",X"01",X"06",X"05",X"8F",X"00",X"1D",
		X"01",X"EB",X"08",X"04",X"01",X"10",X"10",X"AA",X"00",X"81",X"02",X"06",X"05",X"AA",X"00",X"75",
		X"04",X"EB",X"08",X"AA",X"00",X"81",X"02",X"06",X"05",X"AA",X"00",X"35",X"04",X"6B",X"08",X"AA",
		X"00",X"81",X"02",X"06",X"05",X"AA",X"00",X"F9",X"03",X"F2",X"07",X"AA",X"00",X"81",X"02",X"06",
		X"05",X"04",X"10",X"10",X"10",X"00",X"FF",X"AA",X"00",X"AA",X"01",X"06",X"05",X"AA",X"00",X"AA",
		X"01",X"F2",X"07",X"AA",X"00",X"AA",X"01",X"06",X"05",X"04",X"10",X"10",X"10",X"B4",X"00",X"68",
		X"01",X"AE",X"06",X"AA",X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"AE",X"06",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"14",X"07",X"04",
		X"10",X"10",X"10",X"AA",X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"14",X"07",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"80",X"07",X"AA",X"00",X"53",X"01",X"75",
		X"04",X"AA",X"00",X"53",X"01",X"80",X"07",X"AA",X"00",X"53",X"01",X"75",X"04",X"04",X"01",X"01",
		X"10",X"AA",X"00",X"AA",X"01",X"F2",X"07",X"04",X"10",X"10",X"10",X"AA",X"00",X"53",X"01",X"75",
		X"04",X"AA",X"00",X"53",X"01",X"F2",X"07",X"AA",X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",
		X"01",X"6B",X"08",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"01",X"06",X"05",X"04",X"10",X"10",
		X"03",X"00",X"18",X"09",X"04",X"08",X"08",X"10",X"05",X"08",X"F8",X"02",X"52",X"97",X"00",X"2E",
		X"01",X"5D",X"02",X"A0",X"00",X"40",X"01",X"81",X"02",X"97",X"00",X"2E",X"01",X"5D",X"02",X"A0",
		X"00",X"40",X"01",X"81",X"02",X"2E",X"01",X"5D",X"02",X"B9",X"04",X"40",X"01",X"81",X"02",X"06",
		X"05",X"2E",X"01",X"5D",X"02",X"B9",X"04",X"40",X"01",X"81",X"02",X"06",X"05",X"00",X"FF",X"75",
		X"04",X"EB",X"08",X"AA",X"00",X"81",X"02",X"06",X"05",X"AA",X"00",X"35",X"04",X"6B",X"08",X"AA",
		X"00",X"81",X"02",X"06",X"05",X"AA",X"00",X"F9",X"03",X"F2",X"07",X"AA",X"00",X"81",X"02",X"06",
		X"05",X"04",X"10",X"10",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"00",X"09",X"09",X"04",X"10",X"10",X"10",X"05",X"08",X"F8",X"02",X"42",X"97",X"00",X"2E",
		X"01",X"5D",X"02",X"8F",X"00",X"1D",X"01",X"3B",X"02",X"8F",X"00",X"1D",X"01",X"3B",X"02",X"8F",
		X"00",X"1D",X"01",X"3B",X"02",X"2E",X"01",X"5D",X"02",X"B9",X"04",X"1D",X"01",X"3B",X"02",X"75",
		X"04",X"1D",X"01",X"3B",X"02",X"75",X"04",X"1D",X"01",X"3B",X"02",X"75",X"04",X"5D",X"02",X"B9",
		X"04",X"73",X"09",X"3B",X"02",X"75",X"04",X"EB",X"08",X"3B",X"02",X"75",X"04",X"EB",X"08",X"3B",
		X"02",X"75",X"04",X"EB",X"08",X"04",X"01",X"01",X"01",X"3B",X"02",X"75",X"04",X"EB",X"08",X"8F",
		X"00",X"1D",X"01",X"75",X"04",X"8F",X"00",X"1D",X"01",X"F9",X"03",X"8F",X"00",X"1D",X"01",X"8A",
		X"03",X"8F",X"00",X"1D",X"01",X"57",X"03",X"04",X"01",X"01",X"10",X"8F",X"00",X"1D",X"01",X"75",
		X"04",X"04",X"10",X"10",X"10",X"AA",X"00",X"53",X"01",X"57",X"03",X"04",X"01",X"01",X"10",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"04",X"10",X"10",X"10",X"8F",X"00",X"1D",X"01",X"57",X"03",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"04",X"01",X"01",X"10",X"AA",X"00",X"53",X"01",X"57",X"03",X"04",
		X"10",X"10",X"10",X"8F",X"00",X"1D",X"01",X"75",X"04",X"7F",X"00",X"FE",X"00",X"57",X"03",X"AA",
		X"00",X"53",X"01",X"75",X"04",X"AA",X"00",X"53",X"01",X"57",X"03",X"AA",X"00",X"53",X"01",X"75",
		X"04",X"04",X"01",X"01",X"10",X"AA",X"00",X"AA",X"00",X"57",X"03",X"04",X"10",X"10",X"10",X"BE",
		X"04",X"7D",X"01",X"75",X"04",X"D6",X"00",X"AC",X"01",X"57",X"03",X"04",X"01",X"01",X"10",X"D6",
		X"00",X"AC",X"01",X"75",X"04",X"04",X"10",X"10",X"10",X"CA",X"00",X"94",X"01",X"C0",X"03",X"04",
		X"01",X"01",X"10",X"94",X"01",X"E0",X"01",X"75",X"04",X"04",X"10",X"10",X"10",X"1D",X"01",X"3B",
		X"02",X"C0",X"03",X"04",X"01",X"01",X"10",X"1D",X"01",X"3B",X"02",X"75",X"04",X"04",X"10",X"10",
		X"10",X"D6",X"00",X"AC",X"01",X"C0",X"03",X"1D",X"01",X"3B",X"02",X"75",X"04",X"F0",X"00",X"E0",
		X"01",X"C0",X"03",X"D6",X"00",X"AC",X"01",X"75",X"04",X"00",X"00",X"01",X"01",X"01",X"01",X"8F",
		X"00",X"1D",X"01",X"1D",X"01",X"01",X"01",X"01",X"01",X"AA",X"00",X"53",X"01",X"53",X"01",X"01",
		X"01",X"01",X"01",X"D6",X"00",X"AC",X"01",X"AC",X"01",X"01",X"01",X"01",X"01",X"B4",X"00",X"68",
		X"01",X"68",X"01",X"01",X"01",X"01",X"01",X"AA",X"00",X"53",X"01",X"53",X"01",X"01",X"01",X"01",
		X"01",X"B4",X"00",X"68",X"01",X"68",X"01",X"01",X"01",X"01",X"01",X"AA",X"00",X"53",X"01",X"53",
		X"01",X"01",X"01",X"01",X"01",X"02",X"06",X"D6",X"00",X"AC",X"01",X"AC",X"01",X"01",X"01",X"01",
		X"01",X"6B",X"00",X"7F",X"00",X"8F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5C",X"46",X"92",X"92",X"92",X"75",X"75",X"75",X"85",X"FE",X"85",X"85",X"46",X"46",X"75",X"46",
		X"46",X"92",X"92",X"92",X"85",X"75",X"75",X"75",X"5C",X"85",X"5C",X"5C",X"FE",X"5C",X"5C",X"3B",
		X"46",X"46",X"46",X"46",X"75",X"85",X"46",X"85",X"5C",X"FE",X"5C",X"5C",X"5C",X"5C",X"75",X"85",
		X"92",X"75",X"75",X"75",X"75",X"5C",X"46",X"46",X"46",X"5C",X"92",X"92",X"92",X"46",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"9E",X"A9",X"98",X"AE",
		X"92",X"B3",X"8D",X"B7",X"85",X"B7",X"85",X"B3",X"8D",X"AE",X"92",X"A9",X"A8",X"A5",X"9E",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"8E",X"42",X"7E",X"47",X"E6",X"C3",X"28",X"12",
		X"FE",X"80",X"20",X"59",X"78",X"E6",X"18",X"FE",X"18",X"20",X"52",X"3A",X"AF",X"42",X"CB",X"4F",
		X"20",X"4B",X"21",X"9D",X"42",X"35",X"C0",X"36",X"01",X"DD",X"2A",X"91",X"42",X"21",X"8F",X"42",
		X"CB",X"46",X"C2",X"09",X"22",X"3E",X"08",X"32",X"9B",X"42",X"0E",X"00",X"08",X"47",X"08",X"0A",
		X"CB",X"57",X"C2",X"45",X"21",X"CB",X"5F",X"20",X"2A",X"CB",X"6F",X"C2",X"83",X"21",X"57",X"3A",
		X"86",X"42",X"CB",X"5F",X"20",X"08",X"FD",X"E5",X"C1",X"78",X"FE",X"41",X"28",X"07",X"CB",X"72",
		X"C2",X"CC",X"21",X"18",X"08",X"3A",X"00",X"60",X"CB",X"7F",X"C2",X"CC",X"21",X"21",X"CD",X"42",
		X"CB",X"A6",X"C9",X"3A",X"5C",X"42",X"FE",X"E0",X"28",X"F3",X"C6",X"10",X"47",X"3A",X"5F",X"42",
		X"4F",X"CD",X"4A",X"24",X"38",X"E7",X"CD",X"04",X"25",X"DD",X"7E",X"C0",X"EB",X"DD",X"22",X"97",
		X"42",X"DD",X"E5",X"E1",X"01",X"20",X"00",X"A7",X"ED",X"42",X"22",X"99",X"42",X"A7",X"ED",X"42",
		X"22",X"93",X"42",X"DD",X"E5",X"E1",X"01",X"60",X"00",X"A7",X"ED",X"42",X"EB",X"0E",X"11",X"CD",
		X"B8",X"23",X"C3",X"F3",X"22",X"3A",X"5C",X"42",X"FE",X"10",X"CA",X"FD",X"20",X"D6",X"10",X"47",
		X"3A",X"5F",X"42",X"4F",X"CD",X"4A",X"24",X"DA",X"FD",X"20",X"CD",X"04",X"25",X"DD",X"7E",X"20",
		X"EB",X"DD",X"22",X"97",X"42",X"DD",X"E5",X"E1",X"01",X"20",X"00",X"09",X"22",X"99",X"42",X"09",
		X"22",X"93",X"42",X"DD",X"E5",X"E1",X"01",X"20",X"00",X"09",X"EB",X"0E",X"21",X"CD",X"B8",X"23",
		X"C3",X"3E",X"23",X"3A",X"5F",X"42",X"FE",X"20",X"CA",X"FD",X"20",X"D6",X"10",X"4F",X"3A",X"5C",
		X"42",X"47",X"CD",X"4A",X"24",X"DA",X"FD",X"20",X"CD",X"04",X"25",X"DD",X"7E",X"FF",X"EB",X"DD",
		X"22",X"97",X"42",X"DD",X"E5",X"E1",X"2B",X"22",X"99",X"42",X"2B",X"22",X"93",X"42",X"DD",X"E5",
		X"E1",X"01",X"22",X"00",X"A7",X"ED",X"42",X"EB",X"0E",X"81",X"CD",X"B8",X"23",X"3A",X"5F",X"42",
		X"FE",X"30",X"C2",X"5D",X"22",X"CB",X"CE",X"CB",X"D6",X"C3",X"5D",X"22",X"3A",X"5F",X"42",X"FE",
		X"E0",X"CA",X"FD",X"20",X"C6",X"10",X"4F",X"3A",X"5C",X"42",X"47",X"CD",X"4A",X"24",X"DA",X"FD",
		X"20",X"CD",X"04",X"25",X"DD",X"7E",X"02",X"EB",X"DD",X"22",X"97",X"42",X"DD",X"E5",X"E1",X"23",
		X"22",X"99",X"42",X"23",X"22",X"93",X"42",X"DD",X"E5",X"E1",X"01",X"1E",X"00",X"A7",X"ED",X"42",
		X"EB",X"0E",X"41",X"CD",X"B8",X"23",X"C3",X"A8",X"22",X"0E",X"00",X"08",X"47",X"08",X"0A",X"57",
		X"E6",X"2C",X"20",X"19",X"3A",X"86",X"42",X"CB",X"5F",X"20",X"26",X"FD",X"E5",X"C1",X"78",X"FE",
		X"41",X"20",X"1E",X"3A",X"00",X"60",X"CB",X"7F",X"CA",X"FD",X"20",X"18",X"19",X"CB",X"57",X"28",
		X"04",X"CB",X"66",X"18",X"13",X"CB",X"5F",X"28",X"04",X"CB",X"6E",X"18",X"0B",X"CB",X"76",X"18",
		X"07",X"CB",X"72",X"CA",X"FD",X"20",X"CB",X"7E",X"C4",X"35",X"25",X"CD",X"04",X"25",X"CB",X"66",
		X"C2",X"F3",X"22",X"CB",X"6E",X"C2",X"3E",X"23",X"CB",X"76",X"C2",X"A8",X"22",X"21",X"5F",X"42",
		X"35",X"35",X"CD",X"0D",X"24",X"CD",X"5B",X"33",X"78",X"F5",X"A7",X"28",X"0D",X"FE",X"01",X"28",
		X"03",X"CD",X"89",X"22",X"11",X"FF",X"FF",X"CD",X"32",X"24",X"F1",X"FE",X"03",X"28",X"04",X"CB",
		X"4E",X"28",X"03",X"CD",X"89",X"22",X"C3",X"67",X"23",X"DD",X"2A",X"91",X"42",X"E5",X"DD",X"7E",
		X"00",X"21",X"C4",X"24",X"CD",X"3C",X"24",X"DD",X"71",X"00",X"DD",X"7E",X"E0",X"21",X"D4",X"24",
		X"CD",X"3C",X"24",X"DD",X"71",X"E0",X"E1",X"C9",X"21",X"5F",X"42",X"34",X"34",X"CD",X"0D",X"24",
		X"CD",X"5B",X"33",X"78",X"F5",X"A7",X"28",X"0D",X"FE",X"01",X"28",X"03",X"CD",X"D4",X"22",X"11",
		X"01",X"00",X"CD",X"32",X"24",X"F1",X"FE",X"03",X"28",X"04",X"CB",X"4E",X"28",X"03",X"CD",X"D4",
		X"22",X"C3",X"67",X"23",X"DD",X"2A",X"91",X"42",X"E5",X"DD",X"7E",X"01",X"21",X"E4",X"24",X"CD",
		X"3C",X"24",X"DD",X"71",X"01",X"DD",X"7E",X"E1",X"21",X"F4",X"24",X"CD",X"3C",X"24",X"DD",X"71",
		X"E1",X"E1",X"C9",X"21",X"5C",X"42",X"34",X"34",X"CD",X"0D",X"24",X"CD",X"5B",X"33",X"78",X"F5",
		X"A7",X"28",X"0D",X"FE",X"01",X"28",X"03",X"CD",X"1F",X"23",X"11",X"E0",X"FF",X"CD",X"32",X"24",
		X"F1",X"FE",X"03",X"28",X"04",X"CB",X"4E",X"28",X"03",X"CD",X"1F",X"23",X"C3",X"67",X"23",X"DD",
		X"2A",X"91",X"42",X"E5",X"DD",X"7E",X"E0",X"21",X"84",X"24",X"CD",X"3C",X"24",X"DD",X"71",X"E0",
		X"DD",X"7E",X"E1",X"21",X"94",X"24",X"CD",X"3C",X"24",X"DD",X"71",X"E1",X"E1",X"C9",X"21",X"5C",
		X"42",X"35",X"35",X"CD",X"0D",X"24",X"CD",X"5B",X"33",X"78",X"F5",X"A7",X"28",X"0D",X"FE",X"01",
		X"28",X"03",X"CD",X"7F",X"23",X"11",X"20",X"00",X"CD",X"32",X"24",X"F1",X"FE",X"03",X"28",X"04",
		X"CB",X"4E",X"28",X"03",X"CD",X"7F",X"23",X"CB",X"5E",X"28",X"04",X"3E",X"19",X"18",X"02",X"3E",
		X"26",X"32",X"9D",X"42",X"21",X"9B",X"42",X"35",X"C0",X"21",X"8F",X"42",X"CB",X"86",X"C9",X"DD",
		X"2A",X"91",X"42",X"E5",X"DD",X"7E",X"00",X"21",X"A4",X"24",X"CD",X"3C",X"24",X"DD",X"71",X"00",
		X"DD",X"7E",X"01",X"21",X"B4",X"24",X"CD",X"3C",X"24",X"DD",X"71",X"01",X"E1",X"C9",X"06",X"00",
		X"FE",X"10",X"C8",X"FE",X"B4",X"D0",X"04",X"FE",X"50",X"C8",X"04",X"FE",X"4C",X"D0",X"04",X"FE",
		X"4A",X"D0",X"04",X"FE",X"48",X"D0",X"04",X"C9",X"47",X"7E",X"E6",X"08",X"B1",X"77",X"78",X"CD",
		X"9E",X"23",X"78",X"FE",X"00",X"C8",X"FE",X"02",X"28",X"18",X"38",X"32",X"FE",X"05",X"28",X"0E",
		X"79",X"E6",X"30",X"78",X"28",X"05",X"FE",X"04",X"C8",X"18",X"03",X"FE",X"03",X"C8",X"CB",X"D6",
		X"18",X"28",X"3E",X"50",X"12",X"13",X"12",X"EB",X"01",X"1F",X"00",X"09",X"EB",X"12",X"13",X"12",
		X"CB",X"DE",X"E5",X"21",X"BD",X"42",X"CB",X"C6",X"21",X"BC",X"42",X"36",X"03",X"E1",X"C5",X"D5",
		X"01",X"00",X"00",X"16",X"10",X"CD",X"CC",X"06",X"D1",X"C1",X"CB",X"CE",X"C9",X"06",X"00",X"21",
		X"8F",X"42",X"3A",X"9B",X"42",X"FE",X"07",X"28",X"0B",X"FE",X"03",X"28",X"01",X"C9",X"CB",X"4E",
		X"28",X"0E",X"18",X"0B",X"CB",X"4E",X"28",X"08",X"CB",X"56",X"28",X"03",X"CB",X"8E",X"04",X"04",
		X"04",X"C9",X"E5",X"2A",X"91",X"42",X"19",X"22",X"91",X"42",X"E1",X"C9",X"06",X"08",X"4F",X"BE",
		X"20",X"03",X"23",X"4E",X"C9",X"23",X"23",X"10",X"F6",X"C9",X"D5",X"E5",X"DD",X"E5",X"DD",X"2A",
		X"A9",X"42",X"16",X"03",X"DD",X"CB",X"00",X"46",X"20",X"17",X"DD",X"CB",X"00",X"4E",X"20",X"11",
		X"DD",X"66",X"02",X"DD",X"6E",X"01",X"78",X"BE",X"20",X"07",X"23",X"23",X"23",X"79",X"BE",X"28",
		X"0D",X"D5",X"11",X"07",X"00",X"DD",X"19",X"D1",X"15",X"20",X"D9",X"A7",X"18",X"01",X"37",X"DD",
		X"E1",X"E1",X"D1",X"C9",X"3E",X"48",X"50",X"40",X"40",X"42",X"42",X"46",X"46",X"3E",X"44",X"48",
		X"4A",X"10",X"4B",X"10",X"3F",X"49",X"50",X"41",X"41",X"43",X"43",X"47",X"47",X"3F",X"45",X"49",
		X"4A",X"10",X"4B",X"10",X"38",X"48",X"50",X"3A",X"3A",X"3C",X"3C",X"44",X"44",X"38",X"46",X"48",
		X"4A",X"10",X"4B",X"10",X"39",X"49",X"50",X"3B",X"3B",X"3D",X"3D",X"45",X"45",X"39",X"47",X"49",
		X"4A",X"10",X"4B",X"10",X"32",X"4A",X"50",X"34",X"34",X"36",X"36",X"44",X"44",X"32",X"45",X"4A",
		X"48",X"10",X"49",X"10",X"33",X"4B",X"50",X"35",X"35",X"37",X"37",X"46",X"46",X"33",X"47",X"4B",
		X"48",X"10",X"49",X"10",X"2C",X"4A",X"50",X"2E",X"2E",X"30",X"30",X"45",X"45",X"2C",X"44",X"4A",
		X"48",X"10",X"49",X"10",X"2D",X"4B",X"50",X"2F",X"2F",X"31",X"31",X"47",X"47",X"2D",X"46",X"4B",
		X"48",X"10",X"49",X"10",X"F5",X"E5",X"21",X"CD",X"42",X"CB",X"E6",X"FD",X"7E",X"06",X"FE",X"01",
		X"28",X"16",X"3A",X"A6",X"42",X"B7",X"28",X"10",X"3A",X"8F",X"42",X"CB",X"5F",X"20",X"09",X"3A",
		X"7F",X"43",X"E6",X"0F",X"F6",X"40",X"18",X"07",X"3A",X"7F",X"43",X"E6",X"0F",X"F6",X"30",X"32",
		X"7F",X"43",X"E1",X"F1",X"C9",X"E5",X"3A",X"8F",X"42",X"E6",X"08",X"F6",X"01",X"47",X"CD",X"DE",
		X"33",X"28",X"06",X"E6",X"30",X"F6",X"CF",X"18",X"04",X"E6",X"C0",X"F6",X"3F",X"2F",X"B0",X"32",
		X"90",X"42",X"2A",X"91",X"42",X"3A",X"9B",X"42",X"FE",X"06",X"20",X"05",X"2A",X"97",X"42",X"18",
		X"07",X"FE",X"02",X"20",X"03",X"2A",X"99",X"42",X"22",X"95",X"42",X"47",X"3E",X"08",X"90",X"32",
		X"9C",X"42",X"2A",X"97",X"42",X"ED",X"5B",X"93",X"42",X"22",X"93",X"42",X"ED",X"53",X"97",X"42",
		X"CD",X"8A",X"2B",X"3A",X"90",X"42",X"32",X"8F",X"42",X"3A",X"9C",X"42",X"32",X"9B",X"42",X"2A",
		X"95",X"42",X"22",X"91",X"42",X"E1",X"C9",X"3A",X"8E",X"42",X"CB",X"47",X"C0",X"CB",X"77",X"C0",
		X"2A",X"A2",X"42",X"7E",X"A7",X"20",X"12",X"2A",X"A0",X"42",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"CB",X"47",X"20",X"2A",X"E5",X"DD",X"E1",
		X"23",X"47",X"4E",X"79",X"E6",X"0F",X"20",X"24",X"CD",X"D5",X"25",X"DD",X"66",X"07",X"DD",X"6E",
		X"06",X"C3",X"F1",X"25",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"22",X"A2",
		X"42",X"C9",X"06",X"80",X"10",X"FE",X"C9",X"CD",X"E2",X"25",X"18",X"E8",X"CD",X"E2",X"25",X"18",
		X"E4",X"DD",X"35",X"02",X"C0",X"CB",X"50",X"CA",X"F6",X"26",X"CB",X"60",X"C4",X"44",X"26",X"CB",
		X"68",X"C4",X"41",X"26",X"23",X"23",X"23",X"CB",X"70",X"C4",X"44",X"26",X"CB",X"78",X"C4",X"41",
		X"26",X"DD",X"35",X"03",X"20",X"1B",X"DD",X"CB",X"00",X"96",X"CB",X"58",X"28",X"13",X"DD",X"56",
		X"05",X"DD",X"5E",X"04",X"1A",X"FE",X"50",X"28",X"08",X"FE",X"4E",X"28",X"04",X"DD",X"CB",X"00",
		X"9E",X"3A",X"9E",X"42",X"DD",X"CB",X"00",X"5E",X"28",X"03",X"3A",X"9F",X"42",X"DD",X"77",X"02",
		X"C9",X"35",X"35",X"C9",X"34",X"34",X"C9",X"D5",X"E5",X"DD",X"E5",X"01",X"00",X"00",X"DD",X"56",
		X"05",X"DD",X"5E",X"04",X"D5",X"DD",X"E1",X"7E",X"23",X"23",X"23",X"56",X"21",X"B2",X"26",X"DD",
		X"5E",X"E0",X"CD",X"99",X"26",X"21",X"B5",X"26",X"DD",X"5E",X"00",X"CD",X"99",X"26",X"7A",X"21",
		X"BB",X"26",X"DD",X"5E",X"01",X"CD",X"99",X"26",X"FE",X"20",X"20",X"0F",X"F5",X"DD",X"7E",X"02",
		X"FE",X"10",X"28",X"06",X"FE",X"4A",X"28",X"02",X"CB",X"B9",X"F1",X"21",X"B8",X"26",X"DD",X"5E",
		X"00",X"CD",X"99",X"26",X"DD",X"E1",X"E1",X"D1",X"C9",X"F5",X"BE",X"28",X"0F",X"7B",X"23",X"1E",
		X"02",X"BE",X"28",X"06",X"23",X"1D",X"20",X"F9",X"CB",X"C1",X"CB",X"C0",X"CB",X"09",X"CB",X"08",
		X"F1",X"C9",X"E0",X"46",X"4B",X"10",X"44",X"4A",X"20",X"44",X"48",X"E0",X"45",X"49",X"E5",X"1E",
		X"00",X"56",X"23",X"23",X"23",X"FD",X"7E",X"06",X"FE",X"01",X"3A",X"5C",X"42",X"20",X"02",X"3E",
		X"10",X"BA",X"28",X"08",X"38",X"04",X"CB",X"E3",X"18",X"02",X"CB",X"EB",X"56",X"FD",X"7E",X"06",
		X"FE",X"01",X"3A",X"5F",X"42",X"20",X"02",X"3E",X"20",X"BA",X"28",X"08",X"38",X"04",X"CB",X"F3",
		X"18",X"02",X"CB",X"FB",X"E1",X"C9",X"CD",X"47",X"26",X"CD",X"BE",X"26",X"DD",X"CB",X"00",X"5E",
		X"C2",X"65",X"28",X"FD",X"7E",X"06",X"FE",X"01",X"CC",X"B4",X"28",X"DD",X"CB",X"00",X"4E",X"C4",
		X"0D",X"35",X"DD",X"7E",X"00",X"E6",X"30",X"7B",X"CA",X"B1",X"27",X"E6",X"C0",X"5F",X"28",X"05",
		X"CD",X"6A",X"28",X"18",X"18",X"79",X"E6",X"C0",X"20",X"23",X"78",X"E6",X"C0",X"FE",X"C0",X"5F",
		X"20",X"0B",X"CD",X"AC",X"28",X"28",X"04",X"CB",X"BB",X"18",X"02",X"CB",X"B3",X"CD",X"C9",X"28",
		X"E6",X"F0",X"20",X"09",X"7B",X"DD",X"CB",X"00",X"DE",X"CD",X"6C",X"28",X"76",X"DD",X"7E",X"00",
		X"E6",X"0F",X"57",X"DD",X"7E",X"00",X"E6",X"30",X"B2",X"DD",X"77",X"00",X"3A",X"AB",X"42",X"B7",
		X"28",X"11",X"3A",X"AC",X"42",X"BE",X"20",X"0B",X"DD",X"7E",X"00",X"E6",X"30",X"CD",X"6A",X"28",
		X"C3",X"3F",X"28",X"DD",X"7E",X"00",X"E6",X"30",X"A1",X"20",X"1D",X"79",X"E6",X"C0",X"5F",X"28",
		X"14",X"FE",X"C0",X"20",X"0B",X"CD",X"AC",X"28",X"28",X"04",X"CB",X"BB",X"18",X"02",X"CB",X"B3",
		X"7B",X"CD",X"6C",X"28",X"76",X"59",X"18",X"F8",X"79",X"E6",X"C0",X"5F",X"28",X"0B",X"FE",X"C0",
		X"28",X"07",X"CD",X"C9",X"28",X"FE",X"A0",X"30",X"E7",X"DD",X"7E",X"00",X"E6",X"30",X"5F",X"18",
		X"DF",X"E6",X"30",X"5F",X"28",X"05",X"CD",X"6A",X"28",X"18",X"18",X"79",X"E6",X"30",X"20",X"23",
		X"78",X"E6",X"30",X"FE",X"30",X"5F",X"20",X"0B",X"CD",X"AC",X"28",X"28",X"04",X"CB",X"AB",X"18",
		X"02",X"CB",X"A3",X"CD",X"C9",X"28",X"E6",X"F0",X"20",X"09",X"7B",X"DD",X"CB",X"00",X"DE",X"CD",
		X"6C",X"28",X"76",X"DD",X"7E",X"00",X"E6",X"0F",X"57",X"DD",X"7E",X"00",X"E6",X"C0",X"B2",X"DD",
		X"77",X"00",X"3A",X"AB",X"42",X"B7",X"28",X"09",X"3A",X"AC",X"42",X"BE",X"20",X"03",X"C3",X"3F",
		X"28",X"DD",X"7E",X"00",X"E6",X"C0",X"A1",X"20",X"1D",X"79",X"E6",X"30",X"5F",X"28",X"14",X"FE",
		X"30",X"20",X"0B",X"CD",X"AC",X"28",X"28",X"04",X"CB",X"AB",X"18",X"02",X"CB",X"A3",X"7B",X"CD",
		X"6C",X"28",X"76",X"59",X"18",X"F8",X"79",X"E6",X"30",X"5F",X"28",X"0B",X"FE",X"30",X"28",X"07",
		X"CD",X"C9",X"28",X"FE",X"A0",X"30",X"E7",X"DD",X"7E",X"00",X"E6",X"C0",X"5F",X"18",X"DF",X"79",
		X"E6",X"30",X"5F",X"28",X"14",X"FE",X"30",X"20",X"0B",X"CD",X"AC",X"28",X"28",X"04",X"CB",X"AB",
		X"18",X"02",X"CB",X"A3",X"7B",X"CD",X"6C",X"28",X"76",X"79",X"E6",X"C0",X"5F",X"FE",X"C0",X"20",
		X"F3",X"1E",X"40",X"18",X"EF",X"7B",X"CD",X"6C",X"28",X"76",X"A1",X"C8",X"4F",X"DD",X"CB",X"00",
		X"D6",X"DD",X"7E",X"00",X"E6",X"0F",X"B1",X"47",X"F1",X"DD",X"36",X"03",X"08",X"DD",X"70",X"00",
		X"E5",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"40",X"00",X"CB",X"60",X"28",X"03",X"A7",X"ED",
		X"52",X"CB",X"68",X"28",X"01",X"19",X"CB",X"70",X"28",X"02",X"23",X"23",X"CB",X"78",X"28",X"02",
		X"2B",X"2B",X"DD",X"75",X"04",X"DD",X"74",X"05",X"E1",X"C3",X"FA",X"25",X"57",X"CD",X"C9",X"28",
		X"CB",X"7F",X"7A",X"C9",X"7E",X"B7",X"20",X"09",X"FD",X"35",X"06",X"DD",X"CB",X"00",X"C6",X"F1",
		X"C9",X"7B",X"B7",X"C0",X"3E",X"20",X"C3",X"6C",X"28",X"D9",X"2A",X"A7",X"42",X"E5",X"D1",X"29",
		X"29",X"E5",X"C1",X"29",X"09",X"19",X"23",X"22",X"A7",X"42",X"7C",X"D9",X"C9",X"DD",X"2A",X"A9",
		X"42",X"06",X"03",X"DD",X"CB",X"00",X"46",X"20",X"15",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"DD",
		X"56",X"06",X"DD",X"5E",X"05",X"C5",X"DD",X"E5",X"CD",X"06",X"29",X"DD",X"E1",X"C1",X"11",X"07",
		X"00",X"DD",X"19",X"10",X"DE",X"C9",X"DD",X"CB",X"00",X"4E",X"20",X"42",X"3A",X"AB",X"42",X"A7",
		X"C0",X"DD",X"CB",X"00",X"7E",X"3A",X"8F",X"42",X"20",X"17",X"CB",X"47",X"C0",X"3A",X"5C",X"42",
		X"BE",X"C0",X"3A",X"5F",X"42",X"D6",X"10",X"23",X"23",X"23",X"BE",X"C0",X"DD",X"CB",X"00",X"FE",
		X"C9",X"CB",X"47",X"C8",X"3E",X"01",X"32",X"AB",X"42",X"7E",X"32",X"AC",X"42",X"DD",X"36",X"03",
		X"FF",X"DD",X"36",X"04",X"04",X"DD",X"CB",X"00",X"CE",X"DD",X"CB",X"00",X"96",X"C9",X"DD",X"35",
		X"03",X"C0",X"DD",X"CB",X"00",X"56",X"20",X"30",X"DD",X"36",X"03",X"50",X"DD",X"CB",X"04",X"46",
		X"7E",X"06",X"04",X"28",X"03",X"80",X"18",X"01",X"90",X"77",X"DD",X"35",X"04",X"C0",X"DD",X"CB",
		X"00",X"D6",X"DD",X"CB",X"00",X"9E",X"DD",X"CB",X"00",X"E6",X"DD",X"36",X"03",X"80",X"AF",X"32",
		X"AD",X"42",X"21",X"CA",X"42",X"CB",X"DE",X"C9",X"DD",X"CB",X"00",X"5E",X"C2",X"26",X"2A",X"DD",
		X"36",X"03",X"03",X"23",X"23",X"23",X"7E",X"FE",X"E0",X"28",X"63",X"E6",X"0F",X"20",X"17",X"DD",
		X"CB",X"00",X"66",X"20",X"05",X"CD",X"DE",X"2B",X"38",X"54",X"13",X"13",X"DD",X"72",X"06",X"DD",
		X"73",X"05",X"DD",X"CB",X"00",X"A6",X"34",X"34",X"5E",X"2B",X"2B",X"2B",X"56",X"DD",X"E5",X"CD",
		X"10",X"2B",X"AF",X"32",X"AE",X"42",X"CD",X"1F",X"2B",X"38",X"12",X"CB",X"41",X"20",X"09",X"CB",
		X"59",X"20",X"F3",X"CD",X"3C",X"2B",X"18",X"EE",X"CD",X"6C",X"2B",X"18",X"E9",X"21",X"5C",X"42",
		X"3A",X"8E",X"42",X"CB",X"47",X"20",X"10",X"CB",X"4F",X"20",X"09",X"CB",X"77",X"20",X"08",X"CD",
		X"71",X"2B",X"18",X"03",X"CD",X"6C",X"2B",X"DD",X"E1",X"3A",X"AE",X"42",X"A7",X"C8",X"DD",X"CB",
		X"00",X"DE",X"DD",X"CB",X"00",X"F6",X"DD",X"36",X"03",X"FF",X"21",X"CC",X"42",X"CB",X"9E",X"21",
		X"CA",X"42",X"CB",X"9E",X"CB",X"E6",X"3A",X"AD",X"42",X"A7",X"C0",X"3A",X"8E",X"42",X"CB",X"4F",
		X"C0",X"DD",X"CB",X"00",X"EE",X"C9",X"DD",X"CB",X"00",X"6E",X"28",X"2A",X"DD",X"36",X"03",X"8C",
		X"DD",X"CB",X"00",X"76",X"28",X"08",X"DD",X"CB",X"00",X"B6",X"23",X"36",X"22",X"C9",X"23",X"7E",
		X"FE",X"23",X"28",X"03",X"36",X"23",X"C9",X"CD",X"EE",X"2A",X"2B",X"DD",X"CB",X"00",X"C6",X"AF",
		X"77",X"23",X"23",X"23",X"77",X"C9",X"DD",X"CB",X"00",X"76",X"28",X"77",X"3A",X"AD",X"42",X"A7",
		X"20",X"09",X"CD",X"EE",X"2A",X"CD",X"4B",X"2A",X"C3",X"F9",X"2A",X"DD",X"CB",X"00",X"B6",X"DD",
		X"36",X"03",X"FF",X"47",X"FD",X"7E",X"06",X"90",X"FD",X"77",X"06",X"3A",X"8E",X"42",X"CB",X"4F",
		X"C4",X"0A",X"2B",X"E5",X"21",X"10",X"00",X"1E",X"25",X"05",X"28",X"04",X"29",X"1C",X"10",X"FC",
		X"16",X"00",X"E5",X"C1",X"CD",X"CC",X"06",X"E1",X"7E",X"D6",X"08",X"77",X"C6",X"10",X"57",X"23",
		X"73",X"23",X"36",X"07",X"23",X"5E",X"CD",X"10",X"2B",X"AF",X"32",X"AE",X"42",X"CD",X"1F",X"2B",
		X"D8",X"CB",X"41",X"28",X"F8",X"3A",X"AE",X"42",X"A7",X"20",X"0F",X"3C",X"32",X"AE",X"42",X"72",
		X"23",X"36",X"24",X"23",X"36",X"07",X"23",X"73",X"18",X"E3",X"DD",X"CB",X"00",X"C6",X"CD",X"4F",
		X"2A",X"18",X"DA",X"CD",X"F3",X"2A",X"CD",X"4B",X"2A",X"CD",X"EE",X"2A",X"CD",X"10",X"2B",X"CD",
		X"1F",X"2B",X"D8",X"CB",X"41",X"28",X"F8",X"DD",X"CB",X"00",X"C6",X"C3",X"4F",X"2A",X"AF",X"32",
		X"AB",X"42",X"C9",X"3A",X"8E",X"42",X"CB",X"4F",X"C8",X"3A",X"8E",X"42",X"CB",X"F7",X"32",X"8E",
		X"42",X"3E",X"05",X"32",X"9B",X"42",X"AF",X"32",X"9D",X"42",X"3E",X"00",X"32",X"5D",X"42",X"C9",
		X"E5",X"2A",X"A0",X"42",X"01",X"0A",X"00",X"A7",X"ED",X"42",X"E5",X"DD",X"E1",X"E1",X"C9",X"01",
		X"0A",X"00",X"DD",X"09",X"DD",X"7E",X"00",X"A7",X"28",X"10",X"CB",X"47",X"20",X"F4",X"47",X"DD",
		X"4E",X"01",X"DD",X"66",X"07",X"DD",X"6E",X"06",X"A7",X"C9",X"37",X"C9",X"CD",X"B3",X"2B",X"CD",
		X"C1",X"2B",X"D8",X"DD",X"CB",X"01",X"56",X"28",X"09",X"DD",X"CB",X"01",X"66",X"28",X"03",X"CD",
		X"5B",X"33",X"DD",X"CB",X"01",X"4E",X"C4",X"5F",X"36",X"DD",X"CB",X"01",X"C6",X"3A",X"AD",X"42",
		X"3C",X"32",X"AD",X"42",X"79",X"FE",X"E0",X"C0",X"32",X"AE",X"42",X"C9",X"CD",X"B9",X"2B",X"18",
		X"F3",X"CD",X"B3",X"2B",X"CD",X"C1",X"2B",X"D8",X"CD",X"5B",X"33",X"3A",X"8E",X"42",X"CB",X"CF",
		X"32",X"8E",X"42",X"C5",X"CD",X"8A",X"2B",X"C1",X"18",X"DA",X"3A",X"8F",X"42",X"CB",X"47",X"C8",
		X"CB",X"4F",X"C8",X"CB",X"67",X"28",X"05",X"CD",X"F8",X"22",X"18",X"EE",X"CB",X"6F",X"28",X"05",
		X"CD",X"43",X"23",X"18",X"E5",X"CB",X"77",X"28",X"05",X"CD",X"AD",X"22",X"18",X"DC",X"CD",X"62",
		X"22",X"18",X"D7",X"46",X"23",X"23",X"23",X"4E",X"C9",X"46",X"23",X"23",X"23",X"34",X"34",X"4E",
		X"C9",X"7A",X"C5",X"B8",X"30",X"03",X"4F",X"78",X"41",X"90",X"C1",X"FE",X"0D",X"30",X"0D",X"7B",
		X"C6",X"08",X"B9",X"28",X"05",X"C6",X"02",X"B9",X"20",X"02",X"A7",X"C9",X"37",X"C9",X"DD",X"E5",
		X"D5",X"DD",X"E1",X"DD",X"7E",X"02",X"FE",X"50",X"28",X"28",X"FE",X"4E",X"28",X"24",X"CD",X"16",
		X"2C",X"DD",X"77",X"02",X"DD",X"7E",X"E2",X"CD",X"16",X"2C",X"DD",X"77",X"E2",X"DD",X"7E",X"01",
		X"CD",X"16",X"2C",X"DD",X"77",X"01",X"DD",X"7E",X"E1",X"CD",X"16",X"2C",X"DD",X"77",X"E1",X"A7",
		X"18",X"01",X"37",X"DD",X"E1",X"C9",X"E5",X"21",X"29",X"2C",X"06",X"06",X"BE",X"28",X"06",X"23",
		X"23",X"10",X"F9",X"E1",X"C9",X"23",X"7E",X"E1",X"C9",X"44",X"4A",X"45",X"4A",X"46",X"4B",X"47",
		X"4B",X"48",X"10",X"49",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"20",X"35",X"38",X"00",X"00",X"54",X"52",X"55",X"44",X"41",X"54",X"15",X"39",X"00",X"00",
		X"49",X"57",X"44",X"41",X"54",X"41",X"1D",X"39",X"00",X"00",X"4F",X"49",X"4B",X"44",X"41",X"54",
		X"41",X"39",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"16",X"00",X"CD",X"EC",X"00",X"CA",X"26",X"21",X"3A",
		X"89",X"42",X"FE",X"00",X"20",X"59",X"CD",X"DC",X"00",X"CA",X"26",X"21",X"1E",X"01",X"CD",X"EC",
		X"00",X"FE",X"00",X"28",X"24",X"FE",X"01",X"20",X"19",X"21",X"8C",X"42",X"7E",X"B7",X"28",X"04",
		X"36",X"00",X"18",X"15",X"3E",X"01",X"77",X"32",X"89",X"42",X"3E",X"03",X"32",X"8A",X"42",X"C3",
		X"26",X"21",X"21",X"8B",X"42",X"34",X"1C",X"18",X"03",X"21",X"8B",X"42",X"34",X"3E",X"01",X"32",
		X"89",X"42",X"3E",X"04",X"32",X"8A",X"42",X"3A",X"8D",X"42",X"B7",X"20",X"07",X"3A",X"88",X"42",
		X"B7",X"20",X"01",X"14",X"3A",X"88",X"42",X"83",X"27",X"32",X"88",X"42",X"C3",X"26",X"21",X"FE",
		X"01",X"21",X"8A",X"42",X"20",X"0E",X"35",X"C2",X"26",X"21",X"3E",X"02",X"32",X"89",X"42",X"36",
		X"03",X"C3",X"26",X"21",X"35",X"20",X"07",X"AF",X"32",X"89",X"42",X"C3",X"26",X"21",X"CD",X"DC",
		X"00",X"CA",X"26",X"21",X"36",X"03",X"3A",X"00",X"78",X"3A",X"7C",X"42",X"C3",X"B6",X"00",X"3A",
		X"BE",X"42",X"B7",X"C8",X"3A",X"BA",X"42",X"67",X"2E",X"00",X"3A",X"B0",X"42",X"57",X"A7",X"20",
		X"0E",X"CD",X"AD",X"31",X"20",X"0E",X"21",X"B1",X"42",X"35",X"20",X"0F",X"3C",X"18",X"0C",X"CD",
		X"AD",X"31",X"28",X"07",X"06",X"05",X"AF",X"21",X"B1",X"42",X"70",X"32",X"B0",X"42",X"7A",X"32",
		X"AF",X"42",X"3A",X"8E",X"42",X"47",X"E6",X"43",X"C0",X"CB",X"78",X"C0",X"3A",X"AF",X"42",X"FE",
		X"03",X"C0",X"3E",X"14",X"32",X"B2",X"42",X"CD",X"40",X"33",X"06",X"80",X"2A",X"93",X"42",X"22",
		X"B5",X"42",X"3A",X"8F",X"42",X"CB",X"47",X"20",X"10",X"2A",X"91",X"42",X"22",X"B5",X"42",X"CD",
		X"E1",X"32",X"22",X"B5",X"42",X"30",X"0C",X"18",X"08",X"CB",X"4F",X"28",X"06",X"CB",X"57",X"20",
		X"02",X"CB",X"D0",X"78",X"32",X"8E",X"42",X"21",X"CA",X"42",X"CB",X"EE",X"C9",X"CB",X"66",X"C8",
		X"CB",X"CA",X"C9",X"3A",X"8E",X"42",X"47",X"E6",X"43",X"C0",X"21",X"B7",X"42",X"35",X"C0",X"36",
		X"03",X"CB",X"78",X"C8",X"CB",X"50",X"28",X"0D",X"21",X"CA",X"42",X"CB",X"AE",X"21",X"CC",X"42",
		X"CB",X"AE",X"C3",X"5B",X"33",X"CB",X"60",X"C2",X"8E",X"32",X"CD",X"A3",X"32",X"CD",X"7E",X"33",
		X"DD",X"21",X"6C",X"42",X"DD",X"56",X"00",X"DD",X"5E",X"03",X"CD",X"DE",X"33",X"06",X"08",X"28",
		X"0C",X"CB",X"67",X"7A",X"20",X"03",X"90",X"18",X"01",X"80",X"57",X"18",X"0A",X"CB",X"77",X"7B",
		X"20",X"03",X"90",X"18",X"01",X"80",X"5F",X"CD",X"10",X"2B",X"CD",X"1F",X"2B",X"38",X"58",X"CB",
		X"41",X"20",X"F7",X"CB",X"59",X"20",X"F3",X"DD",X"7E",X"08",X"FE",X"05",X"28",X"EC",X"CD",X"B3",
		X"2B",X"7A",X"CD",X"99",X"32",X"30",X"E3",X"7B",X"41",X"CD",X"99",X"32",X"30",X"DC",X"DD",X"CB",
		X"01",X"4E",X"C4",X"5F",X"36",X"DD",X"22",X"B3",X"42",X"DD",X"CB",X"01",X"D6",X"DD",X"CB",X"01",
		X"E6",X"DD",X"34",X"08",X"DD",X"36",X"09",X"80",X"21",X"CA",X"42",X"CB",X"F6",X"3A",X"8E",X"42",
		X"CB",X"DF",X"CB",X"E7",X"32",X"8E",X"42",X"3E",X"14",X"32",X"B2",X"42",X"21",X"CA",X"42",X"CB",
		X"AE",X"21",X"CC",X"42",X"CB",X"AE",X"C9",X"CD",X"DE",X"33",X"28",X"05",X"3A",X"6C",X"42",X"18",
		X"03",X"3A",X"6F",X"42",X"E6",X"0F",X"20",X"0F",X"CD",X"E1",X"32",X"22",X"B5",X"42",X"30",X"07",
		X"3A",X"8E",X"42",X"CB",X"9F",X"18",X"CB",X"21",X"B2",X"42",X"35",X"C0",X"18",X"F2",X"CB",X"58",
		X"C0",X"21",X"B2",X"42",X"35",X"C0",X"C3",X"5B",X"33",X"B8",X"30",X"03",X"67",X"78",X"44",X"90",
		X"FE",X"05",X"C9",X"3A",X"8F",X"42",X"4F",X"21",X"6C",X"42",X"E6",X"30",X"20",X"03",X"21",X"6F",
		X"42",X"DD",X"21",X"6D",X"42",X"06",X"03",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"CD",X"CF",X"32",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"23",X"23",X"23",X"23",X"10",X"E9",X"C9",X"CB",
		X"79",X"C2",X"41",X"26",X"CB",X"71",X"C2",X"44",X"26",X"CB",X"69",X"C2",X"41",X"26",X"C3",X"44",
		X"26",X"C5",X"D5",X"DD",X"E5",X"2A",X"B5",X"42",X"DD",X"21",X"34",X"33",X"3A",X"8F",X"42",X"47",
		X"3A",X"6F",X"42",X"4F",X"3A",X"6C",X"42",X"CB",X"60",X"20",X"1B",X"DD",X"23",X"DD",X"23",X"DD",
		X"23",X"CB",X"68",X"20",X"11",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"79",X"CB",X"70",X"20",X"06",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"BE",X"00",X"28",X"16",X"DD",X"56",X"02",X"DD",X"5E",
		X"01",X"19",X"7E",X"FE",X"50",X"28",X"0A",X"FE",X"4E",X"28",X"06",X"A7",X"DD",X"E1",X"D1",X"C1",
		X"C9",X"37",X"18",X"F8",X"E0",X"C0",X"FF",X"10",X"40",X"00",X"E0",X"02",X"00",X"20",X"FE",X"FF",
		X"21",X"6C",X"42",X"3A",X"5C",X"42",X"57",X"3A",X"5F",X"42",X"5F",X"06",X"03",X"72",X"23",X"36",
		X"00",X"23",X"36",X"07",X"23",X"73",X"23",X"10",X"F4",X"18",X"23",X"F5",X"C5",X"E5",X"21",X"6C",
		X"42",X"06",X"0C",X"36",X"00",X"23",X"10",X"FB",X"3A",X"8E",X"42",X"CB",X"BF",X"CB",X"5F",X"28",
		X"06",X"2A",X"B3",X"42",X"23",X"CB",X"A6",X"32",X"8E",X"42",X"E1",X"C1",X"F1",X"C9",X"DD",X"21",
		X"6D",X"42",X"CD",X"DE",X"33",X"28",X"05",X"21",X"E7",X"33",X"18",X"03",X"21",X"03",X"34",X"3A",
		X"B2",X"42",X"06",X"07",X"BE",X"28",X"08",X"D0",X"23",X"23",X"23",X"23",X"10",X"F6",X"C9",X"23",
		X"4E",X"23",X"56",X"23",X"5E",X"CD",X"DE",X"33",X"28",X"16",X"CB",X"67",X"20",X"26",X"AF",X"B9",
		X"28",X"02",X"CB",X"F9",X"BA",X"28",X"02",X"CB",X"FA",X"BB",X"28",X"18",X"CB",X"FB",X"18",X"14",
		X"CB",X"7F",X"20",X"10",X"AF",X"B9",X"28",X"02",X"CB",X"F1",X"BA",X"28",X"02",X"CB",X"F2",X"BB",
		X"28",X"02",X"CB",X"F3",X"DD",X"71",X"00",X"DD",X"72",X"04",X"DD",X"73",X"08",X"C9",X"3A",X"8F",
		X"42",X"E6",X"30",X"3A",X"8F",X"42",X"C9",X"14",X"01",X"00",X"00",X"11",X"01",X"03",X"00",X"10",
		X"02",X"05",X"00",X"0C",X"01",X"06",X"00",X"09",X"01",X"06",X"03",X"08",X"02",X"04",X"05",X"04",
		X"01",X"06",X"06",X"14",X"07",X"00",X"00",X"11",X"07",X"09",X"00",X"10",X"08",X"0B",X"00",X"0C",
		X"07",X"0C",X"00",X"09",X"07",X"0C",X"09",X"08",X"08",X"0A",X"0B",X"04",X"07",X"0C",X"0C",X"3A",
		X"BE",X"42",X"B7",X"C8",X"21",X"8E",X"42",X"7E",X"E6",X"43",X"C0",X"CD",X"10",X"2B",X"CD",X"1F",
		X"2B",X"D8",X"CB",X"41",X"20",X"F8",X"CB",X"51",X"28",X"F4",X"CB",X"59",X"20",X"59",X"DD",X"7E",
		X"08",X"FE",X"05",X"28",X"68",X"CB",X"61",X"28",X"0B",X"3A",X"AF",X"42",X"FE",X"03",X"28",X"2E",
		X"CB",X"4F",X"20",X"20",X"DD",X"7E",X"09",X"D6",X"03",X"DD",X"77",X"09",X"30",X"D0",X"DD",X"36",
		X"09",X"80",X"DD",X"35",X"08",X"20",X"C7",X"DD",X"CB",X"01",X"96",X"CB",X"61",X"28",X"BF",X"CD",
		X"5B",X"33",X"18",X"BA",X"DD",X"7E",X"09",X"C6",X"04",X"DD",X"77",X"09",X"30",X"B0",X"DD",X"36",
		X"09",X"80",X"DD",X"34",X"08",X"21",X"CA",X"42",X"DD",X"7E",X"08",X"FE",X"05",X"20",X"04",X"CB",
		X"FE",X"18",X"9B",X"CB",X"F6",X"18",X"97",X"DD",X"34",X"09",X"20",X"92",X"DD",X"CB",X"00",X"C6",
		X"FD",X"35",X"06",X"AF",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"18",X"81",X"DD",X"34",X"09",
		X"DD",X"7E",X"09",X"FE",X"8D",X"C2",X"2E",X"34",X"DD",X"36",X"09",X"C8",X"DD",X"CB",X"01",X"DE",
		X"CB",X"61",X"28",X"03",X"CD",X"5B",X"33",X"23",X"E5",X"23",X"36",X"07",X"23",X"7E",X"CB",X"48",
		X"20",X"05",X"21",X"F5",X"34",X"18",X"03",X"21",X"01",X"35",X"06",X"04",X"BE",X"30",X"06",X"23",
		X"23",X"23",X"10",X"F8",X"76",X"23",X"5E",X"23",X"4E",X"E1",X"73",X"06",X"00",X"16",X"00",X"CD",
		X"CC",X"06",X"C3",X"2E",X"34",X"D0",X"32",X"05",X"A0",X"31",X"04",X"70",X"30",X"03",X"00",X"1B",
		X"02",X"D0",X"33",X"10",X"A0",X"32",X"05",X"70",X"31",X"04",X"00",X"30",X"03",X"3A",X"BF",X"42",
		X"B7",X"C0",X"C5",X"D5",X"E5",X"DD",X"E5",X"DD",X"46",X"05",X"DD",X"4E",X"04",X"C5",X"DD",X"E1",
		X"46",X"23",X"7E",X"E6",X"C0",X"4F",X"20",X"1B",X"78",X"FE",X"E0",X"28",X"64",X"3E",X"E0",X"32",
		X"C0",X"42",X"3E",X"10",X"32",X"C1",X"42",X"11",X"C0",X"FF",X"ED",X"53",X"C2",X"42",X"DD",X"7E",
		X"C0",X"18",X"19",X"78",X"FE",X"10",X"28",X"49",X"3E",X"10",X"32",X"C0",X"42",X"3E",X"F0",X"32",
		X"C1",X"42",X"11",X"40",X"00",X"ED",X"53",X"C2",X"42",X"DD",X"7E",X"40",X"FE",X"50",X"28",X"31",
		X"FE",X"4E",X"28",X"2D",X"CD",X"C9",X"28",X"E6",X"03",X"20",X"26",X"3E",X"15",X"B1",X"77",X"23",
		X"36",X"07",X"DD",X"22",X"C4",X"42",X"DD",X"E1",X"DD",X"CB",X"01",X"CE",X"DD",X"36",X"02",X"01",
		X"DD",X"36",X"08",X"02",X"DD",X"36",X"09",X"FF",X"DD",X"22",X"C6",X"42",X"3E",X"01",X"32",X"BF",
		X"42",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"3A",X"BF",X"42",X"B7",X"C8",X"3A",X"8E",X"42",X"E6",
		X"43",X"C0",X"DD",X"2A",X"C6",X"42",X"DD",X"35",X"09",X"C0",X"DD",X"36",X"09",X"78",X"DD",X"35",
		X"08",X"CA",X"5F",X"36",X"DD",X"66",X"07",X"DD",X"6E",X"06",X"46",X"23",X"23",X"23",X"4E",X"DD",
		X"21",X"60",X"42",X"3E",X"1D",X"57",X"3A",X"C1",X"42",X"FE",X"10",X"28",X"02",X"CB",X"FA",X"7A",
		X"32",X"C9",X"42",X"21",X"CB",X"42",X"CB",X"C6",X"AF",X"32",X"C8",X"42",X"ED",X"5B",X"C2",X"42",
		X"CD",X"EB",X"35",X"3A",X"C8",X"42",X"B7",X"C8",X"C3",X"84",X"0C",X"3A",X"C1",X"42",X"80",X"47",
		X"2A",X"C4",X"42",X"19",X"22",X"C4",X"42",X"3A",X"C9",X"42",X"DD",X"70",X"00",X"DD",X"77",X"01",
		X"DD",X"36",X"02",X"07",X"DD",X"71",X"03",X"3C",X"32",X"C9",X"42",X"CD",X"38",X"36",X"3A",X"C9",
		X"42",X"FE",X"20",X"C8",X"FE",X"A0",X"C8",X"3A",X"C0",X"42",X"B8",X"C8",X"19",X"CD",X"2B",X"36",
		X"D8",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"18",X"C0",X"7E",X"FE",X"50",X"28",X"06",
		X"FE",X"4E",X"28",X"02",X"A7",X"C9",X"37",X"C9",X"C5",X"E5",X"3A",X"5C",X"42",X"CD",X"55",X"36",
		X"30",X"10",X"3A",X"5F",X"42",X"41",X"CD",X"55",X"36",X"30",X"07",X"3A",X"C8",X"42",X"3C",X"32",
		X"C8",X"42",X"E1",X"C1",X"C9",X"B8",X"30",X"03",X"67",X"78",X"44",X"90",X"FE",X"09",X"C9",X"C5",
		X"E5",X"DD",X"E5",X"AF",X"32",X"BF",X"42",X"DD",X"2A",X"C6",X"42",X"DD",X"CB",X"01",X"8E",X"DD",
		X"36",X"08",X"00",X"DD",X"66",X"07",X"DD",X"6E",X"06",X"23",X"23",X"36",X"06",X"21",X"6B",X"42",
		X"06",X"0C",X"CD",X"69",X"0A",X"DD",X"E1",X"E1",X"C1",X"C9",X"3A",X"CA",X"42",X"CB",X"47",X"20",
		X"0C",X"3A",X"CC",X"42",X"CB",X"47",X"20",X"05",X"3A",X"8D",X"42",X"B7",X"C8",X"FD",X"21",X"CA",
		X"42",X"DD",X"21",X"D2",X"42",X"16",X"00",X"1E",X"00",X"FD",X"CB",X"00",X"3E",X"38",X"38",X"FD",
		X"CB",X"02",X"3E",X"38",X"1A",X"01",X"0E",X"00",X"DD",X"09",X"14",X"7A",X"FE",X"08",X"20",X"04",
		X"FD",X"23",X"18",X"E5",X"FE",X"10",X"20",X"E1",X"7B",X"FE",X"00",X"CC",X"97",X"37",X"C9",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"DD",X"35",X"04",X"28",X"14",X"01",X"06",X"00",X"A7",X"ED",X"42",
		X"06",X"0B",X"CD",X"C0",X"37",X"18",X"CE",X"FD",X"CB",X"02",X"3E",X"CD",X"8A",X"37",X"7E",X"FE",
		X"06",X"D2",X"7F",X"37",X"FE",X"00",X"20",X"08",X"23",X"7E",X"FE",X"00",X"28",X"B7",X"18",X"EB",
		X"FE",X"01",X"28",X"49",X"FE",X"02",X"20",X"30",X"23",X"7E",X"CB",X"BF",X"FE",X"00",X"28",X"3D",
		X"DD",X"4E",X"05",X"47",X"E6",X"0F",X"28",X"0A",X"78",X"E6",X"F0",X"28",X"0E",X"DD",X"70",X"05",
		X"18",X"2B",X"79",X"E6",X"0F",X"4F",X"78",X"E6",X"F0",X"18",X"07",X"79",X"E6",X"F0",X"4F",X"78",
		X"E6",X"0F",X"B1",X"DD",X"77",X"05",X"18",X"15",X"FE",X"03",X"20",X"14",X"23",X"7E",X"DD",X"77",
		X"0B",X"23",X"7E",X"DD",X"77",X"0C",X"23",X"7E",X"E6",X"0F",X"DD",X"77",X"0D",X"23",X"18",X"9E",
		X"FE",X"04",X"20",X"17",X"23",X"7E",X"E6",X"1F",X"DD",X"77",X"08",X"23",X"7E",X"E6",X"1F",X"DD",
		X"77",X"09",X"23",X"7E",X"E6",X"1F",X"DD",X"77",X"0A",X"18",X"E2",X"23",X"7E",X"E6",X"1F",X"DD",
		X"77",X"06",X"23",X"7E",X"E6",X"3F",X"CB",X"FF",X"CB",X"F7",X"DD",X"77",X"07",X"18",X"CE",X"06",
		X"0E",X"CD",X"C0",X"37",X"CD",X"FF",X"37",X"C3",X"B5",X"36",X"DD",X"6E",X"00",X"DD",X"75",X"02",
		X"DD",X"66",X"01",X"DD",X"74",X"03",X"C9",X"0E",X"08",X"AF",X"CD",X"A4",X"37",X"0C",X"CD",X"A4",
		X"37",X"0C",X"18",X"00",X"F5",X"C5",X"32",X"00",X"48",X"32",X"00",X"4A",X"06",X"49",X"02",X"32",
		X"03",X"48",X"32",X"00",X"48",X"4F",X"02",X"32",X"01",X"48",X"32",X"00",X"48",X"C1",X"F1",X"C9",
		X"7B",X"FE",X"00",X"20",X"2B",X"1C",X"0E",X"00",X"7E",X"CD",X"A4",X"37",X"23",X"0C",X"79",X"FE",
		X"06",X"20",X"F5",X"DD",X"75",X"02",X"DD",X"74",X"03",X"DD",X"E5",X"E1",X"D5",X"11",X"06",X"00",
		X"19",X"D1",X"0E",X"06",X"7E",X"CD",X"A4",X"37",X"0C",X"23",X"79",X"B8",X"20",X"F6",X"18",X"0A",
		X"01",X"06",X"00",X"09",X"DD",X"75",X"02",X"DD",X"74",X"03",X"FD",X"CB",X"02",X"FE",X"C9",X"E5",
		X"DD",X"7E",X"05",X"E6",X"0F",X"21",X"24",X"38",X"06",X"00",X"4F",X"09",X"7E",X"47",X"DD",X"4E",
		X"05",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"0D",X"28",X"04",X"80",X"0D",X"20",X"FC",
		X"DD",X"77",X"04",X"E1",X"C9",X"01",X"02",X"03",X"04",X"06",X"08",X"0C",X"10",X"18",X"20",X"06",
		X"06",X"06",X"06",X"06",X"06",X"00",X"10",X"00",X"10",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",
		X"00",X"05",X"04",X"80",X"10",X"80",X"10",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",
		X"04",X"00",X"11",X"00",X"11",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"80",
		X"11",X"80",X"11",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"12",X"00",
		X"12",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"13",X"00",X"13",X"00",
		X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"14",X"00",X"14",X"00",X"46",X"04",
		X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"15",X"00",X"15",X"00",X"46",X"04",X"B8",X"05",
		X"05",X"05",X"00",X"05",X"04",X"00",X"16",X"00",X"16",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",
		X"00",X"05",X"04",X"80",X"16",X"80",X"16",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",
		X"04",X"E0",X"17",X"E0",X"17",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",
		X"18",X"00",X"18",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"19",X"00",
		X"19",X"00",X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"80",X"1B",X"80",X"1B",X"00",
		X"46",X"04",X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"1C",X"00",X"1C",X"00",X"46",X"04",
		X"B8",X"05",X"05",X"05",X"00",X"05",X"04",X"00",X"1E",X"00",X"1E",X"00",X"46",X"04",X"B8",X"05",
		X"05",X"05",X"00",X"05",X"04",X"CC",X"50",X"18",X"53",X"9A",X"50",X"C8",X"52",X"58",X"42",X"A0",
		X"70",X"6E",X"51",X"78",X"42",X"40",X"A0",X"F4",X"52",X"7C",X"42",X"30",X"40",X"28",X"53",X"58",
		X"42",X"C0",X"60",X"EC",X"50",X"78",X"42",X"90",X"B0",X"B6",X"51",X"7C",X"42",X"40",X"80",X"F0",
		X"52",X"09",X"16",X"04",X"07",X"3C",X"04",X"E8",X"50",X"00",X"40",X"42",X"C0",X"40",X"12",X"F6",
		X"50",X"01",X"44",X"42",X"C0",X"B0",X"80",X"7A",X"52",X"00",X"48",X"42",X"60",X"D0",X"10",X"2E",
		X"53",X"00",X"4C",X"42",X"30",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"09",X"16",X"04",X"07",X"37",X"04",X"AC",X"51",X"01",X"40",X"42",X"90",X"60",X"82",X"38",
		X"51",X"01",X"44",X"42",X"B0",X"C0",X"40",X"F8",X"52",X"00",X"48",X"42",X"40",X"C0",X"12",X"2A",
		X"53",X"00",X"4C",X"42",X"30",X"50",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"11",X"04",X"07",X"32",X"05",X"68",X"51",X"00",X"40",X"42",X"A0",X"40",X"20",X"78",
		X"51",X"01",X"44",X"42",X"A0",X"C0",X"80",X"78",X"52",X"00",X"48",X"42",X"60",X"C0",X"12",X"6C",
		X"52",X"01",X"4C",X"42",X"60",X"60",X"42",X"32",X"53",X"00",X"50",X"42",X"30",X"90",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"07",X"11",X"04",X"07",X"2D",X"05",X"A8",X"51",X"01",X"40",X"42",X"90",X"40",X"82",X"6E",
		X"51",X"00",X"44",X"42",X"A0",X"70",X"20",X"FA",X"51",X"00",X"48",X"42",X"80",X"D0",X"12",X"38",
		X"53",X"01",X"4C",X"42",X"30",X"C0",X"40",X"AA",X"52",X"00",X"50",X"42",X"50",X"50",X"12",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"04",X"07",X"1E",X"06",X"A6",X"51",X"00",X"40",X"42",X"90",X"30",X"12",X"34",
		X"51",X"01",X"44",X"42",X"B0",X"A0",X"80",X"F4",X"51",X"00",X"48",X"42",X"80",X"A0",X"22",X"AA",
		X"52",X"01",X"4C",X"42",X"50",X"50",X"40",X"F0",X"52",X"00",X"50",X"42",X"40",X"80",X"12",X"BA",
		X"52",X"01",X"54",X"42",X"50",X"D0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"06",X"0E",X"04",X"07",X"0F",X"06",X"68",X"51",X"00",X"40",X"42",X"A0",X"40",X"10",X"EE",
		X"51",X"01",X"44",X"42",X"80",X"70",X"82",X"30",X"51",X"00",X"48",X"42",X"B0",X"80",X"22",X"38",
		X"52",X"01",X"4C",X"42",X"70",X"C0",X"40",X"A8",X"52",X"01",X"50",X"42",X"50",X"40",X"42",X"34",
		X"53",X"00",X"54",X"42",X"30",X"A0",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"04",X"07",X"01",X"06",X"6C",X"51",X"00",X"40",X"42",X"A0",X"60",X"10",X"72",
		X"51",X"00",X"44",X"42",X"A0",X"90",X"22",X"F6",X"51",X"01",X"48",X"42",X"80",X"B0",X"82",X"68",
		X"52",X"01",X"4C",X"42",X"60",X"40",X"42",X"AE",X"52",X"00",X"50",X"42",X"50",X"70",X"12",X"B8",
		X"52",X"00",X"54",X"42",X"50",X"C0",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"06",X"0E",X"04",X"07",X"01",X"06",X"E8",X"51",X"01",X"40",X"42",X"80",X"40",X"42",X"70",
		X"51",X"01",X"44",X"42",X"A0",X"80",X"82",X"36",X"51",X"00",X"48",X"42",X"B0",X"B0",X"22",X"6C",
		X"52",X"01",X"4C",X"42",X"60",X"60",X"42",X"F4",X"52",X"00",X"50",X"42",X"40",X"A0",X"12",X"76",
		X"52",X"01",X"54",X"42",X"60",X"B0",X"82",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
