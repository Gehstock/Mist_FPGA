`define BUILD_DATE "190827"
`define BUILD_TIME "181730"
