library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"10",X"10",X"1C",X"1E",X"7E",X"7E",X"1F",X"7F",X"FE",X"FE",X"FE",X"FC",X"D0",X"10",X"00",
		X"00",X"00",X"06",X"1E",X"9E",X"9E",X"9E",X"1E",X"1E",X"0E",X"5E",X"5E",X"5E",X"06",X"00",X"00",
		X"00",X"10",X"10",X"7C",X"7E",X"1E",X"1E",X"7F",X"FF",X"FE",X"FE",X"FE",X"FC",X"D0",X"10",X"00",
		X"00",X"00",X"06",X"1E",X"5E",X"5E",X"5E",X"1E",X"1E",X"0E",X"9E",X"9E",X"9E",X"06",X"00",X"00",
		X"00",X"10",X"10",X"1C",X"DE",X"DE",X"1E",X"1F",X"DF",X"DE",X"1E",X"1E",X"FC",X"10",X"10",X"00",
		X"00",X"00",X"06",X"5E",X"5C",X"5C",X"18",X"1C",X"1C",X"9C",X"9E",X"9E",X"1E",X"06",X"00",X"00",
		X"00",X"10",X"10",X"1C",X"9E",X"9E",X"1E",X"1F",X"9F",X"9E",X"1E",X"1E",X"FC",X"10",X"10",X"00",
		X"00",X"00",X"06",X"9E",X"9D",X"9D",X"18",X"1C",X"1D",X"5D",X"5E",X"5E",X"1E",X"06",X"00",X"00",
		X"00",X"00",X"18",X"7E",X"7E",X"1F",X"7F",X"FE",X"FE",X"FE",X"FC",X"D0",X"10",X"00",X"00",X"00",
		X"00",X"1E",X"9E",X"9E",X"9E",X"1E",X"1E",X"0E",X"5E",X"5E",X"5E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"3E",X"7F",X"7F",X"7F",X"7F",X"7E",X"68",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2F",X"2F",X"0F",X"0F",X"07",X"4F",X"4F",X"4F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"98",X"BE",X"BF",X"BF",X"BF",X"B4",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"03",X"17",X"17",X"17",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"D8",X"DE",X"DF",X"DA",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"13",X"13",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C2",X"C3",X"B2",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"13",X"13",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"84",X"87",X"37",X"37",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"17",X"17",X"17",X"06",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0E",X"CF",X"CF",X"0F",X"0F",X"CE",X"C8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"4F",X"4E",X"4E",X"0C",X"0E",X"0E",X"2E",X"2F",X"00",
		X"00",X"00",X"00",X"10",X"10",X"1C",X"DE",X"DE",X"1E",X"1F",X"DF",X"DE",X"1E",X"18",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"06",X"5E",X"5C",X"5C",X"18",X"1C",X"1C",X"9C",X"9E",X"9E",X"1E",X"00",
		X"00",X"00",X"E1",X"79",X"78",X"38",X"38",X"38",X"18",X"38",X"B8",X"F8",X"79",X"E1",X"00",X"00",
		X"20",X"A0",X"50",X"58",X"B0",X"76",X"36",X"B0",X"70",X"B0",X"31",X"71",X"B0",X"50",X"50",X"88",
		X"00",X"00",X"C0",X"F0",X"F1",X"71",X"71",X"30",X"70",X"71",X"71",X"F1",X"F0",X"C0",X"00",X"00",
		X"40",X"20",X"A1",X"60",X"63",X"63",X"60",X"E0",X"60",X"6C",X"EC",X"60",X"B0",X"21",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"A4",X"B0",X"FC",X"DD",X"FE",X"DE",X"FE",X"FF",X"FE",X"FD",X"F8",X"EA",X"D0",
		X"00",X"10",X"90",X"1D",X"DF",X"DF",X"1F",X"1F",X"DF",X"DF",X"1F",X"1F",X"FF",X"93",X"13",X"00",
		X"00",X"00",X"07",X"1E",X"9C",X"9C",X"98",X"1C",X"1C",X"9C",X"9E",X"9E",X"1E",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"40",X"E0",X"30",X"30",X"30",X"B0",X"70",X"30",X"20",X"60",X"C0",X"00",X"00",
		X"00",X"0D",X"9B",X"7E",X"7C",X"FB",X"F5",X"FA",X"FD",X"FE",X"FE",X"7D",X"FC",X"BC",X"0B",X"00",
		X"00",X"00",X"07",X"1E",X"9C",X"9C",X"98",X"1C",X"1C",X"9C",X"9E",X"9E",X"1E",X"07",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"00",X"00",
		X"00",X"07",X"25",X"0D",X"3F",X"BB",X"7F",X"7B",X"7F",X"FF",X"7F",X"BF",X"1F",X"57",X"0B",X"00",
		X"00",X"A0",X"78",X"C8",X"9C",X"66",X"A6",X"46",X"B6",X"CE",X"C6",X"A4",X"8C",X"98",X"60",X"00",
		X"00",X"01",X"03",X"0F",X"0F",X"1F",X"1E",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"07",X"01",X"00",
		X"00",X"00",X"81",X"00",X"80",X"20",X"00",X"80",X"20",X"00",X"00",X"00",X"81",X"80",X"00",X"00",
		X"00",X"00",X"00",X"1B",X"36",X"14",X"48",X"B0",X"C4",X"28",X"24",X"32",X"0B",X"04",X"00",X"00",
		X"58",X"0E",X"21",X"09",X"1A",X"20",X"00",X"00",X"00",X"00",X"28",X"04",X"06",X"21",X"02",X"18",
		X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"04",X"88",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A4",X"40",X"82",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"01",X"10",X"04",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"02",X"42",X"A6",X"8B",X"D3",X"EE",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"06",X"02",X"00",X"01",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"90",X"48",X"68",X"60",X"A0",X"28",
		X"00",X"F0",X"7C",X"8E",X"3E",X"42",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0C",X"08",X"11",X"12",X"24",X"29",X"31",X"2A",X"26",X"06",X"0A",X"32",X"2A",X"26",
		X"00",X"F0",X"7C",X"8E",X"3E",X"42",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0C",X"08",X"11",X"12",X"24",X"09",X"11",X"2A",X"26",X"26",X"2A",X"32",X"2A",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"2A",X"32",X"0A",X"06",X"26",X"2A",X"32",X"32",X"2A",X"26",X"06",X"0A",X"32",X"2A",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"2A",X"32",X"2A",X"26",X"26",X"2A",X"12",X"12",X"2A",X"26",X"26",X"2A",X"32",X"2A",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"1F",X"FF",X"1F",X"07",X"03",X"03",X"01",X"01",X"01",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"01",X"01",X"01",X"03",X"03",X"07",X"1F",X"FF",X"FF",X"1F",X"07",X"03",X"03",X"01",X"01",X"01",
		X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"00",X"00",X"0C",X"02",X"01",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"E0",X"F8",X"FF",X"FF",X"F8",X"E0",X"C0",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",
		X"00",X"80",X"98",X"B8",X"B9",X"B3",X"A0",X"B0",X"B3",X"B1",X"B8",X"B8",X"BB",X"98",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"00",X"00",X"0C",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1E",X"3E",X"7E",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"B0",X"70",X"F8",X"78",X"78",X"38",
		X"1C",X"1E",X"1E",X"1F",X"0E",X"0D",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FE",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"9C",X"38",X"C0",X"40",X"20",X"A0",X"A0",X"20",X"40",X"C0",X"38",X"9C",X"80",X"00",
		X"3F",X"FF",X"07",X"03",X"00",X"01",X"19",X"3B",X"3B",X"19",X"01",X"00",X"03",X"07",X"FF",X"3F",
		X"F0",X"FC",X"F0",X"C0",X"B8",X"70",X"80",X"80",X"80",X"80",X"70",X"B8",X"C0",X"F0",X"FC",X"F0",
		X"0F",X"67",X"13",X"01",X"0B",X"B3",X"63",X"67",X"67",X"63",X"B3",X"0B",X"01",X"13",X"67",X"0F",
		X"C0",X"E0",X"E7",X"CE",X"30",X"50",X"48",X"E8",X"E8",X"48",X"50",X"30",X"CE",X"E7",X"E0",X"C0",
		X"0F",X"3F",X"01",X"00",X"00",X"00",X"06",X"0E",X"0E",X"06",X"00",X"00",X"00",X"01",X"3F",X"0F",
		X"FC",X"FF",X"FC",X"70",X"EE",X"DC",X"E0",X"E0",X"E0",X"E0",X"DC",X"EE",X"70",X"FC",X"FF",X"FC",
		X"03",X"19",X"04",X"00",X"02",X"2C",X"18",X"19",X"19",X"18",X"2C",X"02",X"00",X"04",X"19",X"03",
		X"00",X"00",X"00",X"00",X"04",X"02",X"82",X"96",X"6E",X"FE",X"92",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"80",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"04",
		X"00",X"00",X"00",X"04",X"06",X"03",X"87",X"CF",X"7B",X"D2",X"84",X"00",X"00",X"00",X"00",X"00",
		X"04",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",
		X"00",X"10",X"08",X"08",X"78",X"9C",X"10",X"44",X"10",X"9C",X"7C",X"18",X"30",X"20",X"60",X"00",
		X"04",X"10",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"80",X"00",X"80",X"00",X"00",
		X"00",X"60",X"20",X"30",X"7C",X"CE",X"88",X"A2",X"88",X"CE",X"7C",X"18",X"08",X"08",X"10",X"00",
		X"00",X"00",X"80",X"00",X"80",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"10",X"04",
		X"0A",X"00",X"08",X"00",X"00",X"80",X"80",X"00",X"80",X"80",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"06",X"04",X"0C",X"7E",X"C7",X"4B",X"1B",X"4B",X"C7",X"7E",X"18",X"10",X"10",X"20",X"00",
		X"00",X"00",X"00",X"01",X"00",X"01",X"80",X"80",X"00",X"80",X"80",X"00",X"00",X"08",X"00",X"0A",
		X"00",X"20",X"10",X"10",X"18",X"7E",X"C7",X"4B",X"1B",X"4B",X"C7",X"7E",X"0C",X"04",X"06",X"00",
		X"00",X"00",X"08",X"04",X"04",X"2C",X"DC",X"FC",X"24",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"02",X"03",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"20",X"08",X"00",X"00",
		X"00",X"00",X"80",X"CE",X"7B",X"D2",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"30",X"7E",X"49",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"08",X"0C",X"1E",X"70",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"04",X"3C",X"CE",X"88",X"20",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"20",X"30",X"7C",X"CE",X"88",X"A2",X"88",X"C8",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"01",X"01",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"20",X"10",X"10",X"F0",X"38",X"20",X"88",X"20",X"38",X"F8",X"30",X"40",X"00",
		X"00",X"00",X"08",X"20",X"00",X"00",X"00",X"03",X"02",X"00",X"02",X"03",X"00",X"80",X"00",X"00",
		X"80",X"A0",X"00",X"40",X"80",X"10",X"04",X"00",X"00",X"C0",X"20",X"30",X"20",X"80",X"00",X"80",
		X"01",X"0F",X"03",X"6E",X"3E",X"7F",X"5D",X"5C",X"45",X"76",X"5F",X"4C",X"0F",X"0B",X"15",X"0B",
		X"00",X"00",X"00",X"60",X"C4",X"A0",X"80",X"20",X"80",X"60",X"E0",X"C0",X"80",X"10",X"40",X"80",
		X"04",X"2E",X"43",X"08",X"03",X"04",X"80",X"12",X"18",X"DC",X"62",X"D6",X"45",X"88",X"08",X"14",
		X"00",X"C0",X"40",X"60",X"F8",X"9C",X"10",X"44",X"10",X"9C",X"F8",X"30",X"10",X"10",X"20",X"00",
		X"00",X"20",X"40",X"48",X"D0",X"03",X"B3",X"09",X"03",X"93",X"58",X"D0",X"48",X"A8",X"20",X"10",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"80",X"60",X"80",X"20",X"30",X"10",X"10",X"00",X"00",X"10",X"10",X"A0",X"60",X"00",X"E0",X"80",
		X"0F",X"05",X"03",X"0F",X"2C",X"5F",X"56",X"44",X"56",X"5F",X"7F",X"2E",X"2E",X"03",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"58",X"E0",X"C8",X"0C",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"03",X"0B",X"17",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"18",X"40",X"90",X"20",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"18",X"1B",X"33",X"3E",X"36",X"34",X"00",
		X"00",X"00",X"00",X"00",X"80",X"60",X"80",X"20",X"30",X"10",X"10",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"05",X"03",X"0F",X"2C",X"5F",X"56",X"44",X"56",X"5F",X"7F",X"00",
		X"00",X"00",X"00",X"80",X"60",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"3C",X"61",X"6E",X"CC",X"F9",X"D9",X"D0",X"C4",X"D4",X"DA",X"68",X"00",
		X"80",X"60",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"20",X"40",X"80",X"C0",X"E0",X"C0",X"80",
		X"0F",X"1C",X"20",X"66",X"68",X"DA",X"D4",X"C4",X"D0",X"D9",X"F9",X"ED",X"6F",X"77",X"3F",X"0F",
		X"80",X"60",X"00",X"40",X"80",X"00",X"20",X"00",X"00",X"00",X"10",X"80",X"E0",X"60",X"E0",X"80",
		X"0F",X"3C",X"61",X"6E",X"CC",X"F9",X"D9",X"D0",X"C4",X"D4",X"DB",X"6F",X"67",X"3E",X"1C",X"0F",
		X"00",X"30",X"00",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"30",X"00",
		X"06",X"12",X"30",X"30",X"02",X"04",X"0C",X"08",X"62",X"62",X"48",X"34",X"33",X"10",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"12",X"10",X"10",X"00",X"00",X"00",X"00",X"40",X"60",X"40",X"20",X"01",X"00",X"08",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"04",X"20",X"20",X"00",X"00",X"04",X"30",X"80",X"C0",X"80",X"40",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"04",X"07",X"04",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"18",X"38",X"18",X"38",X"18",X"1C",X"1E",X"0F",X"1F",X"08",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"07",X"04",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"08",X"18",X"08",X"18",X"18",X"1C",X"3E",X"1F",X"3F",X"18",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"64",X"07",X"04",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"08",X"18",X"08",X"1A",X"18",X"1C",X"3E",X"1F",X"3F",X"18",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"67",X"04",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"18",X"38",X"18",X"3A",X"18",X"1C",X"1E",X"0F",X"1F",X"08",X"10",X"00",X"00",
		X"00",X"00",X"0C",X"18",X"FC",X"F8",X"3C",X"18",X"58",X"18",X"18",X"3C",X"28",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"20",X"E8",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"18",X"1C",X"38",X"7C",X"18",X"1D",X"0D",X"06",X"27",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"21",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"07",X"04",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"38",X"18",X"38",X"18",X"1C",X"1E",X"0F",X"1F",X"08",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"02",X"00",X"C0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0C",X"0C",X"0E",X"1F",X"0F",X"1F",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"07",X"07",X"03",X"07",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"03",X"07",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"07",X"03",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"98",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"06",X"02",X"06",X"06",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"33",X"02",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"0C",X"1C",X"0C",X"1D",X"0C",X"0E",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"64",X"07",X"04",X"00",X"80",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"08",X"18",X"08",X"1A",X"18",X"1C",X"3E",X"1F",X"3F",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"9C",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"10",X"00",X"00",X"01",X"01",X"00",X"00",X"10",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"67",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"12",X"0C",X"02",X"04",X"04",X"00",X"00",X"08",X"0A",X"04",X"0E",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"64",X"07",X"04",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"18",X"1C",X"08",X"0A",X"10",X"0C",X"06",X"0F",X"0F",X"18",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"67",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"CE",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"73",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"14",X"74",X"13",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"19",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"50",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"FC",X"FE",X"E0",X"C0",X"80",X"80",X"00",X"80",X"C0",X"E0",X"FE",X"FC",X"E0",X"00",X"00",
		X"3F",X"FF",X"07",X"0F",X"07",X"03",X"03",X"00",X"03",X"07",X"0F",X"07",X"FF",X"3F",X"00",X"00",
		X"00",X"E0",X"FC",X"E2",X"C0",X"80",X"80",X"00",X"80",X"C0",X"E2",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"3F",X"FF",X"0F",X"07",X"03",X"03",X"00",X"03",X"07",X"0F",X"FF",X"3F",X"00",X"00",X"00",
		X"60",X"7C",X"BE",X"A0",X"00",X"04",X"10",X"10",X"04",X"00",X"A0",X"7E",X"FC",X"E0",X"00",X"00",
		X"3F",X"FF",X"07",X"0F",X"07",X"00",X"00",X"00",X"00",X"07",X"0F",X"07",X"FC",X"3F",X"00",X"00",
		X"00",X"E0",X"7C",X"A2",X"00",X"04",X"10",X"10",X"04",X"00",X"A2",X"BC",X"60",X"00",X"00",X"00",
		X"00",X"3F",X"FC",X"0F",X"07",X"00",X"00",X"00",X"00",X"07",X"0F",X"FF",X"3F",X"00",X"00",X"00",
		X"F8",X"FE",X"E0",X"40",X"E0",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"60",X"B9",X"5C",X"00",
		X"00",X"0D",X"1C",X"3F",X"60",X"00",X"00",X"10",X"04",X"04",X"10",X"00",X"06",X"70",X"0F",X"00",
		X"00",X"5C",X"BB",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"40",X"E0",X"FE",X"F8",
		X"00",X"0F",X"73",X"01",X"00",X"10",X"04",X"04",X"10",X"00",X"00",X"60",X"3F",X"1C",X"0D",X"00",
		X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"C0",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"0F",X"07",X"07",X"00",X"07",X"0F",X"1F",X"0F",X"FF",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"00",X"80",X"C0",X"E2",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"00",X"03",X"07",X"0F",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"F0",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"03",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"1F",X"E8",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"3F",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"BE",X"DE",X"D0",X"80",X"02",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"7C",X"A2",X"00",X"04",X"10",X"10",X"04",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"FC",X"0F",X"07",X"00",X"00",X"00",X"00",X"07",X"0F",X"00",
		X"00",X"00",X"C0",X"F8",X"7C",X"40",X"00",X"08",X"20",X"20",X"08",X"00",X"40",X"F8",X"C0",X"00",
		X"00",X"00",X"7E",X"FE",X"0F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"0E",X"1F",X"0E",X"F9",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"10",X"10",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"00",X"00",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"F8",X"BC",X"02",X"04",X"10",X"10",X"06",X"FE",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"7F",X"CF",X"07",X"00",X"00",X"00",X"00",X"FF",X"7F",X"1F",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
