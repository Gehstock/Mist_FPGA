library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gravitar_pgm_rom6 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gravitar_pgm_rom6 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"00",X"00",X"A0",X"01",X"FE",X"08",X"A0",X"01",X"FE",X"04",X"98",X"10",X"04",X"10",X"00",
		X"00",X"82",X"02",X"01",X"04",X"8C",X"08",X"FF",X"03",X"80",X"04",X"00",X"01",X"8C",X"20",X"FF",
		X"01",X"86",X"40",X"FF",X"01",X"82",X"40",X"FF",X"01",X"81",X"40",X"FF",X"01",X"00",X"00",X"C0",
		X"10",X"04",X"10",X"00",X"00",X"86",X"50",X"FE",X"03",X"00",X"00",X"98",X"07",X"00",X"01",X"00",
		X"00",X"84",X"07",X"00",X"01",X"00",X"00",X"A1",X"11",X"01",X"03",X"A3",X"11",X"FF",X"01",X"66",
		X"00",X"FF",X"08",X"00",X"05",X"6B",X"00",X"A1",X"08",X"01",X"03",X"A3",X"08",X"FF",X"01",X"6E",
		X"00",X"FF",X"08",X"00",X"05",X"73",X"00",X"A2",X"10",X"00",X"16",X"00",X"00",X"F6",X"10",X"F7",
		X"0A",X"93",X"10",X"09",X"0B",X"00",X"00",X"A7",X"A1",X"00",X"03",X"00",X"00",X"FF",X"A1",X"00",
		X"03",X"00",X"00",X"A7",X"A1",X"00",X"03",X"00",X"00",X"FD",X"A1",X"00",X"03",X"00",X"00",X"A4",
		X"11",X"00",X"05",X"8A",X"00",X"FF",X"11",X"F8",X"05",X"8D",X"00",X"A4",X"11",X"00",X"05",X"90",
		X"00",X"FE",X"11",X"F8",X"05",X"93",X"00",X"F6",X"08",X"F7",X"0A",X"93",X"08",X"09",X"0B",X"96",
		X"00",X"A2",X"08",X"00",X"15",X"9B",X"00",X"80",X"08",X"F8",X"03",X"70",X"08",X"F8",X"03",X"60",
		X"08",X"F8",X"03",X"50",X"08",X"F8",X"03",X"40",X"08",X"F8",X"03",X"00",X"00",X"A4",X"08",X"00",
		X"14",X"00",X"00",X"A9",X"8F",X"D0",X"38",X"A9",X"BF",X"D0",X"34",X"A9",X"0F",X"D0",X"30",X"A9",
		X"1F",X"D0",X"2C",X"A9",X"2F",X"D0",X"28",X"A9",X"5F",X"D0",X"24",X"A9",X"6F",X"D0",X"20",X"A9",
		X"7F",X"D0",X"1C",X"A9",X"3F",X"D0",X"18",X"A9",X"4F",X"D0",X"14",X"A9",X"9F",X"D0",X"10",X"A9",
		X"AF",X"D0",X"11",X"A9",X"CF",X"D0",X"08",X"A9",X"DF",X"D0",X"04",X"A9",X"EF",X"D0",X"00",X"24",
		X"D0",X"D0",X"01",X"60",X"86",X"25",X"84",X"26",X"A8",X"A2",X"0F",X"B9",X"8D",X"DE",X"F0",X"0E",
		X"86",X"8C",X"95",X"8E",X"A9",X"01",X"95",X"AE",X"95",X"BE",X"A9",X"FF",X"85",X"8C",X"88",X"CA",
		X"10",X"E9",X"A6",X"25",X"A4",X"26",X"60",X"A2",X"0F",X"B5",X"8E",X"F0",X"7E",X"E4",X"8C",X"F0",
		X"7A",X"D6",X"AE",X"D0",X"76",X"D6",X"BE",X"D0",X"38",X"F6",X"8E",X"F6",X"8E",X"B5",X"8E",X"0A",
		X"A8",X"B0",X"10",X"B9",X"77",X"DF",X"95",X"9E",X"B9",X"7A",X"DF",X"95",X"BE",X"B9",X"78",X"DF",
		X"4C",X"70",X"E1",X"B9",X"77",X"E0",X"95",X"9E",X"B9",X"7A",X"E0",X"95",X"BE",X"B9",X"78",X"E0",
		X"95",X"AE",X"D0",X"0A",X"95",X"8E",X"B5",X"9E",X"F0",X"04",X"95",X"8E",X"D0",X"CB",X"4C",X"AC",
		X"E1",X"0A",X"A8",X"B0",X"0B",X"B9",X"78",X"DF",X"95",X"AE",X"B9",X"79",X"DF",X"4C",X"98",X"E1",
		X"B9",X"78",X"E0",X"95",X"AE",X"B9",X"79",X"E0",X"B4",X"9E",X"18",X"75",X"9E",X"95",X"9E",X"8A",
		X"4A",X"90",X"09",X"98",X"55",X"9E",X"29",X"F0",X"55",X"9E",X"95",X"9E",X"B5",X"9E",X"E0",X"08",
		X"90",X"06",X"9D",X"F8",X"67",X"4C",X"BB",X"E1",X"9D",X"00",X"60",X"CA",X"30",X"03",X"4C",X"39",
		X"E1",X"60",X"A9",X"00",X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"A9",X"07",X"8D",X"0F",X"60",X"8D",
		X"0F",X"68",X"A2",X"0F",X"A9",X"00",X"9D",X"00",X"60",X"9D",X"00",X"68",X"95",X"8E",X"95",X"9E",
		X"CA",X"10",X"F3",X"A9",X"00",X"8D",X"08",X"60",X"A2",X"00",X"8E",X"08",X"68",X"60",X"48",X"8A",
		X"48",X"20",X"66",X"E4",X"68",X"AA",X"68",X"A0",X"00",X"4C",X"8A",X"E4",X"84",X"22",X"A9",X"00",
		X"A0",X"03",X"20",X"5F",X"E4",X"A4",X"22",X"A9",X"00",X"0A",X"0A",X"C0",X"1D",X"90",X"0A",X"69",
		X"01",X"AA",X"98",X"38",X"E9",X"1D",X"A8",X"10",X"01",X"AA",X"BD",X"7B",X"E2",X"85",X"20",X"BD",
		X"7A",X"E2",X"85",X"1F",X"18",X"71",X"1F",X"85",X"1F",X"90",X"02",X"E6",X"20",X"A0",X"00",X"A2",
		X"00",X"A1",X"1F",X"85",X"22",X"4A",X"4A",X"20",X"56",X"E2",X"A1",X"1F",X"2A",X"26",X"22",X"2A",
		X"A5",X"22",X"2A",X"0A",X"20",X"5C",X"E2",X"A1",X"1F",X"85",X"22",X"20",X"56",X"E2",X"46",X"22",
		X"90",X"DF",X"88",X"4C",X"72",X"E4",X"E6",X"1F",X"D0",X"02",X"E6",X"20",X"29",X"3E",X"D0",X"04",
		X"68",X"68",X"D0",X"EE",X"C9",X"0A",X"90",X"02",X"69",X"0D",X"AA",X"BD",X"46",X"4D",X"91",X"08",
		X"C8",X"BD",X"47",X"4D",X"91",X"08",X"C8",X"A2",X"00",X"60",X"7E",X"E2",X"71",X"E3",X"1D",X"25",
		X"2B",X"33",X"37",X"3B",X"3F",X"47",X"4B",X"57",X"61",X"65",X"6F",X"79",X"87",X"95",X"A1",X"AD",
		X"AD",X"B1",X"B5",X"BB",X"BF",X"C5",X"CD",X"D7",X"E1",X"E5",X"EB",X"A5",X"92",X"BD",X"C2",X"BE",
		X"0A",X"B6",X"00",X"59",X"62",X"48",X"66",X"D2",X"6D",X"9E",X"70",X"0C",X"D4",X"0A",X"B2",X"4C",
		X"00",X"B9",X"E6",X"B2",X"40",X"56",X"52",X"80",X"00",X"83",X"74",X"4D",X"C0",X"4D",X"CE",X"2D",
		X"12",X"0E",X"1A",X"8A",X"40",X"83",X"64",X"78",X"00",X"8B",X"6E",X"BB",X"66",X"90",X"4E",X"9C",
		X"68",X"82",X"70",X"48",X"00",X"BB",X"26",X"9E",X"02",X"B2",X"4A",X"3E",X"26",X"B0",X"00",X"34",
		X"E4",X"CD",X"C0",X"83",X"64",X"78",X"4A",X"3E",X"1A",X"D1",X"70",X"4A",X"00",X"3C",X"E4",X"5D",
		X"8A",X"C6",X"60",X"2E",X"1A",X"9C",X"AF",X"4C",X"B0",X"4D",X"82",X"EC",X"F2",X"B0",X"5A",X"93",
		X"70",X"69",X"60",X"B8",X"00",X"A5",X"92",X"BD",X"C2",X"B4",X"F0",X"2E",X"12",X"09",X"B2",X"C6",
		X"26",X"95",X"C0",X"C4",X"C2",X"3B",X"0A",X"92",X"D2",X"0C",X"12",X"C6",X"12",X"B5",X"C0",X"C5",
		X"8A",X"3E",X"26",X"B0",X"70",X"98",X"6E",X"4C",X"12",X"3E",X"00",X"54",X"32",X"93",X"FB",X"5E",
		X"64",X"92",X"6D",X"3C",X"C2",X"A3",X"60",X"9E",X"00",X"A3",X"60",X"9E",X"00",X"29",X"D2",X"0D",
		X"1A",X"84",X"F1",X"7B",X"60",X"82",X"6C",X"0D",X"1A",X"84",X"F1",X"A4",X"E4",X"C3",X"72",X"B8",
		X"68",X"6C",X"0A",X"C2",X"40",X"5C",X"F0",X"C1",X"42",X"32",X"42",X"86",X"4E",X"7F",X"40",X"0C",
		X"1A",X"BE",X"00",X"A4",X"0A",X"EA",X"6C",X"08",X"00",X"6C",X"AE",X"4D",X"B0",X"09",X"E6",X"6C",
		X"80",X"10",X"1A",X"24",X"2A",X"2E",X"38",X"40",X"48",X"4E",X"58",X"62",X"68",X"6E",X"7E",X"86",
		X"8E",X"18",X"4E",X"9B",X"64",X"08",X"C2",X"A4",X"0A",X"E8",X"00",X"2E",X"0A",X"B3",X"42",X"89",
		X"E2",X"87",X"38",X"E3",X"5B",X"3D",X"92",X"43",X"70",X"B8",X"40",X"41",X"64",X"5A",X"6D",X"BB",
		X"26",X"9E",X"02",X"36",X"64",X"7A",X"6C",X"B8",X"00",X"C5",X"8A",X"3E",X"26",X"B0",X"54",X"CA",
		X"61",X"BE",X"68",X"4D",X"82",X"34",X"E4",X"CD",X"C0",X"92",X"78",X"C0",X"6E",X"63",X"69",X"18",
		X"4E",X"9B",X"64",X"09",X"02",X"A4",X"0A",X"ED",X"C0",X"20",X"4E",X"9B",X"64",X"B8",X"46",X"0D",
		X"20",X"2F",X"40",X"4D",X"8A",X"BB",X"64",X"58",X"00",X"54",X"EC",X"0E",X"12",X"BE",X"00",X"A5",
		X"92",X"BD",X"C2",X"BE",X"0A",X"B6",X"02",X"18",X"4A",X"92",X"02",X"53",X"6C",X"48",X"00",X"3C",
		X"12",X"2D",X"82",X"B9",X"E6",X"B2",X"6F",X"3C",X"12",X"2D",X"82",X"C3",X"62",X"4D",X"C0",X"3C",
		X"12",X"2D",X"82",X"C3",X"62",X"4D",X"C2",X"2C",X"90",X"0D",X"CE",X"9D",X"92",X"B8",X"00",X"A9",
		X"C0",X"D0",X"05",X"20",X"66",X"E4",X"A9",X"20",X"A0",X"00",X"91",X"08",X"4C",X"C3",X"E4",X"90",
		X"04",X"29",X"0F",X"F0",X"05",X"29",X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",
		X"48",X"4D",X"91",X"08",X"BD",X"49",X"4D",X"C8",X"91",X"08",X"20",X"72",X"E4",X"28",X"60",X"38",
		X"E9",X"20",X"4A",X"29",X"1F",X"09",X"E0",X"A0",X"01",X"91",X"08",X"88",X"8A",X"6A",X"91",X"08",
		X"C8",X"D0",X"1F",X"38",X"E9",X"20",X"4A",X"29",X"1F",X"09",X"A0",X"D0",X"EA",X"A4",X"0A",X"09",
		X"60",X"AA",X"98",X"4C",X"6A",X"E4",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"08",X"C8",X"8A",
		X"91",X"08",X"98",X"38",X"65",X"08",X"85",X"08",X"90",X"02",X"E6",X"09",X"60",X"A0",X"00",X"09",
		X"70",X"AA",X"98",X"4C",X"6A",X"E4",X"A8",X"A9",X"00",X"AA",X"84",X"0A",X"A0",X"00",X"0A",X"90",
		X"01",X"88",X"84",X"05",X"0A",X"26",X"05",X"85",X"04",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",
		X"84",X"07",X"0A",X"26",X"07",X"85",X"06",X"A2",X"04",X"A0",X"00",X"B5",X"02",X"91",X"08",X"B5",
		X"03",X"29",X"1F",X"C8",X"91",X"08",X"B5",X"00",X"C8",X"91",X"08",X"B5",X"01",X"45",X"0A",X"29",
		X"1F",X"45",X"0A",X"C8",X"91",X"08",X"D0",X"AA",X"00",X"09",X"0A",X"13",X"14",X"24",X"63",X"04",
		X"5A",X"04",X"50",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",X"02",X"A9",X"07",X"A0",X"FF",
		X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",X"70",X"01",X"48",X"0D",X"71",
		X"01",X"8D",X"71",X"01",X"68",X"0D",X"72",X"01",X"8D",X"72",X"01",X"60",X"A9",X"07",X"8D",X"71",
		X"01",X"A9",X"00",X"8D",X"72",X"01",X"AD",X"74",X"01",X"D0",X"4B",X"AD",X"71",X"01",X"F0",X"46",
		X"A2",X"00",X"8E",X"75",X"01",X"8E",X"79",X"01",X"8E",X"78",X"01",X"A2",X"08",X"38",X"6E",X"78",
		X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"78",X"01",X"2D",X"72",X"01",X"D0",X"02",X"A0",
		X"20",X"8C",X"74",X"01",X"AD",X"78",X"01",X"4D",X"71",X"01",X"8D",X"71",X"01",X"8A",X"0A",X"AA",
		X"BD",X"C8",X"E4",X"8D",X"76",X"01",X"BD",X"C9",X"E4",X"8D",X"77",X"01",X"BD",X"CE",X"E4",X"85",
		X"E1",X"BD",X"CF",X"E4",X"85",X"E2",X"A0",X"00",X"8C",X"00",X"89",X"AD",X"74",X"01",X"D0",X"01",
		X"60",X"AC",X"75",X"01",X"AE",X"76",X"01",X"0A",X"90",X"0D",X"9D",X"40",X"89",X"A9",X"40",X"8D",
		X"74",X"01",X"A0",X"0E",X"4C",X"EA",X"E5",X"10",X"25",X"A9",X"80",X"8D",X"74",X"01",X"AD",X"70",
		X"01",X"F0",X"04",X"A9",X"00",X"91",X"E1",X"B1",X"E1",X"EC",X"77",X"01",X"90",X"08",X"A9",X"00",
		X"8D",X"74",X"01",X"AD",X"79",X"01",X"9D",X"40",X"89",X"A0",X"0C",X"4C",X"DD",X"E5",X"A9",X"08",
		X"8D",X"00",X"89",X"9D",X"40",X"89",X"A9",X"09",X"8D",X"00",X"89",X"EA",X"A9",X"08",X"8D",X"00",
		X"89",X"EC",X"77",X"01",X"AD",X"00",X"70",X"90",X"20",X"4D",X"79",X"01",X"F0",X"13",X"A9",X"00",
		X"AC",X"75",X"01",X"91",X"E1",X"88",X"10",X"FB",X"AD",X"78",X"01",X"0D",X"73",X"01",X"8D",X"73",
		X"01",X"A9",X"00",X"8D",X"74",X"01",X"4C",X"DB",X"E5",X"91",X"E1",X"A0",X"00",X"18",X"6D",X"79",
		X"01",X"8D",X"79",X"01",X"EE",X"75",X"01",X"EE",X"76",X"01",X"8C",X"00",X"89",X"98",X"D0",X"03",
		X"4C",X"06",X"E5",X"60",X"78",X"D8",X"A9",X"FF",X"85",X"02",X"D0",X"11",X"A5",X"00",X"F0",X"0D",
		X"AD",X"00",X"78",X"29",X"40",X"F0",X"06",X"8D",X"80",X"88",X"8D",X"40",X"88",X"8D",X"80",X"89",
		X"AD",X"00",X"78",X"29",X"10",X"F0",X"03",X"4C",X"3A",X"E8",X"AD",X"00",X"80",X"18",X"2A",X"2A",
		X"2A",X"2A",X"49",X"FF",X"29",X"07",X"85",X"00",X"A5",X"00",X"C5",X"02",X"F0",X"CE",X"85",X"02",
		X"AA",X"F0",X"21",X"A9",X"C7",X"8D",X"00",X"20",X"A9",X"60",X"8D",X"01",X"20",X"BC",X"A8",X"E6",
		X"BD",X"B0",X"E6",X"AA",X"B9",X"B8",X"E6",X"9D",X"02",X"20",X"88",X"CA",X"10",X"F6",X"8D",X"80",
		X"88",X"4C",X"FC",X"E5",X"A9",X"20",X"85",X"04",X"A9",X"00",X"85",X"03",X"85",X"01",X"A8",X"A9",
		X"08",X"85",X"00",X"18",X"A5",X"01",X"91",X"03",X"69",X"05",X"85",X"01",X"C8",X"D0",X"F4",X"E6",
		X"04",X"C6",X"00",X"D0",X"EE",X"A0",X"07",X"A2",X"00",X"A9",X"11",X"9D",X"80",X"27",X"9D",X"80",
		X"26",X"48",X"8A",X"18",X"69",X"10",X"AA",X"68",X"88",X"10",X"F0",X"8D",X"B2",X"26",X"8D",X"B2",
		X"27",X"8D",X"DE",X"26",X"8D",X"EE",X"26",X"8D",X"DE",X"27",X"8D",X"EE",X"27",X"A9",X"80",X"8D",
		X"FE",X"26",X"8D",X"FE",X"27",X"4C",X"4E",X"E6",X"01",X"01",X"15",X"2B",X"45",X"71",X"01",X"01",
		X"01",X"01",X"13",X"15",X"19",X"2B",X"01",X"01",X"00",X"20",X"40",X"80",X"00",X"71",X"80",X"01",
		X"00",X"22",X"40",X"80",X"00",X"60",X"80",X"1E",X"00",X"3E",X"40",X"80",X"00",X"20",X"40",X"80",
		X"00",X"71",X"80",X"01",X"00",X"22",X"07",X"E0",X"00",X"20",X"40",X"80",X"80",X"1E",X"00",X"3E",
		X"40",X"80",X"00",X"20",X"40",X"80",X"00",X"71",X"80",X"01",X"00",X"22",X"07",X"E0",X"00",X"20",
		X"40",X"80",X"80",X"1E",X"00",X"3E",X"40",X"80",X"2F",X"51",X"40",X"80",X"00",X"20",X"40",X"80",
		X"00",X"71",X"80",X"01",X"00",X"22",X"07",X"E0",X"00",X"20",X"40",X"80",X"80",X"1E",X"00",X"3E",
		X"40",X"80",X"2F",X"51",X"40",X"80",X"11",X"A0",X"20",X"51",X"40",X"80",X"00",X"20",X"13",X"A0",
		X"00",X"C0",X"15",X"A0",X"00",X"C0",X"2F",X"40",X"00",X"C0",X"A2",X"02",X"AD",X"00",X"78",X"E0",
		X"01",X"F0",X"03",X"B0",X"02",X"4A",X"4A",X"4A",X"B5",X"DB",X"29",X"1F",X"B0",X"37",X"F0",X"10",
		X"C9",X"1B",X"B0",X"0A",X"A8",X"A5",X"E0",X"29",X"07",X"C9",X"07",X"98",X"90",X"02",X"E9",X"01",
		X"95",X"DB",X"AD",X"00",X"78",X"29",X"08",X"D0",X"04",X"A9",X"F0",X"85",X"DE",X"A5",X"DE",X"F0",
		X"08",X"C6",X"DE",X"A9",X"00",X"95",X"DB",X"95",X"D8",X"18",X"B5",X"D8",X"F0",X"23",X"D6",X"D8",
		X"D0",X"1F",X"38",X"B0",X"1C",X"C9",X"1B",X"B0",X"09",X"B5",X"DB",X"69",X"20",X"90",X"D1",X"F0",
		X"01",X"18",X"A9",X"1F",X"B0",X"CA",X"95",X"DB",X"B5",X"D8",X"F0",X"01",X"38",X"A9",X"78",X"95",
		X"D8",X"90",X"2A",X"A9",X"00",X"E0",X"01",X"90",X"16",X"F0",X"0C",X"A5",X"DF",X"29",X"0C",X"4A",
		X"4A",X"F0",X"0C",X"69",X"02",X"D0",X"08",X"A5",X"DF",X"29",X"10",X"F0",X"02",X"A9",X"01",X"38",
		X"48",X"65",X"D1",X"85",X"D1",X"68",X"38",X"65",X"D7",X"85",X"D7",X"F6",X"D3",X"CA",X"30",X"03",
		X"4C",X"2C",X"E7",X"A5",X"DF",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"A5",X"D1",X"38",X"F9",X"DF",
		X"E7",X"30",X"14",X"85",X"D1",X"E6",X"D2",X"C0",X"03",X"D0",X"0C",X"E6",X"D2",X"D0",X"08",X"7F",
		X"02",X"04",X"04",X"05",X"03",X"7F",X"7F",X"A5",X"DF",X"29",X"03",X"A8",X"F0",X"1A",X"4A",X"69",
		X"00",X"49",X"FF",X"38",X"65",X"D7",X"B0",X"08",X"65",X"D2",X"30",X"0E",X"85",X"D2",X"A9",X"00",
		X"C0",X"02",X"B0",X"02",X"E6",X"D6",X"E6",X"D6",X"85",X"D7",X"E6",X"E0",X"A5",X"E0",X"4A",X"B0",
		X"27",X"A0",X"00",X"A2",X"02",X"B5",X"D3",X"F0",X"09",X"C9",X"10",X"90",X"05",X"69",X"EF",X"C8",
		X"95",X"D3",X"CA",X"10",X"F0",X"98",X"D0",X"10",X"A2",X"02",X"B5",X"D3",X"F0",X"07",X"18",X"69",
		X"EF",X"95",X"D3",X"30",X"03",X"CA",X"10",X"F2",X"60",X"CD",X"78",X"A2",X"FE",X"9A",X"A9",X"00",
		X"8D",X"80",X"88",X"D8",X"AA",X"95",X"00",X"9D",X"00",X"01",X"9D",X"00",X"02",X"9D",X"00",X"03",
		X"9D",X"00",X"04",X"9D",X"00",X"05",X"9D",X"00",X"06",X"9D",X"00",X"07",X"9D",X"00",X"20",X"9D",
		X"00",X"21",X"9D",X"00",X"22",X"9D",X"00",X"23",X"9D",X"00",X"24",X"9D",X"00",X"25",X"9D",X"00",
		X"26",X"9D",X"00",X"27",X"9D",X"00",X"60",X"9D",X"00",X"68",X"8D",X"80",X"89",X"E8",X"D0",X"C5",
		X"A9",X"C0",X"8D",X"00",X"88",X"A9",X"07",X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"AD",X"00",X"78",
		X"29",X"10",X"D0",X"03",X"4C",X"D2",X"E8",X"A9",X"01",X"8D",X"00",X"20",X"A9",X"E2",X"8D",X"01",
		X"20",X"A9",X"20",X"8D",X"03",X"20",X"8D",X"03",X"24",X"A9",X"24",X"85",X"09",X"A9",X"02",X"85",
		X"08",X"58",X"E6",X"FB",X"A5",X"FB",X"8D",X"80",X"89",X"D0",X"F9",X"20",X"FC",X"E4",X"AD",X"74",
		X"01",X"8D",X"80",X"89",X"D0",X"F8",X"AD",X"73",X"01",X"4A",X"B0",X"03",X"20",X"9E",X"CB",X"4C",
		X"00",X"90",X"A2",X"11",X"9A",X"8A",X"86",X"00",X"A0",X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",
		X"D0",X"21",X"E8",X"D0",X"F7",X"BA",X"8A",X"8D",X"80",X"89",X"C8",X"59",X"00",X"00",X"D0",X"13",
		X"8A",X"A2",X"00",X"96",X"00",X"C8",X"D0",X"05",X"0A",X"A2",X"00",X"B0",X"4B",X"AA",X"9A",X"96",
		X"00",X"D0",X"D7",X"AA",X"8A",X"A0",X"82",X"29",X"0F",X"F0",X"02",X"A0",X"12",X"8A",X"A2",X"82",
		X"29",X"F0",X"F0",X"02",X"A2",X"12",X"98",X"9A",X"AA",X"8E",X"00",X"60",X"A2",X"A8",X"8E",X"01",
		X"60",X"A0",X"0C",X"A2",X"64",X"2C",X"00",X"78",X"30",X"FB",X"2C",X"00",X"78",X"10",X"FB",X"8D",
		X"80",X"89",X"CA",X"D0",X"F0",X"C0",X"05",X"D0",X"03",X"8E",X"01",X"60",X"88",X"D0",X"E4",X"4A",
		X"B0",X"03",X"BA",X"D0",X"D4",X"4C",X"FF",X"E9",X"A2",X"FF",X"9A",X"A2",X"00",X"8A",X"95",X"00",
		X"E8",X"D0",X"FB",X"A8",X"A9",X"01",X"85",X"01",X"A2",X"11",X"B1",X"00",X"D0",X"27",X"8A",X"91",
		X"00",X"51",X"00",X"D0",X"20",X"8A",X"0A",X"AA",X"90",X"F5",X"C8",X"D0",X"EB",X"8D",X"80",X"89",
		X"E6",X"01",X"A6",X"01",X"E0",X"04",X"90",X"E0",X"A9",X"20",X"E0",X"20",X"90",X"D8",X"E0",X"28",
		X"90",X"D6",X"4C",X"06",X"EA",X"A6",X"01",X"E0",X"20",X"85",X"02",X"90",X"03",X"8A",X"E9",X"1C",
		X"4A",X"4A",X"29",X"07",X"A8",X"A5",X"02",X"84",X"00",X"85",X"01",X"A9",X"01",X"85",X"02",X"A2",
		X"A8",X"A0",X"82",X"A5",X"00",X"D0",X"08",X"A5",X"01",X"29",X"0F",X"F0",X"02",X"A0",X"12",X"8E",
		X"01",X"60",X"8C",X"00",X"60",X"A9",X"09",X"C0",X"12",X"F0",X"02",X"A9",X"01",X"A8",X"A2",X"00",
		X"2C",X"00",X"78",X"30",X"FB",X"2C",X"00",X"78",X"10",X"FB",X"8D",X"80",X"89",X"CA",X"D0",X"F0",
		X"88",X"D0",X"ED",X"8E",X"01",X"60",X"A0",X"09",X"2C",X"00",X"78",X"30",X"FB",X"2C",X"00",X"78",
		X"10",X"FB",X"8D",X"80",X"89",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"A5",X"00",X"D0",X"08",X"A5",
		X"01",X"4A",X"4A",X"4A",X"4A",X"85",X"01",X"C6",X"02",X"F0",X"A4",X"C6",X"00",X"10",X"9C",X"8D",
		X"80",X"89",X"A9",X"FF",X"85",X"74",X"A9",X"00",X"AA",X"9D",X"00",X"01",X"9D",X"00",X"02",X"9D",
		X"00",X"03",X"CA",X"D0",X"F4",X"A8",X"85",X"21",X"A9",X"30",X"85",X"22",X"A9",X"10",X"85",X"23",
		X"8A",X"51",X"21",X"C8",X"D0",X"FB",X"E6",X"22",X"8D",X"80",X"89",X"C6",X"23",X"D0",X"F2",X"95",
		X"6B",X"E8",X"F0",X"18",X"A5",X"22",X"C9",X"60",X"D0",X"04",X"A9",X"90",X"85",X"22",X"C9",X"F0",
		X"90",X"D8",X"A2",X"FF",X"A9",X"28",X"85",X"22",X"A9",X"08",X"D0",X"D2",X"A5",X"6A",X"05",X"6B",
		X"F0",X"0A",X"A9",X"F0",X"A2",X"A2",X"8D",X"04",X"60",X"8E",X"05",X"60",X"A2",X"05",X"AD",X"0A",
		X"68",X"CD",X"0A",X"68",X"D0",X"05",X"CA",X"10",X"F8",X"85",X"75",X"A2",X"05",X"AD",X"0A",X"60",
		X"CD",X"0A",X"60",X"D0",X"05",X"CA",X"10",X"F8",X"85",X"76",X"58",X"20",X"FC",X"E4",X"A0",X"02",
		X"AD",X"73",X"01",X"F0",X"0A",X"85",X"77",X"20",X"DC",X"E4",X"A0",X"00",X"8C",X"73",X"01",X"84",
		X"69",X"4C",X"D7",X"EC",X"AD",X"74",X"01",X"0D",X"71",X"01",X"D0",X"0C",X"20",X"FC",X"E4",X"AD",
		X"73",X"01",X"85",X"77",X"A9",X"02",X"85",X"69",X"60",X"A0",X"A7",X"A9",X"04",X"20",X"5F",X"E4",
		X"A2",X"8E",X"A9",X"4A",X"20",X"53",X"E4",X"A9",X"48",X"A2",X"40",X"A0",X"00",X"20",X"8A",X"E4",
		X"20",X"41",X"EC",X"A9",X"01",X"20",X"7F",X"E4",X"A2",X"46",X"86",X"23",X"A2",X"09",X"B5",X"6A",
		X"F0",X"1B",X"86",X"22",X"20",X"66",X"E4",X"A6",X"23",X"8A",X"38",X"E9",X"08",X"85",X"23",X"A9",
		X"F6",X"A0",X"00",X"20",X"8A",X"E4",X"A5",X"22",X"20",X"54",X"DE",X"A6",X"22",X"CA",X"10",X"DE",
		X"20",X"66",X"E4",X"A9",X"F6",X"A2",X"58",X"A0",X"00",X"20",X"8A",X"E4",X"A2",X"03",X"86",X"22",
		X"A6",X"22",X"A0",X"00",X"B5",X"74",X"F0",X"03",X"BC",X"C9",X"EB",X"B9",X"48",X"4D",X"BE",X"49",
		X"4D",X"20",X"6A",X"E4",X"C6",X"22",X"10",X"E8",X"20",X"A7",X"EC",X"60",X"A2",X"5C",X"A9",X"4B",
		X"4C",X"53",X"E4",X"E6",X"30",X"10",X"06",X"A9",X"00",X"85",X"30",X"E6",X"23",X"A5",X"23",X"29",
		X"07",X"AA",X"BC",X"68",X"EB",X"A9",X"00",X"99",X"F1",X"67",X"BC",X"69",X"EB",X"BD",X"72",X"EB",
		X"99",X"F0",X"67",X"A9",X"A8",X"99",X"F1",X"67",X"A2",X"62",X"A9",X"4B",X"20",X"53",X"E4",X"20",
		X"66",X"E4",X"A4",X"30",X"A5",X"23",X"29",X"07",X"D0",X"04",X"A9",X"01",X"85",X"23",X"20",X"7F",
		X"E4",X"A2",X"90",X"A9",X"4A",X"4C",X"53",X"E4",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",
		X"16",X"00",X"10",X"10",X"40",X"40",X"90",X"90",X"FF",X"FF",X"A2",X"8E",X"A9",X"4A",X"20",X"53",
		X"E4",X"A0",X"06",X"84",X"23",X"20",X"66",X"E4",X"A4",X"23",X"B9",X"BB",X"EB",X"BE",X"C2",X"EB",
		X"20",X"8A",X"E4",X"A5",X"23",X"49",X"FF",X"29",X"07",X"A8",X"20",X"5F",X"E4",X"A5",X"23",X"D0",
		X"07",X"A2",X"1E",X"A9",X"4B",X"4C",X"AC",X"EB",X"A2",X"18",X"A9",X"4B",X"20",X"53",X"E4",X"C6",
		X"23",X"10",X"D2",X"A2",X"3C",X"A9",X"4B",X"20",X"53",X"E4",X"60",X"DE",X"9D",X"1F",X"9D",X"DE",
		X"1F",X"DE",X"F4",X"D8",X"D8",X"10",X"D8",X"10",X"10",X"38",X"34",X"36",X"1E",X"20",X"66",X"E4",
		X"A9",X"01",X"20",X"7D",X"E4",X"A2",X"06",X"86",X"22",X"A4",X"22",X"A9",X"98",X"BE",X"1C",X"EC",
		X"20",X"8A",X"E4",X"A2",X"54",X"A9",X"4B",X"20",X"53",X"E4",X"C6",X"22",X"10",X"EB",X"A2",X"06",
		X"86",X"22",X"A4",X"22",X"B9",X"23",X"EC",X"A2",X"60",X"20",X"8A",X"E4",X"A2",X"4C",X"A9",X"4B",
		X"20",X"53",X"E4",X"C6",X"22",X"10",X"EB",X"AD",X"00",X"88",X"29",X"20",X"D0",X"09",X"06",X"21",
		X"90",X"02",X"E6",X"38",X"4C",X"1B",X"EC",X"A9",X"20",X"85",X"21",X"60",X"B8",X"D0",X"E8",X"00",
		X"18",X"30",X"48",X"B2",X"CC",X"E6",X"00",X"1A",X"34",X"4E",X"A2",X"CE",X"A9",X"4B",X"20",X"53",
		X"E4",X"A9",X"20",X"85",X"21",X"A2",X"C2",X"A9",X"4B",X"20",X"53",X"E4",X"C6",X"21",X"10",X"F5",
		X"60",X"A2",X"0F",X"86",X"22",X"8D",X"0B",X"60",X"EA",X"AD",X"08",X"60",X"85",X"24",X"8D",X"0B",
		X"68",X"EA",X"AD",X"08",X"68",X"48",X"29",X"01",X"18",X"20",X"54",X"DE",X"46",X"24",X"68",X"6A",
		X"C6",X"22",X"10",X"F1",X"A9",X"D0",X"A0",X"00",X"A2",X"F8",X"20",X"8A",X"E4",X"A2",X"07",X"86",
		X"22",X"A9",X"78",X"85",X"39",X"A9",X"07",X"85",X"3A",X"A9",X"00",X"85",X"38",X"A8",X"B1",X"38",
		X"49",X"FF",X"29",X"7F",X"48",X"29",X"01",X"18",X"20",X"54",X"DE",X"68",X"6A",X"C8",X"C6",X"3A",
		X"10",X"F2",X"A9",X"D0",X"A0",X"00",X"A2",X"F8",X"20",X"8A",X"E4",X"A5",X"39",X"18",X"69",X"08",
		X"85",X"39",X"C9",X"90",X"90",X"CF",X"60",X"84",X"24",X"AD",X"00",X"78",X"29",X"0F",X"85",X"21",
		X"AD",X"00",X"80",X"29",X"1F",X"85",X"22",X"AD",X"00",X"88",X"29",X"7F",X"85",X"23",X"A5",X"21",
		X"09",X"10",X"25",X"22",X"09",X"60",X"25",X"23",X"49",X"7F",X"F0",X"07",X"69",X"40",X"8D",X"00",
		X"60",X"A0",X"A4",X"8C",X"01",X"60",X"60",X"A2",X"18",X"2C",X"00",X"78",X"10",X"FB",X"2C",X"00",
		X"78",X"30",X"FB",X"CA",X"10",X"F3",X"E6",X"4F",X"2C",X"00",X"78",X"50",X"FB",X"A9",X"00",X"85",
		X"08",X"A9",X"20",X"85",X"09",X"AD",X"00",X"78",X"49",X"FF",X"29",X"24",X"F0",X"26",X"06",X"7B",
		X"90",X"1F",X"AD",X"00",X"88",X"29",X"40",X"D0",X"06",X"20",X"C2",X"E1",X"20",X"F4",X"E5",X"E6",
		X"69",X"E6",X"69",X"A9",X"00",X"A2",X"06",X"9D",X"00",X"60",X"9D",X"00",X"68",X"CA",X"CA",X"10",
		X"F6",X"4C",X"28",X"ED",X"A9",X"20",X"85",X"7B",X"A5",X"69",X"C9",X"0C",X"D0",X"0E",X"A5",X"38",
		X"29",X"07",X"D0",X"02",X"A9",X"01",X"09",X"C0",X"A8",X"4C",X"3E",X"ED",X"A0",X"A7",X"A9",X"04",
		X"20",X"5F",X"E4",X"A2",X"8E",X"A9",X"4A",X"20",X"53",X"E4",X"20",X"78",X"ED",X"20",X"66",X"E4",
		X"20",X"13",X"E4",X"A9",X"C0",X"85",X"F8",X"8D",X"40",X"88",X"8D",X"80",X"89",X"AD",X"00",X"78",
		X"29",X"10",X"D0",X"03",X"4C",X"D7",X"EC",X"4C",X"3A",X"E8",X"93",X"EA",X"A8",X"EA",X"1B",X"EB",
		X"22",X"EB",X"29",X"EC",X"79",X"EB",X"CC",X"EB",X"A6",X"69",X"E0",X"0E",X"90",X"04",X"A2",X"02",
		X"86",X"69",X"BD",X"6B",X"ED",X"48",X"BD",X"6A",X"ED",X"48",X"60",X"A9",X"00",X"85",X"00",X"8D",
		X"13",X"E4",X"20",X"C2",X"E1",X"20",X"FC",X"E4",X"AD",X"74",X"01",X"30",X"32",X"A6",X"35",X"AD",
		X"00",X"88",X"29",X"20",X"85",X"35",X"D0",X"27",X"AD",X"00",X"80",X"29",X"02",X"D0",X"0D",X"A5",
		X"00",X"D0",X"03",X"4C",X"3A",X"E8",X"20",X"DF",X"ED",X"4C",X"CF",X"ED",X"8A",X"29",X"20",X"F0",
		X"0E",X"E6",X"00",X"E6",X"00",X"A5",X"00",X"C9",X"08",X"90",X"04",X"A9",X"00",X"85",X"00",X"20",
		X"03",X"EE",X"20",X"11",X"EE",X"AD",X"00",X"78",X"29",X"10",X"F0",X"BC",X"4C",X"3A",X"E8",X"A6",
		X"00",X"E0",X"08",X"90",X"04",X"A2",X"00",X"86",X"00",X"BD",X"F3",X"ED",X"48",X"BD",X"F2",X"ED",
		X"48",X"60",X"F9",X"ED",X"F9",X"ED",X"FC",X"ED",X"FF",X"ED",X"4C",X"D8",X"E4",X"4C",X"D4",X"E4",
		X"4C",X"DC",X"E4",X"A5",X"1D",X"29",X"1F",X"C9",X"1F",X"D0",X"05",X"68",X"68",X"4C",X"E1",X"90",
		X"60",X"2C",X"00",X"78",X"50",X"FB",X"A9",X"20",X"85",X"09",X"A9",X"00",X"85",X"08",X"A2",X"A6",
		X"A9",X"4B",X"20",X"53",X"E4",X"A9",X"01",X"A0",X"40",X"20",X"7F",X"E4",X"20",X"32",X"EF",X"20",
		X"49",X"EF",X"20",X"68",X"EF",X"20",X"A1",X"EF",X"A2",X"40",X"A9",X"B0",X"20",X"EE",X"E1",X"A0",
		X"29",X"20",X"FC",X"E1",X"A5",X"00",X"4A",X"A8",X"B9",X"98",X"EE",X"AA",X"B9",X"94",X"EE",X"48",
		X"A9",X"E0",X"20",X"EE",X"E1",X"68",X"A8",X"20",X"FC",X"E1",X"20",X"ED",X"EE",X"A9",X"F0",X"A2",
		X"D0",X"20",X"EE",X"E1",X"20",X"9C",X"EE",X"20",X"AD",X"EE",X"A2",X"C0",X"A9",X"F0",X"20",X"EE",
		X"E1",X"18",X"A5",X"22",X"20",X"47",X"DE",X"A5",X"21",X"20",X"47",X"DE",X"AD",X"74",X"01",X"10",
		X"0C",X"A9",X"F0",X"A2",X"50",X"20",X"EE",X"E1",X"A0",X"27",X"20",X"FC",X"E1",X"20",X"13",X"E4",
		X"8D",X"40",X"88",X"60",X"28",X"2A",X"2B",X"2C",X"30",X"30",X"30",X"30",X"A5",X"3A",X"18",X"20",
		X"47",X"DE",X"A5",X"39",X"20",X"47",X"DE",X"A5",X"38",X"20",X"47",X"DE",X"60",X"A9",X"00",X"85",
		X"21",X"85",X"22",X"AD",X"54",X"04",X"85",X"38",X"AD",X"55",X"04",X"85",X"39",X"AD",X"56",X"04",
		X"85",X"3A",X"A5",X"23",X"05",X"24",X"F0",X"24",X"F8",X"A5",X"21",X"18",X"69",X"01",X"85",X"21",
		X"A5",X"22",X"69",X"00",X"85",X"22",X"D8",X"A5",X"38",X"38",X"E5",X"23",X"85",X"38",X"A5",X"39",
		X"E5",X"24",X"85",X"39",X"A5",X"3A",X"E9",X"00",X"85",X"3A",X"10",X"DC",X"60",X"AD",X"52",X"04",
		X"0A",X"85",X"21",X"AD",X"53",X"04",X"2A",X"85",X"22",X"AD",X"50",X"04",X"18",X"65",X"21",X"85",
		X"21",X"85",X"23",X"AD",X"51",X"04",X"65",X"22",X"85",X"22",X"85",X"24",X"A0",X"0F",X"A9",X"00",
		X"85",X"38",X"85",X"39",X"85",X"3A",X"F8",X"06",X"21",X"26",X"22",X"A5",X"38",X"65",X"38",X"85",
		X"38",X"A5",X"39",X"65",X"39",X"85",X"39",X"A5",X"3A",X"65",X"3A",X"85",X"3A",X"88",X"10",X"E7",
		X"D8",X"60",X"A2",X"68",X"A9",X"FC",X"20",X"EE",X"E1",X"A5",X"F0",X"29",X"10",X"F0",X"05",X"A9",
		X"1C",X"4C",X"46",X"EF",X"A9",X"22",X"4C",X"F8",X"D9",X"A9",X"F0",X"A2",X"58",X"20",X"EE",X"E1",
		X"A5",X"F1",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"B9",X"60",X"EF",X"18",X"20",X"47",X"DE",X"60",
		X"00",X"00",X"14",X"24",X"15",X"13",X"00",X"00",X"A9",X"F0",X"A2",X"60",X"20",X"EE",X"E1",X"A5",
		X"F1",X"29",X"03",X"A8",X"B9",X"9D",X"EF",X"18",X"20",X"54",X"DE",X"A5",X"F1",X"29",X"0C",X"4A",
		X"4A",X"A8",X"B9",X"99",X"EF",X"20",X"54",X"DE",X"A5",X"F1",X"29",X"10",X"D0",X"05",X"A9",X"01",
		X"4C",X"95",X"EF",X"A9",X"02",X"20",X"54",X"DE",X"60",X"01",X"04",X"05",X"06",X"00",X"02",X"01",
		X"00",X"A9",X"C0",X"A2",X"D0",X"20",X"EE",X"E1",X"A5",X"F0",X"4A",X"4A",X"29",X"03",X"A8",X"B9",
		X"F0",X"EF",X"85",X"21",X"AD",X"C6",X"45",X"AE",X"C7",X"45",X"20",X"6A",X"E4",X"A2",X"FB",X"A9",
		X"F8",X"A0",X"00",X"20",X"8A",X"E4",X"C6",X"21",X"10",X"EA",X"AD",X"00",X"88",X"30",X"20",X"A9",
		X"C0",X"A2",X"B0",X"20",X"EE",X"E1",X"A9",X"18",X"20",X"F8",X"D9",X"A6",X"18",X"AD",X"00",X"88",
		X"29",X"40",X"85",X"18",X"D0",X"09",X"8A",X"F0",X"06",X"A5",X"F8",X"49",X"C0",X"85",X"F8",X"60",
		X"02",X"03",X"04",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"E8",X"3A",X"E8",X"EA",X"CB");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
