library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpe_13l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpe_13l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"33",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"F7",X"F1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F1",X"33",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",
		X"80",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"F6",X"F3",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F1",X"77",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F6",
		X"C0",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F1",X"FF",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F7",
		X"D1",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"10",X"F1",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",
		X"F3",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"FF",X"FE",X"00",X"00",
		X"00",X"00",X"00",X"10",X"F3",X"FB",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"10",X"FF",
		X"F1",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"30",X"F3",X"F9",X"FE",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"0F",X"10",X"FE",
		X"F3",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"FF",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"F3",X"FD",X"FA",X"00",X"00",X"00",X"00",X"11",X"98",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"08",X"0F",X"30",X"FE",
		X"F7",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"71",X"FF",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"F0",X"F1",X"FF",X"F0",X"00",X"00",X"00",X"00",X"33",X"B8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"88",X"00",X"00",X"08",X"09",X"30",X"FF",
		X"F3",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"F8",X"FF",X"FC",X"C0",X"00",
		X"00",X"00",X"00",X"F0",X"F1",X"FF",X"F0",X"00",X"00",X"00",X"00",X"33",X"E8",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"A8",X"00",X"00",X"09",X"0C",X"30",X"FF",
		X"F3",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F8",X"FF",X"FE",X"C0",X"00",
		X"00",X"00",X"10",X"F0",X"F3",X"FF",X"F0",X"00",X"00",X"00",X"00",X"77",X"F8",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"EC",X"00",X"00",X"09",X"08",X"71",X"FF",
		X"FB",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FC",X"F7",X"FC",X"E0",X"00",
		X"00",X"00",X"30",X"F0",X"F1",X"FF",X"F8",X"00",X"00",X"00",X"00",X"77",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"FC",X"00",X"00",X"09",X"08",X"71",X"FF",
		X"FB",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FC",X"F7",X"F8",X"E0",X"00",
		X"00",X"10",X"30",X"F0",X"F1",X"FF",X"F8",X"80",X"00",X"00",X"00",X"77",X"F0",X"E0",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"FC",X"80",X"00",X"0B",X"08",X"70",X"FE",
		X"FF",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FE",X"FF",X"F8",X"E0",X"00",
		X"00",X"30",X"B0",X"F0",X"F3",X"FF",X"F8",X"80",X"00",X"00",X"00",X"FF",X"F8",X"E0",X"00",X"00",
		X"00",X"33",X"88",X"00",X"00",X"00",X"00",X"00",X"F7",X"F8",X"80",X"00",X"0B",X"0C",X"70",X"FE",
		X"FF",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FE",X"FF",X"FC",X"E0",X"00",
		X"00",X"30",X"F0",X"FD",X"FB",X"FF",X"FC",X"80",X"00",X"00",X"00",X"FF",X"F8",X"E0",X"00",X"00",
		X"00",X"33",X"88",X"00",X"00",X"00",X"00",X"00",X"F3",X"F8",X"80",X"00",X"06",X"0C",X"71",X"FE",
		X"F7",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"EE",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FC",X"FF",X"FC",X"E0",X"00",
		X"00",X"F0",X"F0",X"FF",X"FD",X"FF",X"FC",X"C4",X"00",X"11",X"11",X"FF",X"F8",X"E0",X"00",X"00",
		X"00",X"77",X"C0",X"00",X"00",X"00",X"00",X"00",X"F7",X"FC",X"C0",X"80",X"00",X"04",X"71",X"FF",
		X"F6",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F7",X"C4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"FE",X"FF",X"F8",X"E0",X"00",
		X"00",X"F0",X"F0",X"F7",X"FE",X"FF",X"FC",X"C4",X"00",X"33",X"BB",X"FB",X"F0",X"E0",X"00",X"00",
		X"00",X"FF",X"C0",X"00",X"00",X"00",X"00",X"D0",X"F3",X"FD",X"D0",X"80",X"00",X"02",X"70",X"FF",
		X"F6",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F7",X"C4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"FF",X"FF",X"F0",X"E0",X"00",
		X"30",X"F0",X"F0",X"FB",X"FF",X"FF",X"FF",X"E0",X"00",X"33",X"FF",X"F7",X"F0",X"F4",X"00",X"00",
		X"00",X"FF",X"C8",X"00",X"00",X"00",X"10",X"F0",X"F3",X"FD",X"F8",X"80",X"00",X"00",X"70",X"FF",
		X"F6",X"DD",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"F7",X"FF",X"FF",X"F0",X"F0",X"00",
		X"70",X"F0",X"F3",X"FD",X"FF",X"FF",X"FF",X"E8",X"00",X"77",X"FF",X"FF",X"F8",X"FC",X"00",X"00",
		X"11",X"FE",X"C0",X"00",X"00",X"00",X"10",X"F4",X"F7",X"FF",X"FC",X"80",X"00",X"00",X"78",X"FF",
		X"FE",X"FF",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FB",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"F7",X"F7",X"FE",X"F0",X"F0",X"80",
		X"71",X"F8",X"F7",X"FF",X"FF",X"FF",X"FF",X"F0",X"33",X"FF",X"FF",X"FD",X"F0",X"F8",X"00",X"00",
		X"11",X"FC",X"E0",X"C0",X"00",X"00",X"10",X"FC",X"FF",X"FF",X"FC",X"C0",X"00",X"00",X"F3",X"FE",
		X"FE",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FB",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"F7",X"F7",X"FE",X"F0",X"F0",X"E0",
		X"FF",X"FA",X"F7",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"FD",X"FF",X"FC",X"F1",X"F0",X"C0",X"00",
		X"33",X"F8",X"E0",X"C0",X"00",X"00",X"11",X"FE",X"FF",X"FF",X"FD",X"C4",X"00",X"00",X"F3",X"FE",
		X"FF",X"FF",X"EE",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"33",X"FF",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"F7",X"F7",X"FF",X"F0",X"F1",X"F1",
		X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FE",X"F3",X"FF",X"F0",X"FF",X"FE",X"F0",X"F0",X"C0",X"00",
		X"33",X"F8",X"E0",X"E0",X"00",X"00",X"33",X"FF",X"F7",X"FF",X"FF",X"F8",X"00",X"33",X"F3",X"FE",
		X"FF",X"FF",X"FF",X"88",X"00",X"00",X"77",X"66",X"00",X"00",X"33",X"FF",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"FF",X"F3",X"F3",X"FD",
		X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FC",X"F7",X"FE",X"F0",X"FF",X"FF",X"F0",X"F0",X"E0",X"00",
		X"BB",X"FE",X"E0",X"E0",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"88",X"00",X"00",X"77",X"EC",X"00",X"00",X"33",X"FF",X"FF",X"CC",X"00",X"00",
		X"00",X"11",X"CC",X"00",X"00",X"00",X"00",X"00",X"11",X"FD",X"FF",X"FB",X"FE",X"F7",X"F7",X"FB",
		X"FE",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"F7",X"FE",X"F0",X"F0",X"E0",X"11",
		X"FF",X"FC",X"F0",X"E0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"88",X"FF",X"F7",X"FF",
		X"FF",X"FC",X"FF",X"88",X"00",X"11",X"FF",X"EC",X"00",X"00",X"33",X"FF",X"FD",X"CC",X"00",X"00",
		X"00",X"11",X"CC",X"00",X"00",X"00",X"00",X"00",X"11",X"FC",X"FF",X"FF",X"FD",X"FE",X"FF",X"F7",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FC",X"F8",X"FF",X"F8",X"F0",X"F1",X"F0",X"11",
		X"FF",X"FC",X"FC",X"F1",X"00",X"00",X"FF",X"FF",X"FD",X"FF",X"FF",X"F2",X"88",X"FF",X"F7",X"FF",
		X"FF",X"F8",X"F3",X"88",X"00",X"11",X"FF",X"EA",X"00",X"00",X"77",X"FF",X"FF",X"EC",X"00",X"00",
		X"00",X"11",X"FE",X"00",X"00",X"00",X"00",X"00",X"11",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FD",X"F9",X"FF",X"FE",X"F6",X"F3",X"F8",X"11",
		X"FF",X"F9",X"F9",X"F9",X"80",X"11",X"FF",X"F7",X"FD",X"FF",X"FE",X"F5",X"99",X"FF",X"FB",X"FF",
		X"FF",X"F0",X"F3",X"88",X"00",X"30",X"FF",X"EE",X"00",X"00",X"77",X"FB",X"FF",X"E8",X"00",X"00",
		X"00",X"11",X"FE",X"C0",X"00",X"00",X"00",X"00",X"11",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"F3",X"FC",X"33",
		X"FF",X"F7",X"F9",X"FB",X"80",X"11",X"FF",X"F1",X"FF",X"F8",X"FE",X"F5",X"99",X"FF",X"FF",X"FF",
		X"FE",X"F0",X"F0",X"EE",X"00",X"31",X"FF",X"EE",X"00",X"00",X"77",X"FB",X"FF",X"EA",X"00",X"00",
		X"00",X"11",X"FE",X"C0",X"00",X"00",X"00",X"00",X"11",X"F9",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"F9",X"FF",X"F7",X"FE",X"B3",
		X"FE",X"FF",X"FF",X"FB",X"80",X"11",X"FE",X"F0",X"F3",X"FF",X"FE",X"FF",X"99",X"FF",X"FF",X"FF",
		X"FF",X"F1",X"F5",X"EE",X"00",X"31",X"FF",X"FE",X"00",X"00",X"FF",X"FE",X"F7",X"E6",X"00",X"00",
		X"10",X"F3",X"FD",X"F0",X"00",X"00",X"00",X"00",X"17",X"FD",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",
		X"FF",X"FF",X"FF",X"F3",X"C0",X"73",X"FE",X"F0",X"F3",X"FF",X"FC",X"FF",X"BB",X"FF",X"FC",X"F7",
		X"FF",X"F1",X"FF",X"EE",X"00",X"F1",X"FF",X"FC",X"00",X"00",X"FF",X"FE",X"FF",X"FF",X"00",X"00",
		X"10",X"F3",X"FB",X"F0",X"00",X"00",X"00",X"11",X"F9",X"FF",X"FF",X"FD",X"FC",X"F3",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",
		X"FF",X"FF",X"FE",X"FF",X"C0",X"73",X"FC",X"F4",X"FB",X"FF",X"FB",X"FF",X"BB",X"FF",X"FF",X"F7",
		X"FF",X"FB",X"FF",X"FF",X"88",X"F3",X"FF",X"FC",X"00",X"10",X"FF",X"FE",X"FF",X"FF",X"C0",X"00",
		X"10",X"F7",X"FF",X"F4",X"80",X"00",X"00",X"32",X"F8",X"FF",X"FF",X"F9",X"FE",X"F1",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"C8",X"F7",X"FC",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"FF",X"FB",X"FF",X"FF",X"98",X"FD",X"FF",X"F0",X"00",X"30",X"FF",X"FE",X"F7",X"FF",X"C0",X"00",
		X"70",X"FF",X"FF",X"FC",X"80",X"00",X"00",X"74",X"F9",X"F7",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FD",X"FF",X"E8",X"F7",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"FB",X"FF",X"FF",X"F8",X"FE",X"FE",X"FC",X"E0",X"30",X"FF",X"F7",X"FF",X"FF",X"C0",X"00",
		X"70",X"FF",X"F7",X"FC",X"80",X"00",X"00",X"F8",X"FB",X"F7",X"FF",X"FF",X"FF",X"FA",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"FF",X"FC",X"F7",X"F2",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FD",X"FE",X"E0",X"30",X"FF",X"F7",X"FF",X"FE",X"C4",X"00",
		X"71",X"F7",X"F7",X"FD",X"80",X"10",X"CC",X"F2",X"FB",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F9",X"FB",X"FF",X"FC",X"F7",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"F0",X"74",X"FF",X"F3",X"FF",X"FE",X"F7",X"00",
		X"F1",X"F3",X"FB",X"FB",X"80",X"10",X"FF",X"FF",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FB",X"FF",X"FC",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"F0",X"F8",X"FF",X"F7",X"FF",X"FC",X"F7",X"CC",
		X"F3",X"F7",X"FF",X"FB",X"C0",X"30",X"FF",X"FF",X"F3",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"F0",X"F0",X"FF",X"F7",X"FF",X"FB",X"FF",X"FF",
		X"FB",X"FB",X"FF",X"F7",X"FB",X"F9",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"F0",X"FC",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F4",X"F5",X"FC",X"F7",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F6",X"F7",X"FC",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FC",X"F7",X"FF",X"FF",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F8",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"F8",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
