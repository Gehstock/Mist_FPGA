library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GAL_HIT is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GAL_HIT is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"65",X"75",X"88",X"90",X"93",X"9B",X"A3",X"A3",X"A3",X"A6",X"9E",X"9B",X"9B",X"A3",X"AB",X"B6",
		X"B9",X"B9",X"BE",X"B9",X"AE",X"A6",X"9E",X"98",X"88",X"78",X"68",X"65",X"65",X"65",X"62",X"68",
		X"68",X"65",X"5D",X"52",X"47",X"47",X"4A",X"4D",X"4D",X"4D",X"52",X"65",X"7D",X"88",X"90",X"9B",
		X"A3",X"AE",X"AE",X"AB",X"AB",X"9E",X"98",X"88",X"70",X"52",X"37",X"1F",X"17",X"1F",X"27",X"3A",
		X"5A",X"68",X"78",X"83",X"93",X"A3",X"AB",X"AE",X"A3",X"93",X"88",X"88",X"83",X"88",X"8B",X"88",
		X"78",X"62",X"4A",X"42",X"3A",X"42",X"4D",X"55",X"65",X"78",X"83",X"8B",X"93",X"90",X"88",X"88",
		X"98",X"A6",X"A6",X"AB",X"9E",X"8B",X"7D",X"68",X"70",X"88",X"AB",X"CE",X"E9",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"DC",X"9B",X"4D",X"14",X"01",X"04",X"2F",X"52",X"5D",X"68",X"78",X"80",X"78",X"70",
		X"5D",X"47",X"32",X"1F",X"14",X"09",X"11",X"1C",X"32",X"52",X"83",X"B9",X"D1",X"C9",X"AB",X"8B",
		X"70",X"68",X"75",X"78",X"80",X"8B",X"8B",X"98",X"AB",X"BE",X"C1",X"AB",X"83",X"5D",X"3A",X"17",
		X"11",X"17",X"27",X"3A",X"65",X"90",X"AE",X"B6",X"9B",X"78",X"55",X"4A",X"4D",X"5A",X"5D",X"52",
		X"4A",X"4A",X"52",X"78",X"AB",X"D4",X"FC",X"FC",X"F7",X"E9",X"E1",X"D1",X"C9",X"BE",X"AB",X"90",
		X"52",X"14",X"01",X"01",X"01",X"01",X"01",X"01",X"2F",X"4A",X"52",X"47",X"47",X"62",X"70",X"7D",
		X"7D",X"78",X"7D",X"90",X"B3",X"CE",X"EC",X"FC",X"FC",X"FC",X"FC",X"F4",X"E9",X"F4",X"FC",X"FC",
		X"FC",X"FC",X"CE",X"98",X"65",X"2C",X"01",X"01",X"01",X"01",X"01",X"32",X"6D",X"7D",X"68",X"4A",
		X"27",X"11",X"1C",X"3A",X"4D",X"62",X"68",X"65",X"68",X"70",X"80",X"9B",X"D1",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"DC",X"A3",X"75",X"55",X"62",X"80",X"A3",X"BE",X"CE",X"C1",X"90",X"4A",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"37",X"88",X"C9",X"FC",X"FC",X"FC",X"FC",X"FC",X"DC",
		X"B6",X"90",X"68",X"3F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1F",X"83",X"BE",X"D1",X"CE",
		X"D4",X"F4",X"FC",X"FC",X"FC",X"F7",X"D1",X"CE",X"DC",X"F7",X"FC",X"FC",X"FC",X"FC",X"D1",X"8B",
		X"68",X"68",X"88",X"A6",X"C1",X"D9",X"D4",X"BE",X"A3",X"88",X"75",X"68",X"62",X"5D",X"62",X"68",
		X"6D",X"78",X"75",X"55",X"2C",X"11",X"11",X"2F",X"55",X"75",X"83",X"93",X"9E",X"B9",X"E9",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BE",X"68",X"32",X"11",X"17",X"32",X"52",X"7D",
		X"AE",X"E1",X"F7",X"E1",X"A3",X"62",X"17",X"01",X"01",X"01",X"01",X"01",X"1C",X"4D",X"7D",X"90",
		X"9B",X"A6",X"B6",X"BE",X"A6",X"70",X"37",X"14",X"14",X"1C",X"14",X"1C",X"2F",X"3A",X"3A",X"3A",
		X"4A",X"52",X"4A",X"47",X"3A",X"24",X"11",X"14",X"27",X"3A",X"65",X"9E",X"D4",X"FC",X"FC",X"F7",
		X"D4",X"AB",X"93",X"93",X"93",X"83",X"68",X"4D",X"37",X"37",X"5D",X"9B",X"EC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"F7",X"CE",X"AB",X"93",X"7D",X"65",X"65",X"75",X"88",X"93",X"98",X"98",X"93",
		X"93",X"90",X"93",X"8B",X"90",X"90",X"90",X"8B",X"8B",X"90",X"8B",X"90",X"90",X"90",X"90",X"8B",
		X"8B",X"8B",X"8B",X"8B",X"88",X"88",X"88",X"88",X"88",X"83",X"83",X"80",X"83",X"80",X"80",X"80",
		X"80",X"7D",X"7D",X"7D",X"80",X"80",X"80",X"78",X"78",X"78",X"7D",X"78",X"75",X"78",X"75",X"78",
		X"78",X"78",X"75",X"78",X"75",X"70",X"75",X"75",X"75",X"75",X"70",X"6D",X"68",X"6D",X"70",X"6D",
		X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"70",X"70",X"70",X"75",X"75",X"75",X"75",
		X"75",X"70",X"62",X"4D",X"4D",X"4D",X"47",X"4A",X"68",X"98",X"B6",X"B3",X"9B",X"78",X"5A",X"3F",
		X"32",X"2F",X"32",X"3F",X"5A",X"90",X"D1",X"FC",X"FC",X"FC",X"FC",X"FC",X"E9",X"90",X"4D",X"3A",
		X"47",X"5D",X"5D",X"4D",X"3A",X"27",X"1C",X"14",X"11",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"04",X"4A",X"9E",X"F7",X"FC",X"FC",X"FC",X"FC",X"EC",X"E4",X"E4",X"D1",X"AB",X"80",X"62",X"47",
		X"37",X"2F",X"2C",X"24",X"04",X"01",X"24",X"52",X"70",X"70",X"62",X"4D",X"3F",X"37",X"37",X"3A",
		X"4D",X"62",X"78",X"93",X"AE",X"D1",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"B6",X"68",
		X"2C",X"01",X"01",X"01",X"01",X"01",X"01",X"09",X"47",X"65",X"68",X"68",X"62",X"5A",X"52",X"4D",
		X"52",X"4D",X"52",X"52",X"5A",X"5D",X"65",X"68",X"6D",X"70",X"75",X"75",X"75",X"65",X"37",X"1C",
		X"09",X"09",X"1C",X"32",X"4D",X"70",X"93",X"AB",X"C9",X"D9",X"E9",X"EF",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"F7",X"6D",X"0C",X"01",X"01",X"01",X"01",X"01",X"17",X"62",X"83",X"78",
		X"5A",X"37",X"14",X"04",X"01",X"01",X"01",X"01",X"04",X"11",X"1C",X"1C",X"01",X"01",X"0C",X"3F",
		X"6D",X"7D",X"78",X"68",X"65",X"83",X"B3",X"E1",X"F4",X"E4",X"C6",X"A3",X"8B",X"75",X"68",X"65",
		X"5D",X"62",X"65",X"62",X"5A",X"3F",X"27",X"17",X"1F",X"5A",X"9E",X"CE",X"D4",X"C9",X"AE",X"A6",
		X"AE",X"AB",X"9B",X"83",X"80",X"98",X"9B",X"9B",X"9B",X"B6",X"D9",X"E4",X"E1",X"DC",X"E1",X"D4",
		X"B3",X"83",X"5A",X"3A",X"1F",X"11",X"0C",X"11",X"14",X"1C",X"1F",X"2C",X"2C",X"1F",X"27",X"32",
		X"3F",X"5D",X"83",X"9B",X"93",X"93",X"88",X"7D",X"7D",X"75",X"70",X"70",X"6D",X"68",X"68",X"68",
		X"5A",X"5A",X"75",X"88",X"93",X"93",X"90",X"90",X"88",X"83",X"80",X"80",X"7D",X"7D",X"7D",X"80",
		X"7D",X"80",X"80",X"80",X"80",X"83",X"80",X"80",X"7D",X"7D",X"80",X"80",X"83",X"83",X"80",X"80",
		X"80",X"7D",X"7D",X"70",X"70",X"6D",X"75",X"83",X"90",X"93",X"90",X"88",X"88",X"80",X"78",X"7D",
		X"70",X"68",X"70",X"78",X"78",X"7D",X"78",X"78",X"78",X"75",X"78",X"75",X"70",X"68",X"4D",X"3A",
		X"4A",X"70",X"93",X"A3",X"B6",X"B9",X"B3",X"A3",X"90",X"80",X"75",X"70",X"68",X"68",X"68",X"65",
		X"68",X"68",X"68",X"68",X"68",X"6D",X"6D",X"70",X"70",X"75",X"75",X"75",X"75",X"78",X"75",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"70",X"55",X"37",X"1F",X"24",X"47",X"68",X"7D",X"88",X"8B",
		X"88",X"88",X"88",X"8B",X"AB",X"CE",X"E9",X"FC",X"FC",X"FC",X"FC",X"EF",X"C9",X"AB",X"80",X"5A",
		X"4A",X"47",X"37",X"2C",X"32",X"4D",X"70",X"78",X"7D",X"8B",X"90",X"88",X"68",X"4A",X"2C",X"1C",
		X"11",X"09",X"01",X"01",X"01",X"01",X"14",X"27",X"47",X"70",X"AE",X"E1",X"F4",X"E4",X"D1",X"AE",
		X"93",X"80",X"70",X"68",X"62",X"62",X"65",X"68",X"6D",X"75",X"78",X"78",X"65",X"4A",X"4D",X"5A",
		X"62",X"65",X"68",X"88",X"B9",X"EC",X"FC",X"F4",X"D1",X"B6",X"B3",X"AE",X"A3",X"98",X"A3",X"C6",
		X"D9",X"D4",X"D4",X"E1",X"E1",X"C9",X"9E",X"78",X"62",X"3F",X"32",X"2C",X"27",X"2C",X"32",X"37",
		X"3F",X"47",X"4A",X"52",X"55",X"5A",X"5D",X"5D",X"5A",X"3F",X"27",X"14",X"11",X"14",X"24",X"4A",
		X"80",X"A6",X"BE",X"C6",X"CE",X"E4",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"DC",X"BE",X"AB",X"8B",
		X"5D",X"2F",X"14",X"01",X"01",X"01",X"01",X"01",X"01",X"17",X"3F",X"65",X"70",X"6D",X"5D",X"4D",
		X"4D",X"68",X"9B",X"BE",X"C9",X"B9",X"B3",X"AB",X"9B",X"A3",X"B3",X"C6",X"D1",X"B6",X"8B",X"52",
		X"1C",X"11",X"11",X"14",X"37",X"62",X"90",X"9E",X"9B",X"83",X"75",X"5D",X"47",X"32",X"2F",X"24",
		X"17",X"11",X"11",X"17",X"27",X"5D",X"A3",X"E1",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"EF",X"CE",
		X"9B",X"7D",X"68",X"62",X"62",X"7D",X"98",X"9E",X"93",X"7D",X"6D",X"5D",X"55",X"52",X"52",X"52",
		X"55",X"55",X"5D",X"62",X"65",X"68",X"6D",X"70",X"75",X"7D",X"78",X"7D",X"80",X"83",X"78",X"62",
		X"3A",X"27",X"14",X"17",X"27",X"3F",X"5A",X"78",X"98",X"AE",X"C6",X"DC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"F7",X"A6",X"80",X"70",X"62",X"65",X"7D",X"98",X"A6",X"9B",X"80",X"62",X"32",
		X"04",X"01",X"01",X"01",X"01",X"01",X"11",X"3A",X"5D",X"83",X"98",X"93",X"88",X"83",X"88",X"78",
		X"5D",X"4A",X"37",X"2C",X"24",X"27",X"24",X"17",X"14",X"32",X"5D",X"80",X"90",X"90",X"93",X"93",
		X"93",X"90",X"8B",X"8B",X"8B",X"8B",X"90",X"93",X"93",X"98",X"98",X"9B",X"9B",X"9B",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9B",X"9E",X"9B",X"98",X"98",X"98",X"93",X"93",X"90",X"93",X"8B",
		X"88",X"75",X"52",X"37",X"1F",X"1C",X"27",X"37",X"4D",X"68",X"83",X"AE",X"E4",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"D1",X"9B",X"65",X"42",X"3A",X"52",X"80",X"AE",X"D4",X"E9",X"E4",X"C6",
		X"80",X"3A",X"11",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"32",X"88",X"C6",X"F7",X"FC",
		X"E4",X"CE",X"B9",X"A3",X"80",X"62",X"47",X"37",X"2F",X"2C",X"2F",X"37",X"3F",X"3A",X"32",X"3A",
		X"37",X"32",X"37",X"3A",X"52",X"7D",X"B3",X"DC",X"E4",X"E1",X"D1",X"D1",X"E1",X"FC",X"FC",X"FC",
		X"FC",X"F4",X"CE",X"A3",X"83",X"75",X"7D",X"83",X"83",X"88",X"98",X"A6",X"A6",X"98",X"88",X"75",
		X"68",X"5D",X"5A",X"5A",X"5A",X"62",X"65",X"68",X"6D",X"70",X"75",X"75",X"75",X"7D",X"83",X"83",
		X"80",X"75",X"68",X"70",X"80",X"8B",X"93",X"98",X"98",X"90",X"90",X"8B",X"90",X"98",X"A3",X"AE",
		X"B6",X"C9",X"C9",X"C1",X"B3",X"A3",X"98",X"8B",X"78",X"75",X"70",X"6D",X"65",X"68",X"70",X"80",
		X"83",X"83",X"88",X"8B",X"83",X"78",X"68",X"5D",X"52",X"42",X"2C",X"27",X"2C",X"3A",X"47",X"42",
		X"42",X"52",X"70",X"8B",X"A6",X"AB",X"A3",X"9E",X"9E",X"B3",X"B9",X"B9",X"BE",X"BE",X"B9",X"A3",
		X"88",X"68",X"5D",X"5A",X"5A",X"52",X"52",X"68",X"70",X"65",X"62",X"62",X"68",X"7D",X"8B",X"8B",
		X"83",X"75",X"65",X"68",X"75",X"80",X"9B",X"C1",X"EC",X"FC",X"FC",X"F7",X"EF",X"E9",X"D1",X"A3",
		X"78",X"5D",X"42",X"2C",X"14",X"0C",X"09",X"0C",X"0C",X"17",X"2C",X"47",X"62",X"75",X"75",X"68",
		X"62",X"52",X"4A",X"4A",X"42",X"3F",X"4A",X"55",X"68",X"90",X"A3",X"B9",X"C6",X"CE",X"E4",X"FC",
		X"FC",X"EC",X"E9",X"E9",X"DC",X"C1",X"B3",X"A6",X"98",X"75",X"52",X"3A",X"2C",X"1C",X"11",X"01",
		X"0C",X"1F",X"37",X"52",X"70",X"78",X"78",X"68",X"62",X"62",X"75",X"98",X"B6",X"BE",X"B3",X"AB",
		X"A6",X"9B",X"9E",X"AE",X"B9",X"C1",X"AE",X"90",X"5D",X"32",X"2C",X"27",X"2C",X"3F",X"62",X"83",
		X"93",X"90",X"88",X"80",X"70",X"5D",X"52",X"47",X"3A",X"2F",X"24",X"1F",X"2C",X"3A",X"68",X"A3",
		X"D4",X"F4",X"FC",X"FC",X"F4",X"E9",X"E9",X"DC",X"B9",X"90",X"78",X"68",X"5D",X"62",X"7D",X"93",
		X"9B",X"90",X"7D",X"70",X"5D",X"5A",X"52",X"52",X"52",X"55",X"5A",X"5D",X"65",X"68",X"68",X"70",
		X"70",X"75",X"78",X"78",X"7D",X"80",X"80",X"78",X"65",X"3F",X"27",X"17",X"1C",X"2C",X"3F",X"5D",
		X"78",X"93",X"AE",X"C6",X"DC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F7",X"A6",X"80",X"70",
		X"62",X"65",X"7D",X"98",X"A6",X"9B",X"80",X"62",X"32",X"04",X"01",X"01",X"01",X"01",X"01",X"11",
		X"3A",X"5D",X"83",X"98",X"93",X"88",X"83",X"88",X"78",X"5D",X"4A",X"37",X"2C",X"24",X"27",X"24",
		X"17",X"14",X"32",X"5D",X"80",X"90",X"90",X"93",X"93",X"93",X"90",X"8B",X"8B",X"8B",X"8B",X"90",
		X"93",X"93",X"98",X"98",X"9B",X"9B",X"9B",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9B",X"9E",
		X"9B",X"98",X"98",X"98",X"93",X"93",X"90",X"93",X"8B",X"88",X"75",X"52",X"37",X"1F",X"1C",X"24",
		X"37",X"4D",X"68",X"88",X"AE",X"E4",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"D4",X"9B",X"65",
		X"3F",X"37",X"52",X"80",X"B3",X"D9",X"EC",X"EC",X"C9",X"7D",X"37",X"04",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"27",X"88",X"D1",X"FC",X"FC",X"EC",X"D1",X"BE",X"A3",X"7D",X"62",X"3A",
		X"2C",X"1F",X"1F",X"24",X"2C",X"32",X"2C",X"27",X"2F",X"27",X"27",X"27",X"2C",X"47",X"7D",X"C1",
		X"F7",X"FC",X"FC",X"E9",X"E1",X"EC",X"FC",X"FC",X"FC",X"FC",X"FC",X"E4",X"AE",X"88",X"78",X"83",
		X"8B",X"8B",X"93",X"A3",X"B9",X"BE",X"A6",X"90",X"75",X"65",X"52",X"52",X"52",X"4D",X"55",X"5D",
		X"62",X"68",X"70",X"70",X"70",X"75",X"80",X"8B",X"90",X"90",X"8B",X"83",X"90",X"98",X"9B",X"9E",
		X"9E",X"9B",X"93",X"93",X"8B",X"90",X"8B",X"8B",X"8B",X"88",X"8B",X"8B",X"8B",X"8B",X"88",X"8B",
		X"8B",X"8B",X"8B",X"8B",X"8B",X"88",X"8B",X"88",X"88",X"88",X"88",X"83",X"83",X"80",X"80",X"80",
		X"80",X"7D",X"65",X"47",X"52",X"68",X"78",X"78",X"65",X"5A",X"5D",X"6D",X"75",X"78",X"70",X"68",
		X"70",X"90",X"C9",X"EC",X"FC",X"FC",X"FC",X"FC",X"E1",X"A6",X"68",X"42",X"3A",X"37",X"3A",X"5D",
		X"7D",X"83",X"68",X"55",X"52",X"47",X"32",X"17",X"09",X"01",X"01",X"09",X"17",X"2C",X"52",X"9B",
		X"E1",X"FC",X"FC",X"FC",X"FC",X"FC",X"F4",X"DC",X"A6",X"78",X"62",X"47",X"1F",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"3F",X"7D",X"A3",X"9B",X"80",X"5D",X"4A",X"5A",X"7D",X"90",X"9B",X"AB",
		X"A6",X"AB",X"AB",X"9E",X"A6",X"BE",X"D4",X"E4",X"D4",X"A6",X"88",X"7D",X"88",X"88",X"83",X"90",
		X"A3",X"AB",X"A6",X"9E",X"98",X"8B",X"83",X"80",X"80",X"80",X"83",X"83",X"88",X"8B",X"8B",X"90",
		X"90",X"90",X"93",X"98",X"98",X"9B",X"93",X"98",X"93",X"93",X"93",X"93",X"93",X"93",X"90",X"90",
		X"90",X"8B",X"8B",X"83",X"80",X"7D",X"68",X"52",X"52",X"62",X"68",X"88",X"AB",X"C6",X"C9",X"C9",
		X"B6",X"A6",X"9E",X"8B",X"83",X"8B",X"A3",X"B3",X"AE",X"98",X"80",X"6D",X"5D",X"52",X"47",X"42",
		X"47",X"3F",X"47",X"42",X"42",X"4D",X"62",X"65",X"68",X"68",X"68",X"68",X"68",X"68",X"68",X"68",
		X"65",X"68",X"68",X"68",X"6D",X"70",X"6D",X"6D",X"70",X"75",X"70",X"75",X"78",X"75",X"78",X"75",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"7D",X"80",X"80",X"6D",X"65",X"70",X"80",X"80",X"68",
		X"52",X"32",X"2C",X"37",X"68",X"9B",X"B6",X"B6",X"B6",X"C1",X"D4",X"D9",X"C6",X"A3",X"78",X"5A",
		X"3F",X"32",X"32",X"3A",X"55",X"8B",X"CE",X"FC",X"FC",X"FC",X"FC",X"FC",X"E1",X"A3",X"62",X"2F",
		X"1C",X"09",X"01",X"01",X"1C",X"47",X"5D",X"68",X"80",X"93",X"90",X"80",X"70",X"5A",X"4D",X"52",
		X"68",X"78",X"7D",X"70",X"5D",X"4A",X"3A",X"32",X"32",X"2F",X"27",X"27",X"1C",X"11",X"09",X"0C",
		X"14",X"2C",X"42",X"75",X"AB",X"DC",X"F7",X"FC",X"FC",X"F7",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"BE",X"88",X"4D",X"11",X"01",X"01",X"0C",X"3F",X"75",X"9E",X"B6",X"B3",
		X"93",X"70",X"52",X"3A",X"1F",X"11",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"24",X"3F",
		X"52",X"62",X"68",X"7D",X"9E",X"C1",X"E4",X"FC",X"FC",X"F7",X"E1",X"BE",X"A3",X"90",X"80",X"88",
		X"AB",X"E1",X"FC",X"FC",X"FC",X"FC",X"F7",X"BE",X"7D",X"3F",X"0C",X"01",X"01",X"01",X"01",X"27",
		X"70",X"B6",X"E9",X"FC",X"FC",X"E9",X"AE",X"83",X"62",X"4D",X"2F",X"04",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"3F",X"98",X"CE",X"D1",X"BE",X"B6",X"C1",X"D4",X"E9",X"FC",X"E9",X"C9",X"AB",
		X"9B",X"88",X"5D",X"37",X"27",X"27",X"1F",X"1C",X"1C",X"1F",X"37",X"70",X"B6",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"F4",X"F4",X"E4",X"C6",X"98",X"70",X"5A",X"3A",X"37",X"47",X"6D",X"AE",X"F7",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"CE",X"93",X"55",X"17",X"01",X"01",X"01",X"1C",X"4A",X"80",X"AB",
		X"B3",X"A6",X"A3",X"A3",X"A3",X"A6",X"9B",X"78",X"42",X"11",X"04",X"11",X"1C",X"1F",X"37",X"55",
		X"7D",X"8B",X"80",X"5D",X"47",X"4D",X"65",X"6D",X"5D",X"4A",X"3F",X"4D",X"7D",X"B6",X"EC",X"FC",
		X"FC",X"FC",X"E4",X"C6",X"9E",X"98",X"9B",X"90",X"75",X"5D",X"62",X"7D",X"9B",X"C6",X"E1",X"E9",
		X"D9",X"B3",X"93",X"83",X"70",X"68",X"5D",X"5A",X"52",X"52",X"52",X"55",X"5D",X"65",X"65",X"68",
		X"5A",X"37",X"2F",X"4A",X"65",X"6D",X"68",X"75",X"93",X"BE",X"E4",X"EC",X"D1",X"B3",X"9E",X"AB",
		X"AB",X"9E",X"80",X"65",X"42",X"32",X"32",X"4A",X"75",X"90",X"A3",X"BE",X"E4",X"FC",X"FC",X"FC",
		X"FC",X"D1",X"93",X"5A",X"3A",X"3A",X"47",X"5A",X"7D",X"A6",X"CE",X"CE",X"B9",X"A6",X"9B",X"80",
		X"52",X"1C",X"01",X"01",X"01",X"11",X"47",X"78",X"9E",X"AB",X"9B",X"78",X"5A",X"2C",X"14",X"1C",
		X"27",X"1F",X"11",X"01",X"01",X"01",X"1C",X"3F",X"75",X"AB",X"C9",X"D4",X"DC",X"CE",X"C9",X"D1",
		X"E1",X"F4",X"FC",X"FC",X"FC",X"E4",X"BE",X"90",X"70",X"4A",X"11",X"01",X"01",X"01",X"01",X"09",
		X"17",X"4A",X"90",X"D4",X"FC",X"FC",X"FC",X"F4",X"E9",X"E9",X"FC",X"FC",X"E4",X"B3",X"80",X"52",
		X"2F",X"1C",X"1F",X"32",X"68",X"AE",X"F4",X"FC",X"FC",X"FC",X"E4",X"C9",X"AB",X"80",X"5D",X"47",
		X"37",X"42",X"75",X"AB",X"DC",X"FC",X"FC",X"FC",X"D9",X"93",X"55",X"37",X"2F",X"3A",X"52",X"62",
		X"68",X"68",X"55",X"27",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1C",X"32",X"4D",X"68",
		X"9B",X"CE",X"E4",X"F4",X"EC",X"E4",X"E4",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"D9",
		X"88",X"4A",X"17",X"04",X"11",X"42",X"75",X"88",X"9B",X"B6",X"BE",X"A6",X"7D",X"4D",X"1C",X"01",
		X"01",X"17",X"27",X"32",X"4D",X"7D",X"A6",X"B3",X"B9",X"C6",X"D1",X"D9",X"D9",X"CE",X"BE",X"A6",
		X"90",X"65",X"27",X"01",X"01",X"01",X"01",X"01",X"01",X"14",X"68",X"93",X"98",X"83",X"75",X"7D",
		X"9E",X"BE",X"C9",X"BE",X"A6",X"9E",X"B6",X"D9",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"D9",X"C1",
		X"B3",X"9B",X"75",X"5D",X"47",X"2F",X"2F",X"4A",X"68",X"7D",X"7D",X"78",X"83",X"90",X"9E",X"AE",
		X"A3",X"83",X"75",X"52",X"3F",X"4A",X"5D",X"62",X"55",X"3F",X"2F",X"24",X"32",X"5A",X"7D",X"90",
		X"AB",X"CE",X"E4",X"FC",X"FC",X"FC",X"E9",X"CE",X"B3",X"98",X"88",X"83",X"83",X"90",X"B3",X"EC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"CE",X"75",X"42",X"27",X"14",X"01",X"01",X"1C",X"3F",X"52",X"5A",
		X"68",X"78",X"68",X"47",X"17",X"01",X"01",X"09",X"27",X"37",X"4A",X"65",X"75",X"6D",X"65",X"68",
		X"68",X"5D",X"4D",X"42",X"27",X"0C",X"0C",X"14",X"1C",X"1F",X"3A",X"68",X"9E",X"CE",X"E1",X"DC",
		X"DC",X"DC",X"DC",X"CE",X"A6",X"75",X"5A",X"4A",X"3A",X"4A",X"70",X"98",X"BE",X"E1",X"E9",X"E4",
		X"B9",X"9E",X"90",X"8B",X"88",X"75",X"52",X"2F",X"2F",X"4A",X"5D",X"68",X"78",X"80",X"70",X"70",
		X"7D",X"8B",X"9E",X"B6",X"BE",X"B6",X"AE",X"9B",X"98",X"AE",X"CE",X"E4",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"E4",X"B9",X"9E",X"88",X"65",X"4D",X"47",X"3F",X"2F",X"11",X"01",X"04",
		X"1F",X"2F",X"2F",X"1F",X"11",X"01",X"0C",X"2C",X"4D",X"62",X"78",X"98",X"AB",X"BE",X"DC",X"F4",
		X"F7",X"E4",X"E1",X"DC",X"C1",X"9E",X"88",X"62",X"3A",X"14",X"01",X"11",X"17",X"27",X"32",X"55",
		X"88",X"B6",X"E4",X"F7",X"E4",X"C6",X"A3",X"75",X"5A",X"52",X"5A",X"68",X"78",X"80",X"80",X"5A",
		X"27",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"11",X"3F",X"70",X"A3",X"C9",X"E1",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"DC",X"C6",X"B3",X"98",X"93",X"9B",X"AB",X"B9",X"AB",X"98",X"83",X"68",X"52",
		X"4A",X"2F",X"17",X"04",X"01",X"0C",X"37",X"75",X"A3",X"B9",X"D1",X"CE",X"B3",X"A3",X"9B",X"93",
		X"93",X"A6",X"BE",X"B9",X"9E",X"7D",X"55",X"37",X"27",X"27",X"4A",X"80",X"A6",X"B3",X"AE",X"AB",
		X"B9",X"C6",X"B9",X"B3",X"A3",X"80",X"5D",X"4A",X"47",X"3A",X"32",X"3A",X"5A",X"7D",X"83",X"90",
		X"8B",X"83",X"7D",X"70",X"65",X"6D",X"7D",X"78",X"65",X"47",X"1F",X"0C",X"01",X"01",X"09",X"2C",
		X"68",X"AE",X"CE",X"D1",X"CE",X"D4",X"E4",X"E4",X"CE",X"A6",X"98",X"9B",X"AB",X"BE",X"CE",X"CE",
		X"B9",X"90",X"52",X"14",X"01",X"01",X"01",X"01",X"09",X"3A",X"78",X"9E",X"AE",X"B9",X"CE",X"CE",
		X"B9",X"A6",X"90",X"7D",X"7D",X"83",X"80",X"68",X"55",X"52",X"4A",X"42",X"37",X"32",X"47",X"75",
		X"A6",X"C1",X"D1",X"D9",X"CE",X"C9",X"B6",X"9B",X"7D",X"62",X"4D",X"4D",X"6D",X"9E",X"D4",X"F4",
		X"EC",X"E4",X"CE",X"A3",X"78",X"65",X"5A",X"4A",X"37",X"2C",X"37",X"5D",X"93",X"C6",X"E9",X"FC",
		X"FC",X"D4",X"A6",X"88",X"75",X"68",X"52",X"27",X"01",X"01",X"01",X"01",X"01",X"11",X"5D",X"9B",
		X"C9",X"D1",X"C9",X"BE",X"B9",X"B9",X"B9",X"B6",X"AE",X"A3",X"98",X"83",X"70",X"4D",X"17",X"01",
		X"01",X"01",X"01",X"01",X"01",X"24",X"47",X"68",X"9B",X"DC",X"FC",X"FC",X"FC",X"FC",X"E9",X"F4",
		X"FC",X"FC",X"FC",X"E4",X"D4",X"C9",X"B3",X"9B",X"98",X"98",X"90",X"83",X"88",X"A6",X"C9",X"DC",
		X"D9",X"BE",X"AB",X"7D",X"52",X"2F",X"27",X"1F",X"11",X"17",X"27",X"2F",X"2F",X"3F",X"52",X"5D",
		X"5A",X"65",X"70",X"75",X"80",X"88",X"8B",X"9B",X"AB",X"BE",X"C6",X"AE",X"83",X"55",X"27",X"09",
		X"09",X"27",X"52",X"83",X"93",X"98",X"93",X"88",X"83",X"80",X"70",X"55",X"3F",X"2C",X"27",X"32",
		X"47",X"65",X"8B",X"AE",X"D4",X"E9",X"D9",X"B3",X"98",X"90",X"93",X"88",X"68",X"4D",X"4A",X"5A",
		X"68",X"6D",X"7D",X"8B",X"90",X"8B",X"88",X"8B",X"98",X"9E",X"9B",X"83",X"62",X"2F",X"09",X"04",
		X"1F",X"47",X"6D",X"98",X"AE",X"B6",X"B3",X"AB",X"9B",X"9B",X"A3",X"B6",X"C6",X"B9",X"9B",X"83",
		X"78",X"6D",X"65",X"5A",X"5A",X"68",X"88",X"A6",X"B6",X"A3",X"8B",X"75",X"68",X"6D",X"6D",X"65",
		X"5D",X"5D",X"68",X"80",X"A3",X"CE",X"DC",X"D4",X"CE",X"CE",X"C9",X"C6",X"CE",X"BE",X"AB",X"90",
		X"80",X"80",X"8B",X"98",X"9E",X"B6",X"DC",X"E4",X"E4",X"E1",X"CE",X"C6",X"B6",X"98",X"80",X"7D",
		X"75",X"70",X"68",X"68",X"62",X"3F",X"11",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"11",X"47",X"68",X"90",X"B6",X"CE",X"D4",X"E1",X"E9",X"E9",X"E4",X"E4",X"E9",X"E4",X"D4",X"C6",
		X"A6",X"78",X"42",X"14",X"01",X"01",X"01",X"01",X"14",X"42",X"78",X"AB",X"D1",X"E1",X"D9",X"C6",
		X"9B",X"7D",X"75",X"78",X"88",X"93",X"8B",X"88",X"70",X"4D",X"2F",X"24",X"1C",X"24",X"27",X"24",
		X"27",X"3A",X"62",X"88",X"B3",X"CE",X"DC",X"EC",X"EF",X"E1",X"CE",X"BE",X"A3",X"83",X"68",X"52",
		X"4D",X"55",X"65",X"78",X"78",X"80",X"90",X"90",X"90",X"8B",X"75",X"5D",X"4D",X"52",X"62",X"80",
		X"A3",X"B6",X"B6",X"B6",X"A6",X"90",X"83",X"88",X"93",X"9E",X"BE",X"D1",X"C9",X"AE",X"8B",X"62",
		X"3F",X"27",X"1C",X"32",X"62",X"88",X"9B",X"A3",X"AB",X"C1",X"CE",X"C1",X"B6",X"A6",X"90",X"6D",
		X"5D",X"55",X"3F",X"2F",X"2F",X"47",X"5D",X"65",X"6D",X"75",X"78",X"83",X"7D",X"75",X"7D",X"83",
		X"80",X"68",X"4D",X"2F",X"14",X"04",X"04",X"17",X"37",X"70",X"A6",X"C1",X"C1",X"B9",X"BE",X"D1",
		X"D4",X"C1",X"A3",X"98",X"9E",X"AE",X"C9",X"D4",X"D4",X"C6",X"98",X"5D",X"24",X"01",X"01",X"01",
		X"01",X"17",X"4A",X"7D",X"A3",X"AE",X"B9",X"C9",X"C6",X"B6",X"A3",X"8B",X"7D",X"80",X"83",X"83",
		X"6D",X"55",X"52",X"4A",X"42",X"37",X"32",X"47",X"75",X"A6",X"C1",X"D1",X"D9",X"CE",X"C9",X"B6",
		X"9B",X"7D",X"62",X"4D",X"4D",X"6D",X"9E",X"D4",X"F4",X"EC",X"E4",X"CE",X"A3",X"78",X"65",X"5A",
		X"4A",X"37",X"2C",X"37",X"5D",X"93",X"C6",X"E9",X"FC",X"FC",X"D4",X"A6",X"88",X"75",X"68",X"52",
		X"27",X"01",X"01",X"01",X"01",X"01",X"11",X"5D",X"9B",X"C9",X"D1",X"C9",X"BE",X"B9",X"B9",X"B9",
		X"B6",X"AE",X"A3",X"98",X"83",X"70",X"4D",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"24",X"47",
		X"68",X"9B",X"DC",X"FC",X"FC",X"FC",X"FC",X"E9",X"F4",X"FC",X"FC",X"FC",X"E4",X"D4",X"C9",X"B3",
		X"9B",X"98",X"98",X"8B",X"83",X"8B",X"A6",X"C9",X"E1",X"DC",X"C1",X"A6",X"7D",X"4D",X"2C",X"24",
		X"17",X"0C",X"11",X"1F",X"2C",X"2C",X"3A",X"52",X"5D",X"5A",X"65",X"70",X"78",X"88",X"90",X"90",
		X"9E",X"AB",X"C1",X"C6",X"A6",X"78",X"3F",X"11",X"01",X"01",X"14",X"47",X"80",X"93",X"98",X"93",
		X"83",X"70",X"65",X"4D",X"2F",X"14",X"04",X"04",X"27",X"47",X"70",X"A3",X"D1",X"FC",X"FC",X"F7",
		X"C9",X"A6",X"9B",X"9B",X"8B",X"70",X"5A",X"5D",X"75",X"7D",X"80",X"8B",X"9E",X"9B",X"93",X"8B",
		X"98",X"A3",X"AE",X"AE",X"93",X"68",X"32",X"04",X"04",X"24",X"52",X"88",X"B6",X"C9",X"B9",X"AB",
		X"98",X"80",X"80",X"90",X"A6",X"B9",X"BE",X"A6",X"93",X"8B",X"80",X"70",X"4D",X"37",X"3F",X"62",
		X"88",X"9E",X"98",X"80",X"65",X"55",X"62",X"68",X"68",X"70",X"75",X"78",X"93",X"C6",X"FC",X"FC",
		X"FC",X"FC",X"F7",X"E9",X"DC",X"D4",X"BE",X"A3",X"80",X"68",X"70",X"75",X"75",X"70",X"80",X"A3",
		X"B3",X"B3",X"AE",X"98",X"83",X"75",X"5D",X"52",X"5A",X"68",X"78",X"83",X"83",X"78",X"4A",X"11",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"37",X"78",X"A6",X"D1",X"E9",X"E4",
		X"E1",X"E1",X"DC",X"D9",X"E9",X"FC",X"FC",X"FC",X"FC",X"EF",X"B9",X"75",X"2F",X"01",X"01",X"01",
		X"01",X"01",X"01",X"27",X"5D",X"9B",X"D4",X"F4",X"EC",X"CE",X"A6",X"93",X"9E",X"B6",X"B6",X"A3",
		X"93",X"8B",X"83",X"70",X"68",X"78",X"93",X"A6",X"9E",X"90",X"83",X"98",X"AE",X"C9",X"D4",X"DC",
		X"CE",X"A6",X"7D",X"65",X"52",X"2C",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"11",X"4D",X"9E",
		X"E4",X"FC",X"FC",X"FC",X"EC",X"EC",X"FC",X"FC",X"FC",X"FC",X"E9",X"AE",X"78",X"4A",X"2F",X"2F",
		X"52",X"8B",X"C6",X"F4",X"FC",X"F7",X"DC",X"B3",X"80",X"4D",X"17",X"01",X"01",X"01",X"1C",X"3F",
		X"70",X"A6",X"D1",X"E9",X"E1",X"CE",X"B9",X"B3",X"AE",X"A6",X"88",X"5A",X"1F",X"01",X"01",X"01",
		X"01",X"01",X"14",X"52",X"8B",X"B9",X"C6",X"B6",X"A6",X"9E",X"90",X"75",X"68",X"52",X"4A",X"52",
		X"68",X"88",X"93",X"83",X"62",X"3F",X"1F",X"17",X"2F",X"4D",X"68",X"75",X"83",X"9E",X"D1",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"D4",X"BE",X"B3",X"A3",X"A6",X"BE",X"D4",X"E1",X"CE",X"B3",X"A6",X"98",
		X"75",X"4A",X"27",X"1C",X"2F",X"4D",X"68",X"7D",X"68",X"47",X"17",X"01",X"01",X"01",X"01",X"01",
		X"04",X"0C",X"1F",X"32",X"4A",X"5D",X"80",X"B3",X"F7",X"FC",X"FC",X"FC",X"EC",X"D4",X"CE",X"BE",
		X"C1",X"CE",X"D9",X"C9",X"A3",X"83",X"70",X"5A",X"3F",X"32",X"3F",X"5D",X"68",X"65",X"47",X"2C",
		X"17",X"04",X"09",X"27",X"4A",X"68",X"90",X"9E",X"98",X"88",X"7D",X"83",X"9E",X"CE",X"E9",X"F7",
		X"E4",X"BE",X"9E",X"68",X"37",X"09",X"01",X"01",X"01",X"04",X"14",X"37",X"55",X"65",X"70",X"88",
		X"AE",X"DC",X"FC",X"F4",X"D1",X"AE",X"93",X"80",X"78",X"83",X"9B",X"B3",X"B3",X"98",X"70",X"47",
		X"24",X"17",X"32",X"62",X"9B",X"C9",X"CE",X"B9",X"A3",X"9B",X"88",X"70",X"5D",X"55",X"68",X"93",
		X"B6",X"BE",X"B3",X"AE",X"AE",X"A3",X"90",X"90",X"98",X"9B",X"AB",X"AB",X"AE",X"B3",X"AB",X"93",
		X"78",X"65",X"68",X"78",X"75",X"70",X"68",X"78",X"8B",X"93",X"93",X"9E",X"B9",X"DC",X"FC",X"FC",
		X"FC",X"D4",X"93",X"62",X"42",X"1C",X"01",X"01",X"04",X"0C",X"0C",X"1F",X"4A",X"78",X"AB",X"C9",
		X"DC",X"E1",X"D9",X"C6",X"AB",X"90",X"70",X"47",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"1C",X"47",X"62",X"75",X"88",X"AB",X"D1",X"E9",X"EC",X"E9",X"E4",X"DC",X"F7",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"E4",X"9E",X"80",X"75",X"7D",X"70",X"6D",X"75",X"80",X"8B",X"80",X"65",
		X"4A",X"2C",X"04",X"01",X"01",X"01",X"04",X"2C",X"52",X"62",X"5A",X"4D",X"5A",X"78",X"9B",X"B3",
		X"C1",X"AB",X"93",X"83",X"78",X"62",X"4D",X"4A",X"52",X"4A",X"3F",X"4D",X"5D",X"7D",X"90",X"9B",
		X"9E",X"83",X"68",X"62",X"5D",X"68",X"78",X"88",X"88",X"8B",X"8B",X"80",X"62",X"47",X"3F",X"3A",
		X"32",X"37",X"37",X"37",X"4D",X"70",X"88",X"8B",X"80",X"70",X"70",X"8B",X"B6",X"D4",X"D4",X"CE",
		X"B9",X"B9",X"C9",X"C9",X"C6",X"B6",X"B9",X"D4",X"FC",X"FC",X"FC",X"FC",X"EC",X"B6",X"80",X"52",
		X"37",X"2F",X"2C",X"37",X"62",X"98",X"D1",X"FC",X"FC",X"EC",X"D1",X"A3",X"68",X"4A",X"32",X"27",
		X"27",X"3A",X"55",X"68",X"62",X"52",X"3F",X"1C",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"37",
		X"5A",X"70",X"88",X"88",X"7D",X"65",X"52",X"47",X"52",X"68",X"83",X"9E",X"AE",X"B6",X"C1",X"B9",
		X"B6",X"AE",X"98",X"78",X"5D",X"42",X"32",X"2C",X"2F",X"4D",X"7D",X"B9",X"F7",X"FC",X"FC",X"FC",
		X"E1",X"AB",X"83",X"65",X"52",X"5A",X"68",X"65",X"52",X"3F",X"3F",X"3F",X"37",X"37",X"52",X"7D",
		X"A6",X"C1",X"BE",X"9E",X"88",X"7D",X"68",X"5A",X"47",X"47",X"62",X"90",X"B3",X"C6",X"D9",X"EF",
		X"FC",X"FC",X"E4",X"CE",X"B9",X"B3",X"B3",X"AE",X"AB",X"9B",X"75",X"55",X"37",X"11",X"01",X"01",
		X"01",X"01",X"04",X"4D",X"88",X"AB",X"B3",X"AE",X"A3",X"9B",X"AE",X"C6",X"CE",X"C9",X"BE",X"B6",
		X"B3",X"AB",X"AE",X"C6",X"EF",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"CE",X"88",X"4A",X"14",X"01",
		X"09",X"2C",X"52",X"78",X"93",X"93",X"78",X"47",X"0C",X"01",X"01",X"01",X"01",X"09",X"09",X"11",
		X"27",X"4D",X"62",X"68",X"7D",X"90",X"9E",X"AE",X"AB",X"8B",X"70",X"62",X"52",X"3A",X"1C",X"04",
		X"11",X"2F",X"5A",X"83",X"9E",X"B3",X"B9",X"B9",X"AB",X"80",X"62",X"4D",X"4D",X"5A",X"65",X"75",
		X"7D",X"83",X"83",X"70",X"4D",X"1F",X"0C",X"14",X"32",X"5D",X"70",X"68",X"65",X"68",X"83",X"9E",
		X"9E",X"93",X"88",X"83",X"9B",X"BE",X"D9",X"E1",X"D1",X"B6",X"A3",X"93",X"88",X"88",X"8B",X"98",
		X"A3",X"C6",X"FC",X"FC",X"FC",X"FC",X"FC",X"F4",X"D4",X"B3",X"88",X"65",X"4A",X"32",X"3A",X"5D",
		X"88",X"B3",X"D4",X"E4",X"E1",X"B9",X"78",X"37",X"11",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"14",X"37",X"42",X"4A",X"5A",X"68",X"78",X"90",X"AE",X"C9",X"E1",X"E1",
		X"C9",X"93",X"65",X"4D",X"32",X"1F",X"17",X"27",X"37",X"3F",X"42",X"4D",X"68",X"88",X"98",X"A3",
		X"B6",X"C9",X"D4",X"E4",X"E4",X"D4",X"BE",X"A6",X"AE",X"C6",X"E4",X"FC",X"FC",X"FC",X"E4",X"AB",
		X"6D",X"3F",X"27",X"2F",X"52",X"83",X"AB",X"AB",X"AE",X"AE",X"AE",X"98",X"70",X"5A",X"5A",X"65",
		X"7D",X"88",X"80",X"5D",X"3A",X"24",X"11",X"11",X"2F",X"52",X"75",X"83",X"93",X"A3",X"C9",X"EF",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"D4",X"98",X"5A",X"1F",X"01",X"01",X"01",X"11",X"2F",
		X"5D",X"90",X"BE",X"E4",X"FC",X"FC",X"D9",X"A3",X"78",X"65",X"68",X"75",X"70",X"65",X"5A",X"4A",
		X"2C",X"14",X"04",X"11",X"37",X"68",X"9B",X"A6",X"9B",X"88",X"83",X"90",X"93",X"90",X"8B",X"83",
		X"7D",X"83",X"93",X"A6",X"B6",X"BE",X"B9",X"9E",X"68",X"42",X"2C",X"2F",X"47",X"5D",X"78",X"88",
		X"90",X"93",X"90",X"70",X"52",X"37",X"17",X"11",X"17",X"2C",X"37",X"3F",X"4D",X"4A",X"3F",X"32",
		X"2F",X"37",X"5A",X"7D",X"9B",X"9E",X"A6",X"AE",X"B6",X"D4",X"FC",X"FC",X"FC",X"FC",X"FC",X"EC",
		X"E1",X"B9",X"93",X"6D",X"5A",X"5A",X"5D",X"68",X"75",X"78",X"83",X"83",X"83",X"83",X"70",X"5D",
		X"4A",X"4D",X"62",X"7D",X"90",X"98",X"88",X"62",X"2F",X"01",X"01",X"01",X"01",X"1C",X"37",X"52",
		X"65",X"68",X"5A",X"52",X"5D",X"75",X"7D",X"75",X"5D",X"4A",X"4D",X"65",X"88",X"AB",X"C6",X"D9",
		X"D4",X"B6",X"93",X"83",X"70",X"5A",X"47",X"47",X"4A",X"3F",X"3A",X"3F",X"32",X"27",X"17",X"1F",
		X"3F",X"68",X"93",X"9E",X"9B",X"93",X"98",X"A6",X"AB",X"AB",X"A3",X"A6",X"BE",X"E1",X"F7",X"FC",
		X"FC",X"EC",X"D1",X"AE",X"93",X"8B",X"9B",X"B3",X"B6",X"B6",X"C6",X"C6",X"B6",X"A6",X"9E",X"93",
		X"7D",X"5D",X"37",X"1C",X"1F",X"27",X"2C",X"37",X"52",X"75",X"93",X"98",X"8B",X"7D",X"65",X"5D",
		X"65",X"75",X"88",X"9B",X"9E",X"9B",X"8B",X"80",X"83",X"8B",X"8B",X"83",X"93",X"AB",X"C9",X"DC",
		X"CE",X"B9",X"A6",X"83",X"5D",X"32",X"17",X"01",X"01",X"04",X"1C",X"4A",X"80",X"B6",X"DC",X"E1",
		X"D4",X"BE",X"A6",X"98",X"90",X"88",X"6D",X"4D",X"2C",X"11",X"04",X"04",X"1C",X"4D",X"83",X"B6",
		X"DC",X"E4",X"D1",X"C1",X"B3",X"9B",X"80",X"68",X"68",X"68",X"75",X"7D",X"7D",X"70",X"52",X"2C",
		X"04",X"01",X"01",X"01",X"11",X"2F",X"47",X"5D",X"78",X"A3",X"D4",X"EC",X"FC",X"FC",X"F7",X"EC",
		X"EF",X"EC",X"D4",X"C9",X"C6",X"B9",X"9E",X"80",X"65",X"68",X"70",X"78",X"7D",X"80",X"93",X"9E",
		X"AB",X"AE",X"AE",X"A3",X"8B",X"68",X"52",X"42",X"32",X"27",X"1C",X"14",X"09",X"01",X"01",X"01",
		X"14",X"3F",X"78",X"A3",X"AE",X"AE",X"A3",X"A6",X"BE",X"D4",X"D9",X"D9",X"D9",X"C6",X"B9",X"AB",
		X"93",X"78",X"65",X"62",X"68",X"70",X"80",X"8B",X"88",X"7D",X"70",X"6D",X"78",X"7D",X"78",X"70",
		X"6D",X"83",X"9E",X"C1",X"CE",X"C1",X"B3",X"98",X"75",X"52",X"3F",X"47",X"5A",X"68",X"7D",X"88",
		X"7D",X"62",X"47",X"2F",X"11",X"01",X"01",X"01",X"01",X"01",X"17",X"3F",X"65",X"78",X"93",X"9B",
		X"9E",X"93",X"98",X"9B",X"98",X"A3",X"A6",X"AB",X"B3",X"C1",X"D1",X"CE",X"BE",X"AE",X"98",X"7D",
		X"75",X"65",X"52",X"4A",X"3F",X"3A",X"3F",X"52",X"68",X"80",X"93",X"AB",X"B6",X"C9",X"E1",X"E4",
		X"D4",X"CE",X"CE",X"C9",X"BE",X"9E",X"7D",X"5A",X"37",X"27",X"1C",X"1F",X"37",X"5A",X"75",X"80",
		X"8B",X"93",X"90",X"8B",X"88",X"88",X"80",X"80",X"83",X"80",X"88",X"A3",X"C6",X"E1",X"FC",X"FC",
		X"F4",X"CE",X"A3",X"80",X"65",X"4A",X"37",X"37",X"3F",X"47",X"52",X"62",X"70",X"7D",X"70",X"62",
		X"52",X"55",X"68",X"78",X"80",X"75",X"65",X"65",X"5D",X"55",X"5A",X"5A",X"65",X"80",X"98",X"A3",
		X"9B",X"8B",X"7D",X"80",X"88",X"90",X"98",X"9B",X"93",X"93",X"9E",X"AE",X"B9",X"B6",X"AE",X"AE",
		X"A6",X"93",X"78",X"65",X"52",X"4D",X"4A",X"52",X"68",X"78",X"88",X"93",X"90",X"83",X"80",X"6D",
		X"5D",X"5D",X"62",X"68",X"6D",X"6D",X"5D",X"4A",X"37",X"2F",X"32",X"52",X"75",X"93",X"A6",X"AE",
		X"AB",X"AE",X"B6",X"C6",X"BE",X"C1",X"B9",X"A6",X"98",X"8B",X"70",X"52",X"3A",X"2C",X"37",X"42",
		X"5A",X"68",X"70",X"78",X"7D",X"88",X"93",X"98",X"90",X"7D",X"7D",X"88",X"90",X"98",X"93",X"7D",
		X"52",X"2C",X"09",X"01",X"01",X"09",X"32",X"52",X"70",X"88",X"9B",X"93",X"90",X"93",X"98",X"90",
		X"83",X"70",X"65",X"62",X"78",X"93",X"AE",X"BE",X"C6",X"B9",X"9E",X"83",X"70",X"65",X"5D",X"5A",
		X"5A",X"5D",X"5A",X"55",X"55",X"47",X"37",X"27",X"1F",X"37",X"5A",X"78",X"88",X"8B",X"8B",X"93",
		X"A3",X"A6",X"AB",X"A6",X"AB",X"BE",X"D4",X"E4",X"EC",X"EC",X"E1",X"C9",X"A6",X"90",X"83",X"90",
		X"98",X"9B",X"9E",X"AE",X"AB",X"A6",X"9E",X"9B",X"9B",X"90",X"78",X"5A",X"3F",X"37",X"37",X"37",
		X"3F",X"52",X"68",X"88",X"83",X"78",X"68",X"5A",X"55",X"65",X"78",X"8B",X"9E",X"A3",X"9B",X"90",
		X"83",X"88",X"8B",X"88",X"80",X"8B",X"9E",X"B9",X"C9",X"B9",X"A6",X"93",X"75",X"52",X"32",X"1C",
		X"11",X"0C",X"14",X"2C",X"5A",X"8B",X"BE",X"DC",X"E1",X"D9",X"C6",X"AE",X"9E",X"98",X"8B",X"75",
		X"55",X"32",X"1C",X"11",X"11",X"24",X"52",X"88",X"B6",X"D9",X"E4",X"CE",X"BE",X"AE",X"98",X"7D",
		X"68",X"65",X"68",X"75",X"78",X"7D",X"70",X"52",X"2F",X"09",X"01",X"01",X"01",X"11",X"2F",X"47",
		X"5A",X"78",X"A3",X"D4",X"EC",X"FC",X"FC",X"F7",X"EC",X"EF",X"EC",X"D4",X"C9",X"C6",X"B9",X"9E",
		X"80",X"65",X"68",X"70",X"78",X"7D",X"80",X"93",X"9E",X"AB",X"AE",X"AE",X"A3",X"8B",X"68",X"52",
		X"42",X"32",X"27",X"1C",X"14",X"09",X"01",X"01",X"01",X"14",X"3F",X"78",X"A3",X"AE",X"AE",X"A3",
		X"A6",X"BE",X"D4",X"D9",X"D9",X"D9",X"C6",X"B9",X"AB",X"93",X"78",X"65",X"62",X"68",X"70",X"80",
		X"8B",X"88",X"7D",X"70",X"6D",X"78",X"7D",X"78",X"70",X"6D",X"83",X"9E",X"C1",X"CE",X"C1",X"B3",
		X"98",X"75",X"52",X"3F",X"47",X"5A",X"68",X"7D",X"88",X"7D",X"62",X"47",X"2C",X"0C",X"01",X"01",
		X"01",X"01",X"01",X"14",X"3A",X"65",X"7D",X"98",X"A3",X"A3",X"98",X"9B",X"9E",X"9E",X"A6",X"AB",
		X"AB",X"B6",X"C6",X"D4",X"CE",X"BE",X"AB",X"90",X"78",X"68",X"5A",X"47",X"32",X"27",X"1F",X"24",
		X"3A",X"62",X"80",X"9E",X"B9",X"CE",X"D4",X"E9",X"EC",X"E1",X"D1",X"D1",X"CE",X"C6",X"A6",X"80",
		X"55",X"2F",X"17",X"04",X"11",X"2F",X"62",X"83",X"9B",X"A6",X"AB",X"9B",X"90",X"8B",X"88",X"78",
		X"70",X"65",X"5A",X"65",X"88",X"A6",X"CE",X"EF",X"FC",X"FC",X"E1",X"B6",X"9E",X"88",X"68",X"52",
		X"4A",X"47",X"3F",X"37",X"3A",X"47",X"47",X"3A",X"2F",X"2F",X"4A",X"68",X"80",X"83",X"75",X"65",
		X"65",X"65",X"68",X"75",X"7D",X"88",X"9E",X"AB",X"AB",X"98",X"80",X"78",X"7D",X"80",X"8B",X"9E",
		X"9E",X"9B",X"9E",X"AE",X"BE",X"C1",X"B3",X"A6",X"A3",X"A6",X"AB",X"9B",X"83",X"68",X"52",X"42",
		X"3F",X"52",X"68",X"80",X"93",X"A3",X"A6",X"B3",X"A6",X"93",X"88",X"88",X"93",X"90",X"83",X"68",
		X"4D",X"37",X"2C",X"2F",X"47",X"68",X"90",X"AB",X"AE",X"A6",X"A6",X"9B",X"88",X"75",X"68",X"62",
		X"52",X"42",X"32",X"27",X"11",X"01",X"01",X"11",X"27",X"3F",X"5A",X"65",X"68",X"78",X"8B",X"A6",
		X"C1",X"C6",X"B9",X"B3",X"B3",X"AB",X"A3",X"8B",X"68",X"42",X"24",X"11",X"11",X"11",X"27",X"4D",
		X"70",X"98",X"B9",X"DC",X"E9",X"E9",X"E1",X"CE",X"AB",X"98",X"90",X"83",X"83",X"93",X"A3",X"B6",
		X"AE",X"A3",X"90",X"78",X"5D",X"4A",X"4D",X"62",X"78",X"83",X"80",X"80",X"83",X"7D",X"68",X"52",
		X"37",X"1F",X"1F",X"2F",X"47",X"55",X"65",X"7D",X"90",X"93",X"98",X"A3",X"AE",X"B3",X"B9",X"B6",
		X"B6",X"C1",X"C6",X"B9",X"A6",X"8B",X"80",X"70",X"65",X"52",X"4A",X"52",X"62",X"65",X"68",X"7D",
		X"90",X"AB",X"C6",X"D1",X"CE",X"AE",X"88",X"68",X"65",X"62",X"52",X"52",X"4D",X"3F",X"2F",X"27",
		X"27",X"3A",X"62",X"83",X"9E",X"B3",X"A6",X"9E",X"93",X"90",X"8B",X"7D",X"68",X"62",X"65",X"65",
		X"65",X"55",X"3F",X"27",X"14",X"11",X"14",X"1C",X"2F",X"4A",X"62",X"78",X"98",X"B6",X"D1",X"E4",
		X"E4",X"E1",X"E4",X"F7",X"FC",X"F7",X"E4",X"D1",X"BE",X"AB",X"98",X"83",X"8B",X"98",X"93",X"90",
		X"93",X"90",X"83",X"78",X"70",X"6D",X"62",X"4A",X"2C",X"17",X"14",X"1C",X"27",X"3F",X"4D",X"5D",
		X"68",X"68",X"68",X"68",X"75",X"8B",X"9E",X"A6",X"9E",X"9B",X"98",X"98",X"93",X"80",X"70",X"62",
		X"52",X"4A",X"42",X"3A",X"2F",X"27",X"2C",X"2F",X"3F",X"5D",X"80",X"90",X"9B",X"A3",X"AE",X"C9",
		X"E1",X"E4",X"DC",X"CE",X"C9",X"CE",X"C6",X"B3",X"98",X"8B",X"83",X"75",X"68",X"6D",X"7D",X"90",
		X"A3",X"B3",X"B9",X"AE",X"98",X"7D",X"70",X"62",X"4A",X"2F",X"17",X"11",X"17",X"24",X"37",X"52",
		X"62",X"75",X"80",X"80",X"80",X"88",X"8B",X"8B",X"98",X"9B",X"9E",X"AB",X"B6",X"AE",X"A3",X"90",
		X"83",X"80",X"7D",X"83",X"90",X"90",X"88",X"75",X"62",X"52",X"47",X"42",X"4A",X"5D",X"75",X"8B",
		X"A3",X"AB",X"AB",X"A3",X"93",X"98",X"9E",X"AE",X"BE",X"BE",X"AB",X"88",X"68",X"52",X"3A",X"37",
		X"47",X"62",X"83",X"98",X"A3",X"9B",X"98",X"98",X"88",X"68",X"52",X"4D",X"52",X"62",X"65",X"62",
		X"62",X"5D",X"4A",X"37",X"27",X"2C",X"3F",X"5D",X"6D",X"75",X"75",X"80",X"90",X"A3",X"B3",X"BE",
		X"C6",X"C1",X"B9",X"AB",X"9E",X"83",X"68",X"52",X"3F",X"27",X"11",X"0C",X"11",X"1C",X"3F",X"68",
		X"9B",X"B6",X"BE",X"B6",X"B3",X"B6",X"BE",X"C9",X"C6",X"AE",X"9B",X"8B",X"80",X"7D",X"83",X"93",
		X"A3",X"AE",X"A3",X"9E",X"9B",X"9E",X"9E",X"9E",X"9E",X"93",X"7D",X"68",X"62",X"5D",X"62",X"5D",
		X"52",X"4D",X"5A",X"52",X"52",X"52",X"52",X"52",X"5A",X"5A",X"5A",X"62",X"68",X"78",X"88",X"90",
		X"98",X"A6",X"B6",X"B9",X"B6",X"B3",X"B6",X"B9",X"B9",X"B6",X"AE",X"AB",X"93",X"78",X"65",X"4D",
		X"32",X"24",X"24",X"32",X"52",X"70",X"83",X"88",X"83",X"7D",X"70",X"65",X"68",X"6D",X"6D",X"6D",
		X"68",X"65",X"68",X"68",X"65",X"5D",X"55",X"5D",X"70",X"8B",X"90",X"93",X"8B",X"80",X"7D",X"7D",
		X"8B",X"9E",X"A6",X"A3",X"9E",X"9E",X"A3",X"A3",X"98",X"88",X"80",X"75",X"68",X"62",X"55",X"4D",
		X"4A",X"4D",X"5D",X"75",X"93",X"AE",X"B6",X"AB",X"93",X"78",X"65",X"52",X"5A",X"5D",X"65",X"78",
		X"88",X"88",X"80",X"75",X"70",X"68",X"5D",X"5A",X"5D",X"62",X"68",X"70",X"75",X"78",X"7D",X"7D",
		X"80",X"78",X"70",X"65",X"5D",X"52",X"5A",X"70",X"8B",X"A3",X"AE",X"AE",X"A6",X"9B",X"90",X"83",
		X"75",X"68",X"55",X"4D",X"4A",X"4A",X"4D",X"5A",X"78",X"93",X"B9",X"D4",X"E4",X"E1",X"CE",X"BE",
		X"AE",X"9B",X"88",X"78",X"78",X"78",X"78",X"68",X"62",X"55",X"4D",X"3A",X"32",X"3A",X"4D",X"68",
		X"7D",X"80",X"7D",X"78",X"75",X"7D",X"88",X"98",X"A3",X"AE",X"AE",X"AB",X"AE",X"B6",X"C6",X"D1",
		X"D4",X"D4",X"C6",X"AB",X"98",X"83",X"78",X"65",X"4D",X"3F",X"3F",X"3F",X"4A",X"5A",X"68",X"70",
		X"68",X"68",X"70",X"80",X"8B",X"93",X"8B",X"7D",X"70",X"6D",X"68",X"70",X"75",X"75",X"78",X"78",
		X"75",X"68",X"65",X"62",X"6D",X"83",X"98",X"AE",X"B6",X"A6",X"98",X"90",X"80",X"75",X"68",X"5D",
		X"62",X"68",X"80",X"93",X"9B",X"93",X"90",X"80",X"6D",X"5A",X"4A",X"42",X"47",X"52",X"5D",X"6D",
		X"83",X"90",X"90",X"83",X"80",X"80",X"75",X"75",X"70",X"68",X"65",X"5A",X"52",X"4D",X"52",X"65",
		X"7D",X"98",X"A6",X"AB",X"AB",X"A6",X"9E",X"9B",X"90",X"80",X"75",X"6D",X"65",X"52",X"52",X"52",
		X"52",X"4D",X"42",X"3F",X"47",X"4A",X"55",X"5D",X"62",X"62",X"62",X"62",X"68",X"7D",X"88",X"93",
		X"A3",X"9E",X"A3",X"98",X"90",X"90",X"98",X"A3",X"B6",X"C1",X"BE",X"B6",X"B3",X"AB",X"9B",X"88",
		X"75",X"70",X"68",X"65",X"70",X"78",X"7D",X"70",X"68",X"68",X"68",X"68",X"65",X"62",X"5D",X"68",
		X"7D",X"90",X"9B",X"9B",X"98",X"98",X"98",X"93",X"98",X"9E",X"9B",X"98",X"93",X"93",X"90",X"83",
		X"80",X"80",X"78",X"68",X"62",X"62",X"65",X"75",X"83",X"88",X"8B",X"90",X"8B",X"7D",X"70",X"68",
		X"65",X"5D",X"55",X"52",X"4D",X"4A",X"4D",X"5A",X"5D",X"65",X"70",X"80",X"8B",X"93",X"9E",X"9E",
		X"9B",X"9E",X"A3",X"9B",X"98",X"90",X"88",X"83",X"83",X"88",X"90",X"A6",X"B9",X"BE",X"C1",X"C6",
		X"C6",X"C6",X"B6",X"9B",X"83",X"65",X"52",X"4A",X"4D",X"5D",X"6D",X"80",X"8B",X"93",X"8B",X"80",
		X"65",X"5A",X"52",X"52",X"52",X"47",X"3F",X"3A",X"47",X"52",X"5D",X"6D",X"83",X"93",X"9B",X"9E",
		X"98",X"8B",X"88",X"80",X"80",X"78",X"6D",X"68",X"68",X"70",X"70",X"68",X"68",X"62",X"5A",X"5A",
		X"5D",X"5A",X"5D",X"65",X"70",X"75",X"8B",X"98",X"9B",X"9B",X"9B",X"93",X"88",X"88",X"83",X"88",
		X"88",X"93",X"9B",X"98",X"8B",X"80",X"78",X"70",X"68",X"68",X"70",X"80",X"88",X"90",X"93",X"9B",
		X"9E",X"98",X"98",X"98",X"98",X"90",X"83",X"78",X"78",X"6D",X"6D",X"78",X"88",X"98",X"A3",X"AB",
		X"AB",X"A6",X"98",X"83",X"70",X"52",X"47",X"37",X"32",X"27",X"27",X"37",X"47",X"4D",X"65",X"75",
		X"88",X"90",X"98",X"90",X"83",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"68",X"62",X"5D",X"4D",X"42",
		X"3A",X"3A",X"3F",X"47",X"52",X"5A",X"68",X"78",X"83",X"90",X"A3",X"AE",X"B6",X"B9",X"B6",X"AE",
		X"B3",X"B6",X"C1",X"C6",X"BE",X"B9",X"B9",X"AE",X"9B",X"88",X"80",X"75",X"68",X"65",X"65",X"70",
		X"78",X"83",X"8B",X"90",X"88",X"7D",X"65",X"5A",X"55",X"5A",X"52",X"4D",X"47",X"42",X"3F",X"47",
		X"4A",X"52",X"65",X"7D",X"93",X"9B",X"98",X"93",X"90",X"93",X"9B",X"A6",X"AE",X"AE",X"A6",X"98",
		X"8B",X"78",X"68",X"5A",X"52",X"52",X"5A",X"65",X"68",X"75",X"75",X"70",X"70",X"7D",X"80",X"83",
		X"83",X"80",X"80",X"80",X"8B",X"98",X"A3",X"A3",X"A6",X"A3",X"9B",X"93",X"90",X"8B",X"88",X"80",
		X"78",X"70",X"62",X"5A",X"5A",X"52",X"52",X"55",X"5A",X"62",X"68",X"75",X"70",X"6D",X"65",X"65",
		X"68",X"6D",X"70",X"70",X"70",X"75",X"75",X"7D",X"83",X"88",X"93",X"9B",X"A3",X"A3",X"A6",X"A6",
		X"A3",X"9E",X"93",X"88",X"80",X"78",X"78",X"78",X"7D",X"80",X"80",X"80",X"7D",X"70",X"68",X"62",
		X"62",X"68",X"70",X"78",X"7D",X"7D",X"78",X"75",X"68",X"68",X"62",X"62",X"68",X"78",X"78",X"7D",
		X"75",X"68",X"6D",X"6D",X"70",X"75",X"7D",X"83",X"80",X"80",X"80",X"83",X"83",X"80",X"80",X"83",
		X"88",X"8B",X"88",X"83",X"80",X"80",X"83",X"8B",X"98",X"9E",X"9E",X"9E",X"9B",X"90",X"83",X"7D",
		X"75",X"6D",X"68",X"75",X"80",X"83",X"88",X"8B",X"90",X"8B",X"83",X"7D",X"75",X"75",X"78",X"7D",
		X"80",X"80",X"75",X"68",X"5D",X"52",X"4A",X"4D",X"52",X"5D",X"68",X"6D",X"78",X"80",X"88",X"8B",
		X"98",X"9B",X"A3",X"A3",X"9B",X"93",X"8B",X"88",X"7D",X"70",X"68",X"65",X"65",X"62",X"62",X"62",
		X"65",X"70",X"78",X"7D",X"80",X"88",X"8B",X"93",X"93",X"90",X"8B",X"88",X"80",X"83",X"88",X"90",
		X"9E",X"9E",X"9B",X"9B",X"93",X"88",X"7D",X"7D",X"7D",X"78",X"7D",X"78",X"75",X"78",X"7D",X"7D",
		X"7D",X"80",X"80",X"80",X"7D",X"78",X"78",X"75",X"70",X"70",X"6D",X"68",X"6D",X"70",X"78",X"80",
		X"80",X"80",X"83",X"88",X"90",X"8B",X"8B",X"8B",X"88",X"80",X"7D",X"78",X"70",X"68",X"68",X"68",
		X"68",X"6D",X"6D",X"70",X"78",X"7D",X"83",X"8B",X"8B",X"90",X"8B",X"88",X"88",X"88",X"88",X"83",
		X"80",X"80",X"83",X"80",X"80",X"7D",X"83",X"83",X"7D",X"7D",X"78",X"75",X"75",X"75",X"78",X"78",
		X"75",X"70",X"70",X"70",X"75",X"78",X"78",X"78",X"75",X"75",X"70",X"70",X"75",X"78",X"75",X"75",
		X"75",X"75",X"78",X"7D",X"80",X"7D",X"7D",X"7D",X"83",X"88",X"8B",X"88",X"88",X"88",X"88",X"88",
		X"8B",X"90",X"90",X"88",X"83",X"7D",X"7D",X"78",X"75",X"75",X"75",X"7D",X"7D",X"80",X"7D",X"78",
		X"75",X"70",X"70",X"78",X"80",X"88",X"88",X"88",X"88",X"83",X"7D",X"78",X"78",X"80",X"83",X"83",
		X"83",X"80",X"78",X"75",X"75",X"75",X"78",X"80",X"80",X"83",X"83",X"80",X"7D",X"78",X"6D",X"68",
		X"65",X"62",X"5D",X"5A",X"62",X"65",X"68",X"75",X"80",X"8B",X"90",X"93",X"90",X"88",X"83",X"80",
		X"78",X"75",X"75",X"70",X"68",X"65",X"5D",X"5D",X"55",X"5A",X"5D",X"65",X"68",X"75",X"75",X"80",
		X"83",X"8B",X"90",X"9B",X"A3",X"A6",X"A6",X"9E",X"9B",X"98",X"98",X"9E",X"9E",X"A3",X"A3",X"A6",
		X"A3",X"9B",X"8B",X"88",X"7D",X"75",X"6D",X"68",X"6D",X"75",X"7D",X"7D",X"83",X"83",X"80",X"75",
		X"6D",X"68",X"68",X"68",X"65",X"62",X"5D",X"5A",X"5A",X"5D",X"62",X"68",X"78",X"80",X"83",X"80",
		X"7D",X"80",X"83",X"8B",X"98",X"9B",X"9B",X"98",X"90",X"8B",X"7D",X"70",X"68",X"62",X"65",X"68",
		X"70",X"78",X"80",X"80",X"80",X"80",X"83",X"83",X"83",X"80",X"7D",X"7D",X"7D",X"83",X"90",X"98",
		X"9B",X"9E",X"9B",X"98",X"90",X"8B",X"83",X"83",X"7D",X"75",X"70",X"65",X"5D",X"5D",X"5A",X"5D",
		X"62",X"65",X"68",X"75",X"75",X"75",X"75",X"68",X"6D",X"6D",X"70",X"70",X"75",X"70",X"75",X"75",
		X"78",X"7D",X"83",X"90",X"98",X"9B",X"9B",X"9E",X"9E",X"9E",X"9E",X"93",X"88",X"83",X"7D",X"7D",
		X"7D",X"80",X"83",X"80",X"80",X"7D",X"75",X"68",X"65",X"65",X"68",X"75",X"78",X"7D",X"78",X"78",
		X"78",X"6D",X"68",X"65",X"68",X"6D",X"78",X"7D",X"7D",X"75",X"6D",X"6D",X"70",X"75",X"78",X"80",
		X"83",X"80",X"80",X"80",X"83",X"83",X"80",X"83",X"83",X"88",X"8B",X"88",X"83",X"80",X"80",X"83",
		X"8B",X"98",X"9E",X"9E",X"9E",X"9B",X"90",X"83",X"7D",X"75",X"6D",X"68",X"75",X"80",X"83",X"88",
		X"8B",X"90",X"8B",X"83",X"7D",X"75",X"75",X"78",X"7D",X"80",X"80",X"75",X"68",X"5D",X"52",X"4A",
		X"4D",X"52",X"5D",X"68",X"6D",X"78",X"80",X"88",X"8B",X"98",X"9B",X"A3",X"A3",X"9B",X"93",X"8B",
		X"88",X"7D",X"70",X"68",X"65",X"65",X"62",X"62",X"62",X"65",X"70",X"78",X"7D",X"80",X"88",X"8B",
		X"93",X"93",X"90",X"8B",X"88",X"80",X"83",X"88",X"90",X"9E",X"9E",X"9B",X"9B",X"93",X"88",X"7D",
		X"7D",X"7D",X"78",X"7D",X"78",X"75",X"78",X"7D",X"7D",X"7D",X"80",X"80",X"80",X"78",X"78",X"75",
		X"75",X"70",X"75",X"6D",X"68",X"6D",X"70",X"78",X"80",X"83",X"80",X"83",X"88",X"90",X"8B",X"8B",
		X"88",X"83",X"7D",X"78",X"75",X"6D",X"68",X"68",X"68",X"65",X"68",X"68",X"68",X"70",X"75",X"7D",
		X"88",X"83",X"88",X"88",X"80",X"83",X"83",X"88",X"8B",X"88",X"88",X"88",X"83",X"80",X"7D",X"80",
		X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"80",X"80",X"80",X"7D",X"75",X"75",X"75",X"75",X"70",
		X"70",X"68",X"68",X"68",X"68",X"70",X"70",X"75",X"75",X"75",X"75",X"78",X"83",X"83",X"83",X"88",
		X"88",X"90",X"98",X"98",X"93",X"90",X"90",X"8B",X"88",X"88",X"8B",X"88",X"80",X"78",X"78",X"75",
		X"70",X"68",X"68",X"65",X"68",X"70",X"78",X"78",X"78",X"75",X"75",X"70",X"78",X"80",X"83",X"83",
		X"80",X"7D",X"70",X"68",X"65",X"68",X"70",X"7D",X"83",X"83",X"83",X"80",X"75",X"70",X"68",X"65",
		X"65",X"65",X"68",X"6D",X"70",X"78",X"7D",X"7D",X"7D",X"83",X"80",X"80",X"80",X"80",X"7D",X"7D",
		X"80",X"83",X"8B",X"90",X"93",X"93",X"8B",X"83",X"7D",X"78",X"70",X"6D",X"68",X"65",X"65",X"62",
		X"65",X"68",X"70",X"7D",X"88",X"88",X"93",X"90",X"90",X"90",X"90",X"93",X"93",X"93",X"98",X"90",
		X"88",X"80",X"78",X"78",X"75",X"78",X"80",X"88",X"90",X"90",X"93",X"8B",X"8B",X"88",X"7D",X"78",
		X"6D",X"65",X"65",X"68",X"6D",X"75",X"80",X"83",X"88",X"88",X"88",X"83",X"83",X"83",X"83",X"80",
		X"7D",X"80",X"7D",X"75",X"6D",X"68",X"5D",X"55",X"52",X"52",X"62",X"68",X"70",X"75",X"75",X"75",
		X"78",X"7D",X"83",X"80",X"83",X"83",X"83",X"83",X"88",X"8B",X"90",X"98",X"98",X"9B",X"9B",X"93",
		X"8B",X"83",X"7D",X"78",X"78",X"70",X"75",X"7D",X"80",X"80",X"83",X"80",X"80",X"75",X"70",X"68",
		X"68",X"68",X"65",X"68",X"68",X"65",X"68",X"70",X"78",X"7D",X"88",X"88",X"88",X"83",X"83",X"80",
		X"80",X"80",X"80",X"7D",X"7D",X"75",X"75",X"68",X"68",X"68",X"68",X"6D",X"6D",X"70",X"70",X"75",
		X"75",X"7D",X"83",X"83",X"88",X"83",X"88",X"83",X"88",X"83",X"83",X"8B",X"88",X"8B",X"88",X"88",
		X"80",X"7D",X"7D",X"75",X"6D",X"68",X"6D",X"70",X"7D",X"80",X"7D",X"83",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"83",X"80",X"80",X"7D",X"7D",X"80",X"80",
		X"83",X"83",X"80",X"80",X"7D",X"78",X"75",X"70",X"68",X"6D",X"75",X"78",X"7D",X"80",X"80",X"80",
		X"7D",X"78",X"7D",X"7D",X"80",X"80",X"80",X"80",X"7D",X"80",X"83",X"88",X"88",X"8B",X"8B",X"8B",
		X"8B",X"88",X"83",X"83",X"80",X"78",X"75",X"75",X"70",X"70",X"75",X"75",X"80",X"83",X"80",X"83",
		X"83",X"83",X"83",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"75",X"75",X"75",X"70",X"70",
		X"75",X"75",X"78",X"7D",X"7D",X"80",X"80",X"83",X"83",X"83",X"83",X"88",X"83",X"83",X"83",X"88",
		X"83",X"83",X"88",X"8B",X"88",X"88",X"80",X"7D",X"7D",X"7D",X"7D",X"80",X"7D",X"80",X"80",X"80",
		X"83",X"83",X"83",X"7D",X"7D",X"75",X"75",X"75",X"75",X"75",X"70",X"75",X"75",X"75",X"78",X"83",
		X"80",X"83",X"80",X"7D",X"80",X"78",X"78",X"80",X"80",X"80",X"7D",X"80",X"80",X"80",X"7D",X"75",
		X"70",X"68",X"68",X"68",X"68",X"68",X"70",X"75",X"7D",X"83",X"8B",X"90",X"90",X"8B",X"83",X"80",
		X"7D",X"7D",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"75",X"75",X"75",X"70",X"70",X"75",X"75",
		X"78",X"7D",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"75",X"78",X"7D",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"78",X"78",X"78",X"7D",X"80",X"80",X"80",X"83",X"83",
		X"8B",X"8B",X"8B",X"88",X"83",X"83",X"80",X"83",X"7D",X"7D",X"7D",X"7D",X"75",X"75",X"78",X"7D",
		X"80",X"80",X"78",X"78",X"78",X"78",X"7D",X"78",X"7D",X"7D",X"78",X"7D",X"78",X"7D",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"78",X"78",X"7D",X"7D",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"78",X"78",
		X"78",X"78",X"78",X"78",X"7D",X"80",X"78",X"80",X"80",X"78",X"78",X"78",X"78",X"7D",X"78",X"7D",
		X"78",X"78",X"7D",X"78",X"78",X"78",X"75",X"78",X"78",X"7D",X"78",X"7D",X"80",X"78",X"7D",X"7D",
		X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"78",X"78",X"78",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"78",X"78",X"7D",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"78",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"80",X"80",X"7D",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"80",
		X"75",X"75",X"75",X"75",X"78",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"75",X"75",X"78",X"80",
		X"80",X"80",X"80",X"80",X"80",X"75",X"75",X"75",X"75",X"83",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7D",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"80",X"88",X"83",
		X"80",X"80",X"7D",X"78",X"75",X"78",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7D",X"7D",X"7D",X"75",X"75",X"75",X"75",X"78",X"83",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"75",X"78",X"75",X"75",X"78",
		X"75",X"78",X"78",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"83",X"83",X"80",X"80",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"83",X"83",X"83",X"83",X"83",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"78",X"78",X"78",X"75",X"75",X"75",X"70",X"75",X"75",X"7D",X"7D",X"80",X"80",X"80",
		X"80",X"80",X"83",X"83",X"83",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"80",X"78",X"78",X"7D",
		X"78",X"7D",X"80",X"80",X"80",X"80",X"80",X"7D",X"80",X"7D",X"7D",X"7D",X"7D",X"78",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"75",X"78",X"78",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"83",
		X"83",X"83",X"88",X"83",X"83",X"83",X"83",X"83",X"83",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"78",
		X"7D",X"78",X"7D",X"80",X"80",X"80",X"80",X"7D",X"7D",X"80",X"7D",X"78",X"78",X"78",X"75",X"75",
		X"75",X"78",X"7D",X"78",X"83",X"80",X"80",X"80",X"80",X"7D",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"78",X"78",X"78",X"78",X"75",X"75",X"75",X"75",X"78",X"7D",X"7D",X"7D",X"80",X"80",X"80",X"80",
		X"83",X"83",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"78",X"78",X"78",X"78",
		X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"7D",X"7D",X"80",X"83",X"83",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"83",X"80",X"83",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"80",X"80",X"80",X"83",X"83",X"83",X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"78",
		X"78",X"78",X"7D",X"78",X"7D",X"7D",X"80",X"80",X"80",X"80",X"7D",X"78",X"7D",X"78",X"78",X"7D",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"78",X"78",X"78",X"7D",X"7D",X"7D",
		X"7D",X"80",X"80",X"80",X"80",X"80",X"83",X"80",X"80",X"83",X"80",X"80",X"83",X"7D",X"7D",X"7D",
		X"7D",X"78",X"78",X"78",X"7D",X"7D",X"7D",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7D",X"80",X"80",X"83",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7D",X"7D",X"7D",X"78",X"7D",X"78",X"78",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7D",X"7D",X"78",X"7D",X"78",X"7D",X"80",X"80",X"80",X"80",X"80",X"7D",X"78",X"7D",
		X"7D",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"78",X"78",X"78",X"7D",X"78",X"78",X"7D",
		X"7D",X"80",X"80",X"80",X"80",X"83",X"83",X"83",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"78",
		X"78",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",X"7D",X"7D",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"78",
		X"7D",X"78",X"7D",X"80",X"80",X"80",X"80",X"7D",X"80",X"83",X"80",X"80",X"80",X"80",X"80",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
