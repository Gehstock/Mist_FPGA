library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps03 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps03 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"10",X"22",X"70",X"20",X"CD",X"42",X"0B",X"23",X"CD",X"1F",X"0B",X"C2",X"26",X"10",X"2A",X"70",
		X"20",X"23",X"22",X"70",X"20",X"21",X"73",X"20",X"11",X"73",X"40",X"06",X"06",X"C3",X"BB",X"04",
		X"35",X"C9",X"21",X"13",X"43",X"C9",X"E5",X"2A",X"70",X"20",X"23",X"22",X"70",X"20",X"E1",X"CD",
		X"3A",X"0B",X"22",X"77",X"20",X"2A",X"77",X"20",X"CD",X"6B",X"10",X"3A",X"77",X"20",X"FE",X"38",
		X"DA",X"15",X"10",X"CD",X"4A",X"0B",X"22",X"75",X"20",X"21",X"75",X"20",X"EF",X"2A",X"77",X"20",
		X"E5",X"7D",X"FE",X"78",X"3E",X"01",X"DA",X"5B",X"10",X"3E",X"02",X"F5",X"FF",X"F1",X"11",X"02",
		X"02",X"DF",X"E1",X"06",X"03",X"11",X"10",X"43",X"C3",X"AC",X"03",X"E5",X"7D",X"FE",X"78",X"D2",
		X"E9",X"08",X"CD",X"C5",X"0F",X"C3",X"E9",X"08",X"CD",X"D2",X"08",X"C0",X"2E",X"7B",X"BE",X"C8",
		X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"C1",X"10",X"34",X"2A",X"79",X"20",X"4E",X"7D",
		X"FE",X"22",X"CC",X"22",X"10",X"22",X"79",X"20",X"CD",X"42",X"0B",X"23",X"CD",X"1F",X"0B",X"C2",
		X"B2",X"10",X"2A",X"79",X"20",X"23",X"22",X"79",X"20",X"21",X"7C",X"20",X"11",X"7C",X"40",X"C3",
		X"1B",X"10",X"E5",X"2A",X"79",X"20",X"23",X"22",X"79",X"20",X"E1",X"CD",X"3A",X"0B",X"22",X"80",
		X"20",X"2A",X"80",X"20",X"CD",X"6B",X"10",X"3A",X"80",X"20",X"FE",X"38",X"DA",X"A9",X"10",X"CD",
		X"4A",X"0B",X"22",X"7E",X"20",X"21",X"7E",X"20",X"EF",X"2A",X"80",X"20",X"C3",X"50",X"10",X"CD",
		X"D2",X"08",X"C0",X"2E",X"84",X"BE",X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"28",
		X"11",X"34",X"2A",X"82",X"20",X"4E",X"7D",X"FE",X"32",X"CC",X"22",X"10",X"22",X"82",X"20",X"CD",
		X"46",X"0B",X"23",X"CD",X"1F",X"0B",X"C2",X"19",X"11",X"2A",X"82",X"20",X"23",X"22",X"82",X"20",
		X"21",X"85",X"20",X"11",X"85",X"40",X"C3",X"1B",X"10",X"E5",X"2A",X"82",X"20",X"23",X"22",X"82",
		X"20",X"E1",X"CD",X"3A",X"0B",X"22",X"89",X"20",X"2A",X"89",X"20",X"CD",X"6B",X"10",X"3A",X"89",
		X"20",X"FE",X"38",X"DA",X"10",X"11",X"CD",X"4A",X"0B",X"22",X"87",X"20",X"21",X"87",X"20",X"EF",
		X"2A",X"89",X"20",X"C3",X"50",X"10",X"CD",X"D2",X"08",X"C0",X"2E",X"8D",X"BE",X"C8",X"23",X"BE",
		X"C2",X"20",X"10",X"23",X"BE",X"C2",X"8F",X"11",X"34",X"2A",X"8B",X"20",X"4E",X"7D",X"FE",X"32",
		X"CC",X"22",X"10",X"22",X"8B",X"20",X"CD",X"46",X"0B",X"23",X"CD",X"1F",X"0B",X"C2",X"80",X"11",
		X"2A",X"8B",X"20",X"23",X"22",X"8B",X"20",X"21",X"8E",X"20",X"11",X"8E",X"40",X"C3",X"1B",X"10",
		X"E5",X"2A",X"8B",X"20",X"23",X"22",X"8B",X"20",X"E1",X"CD",X"3A",X"0B",X"22",X"92",X"20",X"2A",
		X"92",X"20",X"CD",X"6B",X"10",X"3A",X"92",X"20",X"FE",X"38",X"DA",X"77",X"11",X"CD",X"4A",X"0B",
		X"22",X"90",X"20",X"21",X"90",X"20",X"EF",X"2A",X"92",X"20",X"C3",X"50",X"10",X"CD",X"D2",X"08",
		X"C0",X"2E",X"BE",X"BE",X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"CA",X"11",X"34",
		X"CD",X"D8",X"08",X"23",X"CD",X"DC",X"08",X"22",X"C3",X"20",X"CD",X"04",X"12",X"22",X"C1",X"20",
		X"2A",X"C3",X"20",X"CD",X"F0",X"11",X"3A",X"C3",X"20",X"FE",X"74",X"D2",X"FB",X"11",X"21",X"C1",
		X"20",X"EF",X"2A",X"C3",X"20",X"CD",X"D6",X"0F",X"06",X"05",X"11",X"E4",X"44",X"C3",X"AC",X"03",
		X"CD",X"C5",X"0F",X"06",X"05",X"11",X"E4",X"44",X"C3",X"EF",X"08",X"21",X"BF",X"20",X"11",X"BF",
		X"40",X"C3",X"1B",X"10",X"CD",X"ED",X"0E",X"FE",X"22",X"21",X"06",X"00",X"D0",X"FE",X"18",X"2E",
		X"05",X"D0",X"FE",X"13",X"2E",X"04",X"D0",X"FE",X"10",X"2E",X"03",X"D0",X"FE",X"07",X"2E",X"02",
		X"D0",X"2E",X"01",X"C9",X"CD",X"D2",X"08",X"C0",X"2E",X"C5",X"BE",X"C8",X"23",X"BE",X"C2",X"20",
		X"10",X"23",X"BE",X"C2",X"40",X"12",X"34",X"E7",X"2E",X"3D",X"CD",X"DC",X"08",X"22",X"CA",X"20",
		X"CD",X"74",X"12",X"22",X"C8",X"20",X"2A",X"CA",X"20",X"CD",X"F0",X"11",X"3A",X"CA",X"20",X"FE",
		X"74",X"D2",X"5E",X"12",X"21",X"C8",X"20",X"EF",X"2A",X"CA",X"20",X"C3",X"E5",X"11",X"E7",X"2E",
		X"3D",X"AF",X"BE",X"C2",X"6B",X"12",X"21",X"C5",X"20",X"36",X"00",X"21",X"C6",X"20",X"11",X"C6",
		X"40",X"C3",X"1B",X"10",X"CD",X"ED",X"0E",X"FE",X"22",X"21",X"06",X"00",X"D0",X"FE",X"18",X"2E",
		X"05",X"D0",X"FE",X"14",X"2E",X"04",X"D0",X"FE",X"11",X"2E",X"03",X"D0",X"FE",X"08",X"2E",X"02",
		X"D0",X"2E",X"01",X"C9",X"CD",X"D2",X"08",X"C0",X"2E",X"CC",X"BE",X"C8",X"23",X"BE",X"C2",X"20",
		X"10",X"23",X"BE",X"C2",X"B0",X"12",X"34",X"E7",X"2E",X"40",X"CD",X"DC",X"08",X"22",X"D1",X"20",
		X"CD",X"E4",X"12",X"22",X"CF",X"20",X"2A",X"D1",X"20",X"CD",X"F0",X"11",X"3A",X"D1",X"20",X"FE",
		X"74",X"D2",X"CE",X"12",X"21",X"CF",X"20",X"EF",X"2A",X"D1",X"20",X"C3",X"E5",X"11",X"E7",X"2E",
		X"40",X"AF",X"BE",X"C2",X"DB",X"12",X"21",X"CC",X"20",X"36",X"00",X"21",X"CD",X"20",X"11",X"CD",
		X"40",X"C3",X"1B",X"10",X"CD",X"ED",X"0E",X"FE",X"22",X"21",X"06",X"00",X"D0",X"FE",X"18",X"2E",
		X"05",X"D0",X"FE",X"15",X"2E",X"04",X"D0",X"FE",X"12",X"2E",X"03",X"D0",X"FE",X"09",X"2E",X"02",
		X"D0",X"2E",X"01",X"C9",X"21",X"51",X"20",X"AF",X"BE",X"C8",X"2E",X"52",X"BE",X"2E",X"57",X"3A",
		X"05",X"20",X"C2",X"1A",X"13",X"BE",X"DA",X"1F",X"13",X"C9",X"BE",X"D2",X"1F",X"13",X"C9",X"2E",
		X"A9",X"06",X"01",X"70",X"2E",X"B0",X"70",X"2E",X"B7",X"70",X"C9",X"21",X"A9",X"20",X"AF",X"BE",
		X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"42",X"13",X"34",X"CD",X"6B",X"13",X"22",
		X"AE",X"20",X"CD",X"1B",X"14",X"22",X"AC",X"20",X"2A",X"AE",X"20",X"CD",X"7D",X"13",X"CD",X"86",
		X"13",X"3A",X"AE",X"20",X"FE",X"35",X"DA",X"8E",X"13",X"21",X"AC",X"20",X"EF",X"2A",X"AE",X"20",
		X"CD",X"CF",X"0F",X"11",X"E1",X"44",X"06",X"03",X"C3",X"AC",X"03",X"2A",X"56",X"20",X"3A",X"52",
		X"20",X"A7",X"01",X"04",X"12",X"C2",X"7B",X"13",X"01",X"04",X"FB",X"09",X"C9",X"7D",X"FE",X"74",
		X"D2",X"CF",X"0F",X"C3",X"C5",X"0F",X"11",X"E1",X"44",X"06",X"03",X"C3",X"EF",X"08",X"21",X"A9",
		X"20",X"11",X"A9",X"40",X"06",X"07",X"C3",X"BB",X"04",X"21",X"B0",X"20",X"AF",X"BE",X"C8",X"23",
		X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"B0",X"13",X"34",X"CD",X"6B",X"13",X"22",X"B5",X"20",
		X"CD",X"1B",X"14",X"22",X"B3",X"20",X"2A",X"B5",X"20",X"CD",X"7D",X"13",X"CD",X"86",X"13",X"3A",
		X"B5",X"20",X"FE",X"35",X"DA",X"D1",X"13",X"21",X"B3",X"20",X"EF",X"2A",X"B5",X"20",X"C3",X"60",
		X"13",X"21",X"B0",X"20",X"11",X"B0",X"40",X"C3",X"94",X"13",X"21",X"B7",X"20",X"AF",X"BE",X"C8",
		X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"F1",X"13",X"34",X"CD",X"6B",X"13",X"22",X"BC",
		X"20",X"CD",X"1B",X"14",X"22",X"BA",X"20",X"2A",X"BC",X"20",X"CD",X"7D",X"13",X"CD",X"86",X"13",
		X"3A",X"BC",X"20",X"FE",X"35",X"DA",X"12",X"14",X"21",X"BA",X"20",X"EF",X"2A",X"BC",X"20",X"C3",
		X"60",X"13",X"21",X"B7",X"20",X"11",X"B7",X"40",X"C3",X"94",X"13",X"CD",X"ED",X"0E",X"FE",X"23",
		X"21",X"F9",X"00",X"D0",X"FE",X"18",X"2E",X"FA",X"D0",X"FE",X"10",X"2E",X"FB",X"D0",X"FE",X"06",
		X"2E",X"FC",X"D0",X"FE",X"03",X"2E",X"FD",X"D0",X"2E",X"FE",X"C9",X"36",X"00",X"DB",X"02",X"E6",
		X"08",X"C2",X"3E",X"01",X"CD",X"51",X"07",X"21",X"0C",X"23",X"AF",X"BE",X"C2",X"68",X"14",X"CD",
		X"E4",X"08",X"35",X"CA",X"7C",X"02",X"CD",X"33",X"02",X"CD",X"15",X"02",X"CD",X"A0",X"04",X"CD",
		X"85",X"03",X"CD",X"0F",X"4C",X"C3",X"24",X"01",X"E7",X"0F",X"D2",X"97",X"14",X"CD",X"E4",X"08",
		X"35",X"C2",X"BE",X"14",X"CD",X"49",X"02",X"21",X"07",X"39",X"3E",X"1D",X"CD",X"FA",X"14",X"CD",
		X"F7",X"01",X"CD",X"73",X"03",X"21",X"03",X"23",X"36",X"22",X"CD",X"E4",X"08",X"A7",X"C2",X"CD",
		X"14",X"CD",X"F0",X"04",X"C3",X"7F",X"02",X"CD",X"E4",X"08",X"35",X"C2",X"E3",X"14",X"CD",X"49",
		X"02",X"21",X"07",X"39",X"3E",X"1E",X"CD",X"FA",X"14",X"CD",X"F7",X"01",X"CD",X"73",X"03",X"21",
		X"03",X"23",X"36",X"21",X"CD",X"E4",X"08",X"A7",X"C2",X"DB",X"14",X"C3",X"91",X"14",X"CD",X"33",
		X"02",X"21",X"03",X"23",X"36",X"22",X"CD",X"E4",X"08",X"A7",X"CA",X"DB",X"14",X"21",X"03",X"23",
		X"36",X"22",X"CD",X"F0",X"04",X"CD",X"67",X"02",X"C3",X"59",X"14",X"21",X"03",X"23",X"36",X"21",
		X"C3",X"D2",X"14",X"CD",X"33",X"02",X"21",X"03",X"23",X"36",X"21",X"CD",X"E4",X"08",X"A7",X"C2",
		X"DB",X"14",X"21",X"03",X"23",X"36",X"22",X"C3",X"CD",X"14",X"CD",X"F2",X"02",X"21",X"07",X"C8",
		X"11",X"01",X"26",X"3E",X"06",X"DF",X"C9",X"01",X"03",X"00",X"09",X"C9",X"CD",X"ED",X"0E",X"21",
		X"D3",X"20",X"FE",X"18",X"36",X"06",X"D0",X"FE",X"14",X"36",X"0A",X"D0",X"36",X"10",X"FE",X"10",
		X"D0",X"FE",X"07",X"36",X"20",X"D0",X"FE",X"05",X"36",X"30",X"D0",X"FE",X"03",X"36",X"40",X"D0",
		X"36",X"50",X"C9",X"CD",X"48",X"16",X"CD",X"ED",X"0E",X"C6",X"01",X"27",X"77",X"E7",X"2E",X"00",
		X"06",X"4E",X"11",X"00",X"41",X"CD",X"BB",X"04",X"CD",X"15",X"02",X"CD",X"64",X"15",X"CD",X"6E",
		X"03",X"CD",X"CB",X"07",X"CD",X"A0",X"04",X"C3",X"24",X"01",X"06",X"4E",X"C3",X"22",X"02",X"06",
		X"4E",X"C3",X"2D",X"02",X"CD",X"ED",X"0E",X"FE",X"28",X"D2",X"00",X"16",X"FE",X"25",X"CA",X"07",
		X"16",X"FE",X"22",X"CA",X"0E",X"16",X"FE",X"19",X"CA",X"15",X"16",X"FE",X"16",X"CA",X"1C",X"16",
		X"FE",X"13",X"CA",X"23",X"16",X"FE",X"10",X"CA",X"2A",X"16",X"FE",X"07",X"CA",X"31",X"16",X"FE",
		X"04",X"C0",X"3E",X"1D",X"06",X"01",X"C5",X"F5",X"21",X"12",X"CA",X"11",X"01",X"20",X"3E",X"06",
		X"DF",X"CD",X"6E",X"03",X"21",X"12",X"2A",X"11",X"F1",X"15",X"0E",X"06",X"CD",X"54",X"03",X"F1",
		X"CD",X"F2",X"02",X"0E",X"09",X"11",X"F7",X"15",X"CD",X"54",X"03",X"CD",X"85",X"03",X"C1",X"2E",
		X"00",X"60",X"CD",X"F0",X"18",X"06",X"00",X"CD",X"CD",X"07",X"11",X"4F",X"4E",X"CD",X"41",X"4E",
		X"21",X"4A",X"20",X"34",X"2E",X"0A",X"34",X"CD",X"D4",X"01",X"2E",X"4A",X"7E",X"A7",X"D3",X"05",
		X"C2",X"DA",X"15",X"CD",X"D9",X"01",X"21",X"0A",X"20",X"36",X"00",X"CD",X"55",X"16",X"C3",X"6E",
		X"03",X"01",X"0E",X"0D",X"14",X"12",X"1B",X"1C",X"1C",X"1C",X"1B",X"0F",X"0E",X"08",X"0D",X"13",
		X"3E",X"25",X"06",X"09",X"C3",X"96",X"15",X"3E",X"24",X"06",X"08",X"C3",X"96",X"15",X"3E",X"23",
		X"06",X"07",X"C3",X"96",X"15",X"3E",X"22",X"06",X"06",X"C3",X"96",X"15",X"3E",X"21",X"06",X"05",
		X"C3",X"96",X"15",X"3E",X"20",X"06",X"04",X"C3",X"96",X"15",X"3E",X"1F",X"06",X"03",X"C3",X"96",
		X"15",X"3E",X"1E",X"06",X"02",X"C3",X"96",X"15",X"21",X"F1",X"20",X"AF",X"BE",X"06",X"FE",X"CA",
		X"3D",X"09",X"35",X"06",X"01",X"C3",X"2E",X"09",X"CD",X"D9",X"01",X"06",X"A0",X"CD",X"3D",X"09",
		X"06",X"20",X"CD",X"47",X"09",X"CD",X"3E",X"4E",X"C3",X"0E",X"4E",X"21",X"F2",X"20",X"97",X"BE",
		X"06",X"FD",X"CA",X"3D",X"09",X"35",X"06",X"02",X"C3",X"2E",X"09",X"21",X"51",X"20",X"AF",X"BE",
		X"06",X"FB",X"CA",X"3D",X"09",X"06",X"04",X"C3",X"2E",X"09",X"21",X"E5",X"20",X"97",X"BE",X"06",
		X"FC",X"CA",X"47",X"09",X"2E",X"E8",X"7E",X"FE",X"FB",X"06",X"03",X"CA",X"51",X"09",X"A7",X"06",
		X"FE",X"CA",X"47",X"09",X"06",X"02",X"C3",X"51",X"09",X"21",X"F3",X"20",X"AF",X"BE",X"06",X"F7",
		X"CA",X"3D",X"09",X"35",X"06",X"08",X"C3",X"2E",X"09",X"3A",X"0A",X"23",X"FE",X"18",X"06",X"04",
		X"D2",X"56",X"09",X"06",X"FB",X"C3",X"47",X"09",X"06",X"EF",X"C3",X"47",X"09",X"C0",X"23",X"BE",
		X"C0",X"23",X"BE",X"C0",X"06",X"F7",X"C3",X"47",X"09",X"21",X"F4",X"20",X"97",X"BE",X"CA",X"B8",
		X"16",X"35",X"06",X"10",X"C3",X"51",X"09",X"21",X"F5",X"20",X"AF",X"BE",X"CA",X"99",X"16",X"35",
		X"06",X"08",X"C3",X"2E",X"09",X"21",X"F6",X"20",X"97",X"BE",X"CA",X"C4",X"16",X"35",X"06",X"08",
		X"C3",X"51",X"09",X"3A",X"3D",X"20",X"FE",X"12",X"21",X"3E",X"20",X"36",X"40",X"D2",X"39",X"17",
		X"FE",X"0C",X"36",X"50",X"D2",X"47",X"17",X"FE",X"06",X"36",X"60",X"D2",X"59",X"17",X"36",X"7B",
		X"C9",X"21",X"09",X"C4",X"11",X"05",X"02",X"3E",X"00",X"DF",X"C9",X"21",X"09",X"24",X"CD",X"2A",
		X"17",X"21",X"0B",X"24",X"CD",X"2A",X"17",X"21",X"0D",X"24",X"06",X"07",X"11",X"32",X"17",X"C3",
		X"DB",X"03",X"38",X"38",X"38",X"FE",X"7C",X"38",X"10",X"CD",X"11",X"17",X"CD",X"1B",X"17",X"E7",
		X"2E",X"2D",X"36",X"01",X"C3",X"4D",X"17",X"CD",X"11",X"17",X"CD",X"21",X"17",X"E7",X"2E",X"2A",
		X"06",X"01",X"70",X"2E",X"36",X"70",X"C3",X"5F",X"17",X"CD",X"11",X"17",X"CD",X"27",X"17",X"E7",
		X"2E",X"26",X"06",X"01",X"70",X"2E",X"32",X"70",X"C9",X"21",X"23",X"20",X"AF",X"BE",X"C8",X"23",
		X"34",X"7E",X"E6",X"02",X"C2",X"8B",X"17",X"2A",X"25",X"20",X"E5",X"FF",X"3E",X"02",X"11",X"02",
		X"03",X"DF",X"E1",X"11",X"49",X"45",X"06",X"08",X"C3",X"E9",X"03",X"2A",X"25",X"20",X"E5",X"FF",
		X"3E",X"07",X"11",X"02",X"03",X"DF",X"E1",X"01",X"01",X"08",X"CD",X"0F",X"09",X"21",X"00",X"00",
		X"22",X"23",X"20",X"22",X"25",X"20",X"C3",X"6A",X"18",X"21",X"2B",X"20",X"AF",X"BE",X"C8",X"23",
		X"34",X"7E",X"FE",X"03",X"CA",X"D6",X"17",X"11",X"E9",X"44",X"FE",X"02",X"C2",X"C2",X"17",X"11",
		X"01",X"45",X"2A",X"2D",X"20",X"E5",X"D5",X"FF",X"3E",X"06",X"11",X"01",X"07",X"DF",X"D1",X"E1",
		X"01",X"01",X"18",X"C3",X"AB",X"07",X"2A",X"2D",X"20",X"01",X"01",X"18",X"CD",X"0F",X"09",X"21",
		X"00",X"00",X"22",X"2B",X"20",X"22",X"2D",X"20",X"C3",X"6A",X"18",X"21",X"27",X"20",X"AF",X"BE",
		X"C8",X"23",X"34",X"7E",X"FE",X"03",X"CA",X"18",X"18",X"11",X"19",X"45",X"FE",X"02",X"C2",X"04");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
