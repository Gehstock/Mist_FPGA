library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kb_1h is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kb_1h is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",
		X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",
		X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",
		X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",
		X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",
		X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",
		X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",X"C0",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"0F",X"0F",X"0F",X"FE",X"F8",X"E0",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",
		X"00",X"E0",X"F8",X"FE",X"0F",X"0F",X"0F",X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"27",X"07",X"17",X"07",X"03",X"13",X"03",X"23",X"00",X"C0",X"E0",X"F0",X"38",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"C3",X"53",X"FB",X"07",X"07",X"07",X"07",X"03",X"03",X"C3",X"53",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"C3",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"FF",X"44",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"07",X"00",X"00",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"07",X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",X"44",X"07",X"00",X"00",
		X"00",X"07",X"44",X"FF",X"FF",X"44",X"07",X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",X"44",X"07",
		X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",X"44",X"00",X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",
		X"FF",X"57",X"C7",X"07",X"03",X"03",X"03",X"03",X"FF",X"FF",X"57",X"C7",X"03",X"03",X"03",X"03",
		X"57",X"FF",X"FF",X"57",X"C3",X"03",X"03",X"03",X"C7",X"57",X"FF",X"FF",X"53",X"C3",X"03",X"03",
		X"07",X"C7",X"57",X"FF",X"FB",X"53",X"C3",X"03",X"07",X"07",X"C7",X"57",X"FB",X"FB",X"53",X"C3",
		X"07",X"07",X"07",X"C7",X"53",X"FB",X"FB",X"53",X"07",X"07",X"07",X"07",X"C3",X"53",X"FB",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"C7",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"47",X"C7",X"07",X"07",X"03",X"03",X"03",X"03",
		X"03",X"00",X"00",X"08",X"00",X"28",X"44",X"40",X"00",X"82",X"04",X"01",X"92",X"00",X"20",X"04",
		X"00",X"20",X"00",X"00",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"12",X"00",X"60",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"C3",
		X"44",X"FF",X"00",X"00",X"00",X"00",X"FF",X"44",X"57",X"FF",X"07",X"07",X"03",X"03",X"FB",X"53",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"02",X"03",X"02",X"02",X"03",X"02",X"02",X"02",X"07",X"07",X"07",X"07",X"83",X"83",X"83",X"83",
		X"03",X"02",X"03",X"02",X"02",X"03",X"02",X"03",X"87",X"07",X"07",X"07",X"03",X"03",X"03",X"83",
		X"02",X"02",X"02",X"03",X"02",X"02",X"03",X"02",X"87",X"87",X"87",X"87",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"00",X"00",X"00",X"A0",X"D0",X"C8",X"C0",X"C0",
		X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"C0",X"C8",X"D0",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"40",X"B0",X"80",X"80",
		X"3F",X"3F",X"3F",X"1F",X"07",X"00",X"00",X"00",X"80",X"90",X"A0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1F",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"80",X"40",X"20",X"00",X"00",
		X"7F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"1F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"C0",X"A0",X"90",X"80",X"80",
		X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"B0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"90",
		X"05",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"40",X"A0",X"10",X"00",X"00",X"00",X"00",
		X"00",X"02",X"01",X"04",X"02",X"02",X"20",X"12",X"00",X"00",X"20",X"40",X"18",X"98",X"24",X"40",
		X"26",X"0B",X"01",X"02",X"02",X"04",X"00",X"00",X"40",X"20",X"90",X"C0",X"20",X"90",X"00",X"00",
		X"00",X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"62",X"92",X"8A",X"86",X"62",
		X"82",X"7C",X"00",X"8C",X"D2",X"A2",X"82",X"84",X"82",X"7C",X"00",X"08",X"FE",X"48",X"28",X"18",
		X"82",X"7C",X"00",X"9C",X"A2",X"A2",X"A2",X"E4",X"82",X"7C",X"00",X"0C",X"92",X"92",X"52",X"3C",
		X"82",X"7C",X"00",X"C0",X"A0",X"90",X"8E",X"80",X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"00",X"00",
		X"DB",X"DB",X"DF",X"1F",X"00",X"00",X"7F",X"FF",X"FF",X"00",X"00",X"7F",X"FF",X"DB",X"DB",X"DB",
		X"FF",X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"FF",X"C3",X"C3",X"C3",X"FF",X"7E",X"00",X"00",X"7F",
		X"C3",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"C3",X"00",X"00",X"00",X"7E",X"FF",X"C3",X"C3",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"06",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"06",X"06",X"02",X"00",X"00",X"00",
		X"02",X"D9",X"D8",X"DA",X"D9",X"D8",X"D8",X"D8",X"00",X"00",X"80",X"40",X"20",X"80",X"60",X"00",
		X"D8",X"D8",X"D9",X"DA",X"D8",X"D9",X"02",X"00",X"60",X"80",X"20",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1C",X"30",X"40",X"0F",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"40",X"30",X"1C",X"0F",X"03",X"00",X"FE",X"02",X"06",X"00",X"00",X"00",X"80",X"00",
		X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"FE",X"7C",X"00",X"9C",X"A2",X"A2",X"E4",X"00",X"FE",
		X"08",X"08",X"08",X"FF",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",
		X"00",X"00",X"00",X"06",X"36",X"36",X"76",X"76",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",
		X"76",X"76",X"36",X"36",X"06",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",
		X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",X"C0",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",
		X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",
		X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",
		X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",
		X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",
		X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",
		X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",X"C0",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"0F",X"0F",X"0F",X"FE",X"F8",X"E0",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",
		X"00",X"E0",X"F8",X"FE",X"0F",X"0F",X"0F",X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"27",X"07",X"17",X"07",X"03",X"13",X"03",X"23",X"00",X"C0",X"E0",X"F0",X"38",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"C3",X"53",X"FB",X"07",X"07",X"07",X"07",X"03",X"03",X"C3",X"53",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"C3",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"FF",X"44",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"07",X"00",X"00",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"07",X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",X"44",X"07",X"00",X"00",
		X"00",X"07",X"44",X"FF",X"FF",X"44",X"07",X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",X"44",X"07",
		X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",X"44",X"00",X"00",X"00",X"00",X"07",X"44",X"FF",X"FF",
		X"FF",X"57",X"C7",X"07",X"03",X"03",X"03",X"03",X"FF",X"FF",X"57",X"C7",X"03",X"03",X"03",X"03",
		X"57",X"FF",X"FF",X"57",X"C3",X"03",X"03",X"03",X"C7",X"57",X"FF",X"FF",X"53",X"C3",X"03",X"03",
		X"07",X"C7",X"57",X"FF",X"FB",X"53",X"C3",X"03",X"07",X"07",X"C7",X"57",X"FB",X"FB",X"53",X"C3",
		X"07",X"07",X"07",X"C7",X"53",X"FB",X"FB",X"53",X"07",X"07",X"07",X"07",X"C3",X"53",X"FB",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"C7",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"47",X"C7",X"07",X"07",X"03",X"03",X"03",X"03",
		X"03",X"00",X"00",X"08",X"00",X"28",X"44",X"40",X"00",X"82",X"04",X"01",X"92",X"00",X"20",X"04",
		X"00",X"20",X"00",X"00",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"12",X"00",X"60",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"C3",
		X"44",X"FF",X"00",X"00",X"00",X"00",X"FF",X"44",X"57",X"FF",X"07",X"07",X"03",X"03",X"FB",X"53",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"02",X"03",X"02",X"02",X"03",X"02",X"02",X"02",X"07",X"07",X"07",X"07",X"83",X"83",X"83",X"83",
		X"03",X"02",X"03",X"02",X"02",X"03",X"02",X"03",X"87",X"07",X"07",X"07",X"03",X"03",X"03",X"83",
		X"02",X"02",X"02",X"03",X"02",X"02",X"03",X"02",X"87",X"87",X"87",X"87",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"00",X"00",X"00",X"A0",X"D0",X"C8",X"C0",X"C0",
		X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"C0",X"C8",X"D0",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"40",X"B0",X"80",X"80",
		X"3F",X"3F",X"3F",X"1F",X"07",X"00",X"00",X"00",X"80",X"90",X"A0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1F",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"80",X"40",X"20",X"00",X"00",
		X"7F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"1F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"C0",X"A0",X"90",X"80",X"80",
		X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"B0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"90",
		X"05",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"40",X"A0",X"10",X"00",X"00",X"00",X"00",
		X"00",X"02",X"01",X"04",X"02",X"02",X"20",X"12",X"00",X"00",X"20",X"40",X"18",X"98",X"24",X"40",
		X"26",X"0B",X"01",X"02",X"02",X"04",X"00",X"00",X"40",X"20",X"90",X"C0",X"20",X"90",X"00",X"00",
		X"00",X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"62",X"92",X"8A",X"86",X"62",
		X"82",X"7C",X"00",X"8C",X"D2",X"A2",X"82",X"84",X"82",X"7C",X"00",X"08",X"FE",X"48",X"28",X"18",
		X"82",X"7C",X"00",X"9C",X"A2",X"A2",X"A2",X"E4",X"82",X"7C",X"00",X"0C",X"92",X"92",X"52",X"3C",
		X"82",X"7C",X"00",X"C0",X"A0",X"90",X"8E",X"80",X"7C",X"82",X"82",X"7C",X"00",X"7C",X"82",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"00",X"00",
		X"DB",X"DB",X"DF",X"1F",X"00",X"00",X"7F",X"FF",X"FF",X"00",X"00",X"7F",X"FF",X"DB",X"DB",X"DB",
		X"FF",X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"FF",X"C3",X"C3",X"C3",X"FF",X"7E",X"00",X"00",X"7F",
		X"C3",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"C3",X"00",X"00",X"00",X"7E",X"FF",X"C3",X"C3",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"06",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"06",X"06",X"02",X"00",X"00",X"00",
		X"02",X"D9",X"D8",X"DA",X"D9",X"D8",X"D8",X"D8",X"00",X"00",X"80",X"40",X"20",X"80",X"60",X"00",
		X"D8",X"D8",X"D9",X"DA",X"D8",X"D9",X"02",X"00",X"60",X"80",X"20",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1C",X"30",X"40",X"0F",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"40",X"30",X"1C",X"0F",X"03",X"00",X"FE",X"02",X"06",X"00",X"00",X"00",X"80",X"00",
		X"7C",X"00",X"7C",X"82",X"82",X"7C",X"00",X"FE",X"7C",X"00",X"9C",X"A2",X"A2",X"E4",X"00",X"FE",
		X"08",X"08",X"08",X"FF",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",
		X"00",X"00",X"00",X"06",X"36",X"36",X"76",X"76",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",
		X"76",X"76",X"36",X"36",X"06",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",
		X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"C0",X"80",X"80",X"C0",X"80",X"80",X"C0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
