library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"70",X"C3",X"22",X"13",X"00",X"3A",X"2F",X"43",X"11",X"30",X"43",X"18",X"3B",
		X"4F",X"EB",X"21",X"60",X"40",X"C3",X"EF",X"01",X"E1",X"5E",X"23",X"56",X"23",X"C3",X"5D",X"00",
		X"85",X"6F",X"30",X"01",X"24",X"7E",X"C9",X"00",X"87",X"E3",X"E7",X"5F",X"23",X"56",X"EB",X"E9",
		X"E1",X"5E",X"23",X"56",X"23",X"4E",X"23",X"3E",X"C7",X"46",X"23",X"C6",X"59",X"91",X"C5",X"06",
		X"00",X"ED",X"B0",X"4F",X"EB",X"09",X"EB",X"C1",X"10",X"F4",X"E9",X"EB",X"85",X"6F",X"D6",X"2C",
		X"E6",X"7F",X"32",X"2F",X"43",X"71",X"2C",X"70",X"2C",X"73",X"2C",X"72",X"C9",X"ED",X"53",X"00",
		X"43",X"E9",X"2A",X"00",X"43",X"E9",X"08",X"D9",X"DD",X"E5",X"FD",X"E5",X"3A",X"00",X"78",X"AF",
		X"32",X"01",X"70",X"32",X"3E",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"C8",
		X"42",X"11",X"06",X"58",X"06",X"04",X"AF",X"96",X"12",X"1C",X"1C",X"12",X"1C",X"1C",X"2C",X"10",
		X"F5",X"3A",X"D7",X"42",X"ED",X"44",X"11",X"36",X"58",X"06",X"03",X"12",X"1C",X"1C",X"10",X"FB",
		X"3A",X"08",X"43",X"4F",X"3A",X"03",X"43",X"A1",X"4F",X"21",X"70",X"42",X"11",X"40",X"58",X"06",
		X"08",X"2C",X"78",X"FE",X"06",X"3E",X"F0",X"38",X"07",X"3C",X"CB",X"41",X"20",X"02",X"3E",X"EF",
		X"96",X"12",X"1C",X"1C",X"1C",X"2D",X"7E",X"12",X"2C",X"2C",X"1C",X"10",X"E4",X"DD",X"21",X"B0",
		X"42",X"06",X"08",X"1C",X"78",X"FE",X"06",X"3E",X"00",X"30",X"01",X"3D",X"DD",X"96",X"01",X"12",
		X"1C",X"1C",X"3E",X"FB",X"DD",X"96",X"00",X"CB",X"41",X"20",X"03",X"2F",X"D6",X"05",X"12",X"1C",
		X"DD",X"23",X"DD",X"23",X"10",X"DD",X"21",X"E0",X"42",X"11",X"01",X"58",X"06",X"20",X"7E",X"12",
		X"2C",X"1C",X"1C",X"10",X"F9",X"21",X"10",X"42",X"06",X"08",X"7E",X"12",X"2C",X"1C",X"7E",X"12",
		X"2C",X"1C",X"1C",X"1C",X"10",X"F4",X"01",X"28",X"01",X"CF",X"21",X"01",X"70",X"36",X"00",X"36",
		X"01",X"FD",X"E1",X"DD",X"E1",X"D9",X"08",X"C9",X"2A",X"84",X"42",X"23",X"7D",X"B4",X"28",X"03",
		X"22",X"84",X"42",X"CD",X"62",X"00",X"CD",X"86",X"01",X"CD",X"21",X"07",X"CD",X"72",X"04",X"CD",
		X"59",X"05",X"CD",X"44",X"08",X"CD",X"D2",X"08",X"CD",X"46",X"11",X"CD",X"0B",X"02",X"CD",X"30",
		X"02",X"CD",X"6F",X"20",X"CD",X"E2",X"1E",X"CD",X"92",X"1B",X"CD",X"AA",X"1D",X"26",X"40",X"AF",
		X"C6",X"60",X"6F",X"7E",X"D6",X"01",X"38",X"16",X"77",X"20",X"13",X"E5",X"7D",X"D6",X"60",X"87",
		X"87",X"C6",X"80",X"6F",X"4E",X"2C",X"46",X"2C",X"5E",X"2C",X"56",X"EB",X"CF",X"E1",X"7D",X"D6",
		X"5F",X"E6",X"1F",X"20",X"DB",X"C9",X"21",X"18",X"43",X"34",X"7E",X"E6",X"0F",X"C0",X"7E",X"0F",
		X"0F",X"0F",X"0F",X"47",X"3A",X"19",X"43",X"2F",X"B0",X"4F",X"3A",X"15",X"43",X"D6",X"01",X"30",
		X"02",X"AF",X"4F",X"28",X"01",X"79",X"32",X"01",X"60",X"79",X"32",X"00",X"60",X"21",X"20",X"53",
		X"11",X"80",X"50",X"3A",X"03",X"43",X"A7",X"28",X"01",X"EB",X"3C",X"4F",X"3A",X"1A",X"43",X"A0",
		X"CC",X"D1",X"01",X"C4",X"E0",X"01",X"EB",X"3A",X"02",X"43",X"A7",X"28",X"13",X"79",X"EE",X"03",
		X"4F",X"E5",X"FD",X"E1",X"FD",X"36",X"00",X"19",X"FD",X"36",X"20",X"1E",X"FD",X"71",X"40",X"C9",
		X"E5",X"FD",X"E1",X"3E",X"24",X"FD",X"77",X"00",X"FD",X"77",X"20",X"FD",X"77",X"40",X"C9",X"06",
		X"20",X"7E",X"A7",X"28",X"04",X"2C",X"10",X"F9",X"C9",X"71",X"7D",X"D6",X"60",X"87",X"87",X"C6",
		X"80",X"6F",X"C1",X"71",X"2C",X"70",X"2C",X"73",X"2C",X"72",X"C9",X"21",X"1D",X"43",X"11",X"1C",
		X"43",X"01",X"00",X"03",X"1A",X"87",X"38",X"11",X"F0",X"3F",X"7E",X"CE",X"00",X"27",X"FE",X"60",
		X"38",X"02",X"3E",X"00",X"77",X"2C",X"10",X"F1",X"C9",X"71",X"2C",X"10",X"FC",X"0F",X"12",X"C9",
		X"3A",X"15",X"43",X"FE",X"99",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"60",X"2F",X"0F",X"21",X"11",X"43",X"7E",X"17",X"77",X"E6",X"0F",X"D6",X"0C",X"CC",
		X"A0",X"25",X"3A",X"00",X"60",X"2F",X"0F",X"0F",X"21",X"12",X"43",X"7E",X"17",X"77",X"E6",X"0F",
		X"D6",X"0C",X"C0",X"01",X"93",X"02",X"CF",X"21",X"13",X"43",X"34",X"34",X"7E",X"FE",X"02",X"C0",
		X"01",X"85",X"02",X"CF",X"C9",X"3E",X"08",X"D7",X"C3",X"CF",X"25",X"00",X"32",X"04",X"60",X"35",
		X"20",X"F3",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"0C",X"43",
		X"21",X"15",X"43",X"86",X"27",X"30",X"02",X"3E",X"99",X"77",X"21",X"6B",X"22",X"D4",X"22",X"20",
		X"3A",X"16",X"43",X"A7",X"C8",X"11",X"15",X"43",X"21",X"BF",X"52",X"01",X"01",X"01",X"C3",X"5C",
		X"03",X"21",X"05",X"43",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1C",X"2C",X"10",X"F7",X"C9",
		X"1A",X"77",X"1C",X"2C",X"10",X"FA",X"C9",X"47",X"E6",X"F0",X"4F",X"78",X"1F",X"47",X"38",X"06",
		X"1F",X"1F",X"1F",X"E6",X"0F",X"4F",X"3E",X"03",X"90",X"E6",X"07",X"47",X"E7",X"2D",X"7E",X"89",
		X"27",X"77",X"0E",X"00",X"10",X"F7",X"D0",X"36",X"99",X"2C",X"36",X"99",X"2C",X"36",X"90",X"C9",
		X"4F",X"C5",X"79",X"CD",X"0A",X"03",X"C1",X"10",X"F8",X"C9",X"47",X"3A",X"17",X"43",X"A7",X"C0",
		X"78",X"21",X"0D",X"40",X"CD",X"D7",X"02",X"CD",X"4B",X"04",X"CD",X"31",X"03",X"11",X"0D",X"40",
		X"CD",X"C1",X"02",X"11",X"2D",X"40",X"CD",X"C1",X"02",X"11",X"05",X"43",X"21",X"41",X"52",X"18",
		X"28",X"11",X"0D",X"40",X"3A",X"03",X"43",X"A7",X"20",X"1C",X"21",X"A1",X"53",X"18",X"1A",X"11",
		X"0D",X"40",X"21",X"2D",X"40",X"3A",X"03",X"43",X"A7",X"28",X"01",X"EB",X"E5",X"CD",X"3A",X"03",
		X"D1",X"3A",X"02",X"43",X"A7",X"C8",X"21",X"01",X"51",X"01",X"04",X"03",X"3E",X"E0",X"C5",X"47",
		X"1A",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"20",X"07",X"0D",X"FA",X"70",X"03",X"3E",X"24",X"FA",
		X"0E",X"00",X"77",X"1A",X"E6",X"0F",X"20",X"07",X"0D",X"FA",X"7F",X"03",X"3E",X"24",X"FA",X"0E",
		X"00",X"D5",X"58",X"16",X"FF",X"19",X"77",X"19",X"D1",X"1C",X"78",X"E3",X"44",X"E1",X"10",X"CE",
		X"C9",X"C6",X"40",X"6F",X"26",X"27",X"66",X"CD",X"9D",X"03",X"67",X"29",X"C9",X"AF",X"6F",X"57",
		X"CB",X"7C",X"28",X"01",X"93",X"CB",X"7B",X"28",X"01",X"94",X"06",X"08",X"29",X"30",X"01",X"19",
		X"10",X"FA",X"84",X"C9",X"2E",X"00",X"06",X"11",X"AF",X"17",X"BB",X"38",X"01",X"93",X"3F",X"ED",
		X"6A",X"10",X"F6",X"C9",X"01",X"00",X"08",X"11",X"00",X"40",X"7C",X"92",X"79",X"9B",X"38",X"05",
		X"4F",X"7C",X"92",X"67",X"A7",X"3F",X"CB",X"13",X"29",X"CB",X"11",X"29",X"CB",X"11",X"10",X"EA",
		X"C9",X"FD",X"21",X"20",X"43",X"7B",X"95",X"30",X"02",X"2F",X"3C",X"FD",X"CB",X"01",X"16",X"4F",
		X"7A",X"94",X"30",X"02",X"2F",X"3C",X"FD",X"CB",X"03",X"16",X"5F",X"B1",X"F2",X"03",X"04",X"CB",
		X"39",X"CB",X"3B",X"FD",X"71",X"00",X"FD",X"73",X"02",X"63",X"CD",X"9D",X"03",X"E5",X"59",X"63",
		X"CD",X"9D",X"03",X"D1",X"19",X"CD",X"C4",X"03",X"FD",X"66",X"00",X"CD",X"B4",X"03",X"7C",X"A7",
		X"7D",X"28",X"02",X"3E",X"FF",X"A7",X"28",X"09",X"FD",X"CB",X"01",X"1E",X"30",X"02",X"2F",X"3C",
		X"1F",X"4F",X"FD",X"66",X"02",X"CD",X"B4",X"03",X"7C",X"A7",X"7D",X"28",X"02",X"3E",X"FF",X"A7",
		X"C8",X"FD",X"CB",X"03",X"1E",X"30",X"02",X"2F",X"3C",X"1F",X"C9",X"3A",X"10",X"40",X"A7",X"C0",
		X"2A",X"0D",X"40",X"7D",X"6C",X"67",X"29",X"29",X"29",X"29",X"7C",X"21",X"0A",X"43",X"BE",X"D8",
		X"3E",X"01",X"32",X"10",X"40",X"21",X"75",X"22",X"CD",X"1D",X"20",X"21",X"0A",X"40",X"34",X"C3",
		X"77",X"18",X"3A",X"D0",X"42",X"3D",X"C0",X"CD",X"B7",X"04",X"29",X"29",X"29",X"29",X"ED",X"5B",
		X"D2",X"42",X"19",X"22",X"D2",X"42",X"7A",X"47",X"E6",X"F8",X"6F",X"26",X"00",X"29",X"29",X"11",
		X"18",X"50",X"19",X"78",X"E6",X"07",X"C6",X"70",X"11",X"20",X"00",X"77",X"2C",X"C6",X"08",X"77",
		X"19",X"C6",X"10",X"77",X"2D",X"D6",X"08",X"77",X"78",X"FE",X"D0",X"D0",X"E6",X"07",X"C6",X"90",
		X"19",X"77",X"2C",X"C6",X"08",X"77",X"C9",X"3A",X"17",X"43",X"A7",X"20",X"34",X"3A",X"D1",X"42",
		X"47",X"21",X"00",X"00",X"3A",X"08",X"43",X"4F",X"3A",X"03",X"43",X"A1",X"3A",X"00",X"60",X"28",
		X"03",X"3A",X"00",X"68",X"87",X"87",X"87",X"87",X"87",X"38",X"09",X"F0",X"3A",X"D3",X"42",X"FE",
		X"D0",X"D0",X"68",X"C9",X"F8",X"3A",X"D3",X"42",X"FE",X"21",X"D8",X"AF",X"90",X"C8",X"6F",X"25",
		X"C9",X"3A",X"18",X"43",X"E6",X"1F",X"FE",X"10",X"20",X"23",X"01",X"00",X"08",X"DD",X"21",X"20",
		X"42",X"CD",X"2D",X"05",X"DD",X"23",X"DD",X"23",X"10",X"F7",X"06",X"07",X"DD",X"21",X"90",X"42",
		X"CD",X"3A",X"05",X"DD",X"23",X"DD",X"23",X"10",X"F7",X"79",X"32",X"86",X"42",X"3A",X"D1",X"42",
		X"47",X"21",X"00",X"00",X"3A",X"86",X"42",X"87",X"38",X"BB",X"C8",X"18",X"AF",X"DD",X"7E",X"00",
		X"A7",X"C8",X"DD",X"6E",X"50",X"DD",X"66",X"51",X"18",X"0D",X"DD",X"7E",X"00",X"DD",X"B6",X"01",
		X"C8",X"DD",X"6E",X"20",X"DD",X"66",X"21",X"0D",X"3A",X"D3",X"42",X"BC",X"3E",X"A0",X"38",X"04",
		X"BD",X"D0",X"18",X"02",X"BD",X"D8",X"0C",X"0C",X"C9",X"3A",X"80",X"42",X"A7",X"C8",X"3A",X"9E",
		X"42",X"A7",X"20",X"47",X"3A",X"D0",X"42",X"3D",X"28",X"06",X"6F",X"67",X"22",X"BE",X"42",X"C9",
		X"CD",X"78",X"06",X"3A",X"17",X"43",X"A7",X"28",X"08",X"3A",X"18",X"43",X"E6",X"1F",X"C0",X"18",
		X"25",X"3A",X"08",X"43",X"47",X"3A",X"03",X"43",X"A0",X"3A",X"00",X"60",X"28",X"03",X"3A",X"00",
		X"68",X"2F",X"07",X"07",X"07",X"07",X"21",X"83",X"42",X"7E",X"17",X"77",X"E6",X"0F",X"D6",X"0C",
		X"C0",X"3E",X"08",X"CD",X"E7",X"05",X"3E",X"B0",X"32",X"9E",X"42",X"3A",X"9E",X"42",X"26",X"00",
		X"87",X"30",X"01",X"25",X"6F",X"29",X"29",X"29",X"3A",X"AE",X"42",X"85",X"32",X"AE",X"42",X"3A",
		X"BE",X"42",X"8C",X"32",X"BE",X"42",X"2A",X"BE",X"42",X"3A",X"18",X"43",X"E6",X"01",X"87",X"3D",
		X"84",X"67",X"7D",X"FE",X"10",X"DA",X"74",X"06",X"22",X"BE",X"42",X"D6",X"18",X"FE",X"40",X"38",
		X"18",X"3E",X"01",X"32",X"C0",X"42",X"C9",X"47",X"3A",X"17",X"43",X"A7",X"C0",X"3E",X"01",X"32",
		X"05",X"68",X"78",X"D7",X"AF",X"32",X"05",X"68",X"C9",X"6F",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"EB",X"21",X"C8",X"42",X"E7",X"EB",X"ED",X"44",X"84",X"67",X"22",X"24",X"43",X"AF",X"32",X"C0",
		X"42",X"7D",X"E6",X"0F",X"FE",X"0C",X"D0",X"7C",X"E6",X"0F",X"D6",X"02",X"FE",X"0C",X"D0",X"3E",
		X"01",X"32",X"C0",X"42",X"7D",X"E6",X"F0",X"0F",X"0F",X"0F",X"CB",X"04",X"CE",X"00",X"6F",X"7C",
		X"E6",X"E0",X"07",X"07",X"07",X"3C",X"47",X"26",X"40",X"3E",X"80",X"07",X"10",X"FD",X"A6",X"C8",
		X"AE",X"77",X"7D",X"D6",X"00",X"21",X"E3",X"42",X"E7",X"21",X"86",X"06",X"E7",X"CD",X"0A",X"03",
		X"2A",X"24",X"43",X"7D",X"0F",X"0F",X"0F",X"E6",X"1E",X"5F",X"7C",X"07",X"07",X"57",X"E6",X"C0",
		X"B3",X"5F",X"7A",X"E6",X"03",X"57",X"21",X"03",X"50",X"19",X"01",X"E0",X"06",X"CF",X"21",X"4B",
		X"22",X"CD",X"1D",X"20",X"AF",X"32",X"9E",X"42",X"3A",X"18",X"43",X"0F",X"3A",X"D3",X"42",X"CE",
		X"07",X"67",X"2E",X"BC",X"22",X"BE",X"42",X"C9",X"51",X"41",X"31",X"21",X"E5",X"DD",X"E1",X"E5",
		X"DD",X"36",X"F0",X"30",X"E1",X"3E",X"08",X"D7",X"E5",X"DD",X"E1",X"DD",X"36",X"F0",X"31",X"3E",
		X"08",X"D7",X"E5",X"DD",X"E1",X"DD",X"36",X"F0",X"28",X"3E",X"08",X"D7",X"E5",X"DD",X"E1",X"3A",
		X"2E",X"42",X"FE",X"03",X"20",X"1E",X"01",X"07",X"07",X"21",X"20",X"42",X"7E",X"B9",X"28",X"14",
		X"2C",X"2C",X"10",X"F8",X"DD",X"36",X"00",X"07",X"DD",X"36",X"F0",X"3C",X"3A",X"FB",X"42",X"DD",
		X"77",X"F1",X"18",X"48",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"50",X"DD",X"77",X"51",X"18",X"3C",
		X"E5",X"FD",X"E1",X"E5",X"3E",X"C0",X"CD",X"D7",X"19",X"E1",X"3E",X"08",X"D7",X"E5",X"FD",X"E1",
		X"3E",X"C4",X"CD",X"D7",X"19",X"3E",X"08",X"D7",X"E5",X"FD",X"E1",X"3E",X"A0",X"CD",X"D7",X"19",
		X"3E",X"08",X"D7",X"E5",X"FD",X"E1",X"CD",X"C8",X"19",X"06",X"08",X"AF",X"21",X"00",X"40",X"B6",
		X"2C",X"10",X"FC",X"A7",X"20",X"06",X"32",X"C3",X"42",X"CD",X"74",X"08",X"21",X"08",X"40",X"35",
		X"C9",X"3A",X"2E",X"42",X"A7",X"C8",X"3A",X"D7",X"42",X"CD",X"FF",X"07",X"3A",X"2E",X"42",X"3D",
		X"C0",X"3A",X"D5",X"42",X"6F",X"26",X"00",X"ED",X"5B",X"D6",X"42",X"3A",X"D4",X"42",X"BA",X"28",
		X"30",X"30",X"06",X"AF",X"95",X"28",X"02",X"6F",X"25",X"29",X"29",X"29",X"29",X"19",X"22",X"D6",
		X"42",X"7C",X"E6",X"03",X"C0",X"CB",X"54",X"20",X"0C",X"F7",X"1B",X"50",X"03",X"02",X"44",X"45",
		X"46",X"47",X"48",X"49",X"C9",X"F7",X"1B",X"50",X"03",X"02",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",
		X"C9",X"21",X"D4",X"42",X"3A",X"D3",X"42",X"86",X"0F",X"47",X"3A",X"18",X"43",X"80",X"FE",X"20",
		X"30",X"02",X"C6",X"20",X"FE",X"D1",X"38",X"02",X"D6",X"2F",X"77",X"C9",X"21",X"32",X"1B",X"11",
		X"E0",X"42",X"01",X"20",X"00",X"ED",X"B0",X"F7",X"51",X"50",X"0A",X"02",X"30",X"31",X"32",X"33",
		X"34",X"35",X"36",X"5F",X"5F",X"5F",X"24",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"5B",X"6B",X"5B",
		X"F7",X"91",X"53",X"0A",X"02",X"30",X"31",X"32",X"33",X"34",X"3D",X"3E",X"53",X"3F",X"53",X"24",
		X"37",X"38",X"39",X"3A",X"40",X"41",X"5F",X"5F",X"5F",X"21",X"99",X"50",X"11",X"20",X"00",X"01",
		X"98",X"18",X"71",X"19",X"10",X"FC",X"3E",X"20",X"21",X"1B",X"50",X"11",X"1E",X"00",X"06",X"20",
		X"36",X"24",X"2C",X"36",X"24",X"2C",X"36",X"67",X"19",X"10",X"F5",X"32",X"D7",X"42",X"32",X"D4",
		X"42",X"ED",X"44",X"11",X"36",X"58",X"06",X"03",X"12",X"1C",X"1C",X"10",X"FB",X"ED",X"44",X"2F",
		X"C6",X"E4",X"CD",X"08",X"08",X"79",X"C6",X"2C",X"4F",X"E6",X"F8",X"6F",X"26",X"00",X"29",X"29",
		X"11",X"1B",X"50",X"19",X"79",X"E6",X"07",X"C6",X"50",X"11",X"20",X"00",X"77",X"2C",X"77",X"2C",
		X"C6",X"10",X"77",X"19",X"C6",X"0C",X"FE",X"70",X"38",X"02",X"3E",X"6F",X"77",X"2D",X"D6",X"10",
		X"77",X"2D",X"77",X"FE",X"5F",X"C0",X"19",X"79",X"E6",X"07",X"C6",X"54",X"77",X"2C",X"77",X"2C",
		X"C6",X"10",X"77",X"C9",X"3A",X"C0",X"42",X"A7",X"C8",X"2A",X"C2",X"42",X"29",X"6C",X"26",X"00",
		X"30",X"01",X"25",X"29",X"29",X"29",X"29",X"4C",X"7D",X"A7",X"21",X"C1",X"42",X"7E",X"CC",X"7E",
		X"08",X"26",X"00",X"87",X"30",X"01",X"25",X"6F",X"29",X"29",X"ED",X"5B",X"C2",X"42",X"19",X"22",
		X"C2",X"42",X"29",X"7C",X"21",X"C8",X"42",X"06",X"04",X"77",X"2C",X"10",X"FC",X"C9",X"A7",X"C8",
		X"DD",X"21",X"00",X"40",X"DD",X"7E",X"00",X"DD",X"B6",X"02",X"DD",X"B6",X"04",X"DD",X"B6",X"06",
		X"5F",X"DD",X"7E",X"01",X"DD",X"B6",X"03",X"DD",X"B6",X"05",X"DD",X"B6",X"07",X"57",X"B3",X"20",
		X"03",X"33",X"33",X"C9",X"CB",X"7E",X"28",X"15",X"06",X"02",X"7B",X"A7",X"20",X"03",X"06",X"FA",
		X"7A",X"05",X"0F",X"30",X"FC",X"78",X"B9",X"7E",X"F8",X"ED",X"44",X"77",X"C9",X"06",X"FE",X"7A",
		X"A7",X"20",X"03",X"06",X"06",X"7B",X"04",X"07",X"30",X"FC",X"79",X"B8",X"7E",X"F8",X"ED",X"44",
		X"77",X"C9",X"3A",X"02",X"42",X"A7",X"C8",X"CD",X"38",X"0D",X"DD",X"21",X"20",X"42",X"06",X"07",
		X"C5",X"DD",X"7E",X"00",X"21",X"02",X"09",X"EF",X"26",X"00",X"34",X"09",X"47",X"0A",X"CE",X"0A",
		X"26",X"00",X"A8",X"0D",X"EE",X"0E",X"C8",X"0E",X"26",X"00",X"26",X"00",X"50",X"0A",X"EE",X"0E",
		X"EE",X"0E",X"DD",X"7E",X"00",X"21",X"23",X"09",X"EF",X"26",X"00",X"2B",X"09",X"2B",X"09",X"2E",
		X"09",X"26",X"00",X"2B",X"09",X"B2",X"0F",X"26",X"00",X"26",X"00",X"26",X"00",X"2E",X"09",X"03",
		X"10",X"4B",X"10",X"DD",X"23",X"DD",X"23",X"C1",X"10",X"B6",X"C9",X"CD",X"D5",X"11",X"CD",X"4D",
		X"0C",X"C3",X"C4",X"0C",X"DD",X"7E",X"50",X"FE",X"DE",X"38",X"1E",X"DD",X"36",X"00",X"02",X"21",
		X"2D",X"0A",X"3A",X"08",X"40",X"3D",X"BE",X"23",X"38",X"04",X"23",X"23",X"18",X"F8",X"5E",X"23",
		X"56",X"EB",X"CD",X"33",X"1D",X"DD",X"77",X"01",X"C9",X"FE",X"C0",X"38",X"3B",X"3A",X"08",X"40",
		X"3D",X"3A",X"04",X"42",X"20",X"03",X"3A",X"05",X"42",X"47",X"DD",X"7E",X"30",X"CD",X"7F",X"09",
		X"DD",X"77",X"30",X"DD",X"7E",X"31",X"CD",X"87",X"09",X"DD",X"77",X"31",X"C3",X"D4",X"0B",X"A7",
		X"FA",X"85",X"09",X"B8",X"D0",X"78",X"C9",X"A7",X"FA",X"8F",X"09",X"B8",X"D8",X"78",X"C9",X"ED",
		X"44",X"B8",X"38",X"01",X"78",X"ED",X"44",X"C9",X"11",X"80",X"01",X"DD",X"6E",X"20",X"DD",X"66",
		X"21",X"19",X"DD",X"75",X"20",X"DD",X"74",X"21",X"CD",X"AF",X"09",X"CD",X"D4",X"09",X"C9",X"DD",
		X"7E",X"21",X"87",X"1E",X"20",X"CD",X"91",X"03",X"7C",X"DD",X"86",X"30",X"87",X"6F",X"26",X"00",
		X"30",X"01",X"25",X"DD",X"56",X"50",X"DD",X"5E",X"40",X"29",X"29",X"29",X"19",X"DD",X"75",X"40",
		X"DD",X"74",X"50",X"C9",X"DD",X"7E",X"21",X"1E",X"10",X"CD",X"91",X"03",X"7C",X"DD",X"86",X"31",
		X"87",X"6F",X"26",X"00",X"30",X"01",X"25",X"DD",X"56",X"51",X"DD",X"5E",X"41",X"29",X"29",X"29",
		X"19",X"DD",X"75",X"41",X"DD",X"74",X"51",X"DD",X"7E",X"31",X"87",X"38",X"1A",X"C8",X"DD",X"7E",
		X"51",X"C6",X"08",X"FE",X"F8",X"D8",X"DD",X"7E",X"31",X"ED",X"44",X"DD",X"77",X"31",X"DD",X"36",
		X"51",X"EF",X"DD",X"36",X"21",X"80",X"C9",X"DD",X"7E",X"51",X"FE",X"F8",X"D8",X"DD",X"7E",X"31",
		X"ED",X"44",X"DD",X"77",X"31",X"AF",X"DD",X"77",X"51",X"DD",X"77",X"21",X"C9",X"06",X"39",X"0A",
		X"12",X"3B",X"0A",X"1E",X"41",X"0A",X"FF",X"45",X"0A",X"FF",X"B4",X"01",X"78",X"05",X"96",X"FF",
		X"B4",X"03",X"78",X"FF",X"96",X"FF",X"78",X"DD",X"35",X"01",X"C0",X"DD",X"36",X"00",X"03",X"C9",
		X"CD",X"D4",X"0B",X"DD",X"7E",X"50",X"FE",X"08",X"30",X"54",X"AF",X"DD",X"36",X"00",X"03",X"DD",
		X"77",X"50",X"DD",X"77",X"51",X"6F",X"67",X"32",X"2E",X"42",X"22",X"7E",X"42",X"32",X"81",X"42",
		X"32",X"03",X"42",X"32",X"02",X"42",X"32",X"80",X"42",X"32",X"C0",X"42",X"32",X"C5",X"42",X"3E",
		X"02",X"32",X"D0",X"42",X"21",X"65",X"23",X"CD",X"4D",X"20",X"21",X"93",X"22",X"CD",X"4D",X"20",
		X"21",X"85",X"22",X"CD",X"1D",X"20",X"3E",X"03",X"CD",X"06",X"20",X"F7",X"8D",X"51",X"01",X"09",
		X"43",X"24",X"0E",X"22",X"0B",X"24",X"0E",X"22",X"0B",X"01",X"72",X"0B",X"CF",X"C9",X"C6",X"10",
		X"2E",X"DE",X"BD",X"30",X"01",X"6F",X"DD",X"66",X"51",X"22",X"7E",X"42",X"E6",X"07",X"C0",X"CB",
		X"5D",X"2E",X"34",X"28",X"01",X"2C",X"3A",X"FB",X"42",X"67",X"22",X"1E",X"42",X"C9",X"CD",X"D4",
		X"0B",X"DD",X"7E",X"50",X"FE",X"D0",X"38",X"0D",X"3A",X"0A",X"42",X"ED",X"44",X"DD",X"77",X"30",
		X"DD",X"36",X"31",X"00",X"C9",X"2A",X"C2",X"42",X"29",X"6C",X"26",X"00",X"30",X"01",X"25",X"DD",
		X"7E",X"10",X"0F",X"4F",X"E6",X"F0",X"85",X"57",X"7C",X"CE",X"00",X"C0",X"79",X"87",X"87",X"87",
		X"87",X"C6",X"18",X"5F",X"DD",X"6E",X"50",X"DD",X"66",X"51",X"7C",X"92",X"20",X"02",X"7D",X"93",
		X"20",X"24",X"3A",X"08",X"40",X"FE",X"07",X"30",X"0D",X"DD",X"36",X"00",X"01",X"DD",X"6E",X"50",
		X"DD",X"66",X"51",X"C3",X"C8",X"1C",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"50",X"DD",X"77",X"51",
		X"CD",X"B6",X"0B",X"C3",X"0D",X"1F",X"CD",X"E1",X"03",X"67",X"CD",X"4C",X"0B",X"5F",X"CD",X"97",
		X"03",X"DD",X"74",X"31",X"61",X"CD",X"97",X"03",X"DD",X"74",X"30",X"C9",X"7B",X"FE",X"20",X"30",
		X"0C",X"3A",X"C1",X"42",X"A7",X"F2",X"5A",X"0B",X"ED",X"44",X"C6",X"10",X"C9",X"DD",X"7E",X"00",
		X"FE",X"0A",X"3A",X"0A",X"42",X"C0",X"3A",X"08",X"40",X"3D",X"3A",X"07",X"42",X"C0",X"3A",X"08",
		X"42",X"C9",X"3E",X"B4",X"D7",X"AF",X"CD",X"06",X"20",X"06",X"07",X"DD",X"21",X"20",X"42",X"C5",
		X"CD",X"AB",X"0B",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"50",X"DD",X"77",X"51",X"DD",X"23",X"DD",
		X"23",X"C1",X"10",X"EB",X"DD",X"77",X"00",X"DD",X"77",X"50",X"DD",X"77",X"51",X"01",X"00",X"30",
		X"21",X"90",X"42",X"71",X"2C",X"10",X"FC",X"DF",X"39",X"1A",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",
		X"FE",X"04",X"C8",X"FE",X"07",X"C8",X"21",X"00",X"40",X"DD",X"7E",X"10",X"E6",X"1F",X"85",X"6F",
		X"DD",X"7E",X"10",X"E6",X"E0",X"07",X"07",X"07",X"3C",X"4F",X"47",X"3E",X"80",X"07",X"10",X"FD",
		X"AE",X"77",X"41",X"C9",X"CD",X"DB",X"0B",X"CD",X"06",X"0C",X"C9",X"DD",X"7E",X"30",X"DD",X"5E",
		X"40",X"DD",X"56",X"50",X"26",X"00",X"87",X"6F",X"30",X"01",X"25",X"29",X"29",X"29",X"19",X"DD",
		X"75",X"40",X"DD",X"74",X"50",X"7C",X"FE",X"F0",X"D8",X"DD",X"36",X"50",X"00",X"DD",X"7E",X"30",
		X"ED",X"44",X"DD",X"77",X"30",X"C9",X"DD",X"7E",X"31",X"DD",X"5E",X"41",X"DD",X"56",X"51",X"26",
		X"00",X"87",X"6F",X"30",X"01",X"25",X"29",X"29",X"29",X"19",X"DD",X"75",X"41",X"DD",X"74",X"51",
		X"DD",X"7E",X"31",X"87",X"38",X"14",X"C8",X"7C",X"C6",X"08",X"FE",X"F8",X"D8",X"DD",X"7E",X"31",
		X"ED",X"44",X"DD",X"77",X"31",X"DD",X"36",X"51",X"EF",X"C9",X"DD",X"7E",X"51",X"FE",X"F8",X"D8",
		X"DD",X"7E",X"31",X"ED",X"44",X"DD",X"77",X"31",X"DD",X"36",X"51",X"00",X"C9",X"3A",X"9E",X"42",
		X"A7",X"C8",X"3A",X"BE",X"42",X"DD",X"96",X"50",X"FE",X"0C",X"D0",X"3A",X"BF",X"42",X"DD",X"96",
		X"51",X"D6",X"02",X"FE",X"0C",X"D0",X"3E",X"01",X"32",X"C0",X"42",X"CD",X"74",X"06",X"DD",X"7E",
		X"00",X"FE",X"04",X"C8",X"FE",X"0A",X"06",X"02",X"20",X"01",X"04",X"DD",X"7E",X"F1",X"21",X"86",
		X"06",X"E7",X"CD",X"00",X"03",X"CD",X"9A",X"0C",X"DD",X"36",X"00",X"04",X"DD",X"E5",X"E1",X"01",
		X"8C",X"06",X"CF",X"21",X"4B",X"22",X"CD",X"1D",X"20",X"C9",X"DD",X"7E",X"00",X"FE",X"0A",X"C0",
		X"3E",X"03",X"32",X"2E",X"42",X"21",X"93",X"22",X"CD",X"4D",X"20",X"21",X"1D",X"21",X"CD",X"1D",
		X"20",X"3E",X"02",X"CD",X"06",X"20",X"21",X"AD",X"51",X"11",X"20",X"00",X"01",X"24",X"06",X"71",
		X"19",X"10",X"FC",X"C9",X"3A",X"2E",X"42",X"3D",X"C0",X"3E",X"D0",X"DD",X"96",X"50",X"FE",X"E1",
		X"D8",X"3A",X"D7",X"42",X"DD",X"96",X"51",X"C6",X"0C",X"FE",X"19",X"D0",X"DD",X"36",X"00",X"0A",
		X"21",X"93",X"22",X"CD",X"1D",X"20",X"3E",X"01",X"CD",X"06",X"20",X"06",X"07",X"21",X"20",X"42",
		X"7E",X"3D",X"20",X"02",X"36",X"03",X"2C",X"2C",X"10",X"F6",X"3E",X"02",X"32",X"2E",X"42",X"AF",
		X"32",X"03",X"42",X"32",X"81",X"42",X"DD",X"6E",X"50",X"DD",X"66",X"51",X"22",X"7E",X"42",X"7C",
		X"ED",X"44",X"57",X"1E",X"00",X"CD",X"36",X"0B",X"2E",X"34",X"3A",X"FB",X"42",X"67",X"22",X"1E",
		X"42",X"F7",X"1B",X"50",X"03",X"02",X"24",X"24",X"67",X"24",X"24",X"67",X"F7",X"AD",X"51",X"01",
		X"06",X"43",X"24",X"19",X"15",X"0E",X"11",X"C9",X"DD",X"21",X"2E",X"42",X"DD",X"7E",X"00",X"FE",
		X"03",X"C0",X"3A",X"09",X"42",X"87",X"26",X"00",X"30",X"01",X"25",X"6F",X"29",X"29",X"29",X"DD",
		X"5E",X"40",X"DD",X"56",X"50",X"19",X"DD",X"75",X"40",X"DD",X"74",X"50",X"7C",X"FE",X"DD",X"38",
		X"35",X"DD",X"7E",X"51",X"DD",X"36",X"00",X"01",X"DD",X"36",X"50",X"00",X"DD",X"36",X"51",X"00",
		X"01",X"20",X"D0",X"B9",X"30",X"01",X"79",X"B8",X"38",X"01",X"78",X"CD",X"D8",X"07",X"21",X"1D",
		X"21",X"CD",X"4D",X"20",X"AF",X"CD",X"06",X"20",X"3A",X"08",X"40",X"A7",X"C8",X"3E",X"01",X"32",
		X"03",X"42",X"32",X"81",X"42",X"C9",X"E6",X"07",X"C0",X"CB",X"5C",X"2E",X"36",X"28",X"01",X"2C",
		X"3A",X"FB",X"42",X"67",X"22",X"1E",X"42",X"C9",X"CD",X"D4",X"0B",X"21",X"20",X"42",X"01",X"00",
		X"07",X"7E",X"FE",X"05",X"20",X"01",X"0C",X"2C",X"2C",X"10",X"F6",X"79",X"FE",X"03",X"28",X"15",
		X"06",X"07",X"21",X"20",X"42",X"7E",X"FE",X"05",X"20",X"02",X"36",X"03",X"2C",X"2C",X"10",X"F5",
		X"AF",X"32",X"00",X"42",X"C9",X"DD",X"7E",X"50",X"FE",X"58",X"30",X"3D",X"DD",X"E5",X"E1",X"2C",
		X"2C",X"7D",X"FE",X"2E",X"20",X"02",X"2E",X"20",X"7E",X"FE",X"05",X"20",X"F2",X"11",X"50",X"00",
		X"19",X"5E",X"2C",X"56",X"DD",X"6E",X"50",X"DD",X"66",X"51",X"CD",X"E1",X"03",X"67",X"7B",X"FE",
		X"10",X"D8",X"3A",X"04",X"42",X"87",X"5F",X"CD",X"97",X"03",X"DD",X"74",X"31",X"61",X"CD",X"97",
		X"03",X"3A",X"04",X"42",X"84",X"DD",X"77",X"30",X"C9",X"01",X"05",X"07",X"FD",X"21",X"20",X"42",
		X"C5",X"CD",X"60",X"0E",X"C1",X"FD",X"23",X"FD",X"23",X"10",X"F5",X"FD",X"21",X"2E",X"42",X"FD",
		X"2B",X"FD",X"2B",X"FD",X"7E",X"00",X"FE",X"08",X"20",X"F5",X"21",X"2E",X"42",X"2D",X"2D",X"7E",
		X"FE",X"06",X"20",X"F9",X"FD",X"36",X"F0",X"3A",X"11",X"F1",X"FF",X"19",X"7E",X"FD",X"77",X"F1",
		X"11",X"5F",X"00",X"19",X"7E",X"D6",X"10",X"FD",X"77",X"50",X"2C",X"7E",X"FD",X"77",X"51",X"C9",
		X"FD",X"7E",X"00",X"B9",X"C0",X"3A",X"01",X"42",X"87",X"87",X"FD",X"86",X"F1",X"21",X"B6",X"0E",
		X"E7",X"FD",X"77",X"00",X"3A",X"01",X"42",X"2F",X"C6",X"06",X"FD",X"77",X"F1",X"FD",X"7E",X"00",
		X"FE",X"06",X"28",X"0A",X"D6",X"09",X"C0",X"FD",X"77",X"50",X"FD",X"77",X"51",X"C9",X"FD",X"36",
		X"F0",X"3B",X"FD",X"6E",X"50",X"FD",X"66",X"51",X"3A",X"D7",X"42",X"57",X"1E",X"FF",X"FD",X"E5",
		X"CD",X"E1",X"03",X"FD",X"E1",X"67",X"3A",X"06",X"42",X"5F",X"CD",X"97",X"03",X"FD",X"74",X"31",
		X"61",X"CD",X"97",X"03",X"FD",X"74",X"30",X"C9",X"01",X"06",X"09",X"08",X"09",X"01",X"08",X"06",
		X"06",X"08",X"01",X"09",X"08",X"09",X"06",X"01",X"3A",X"2E",X"42",X"FE",X"03",X"28",X"0B",X"AF",
		X"DD",X"77",X"00",X"DD",X"77",X"50",X"DD",X"77",X"51",X"C9",X"2A",X"7E",X"42",X"7D",X"D6",X"10",
		X"DD",X"77",X"50",X"DD",X"74",X"51",X"E6",X"07",X"C0",X"DD",X"36",X"F0",X"3C",X"C9",X"DD",X"7E",
		X"50",X"FE",X"C0",X"30",X"26",X"CD",X"98",X"09",X"01",X"08",X"07",X"FD",X"21",X"20",X"42",X"FD",
		X"7E",X"00",X"B9",X"28",X"07",X"FD",X"23",X"FD",X"23",X"10",X"F4",X"C9",X"DD",X"7E",X"50",X"D6",
		X"10",X"FD",X"77",X"50",X"DD",X"7E",X"51",X"FD",X"77",X"51",X"C9",X"DD",X"7E",X"10",X"E6",X"06",
		X"21",X"E3",X"42",X"E7",X"DD",X"77",X"F1",X"DD",X"36",X"F0",X"2C",X"3A",X"04",X"42",X"DD",X"77",
		X"30",X"DD",X"36",X"00",X"01",X"01",X"09",X"07",X"FD",X"21",X"20",X"42",X"FD",X"7E",X"00",X"B9",
		X"28",X"07",X"FD",X"23",X"FD",X"23",X"10",X"F4",X"C9",X"FD",X"7E",X"10",X"E6",X"06",X"21",X"E3",
		X"42",X"E7",X"FD",X"77",X"F1",X"FD",X"36",X"F0",X"2C",X"DD",X"7E",X"50",X"FD",X"77",X"50",X"DD",
		X"7E",X"51",X"FD",X"77",X"51",X"3A",X"04",X"42",X"FD",X"77",X"30",X"FD",X"77",X"31",X"FD",X"36",
		X"00",X"01",X"01",X"08",X"07",X"FD",X"21",X"20",X"42",X"FD",X"7E",X"00",X"B9",X"28",X"07",X"FD",
		X"23",X"FD",X"23",X"10",X"F4",X"C9",X"FD",X"7E",X"10",X"E6",X"06",X"21",X"E3",X"42",X"E7",X"FD",
		X"77",X"F1",X"FD",X"36",X"F0",X"2C",X"DD",X"7E",X"50",X"FD",X"77",X"50",X"DD",X"7E",X"51",X"FD",
		X"77",X"51",X"3A",X"04",X"42",X"FD",X"77",X"30",X"ED",X"44",X"FD",X"77",X"31",X"FD",X"36",X"00",
		X"01",X"C9",X"3A",X"9E",X"42",X"A7",X"C8",X"3A",X"BE",X"42",X"DD",X"96",X"50",X"FE",X"0C",X"D0",
		X"3A",X"BF",X"42",X"DD",X"96",X"51",X"FE",X"10",X"D0",X"CD",X"74",X"06",X"CD",X"90",X"10",X"DD",
		X"7E",X"F1",X"21",X"3C",X"11",X"E7",X"DD",X"77",X"F1",X"DD",X"36",X"F0",X"3E",X"DD",X"36",X"00",
		X"0B",X"21",X"2E",X"42",X"2D",X"2D",X"7E",X"FE",X"08",X"20",X"F9",X"E5",X"FD",X"E1",X"FD",X"7E",
		X"50",X"C6",X"10",X"FD",X"77",X"50",X"36",X"04",X"01",X"8C",X"06",X"CF",X"21",X"4B",X"22",X"CD",
		X"1D",X"20",X"C9",X"3A",X"9E",X"42",X"A7",X"C8",X"3A",X"BE",X"42",X"DD",X"96",X"50",X"FE",X"0C",
		X"D0",X"3A",X"BF",X"42",X"DD",X"96",X"51",X"D6",X"01",X"FE",X"0E",X"D0",X"CD",X"74",X"06",X"CD",
		X"9D",X"10",X"DD",X"7E",X"F1",X"21",X"40",X"11",X"E7",X"DD",X"77",X"F1",X"DD",X"36",X"F0",X"2C",
		X"DD",X"36",X"00",X"0C",X"21",X"2E",X"42",X"2D",X"2D",X"7E",X"FE",X"09",X"20",X"F9",X"36",X"04",
		X"01",X"8C",X"06",X"CF",X"21",X"4B",X"22",X"CD",X"1D",X"20",X"C9",X"3A",X"9E",X"42",X"A7",X"C8",
		X"3A",X"BE",X"42",X"DD",X"96",X"50",X"FE",X"0C",X"D0",X"3A",X"BF",X"42",X"DD",X"96",X"51",X"D6",
		X"02",X"FE",X"0C",X"D0",X"CD",X"74",X"06",X"CD",X"AA",X"10",X"DD",X"E5",X"E1",X"36",X"04",X"01",
		X"8C",X"06",X"CF",X"21",X"4B",X"22",X"CD",X"1D",X"20",X"AF",X"32",X"03",X"42",X"32",X"81",X"42",
		X"3E",X"F0",X"D7",X"3A",X"80",X"42",X"32",X"81",X"42",X"3A",X"02",X"42",X"32",X"03",X"42",X"C9",
		X"21",X"1A",X"11",X"CD",X"B7",X"10",X"21",X"26",X"11",X"CD",X"EF",X"10",X"C9",X"21",X"1E",X"11",
		X"CD",X"B7",X"10",X"21",X"2E",X"11",X"CD",X"EF",X"10",X"C9",X"21",X"22",X"11",X"CD",X"B7",X"10",
		X"21",X"36",X"11",X"CD",X"EF",X"10",X"C9",X"3A",X"01",X"42",X"E7",X"FE",X"23",X"20",X"07",X"3E",
		X"13",X"CD",X"0A",X"03",X"3E",X"52",X"CD",X"0A",X"03",X"DD",X"7E",X"51",X"E6",X"F8",X"FE",X"18",
		X"30",X"02",X"3E",X"18",X"FE",X"C0",X"38",X"02",X"3E",X"C0",X"6F",X"26",X"00",X"29",X"29",X"DD",
		X"7E",X"50",X"E6",X"F8",X"0F",X"0F",X"0F",X"85",X"6F",X"11",X"21",X"50",X"19",X"EB",X"C9",X"3A",
		X"01",X"42",X"87",X"E7",X"4E",X"23",X"46",X"EB",X"11",X"20",X"00",X"7E",X"FE",X"24",X"20",X"08",
		X"E5",X"19",X"7E",X"E1",X"FE",X"24",X"28",X"03",X"2B",X"18",X"F0",X"71",X"19",X"70",X"3E",X"1E",
		X"D7",X"11",X"E0",X"FF",X"36",X"24",X"19",X"36",X"24",X"C9",X"22",X"32",X"42",X"52",X"32",X"52",
		X"62",X"13",X"52",X"72",X"13",X"23",X"C8",X"C9",X"C8",X"CA",X"C8",X"CB",X"C8",X"CC",X"C8",X"CA",
		X"C8",X"CC",X"C8",X"CD",X"CF",X"F4",X"C8",X"CC",X"C8",X"CE",X"CF",X"F4",X"CF",X"F5",X"03",X"05",
		X"02",X"04",X"05",X"04",X"03",X"02",X"3A",X"80",X"42",X"A7",X"C8",X"DD",X"21",X"90",X"42",X"06",
		X"07",X"C5",X"DD",X"7E",X"00",X"A7",X"C4",X"6B",X"11",X"DD",X"7E",X"01",X"A7",X"C4",X"A4",X"11",
		X"CD",X"EF",X"11",X"DD",X"23",X"DD",X"23",X"C1",X"10",X"E7",X"C9",X"26",X"00",X"87",X"30",X"01",
		X"25",X"6F",X"29",X"29",X"29",X"DD",X"5E",X"10",X"DD",X"56",X"20",X"19",X"DD",X"75",X"10",X"DD",
		X"74",X"20",X"7C",X"D6",X"10",X"FE",X"BD",X"D8",X"DD",X"7E",X"21",X"E6",X"F8",X"6F",X"D6",X"20",
		X"FE",X"C0",X"30",X"2D",X"26",X"00",X"29",X"29",X"11",X"19",X"50",X"19",X"36",X"42",X"01",X"CF",
		X"11",X"CF",X"18",X"1D",X"26",X"00",X"87",X"30",X"01",X"25",X"6F",X"29",X"29",X"29",X"DD",X"5E",
		X"11",X"DD",X"56",X"21",X"19",X"DD",X"75",X"11",X"DD",X"74",X"21",X"7C",X"D6",X"10",X"FE",X"E0",
		X"D8",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"20",X"DD",X"77",X"21",X"C9",X"3E",
		X"08",X"D7",X"36",X"98",X"C9",X"3A",X"D0",X"42",X"3D",X"C0",X"3E",X"B3",X"DD",X"96",X"50",X"FE",
		X"EA",X"D8",X"3A",X"D3",X"42",X"DD",X"96",X"51",X"C6",X"0B",X"FE",X"17",X"D0",X"18",X"19",X"3A",
		X"D0",X"42",X"3D",X"C0",X"3E",X"BF",X"DD",X"96",X"20",X"FE",X"F0",X"D8",X"3A",X"D3",X"42",X"DD",
		X"96",X"21",X"FE",X"F2",X"D8",X"CD",X"C1",X"11",X"AF",X"32",X"D0",X"42",X"01",X"11",X"12",X"CF",
		X"C9",X"3E",X"10",X"CD",X"10",X"13",X"3A",X"D3",X"42",X"FE",X"D0",X"38",X"02",X"3E",X"C8",X"E6",
		X"F8",X"6F",X"26",X"00",X"29",X"29",X"11",X"18",X"50",X"19",X"E5",X"11",X"20",X"00",X"36",X"A4",
		X"2C",X"36",X"A5",X"19",X"36",X"A7",X"2D",X"36",X"A6",X"19",X"36",X"A8",X"2C",X"36",X"A9",X"E1",
		X"3E",X"10",X"D7",X"E5",X"11",X"20",X"00",X"36",X"AA",X"2C",X"36",X"AB",X"19",X"36",X"AD",X"2D",
		X"36",X"AC",X"19",X"36",X"AE",X"2C",X"36",X"AF",X"E1",X"3E",X"10",X"D7",X"11",X"20",X"00",X"3E",
		X"24",X"77",X"2C",X"36",X"98",X"19",X"36",X"98",X"2D",X"77",X"19",X"77",X"2C",X"36",X"98",X"3E",
		X"2D",X"D7",X"3E",X"10",X"D7",X"3A",X"D0",X"42",X"A7",X"C0",X"21",X"2B",X"43",X"77",X"2C",X"77",
		X"2C",X"77",X"06",X"07",X"DD",X"21",X"20",X"42",X"DD",X"7E",X"50",X"D6",X"A0",X"FE",X"30",X"30",
		X"3F",X"DD",X"7E",X"51",X"E6",X"F8",X"0F",X"0F",X"0F",X"C5",X"47",X"11",X"2B",X"43",X"FE",X"0D",
		X"38",X"01",X"1C",X"D6",X"05",X"30",X"01",X"AF",X"FE",X"08",X"38",X"02",X"D6",X"08",X"FE",X"10",
		X"38",X"01",X"AF",X"4F",X"78",X"FE",X"05",X"38",X"0C",X"2F",X"C6",X"1E",X"38",X"01",X"AF",X"FE",
		X"05",X"38",X"02",X"3E",X"05",X"CD",X"EF",X"1B",X"C1",X"1A",X"B5",X"12",X"1C",X"1A",X"B4",X"12",
		X"DD",X"23",X"DD",X"23",X"10",X"B2",X"0E",X"17",X"0D",X"28",X"97",X"79",X"CB",X"2F",X"38",X"03",
		X"2F",X"C6",X"17",X"47",X"11",X"2B",X"43",X"FE",X"0B",X"38",X"03",X"1C",X"D6",X"08",X"21",X"03",
		X"00",X"A7",X"28",X"04",X"29",X"3D",X"20",X"FC",X"1A",X"A5",X"6F",X"1C",X"1A",X"A4",X"B5",X"20",
		X"D7",X"3E",X"04",X"80",X"87",X"87",X"87",X"32",X"D3",X"42",X"3E",X"01",X"32",X"D0",X"42",X"C9",
		X"47",X"3A",X"17",X"43",X"A7",X"C0",X"3E",X"01",X"32",X"03",X"68",X"78",X"D7",X"AF",X"32",X"03",
		X"68",X"C9",X"31",X"F3",X"23",X"3A",X"00",X"78",X"21",X"00",X"60",X"01",X"00",X"03",X"71",X"2C",
		X"7D",X"E6",X"07",X"20",X"F9",X"7C",X"C6",X"08",X"67",X"10",X"F3",X"21",X"00",X"40",X"11",X"00",
		X"04",X"71",X"23",X"1B",X"7B",X"B2",X"20",X"F9",X"3D",X"32",X"28",X"43",X"32",X"00",X"78",X"21",
		X"00",X"50",X"01",X"00",X"04",X"36",X"24",X"23",X"0B",X"79",X"B0",X"20",X"F8",X"AF",X"21",X"C8",
		X"42",X"06",X"04",X"77",X"2C",X"10",X"FC",X"32",X"D7",X"42",X"21",X"10",X"42",X"06",X"70",X"77",
		X"2C",X"10",X"FC",X"21",X"90",X"42",X"06",X"30",X"77",X"2C",X"10",X"FC",X"21",X"00",X"58",X"06",
		X"80",X"77",X"2C",X"10",X"FC",X"3A",X"08",X"43",X"47",X"C3",X"65",X"16",X"00",X"6F",X"67",X"22",
		X"06",X"70",X"C9",X"3A",X"00",X"70",X"4F",X"E6",X"01",X"21",X"D1",X"13",X"E7",X"32",X"0A",X"43",
		X"79",X"0F",X"4F",X"E6",X"01",X"32",X"0B",X"83",X"79",X"0F",X"4F",X"E6",X"01",X"C6",X"02",X"32",
		X"09",X"43",X"79",X"0F",X"E6",X"01",X"32",X"08",X"43",X"3A",X"00",X"68",X"07",X"4F",X"E6",X"01",
		X"26",X"05",X"28",X"02",X"26",X"03",X"79",X"07",X"2F",X"E6",X"01",X"3C",X"6F",X"22",X"0B",X"43",
		X"C9",X"15",X"20",X"00",X"0F",X"0F",X"E6",X"01",X"32",X"0D",X"43",X"C9",X"10",X"12",X"15",X"FF",
		X"31",X"00",X"44",X"CD",X"93",X"13",X"3E",X"01",X"32",X"03",X"70",X"01",X"00",X"28",X"3A",X"00",
		X"78",X"0D",X"20",X"FA",X"10",X"F8",X"00",X"00",X"00",X"00",X"00",X"AF",X"00",X"00",X"32",X"0E",
		X"43",X"AF",X"32",X"03",X"70",X"01",X"00",X"28",X"3A",X"00",X"78",X"AF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"52",X"14",X"3E",X"01",X"32",
		X"02",X"43",X"32",X"88",X"42",X"32",X"89",X"42",X"32",X"8A",X"42",X"32",X"01",X"70",X"32",X"04",
		X"70",X"2A",X"2E",X"43",X"7D",X"BC",X"28",X"F9",X"21",X"30",X"43",X"85",X"6F",X"D6",X"2C",X"E6",
		X"7F",X"32",X"2E",X"43",X"11",X"31",X"14",X"D5",X"5E",X"2C",X"56",X"D5",X"2C",X"5E",X"2C",X"56",
		X"EB",X"C9",X"CD",X"7C",X"14",X"DF",X"59",X"14",X"C9",X"CD",X"80",X"16",X"21",X"7C",X"42",X"35",
		X"28",X"6A",X"7E",X"FE",X"F0",X"D0",X"C6",X"10",X"FE",X"30",X"D8",X"2C",X"2C",X"77",X"E6",X"03",
		X"C0",X"CB",X"56",X"3E",X"34",X"28",X"01",X"3C",X"32",X"1E",X"42",X"C9",X"AF",X"32",X"02",X"42",
		X"32",X"03",X"42",X"32",X"2E",X"42",X"32",X"80",X"42",X"32",X"81",X"42",X"32",X"C0",X"42",X"32",
		X"C5",X"42",X"32",X"D0",X"42",X"32",X"D8",X"42",X"3C",X"32",X"17",X"43",X"CD",X"4F",X"13",X"21",
		X"72",X"1B",X"11",X"E0",X"42",X"01",X"20",X"00",X"ED",X"B0",X"CD",X"9D",X"18",X"CD",X"3F",X"03",
		X"CD",X"4A",X"16",X"CD",X"28",X"02",X"21",X"00",X"C0",X"22",X"7C",X"42",X"22",X"7E",X"42",X"21",
		X"2C",X"02",X"22",X"1C",X"42",X"21",X"34",X"06",X"22",X"1E",X"42",X"C9",X"DF",X"80",X"16",X"F7",
		X"47",X"51",X"01",X"0A",X"43",X"24",X"0E",X"16",X"24",X"0D",X"1B",X"0A",X"1E",X"10",X"3E",X"3C",
		X"D7",X"F7",X"CD",X"50",X"01",X"13",X"0E",X"15",X"0B",X"0A",X"1D",X"24",X"0E",X"0C",X"17",X"0A",
		X"1F",X"0D",X"0A",X"24",X"0E",X"1B",X"18",X"0C",X"1C",X"3E",X"3C",X"D7",X"F7",X"31",X"51",X"01",
		X"0D",X"00",X"00",X"05",X"01",X"24",X"00",X"00",X"00",X"01",X"24",X"00",X"00",X"05",X"F7",X"0F",
		X"53",X"03",X"02",X"E9",X"EC",X"ED",X"EB",X"EE",X"EF",X"3E",X"3C",X"D7",X"F7",X"33",X"51",X"01",
		X"0C",X"00",X"05",X"01",X"24",X"24",X"00",X"00",X"01",X"24",X"24",X"00",X"05",X"F7",X"12",X"53",
		X"02",X"02",X"B0",X"B1",X"B2",X"B3",X"3E",X"3C",X"D7",X"F7",X"35",X"51",X"01",X"0C",X"00",X"02",
		X"01",X"24",X"24",X"00",X"08",X"24",X"24",X"24",X"00",X"04",X"F7",X"14",X"53",X"02",X"02",X"B0",
		X"B1",X"B2",X"B3",X"3E",X"3C",X"D7",X"F7",X"37",X"51",X"01",X"0C",X"00",X"09",X"24",X"24",X"24",
		X"00",X"06",X"24",X"24",X"24",X"00",X"03",X"F7",X"16",X"53",X"02",X"02",X"B0",X"B1",X"B2",X"B3",
		X"3E",X"3C",X"D7",X"F7",X"39",X"51",X"01",X"0C",X"00",X"06",X"24",X"24",X"24",X"00",X"04",X"24",
		X"24",X"24",X"00",X"02",X"F7",X"18",X"53",X"02",X"02",X"B0",X"B1",X"B2",X"B3",X"3E",X"3C",X"D7",
		X"F7",X"9C",X"51",X"01",X"07",X"24",X"24",X"24",X"24",X"12",X"0A",X"1D",X"3E",X"3C",X"D7",X"11",
		X"EF",X"42",X"3E",X"03",X"12",X"1C",X"12",X"1C",X"12",X"F7",X"31",X"51",X"01",X"0D",X"00",X"00",
		X"00",X"01",X"24",X"00",X"00",X"06",X"24",X"24",X"00",X"00",X"04",X"3E",X"3C",X"D7",X"11",X"EF",
		X"42",X"3E",X"04",X"12",X"1C",X"12",X"1C",X"12",X"F7",X"31",X"51",X"01",X"0D",X"00",X"00",X"07",
		X"24",X"24",X"00",X"00",X"05",X"24",X"24",X"00",X"00",X"03",X"3E",X"3C",X"D7",X"11",X"EF",X"42",
		X"3E",X"05",X"12",X"1C",X"12",X"1C",X"12",X"F7",X"31",X"51",X"01",X"0D",X"00",X"00",X"05",X"24",
		X"24",X"00",X"00",X"03",X"24",X"24",X"00",X"00",X"02",X"3E",X"3C",X"D7",X"DF",X"73",X"16",X"CD",
		X"4F",X"13",X"CD",X"8C",X"07",X"CD",X"9D",X"18",X"CD",X"3F",X"03",X"3E",X"06",X"32",X"C1",X"42",
		X"AF",X"32",X"09",X"40",X"32",X"0B",X"40",X"CD",X"D9",X"18",X"AF",X"32",X"D0",X"42",X"3C",X"32",
		X"C0",X"42",X"32",X"C5",X"42",X"32",X"D8",X"42",X"32",X"02",X"42",X"32",X"80",X"42",X"3E",X"78",
		X"D7",X"3E",X"10",X"32",X"D1",X"42",X"CD",X"75",X"12",X"3E",X"08",X"32",X"D5",X"42",X"3E",X"01",
		X"32",X"2E",X"42",X"32",X"03",X"42",X"32",X"81",X"42",X"C9",X"3A",X"0B",X"43",X"A7",X"28",X"14",
		X"F7",X"FF",X"52",X"01",X"06",X"1D",X"12",X"0D",X"0E",X"1B",X"0C",X"3E",X"01",X"32",X"16",X"43",
		X"CD",X"B0",X"02",X"C9",X"C9",X"3A",X"03",X"43",X"A0",X"2F",X"C3",X"8C",X"13",X"00",X"00",X"00",
		X"1B",X"0F",X"C9",X"3A",X"08",X"40",X"A7",X"20",X"04",X"DF",X"52",X"14",X"C9",X"CD",X"23",X"1B",
		X"3A",X"15",X"43",X"A7",X"C8",X"11",X"88",X"02",X"21",X"80",X"40",X"06",X"20",X"4E",X"2C",X"7E",
		X"2C",X"BA",X"20",X"02",X"79",X"BB",X"28",X"06",X"2C",X"2C",X"10",X"F1",X"18",X"0B",X"7D",X"D6",
		X"82",X"0F",X"0F",X"C6",X"60",X"6F",X"7E",X"A7",X"C0",X"21",X"60",X"40",X"01",X"00",X"20",X"71",
		X"2C",X"10",X"FC",X"DF",X"58",X"17",X"AF",X"32",X"17",X"43",X"32",X"10",X"40",X"32",X"09",X"40",
		X"32",X"0B",X"40",X"32",X"02",X"42",X"32",X"03",X"42",X"32",X"2E",X"42",X"32",X"80",X"42",X"32",
		X"81",X"42",X"32",X"C0",X"42",X"32",X"C5",X"42",X"32",X"D0",X"42",X"32",X"D8",X"42",X"3C",X"32",
		X"19",X"43",X"3A",X"09",X"43",X"32",X"0A",X"40",X"CD",X"D9",X"18",X"CD",X"4F",X"13",X"21",X"52",
		X"1B",X"11",X"E0",X"42",X"01",X"20",X"00",X"ED",X"B0",X"CD",X"9D",X"18",X"CD",X"4A",X"16",X"CD",
		X"28",X"02",X"F7",X"ED",X"50",X"01",X"11",X"17",X"18",X"1D",X"1D",X"1E",X"0B",X"24",X"1D",X"1B",
		X"0A",X"1D",X"1C",X"24",X"11",X"1C",X"1E",X"19",X"3A",X"0A",X"43",X"3C",X"28",X"26",X"F7",X"94",
		X"50",X"01",X"18",X"1C",X"1D",X"19",X"24",X"00",X"00",X"00",X"24",X"24",X"24",X"1B",X"18",X"0F",
		X"24",X"10",X"17",X"12",X"14",X"24",X"1C",X"1E",X"17",X"18",X"0B",X"11",X"0A",X"43",X"21",X"94",
		X"51",X"CD",X"BB",X"02",X"F7",X"38",X"51",X"01",X"0E",X"02",X"08",X"09",X"01",X"24",X"1D",X"11",
		X"10",X"12",X"1B",X"22",X"19",X"18",X"0C",X"C9",X"3A",X"15",X"43",X"3D",X"20",X"15",X"F7",X"10",
		X"51",X"01",X"0E",X"24",X"22",X"15",X"17",X"18",X"24",X"1B",X"0E",X"22",X"0A",X"15",X"19",X"24",
		X"01",X"18",X"13",X"F7",X"10",X"51",X"01",X"0E",X"1C",X"1B",X"0E",X"22",X"0A",X"15",X"19",X"24",
		X"02",X"24",X"1B",X"18",X"24",X"01",X"CD",X"3F",X"03",X"21",X"00",X"68",X"AF",X"CB",X"46",X"20",
		X"0A",X"3A",X"15",X"43",X"3D",X"C8",X"CB",X"4E",X"C8",X"3E",X"01",X"32",X"02",X"43",X"DF",X"AF",
		X"18",X"3A",X"0B",X"43",X"A7",X"28",X"0C",X"3A",X"02",X"43",X"2F",X"C6",X"9A",X"21",X"15",X"43",
		X"86",X"27",X"77",X"AF",X"32",X"16",X"43",X"32",X"19",X"43",X"21",X"0D",X"40",X"77",X"2C",X"77",
		X"2C",X"77",X"21",X"2D",X"40",X"77",X"2C",X"77",X"2C",X"77",X"3C",X"32",X"C0",X"42",X"32",X"C5",
		X"42",X"32",X"D8",X"42",X"3E",X"C0",X"32",X"1C",X"43",X"21",X"00",X"40",X"11",X"20",X"40",X"06",
		X"20",X"7E",X"12",X"2C",X"1C",X"10",X"FA",X"3A",X"02",X"43",X"A7",X"20",X"09",X"21",X"20",X"40",
		X"06",X"20",X"77",X"2C",X"10",X"FC",X"21",X"07",X"22",X"CD",X"1D",X"20",X"CD",X"04",X"18",X"3E",
		X"F0",X"D7",X"18",X"45",X"CD",X"4F",X"13",X"CD",X"8C",X"07",X"CD",X"9D",X"18",X"CD",X"3F",X"03",
		X"CD",X"77",X"18",X"CD",X"50",X"19",X"3E",X"06",X"32",X"C1",X"42",X"AF",X"32",X"D0",X"42",X"32",
		X"C3",X"42",X"CD",X"74",X"08",X"3E",X"01",X"32",X"C0",X"42",X"32",X"C5",X"42",X"32",X"D8",X"42",
		X"32",X"1A",X"43",X"21",X"04",X"60",X"00",X"2C",X"77",X"2C",X"77",X"2C",X"77",X"21",X"00",X"68",
		X"77",X"2C",X"77",X"2C",X"77",X"C9",X"CD",X"04",X"18",X"3E",X"3C",X"D7",X"3E",X"10",X"32",X"D1",
		X"42",X"CD",X"75",X"12",X"3E",X"08",X"32",X"D5",X"42",X"3E",X"01",X"32",X"80",X"42",X"32",X"2E",
		X"42",X"21",X"0A",X"40",X"35",X"CD",X"77",X"18",X"3E",X"78",X"D7",X"3E",X"01",X"32",X"02",X"42",
		X"32",X"03",X"42",X"32",X"81",X"42",X"C9",X"3A",X"0A",X"40",X"4F",X"3E",X"05",X"91",X"FD",X"21",
		X"9E",X"52",X"11",X"40",X"00",X"28",X"08",X"47",X"CD",X"C8",X"19",X"FD",X"19",X"10",X"F9",X"79",
		X"A7",X"C8",X"47",X"3E",X"2C",X"CD",X"D7",X"19",X"FD",X"19",X"10",X"F7",X"C9",X"F7",X"60",X"51",
		X"01",X"0A",X"0E",X"1B",X"18",X"0C",X"1C",X"24",X"11",X"10",X"12",X"11",X"C3",X"29",X"03",X"3A",
		X"08",X"40",X"A7",X"C0",X"DF",X"26",X"00",X"AF",X"32",X"03",X"42",X"32",X"81",X"42",X"21",X"65",
		X"23",X"CD",X"4D",X"20",X"3E",X"B4",X"D7",X"DF",X"AF",X"18",X"CD",X"D9",X"18",X"3E",X"78",X"D7",
		X"3E",X"01",X"32",X"03",X"42",X"32",X"81",X"42",X"C9",X"3E",X"2A",X"32",X"08",X"40",X"3E",X"09",
		X"32",X"00",X"42",X"AF",X"32",X"C3",X"42",X"CD",X"74",X"08",X"21",X"C0",X"19",X"11",X"00",X"40",
		X"01",X"08",X"00",X"ED",X"B0",X"21",X"09",X"40",X"7E",X"C6",X"01",X"27",X"FE",X"49",X"30",X"01",
		X"77",X"21",X"0B",X"40",X"7E",X"A7",X"28",X"03",X"3A",X"0D",X"43",X"C6",X"01",X"86",X"38",X"01",
		X"77",X"21",X"E7",X"19",X"CD",X"33",X"1D",X"32",X"04",X"42",X"21",X"F9",X"19",X"CD",X"33",X"1D",
		X"32",X"05",X"42",X"21",X"0B",X"1A",X"CD",X"33",X"1D",X"32",X"06",X"42",X"21",X"0D",X"1A",X"CD",
		X"33",X"1D",X"32",X"07",X"42",X"21",X"21",X"1A",X"CD",X"33",X"1D",X"32",X"08",X"42",X"21",X"35",
		X"1A",X"CD",X"33",X"1D",X"32",X"09",X"42",X"21",X"37",X"1A",X"CD",X"33",X"1D",X"32",X"0A",X"42",
		X"21",X"00",X"00",X"22",X"84",X"42",X"21",X"5E",X"50",X"11",X"20",X"00",X"3A",X"09",X"40",X"E6",
		X"0F",X"28",X"2C",X"FE",X"05",X"28",X"1C",X"38",X"02",X"D6",X"05",X"47",X"36",X"FC",X"2C",X"36",
		X"FD",X"19",X"36",X"FF",X"2D",X"36",X"FE",X"19",X"10",X"F2",X"3A",X"09",X"40",X"E6",X"0F",X"FE",
		X"05",X"38",X"0C",X"36",X"26",X"2C",X"36",X"27",X"19",X"36",X"29",X"2D",X"36",X"28",X"19",X"3A",
		X"09",X"40",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"0F",X"47",X"36",X"2A",X"2C",X"36",X"27",
		X"19",X"36",X"29",X"2D",X"36",X"2B",X"19",X"10",X"F2",X"7C",X"FE",X"52",X"20",X"03",X"7D",X"FE",
		X"5E",X"C8",X"36",X"24",X"2C",X"36",X"24",X"19",X"36",X"24",X"2D",X"36",X"24",X"19",X"18",X"E9",
		X"FC",X"3F",X"FC",X"3F",X"F8",X"1F",X"F0",X"0F",X"3E",X"24",X"FD",X"77",X"00",X"FD",X"77",X"01",
		X"FD",X"77",X"20",X"FD",X"77",X"21",X"C9",X"FD",X"77",X"00",X"3C",X"FD",X"77",X"01",X"3C",X"FD",
		X"77",X"20",X"3C",X"FD",X"77",X"21",X"C9",X"01",X"10",X"02",X"12",X"03",X"14",X"04",X"15",X"06",
		X"16",X"07",X"14",X"0B",X"17",X"0C",X"14",X"FF",X"18",X"01",X"10",X"02",X"12",X"03",X"14",X"04",
		X"15",X"06",X"16",X"07",X"14",X"0B",X"17",X"0C",X"14",X"FF",X"18",X"FF",X"0C",X"01",X"10",X"02",
		X"12",X"03",X"14",X"04",X"15",X"06",X"16",X"07",X"12",X"09",X"17",X"0B",X"18",X"0C",X"14",X"FF",
		X"19",X"01",X"10",X"02",X"12",X"03",X"14",X"04",X"15",X"06",X"16",X"07",X"12",X"09",X"17",X"0B",
		X"18",X"0C",X"14",X"FF",X"19",X"FF",X"0E",X"FF",X"20",X"3A",X"17",X"43",X"A7",X"28",X"04",X"DF",
		X"52",X"14",X"C9",X"DF",X"26",X"00",X"AF",X"32",X"1A",X"43",X"32",X"02",X"42",X"32",X"03",X"42",
		X"32",X"2E",X"42",X"32",X"80",X"42",X"32",X"81",X"42",X"32",X"C0",X"42",X"32",X"C5",X"42",X"32",
		X"D0",X"42",X"32",X"D8",X"42",X"21",X"04",X"60",X"00",X"2C",X"77",X"2C",X"77",X"2C",X"77",X"21",
		X"00",X"68",X"77",X"2C",X"77",X"2C",X"77",X"3A",X"02",X"43",X"A7",X"28",X"2C",X"3A",X"0A",X"40",
		X"A7",X"20",X"15",X"01",X"88",X"1A",X"CF",X"C9",X"CD",X"09",X"1B",X"CD",X"E6",X"1A",X"3E",X"F0",
		X"D7",X"DF",X"95",X"1A",X"C9",X"DF",X"26",X"00",X"3A",X"2A",X"40",X"A7",X"28",X"0B",X"CD",X"CD",
		X"1A",X"01",X"46",X"18",X"CF",X"DF",X"AF",X"18",X"C9",X"3A",X"0A",X"40",X"A7",X"20",X"F2",X"01",
		X"B4",X"1A",X"CF",X"C9",X"AF",X"32",X"D8",X"42",X"CD",X"09",X"1B",X"3E",X"78",X"D7",X"3A",X"03",
		X"43",X"A7",X"C4",X"CD",X"1A",X"AF",X"32",X"1C",X"43",X"DF",X"52",X"14",X"C9",X"06",X"20",X"11",
		X"00",X"40",X"21",X"20",X"40",X"1A",X"4E",X"EB",X"12",X"71",X"1C",X"2C",X"10",X"F7",X"21",X"03",
		X"43",X"7E",X"EE",X"01",X"77",X"C9",X"F7",X"F2",X"51",X"01",X"06",X"1B",X"0E",X"22",X"0A",X"15",
		X"19",X"3A",X"03",X"43",X"A7",X"20",X"09",X"F7",X"72",X"51",X"01",X"03",X"0E",X"17",X"18",X"C9",
		X"F7",X"72",X"51",X"01",X"03",X"18",X"20",X"1D",X"C9",X"21",X"8D",X"51",X"11",X"20",X"00",X"01",
		X"24",X"09",X"71",X"19",X"10",X"FC",X"21",X"72",X"51",X"11",X"20",X"00",X"01",X"24",X"0A",X"71",
		X"19",X"10",X"FC",X"F7",X"94",X"51",X"01",X"09",X"1B",X"0E",X"1F",X"18",X"24",X"0E",X"16",X"0A",
		X"10",X"C9",X"07",X"07",X"07",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"00",X"00",X"03",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"06",X"06",X"06",X"06",
		X"01",X"01",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"04",X"04",X"04",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"01",X"01",X"01",X"01",
		X"01",X"01",X"21",X"89",X"42",X"35",X"C0",X"CD",X"15",X"1D",X"32",X"89",X"42",X"3A",X"03",X"42",
		X"A7",X"C8",X"3A",X"08",X"40",X"A7",X"C8",X"FE",X"0A",X"38",X"0A",X"21",X"00",X"42",X"7E",X"D6",
		X"01",X"DA",X"4A",X"1F",X"77",X"06",X"07",X"DD",X"21",X"20",X"42",X"DD",X"7E",X"00",X"A7",X"28",
		X"42",X"DD",X"23",X"DD",X"23",X"10",X"F4",X"C9",X"3A",X"C3",X"42",X"E6",X"F8",X"0F",X"0F",X"0F",
		X"47",X"2F",X"C6",X"02",X"FE",X"F0",X"38",X"01",X"AF",X"E6",X"0F",X"4F",X"78",X"FE",X"10",X"30",
		X"01",X"2F",X"E6",X"0F",X"3D",X"F2",X"E9",X"1B",X"AF",X"FE",X"0D",X"38",X"02",X"3E",X"0D",X"21",
		X"00",X"00",X"A7",X"28",X"06",X"47",X"37",X"ED",X"6A",X"10",X"FB",X"79",X"A7",X"C8",X"47",X"29",
		X"10",X"FD",X"C9",X"CD",X"C8",X"1B",X"FD",X"21",X"00",X"40",X"FD",X"7E",X"00",X"FD",X"B6",X"02",
		X"FD",X"B6",X"04",X"FD",X"B6",X"06",X"A5",X"5F",X"FD",X"7E",X"01",X"FD",X"B6",X"03",X"FD",X"B6",
		X"05",X"FD",X"B6",X"07",X"A4",X"57",X"21",X"08",X"40",X"3A",X"C1",X"42",X"87",X"38",X"19",X"01",
		X"00",X"01",X"78",X"A3",X"20",X"2C",X"0C",X"CB",X"00",X"30",X"F7",X"2C",X"0E",X"00",X"78",X"A2",
		X"20",X"20",X"0C",X"CB",X"00",X"30",X"F7",X"C9",X"2C",X"01",X"07",X"80",X"78",X"A2",X"20",X"12",
		X"0D",X"CB",X"08",X"30",X"F7",X"2D",X"0E",X"07",X"78",X"A3",X"20",X"06",X"0D",X"CB",X"08",X"30",
		X"F7",X"C9",X"2D",X"2D",X"78",X"A6",X"28",X"FA",X"AE",X"77",X"79",X"0F",X"0F",X"57",X"0F",X"85",
		X"D6",X"00",X"DD",X"77",X"10",X"7A",X"E6",X"C0",X"5F",X"7A",X"E6",X"01",X"57",X"7D",X"D6",X"00",
		X"0F",X"30",X"02",X"14",X"14",X"87",X"83",X"5F",X"FD",X"21",X"03",X"50",X"FD",X"19",X"CD",X"C8",
		X"19",X"DD",X"36",X"F0",X"2C",X"DD",X"7E",X"10",X"E6",X"1E",X"21",X"E3",X"42",X"E7",X"DD",X"77",
		X"F1",X"DD",X"7E",X"10",X"E6",X"E0",X"67",X"DD",X"7E",X"10",X"0F",X"CB",X"1C",X"87",X"87",X"87",
		X"87",X"C6",X"18",X"6F",X"DD",X"7E",X"10",X"E6",X"1E",X"0F",X"C6",X"C8",X"5F",X"16",X"42",X"1A",
		X"84",X"67",X"DD",X"75",X"50",X"DD",X"74",X"51",X"E5",X"21",X"82",X"42",X"7E",X"07",X"07",X"86",
		X"3C",X"77",X"E6",X"7F",X"C6",X"40",X"E1",X"57",X"1E",X"FF",X"CD",X"E1",X"03",X"67",X"3A",X"04",
		X"42",X"5F",X"CD",X"97",X"03",X"DD",X"74",X"31",X"61",X"CD",X"97",X"03",X"DD",X"74",X"30",X"DD",
		X"7E",X"10",X"0F",X"2F",X"E6",X"80",X"DD",X"77",X"21",X"DD",X"36",X"00",X"01",X"21",X"65",X"23",
		X"CD",X"1D",X"20",X"06",X"08",X"AF",X"21",X"00",X"40",X"B6",X"2C",X"10",X"FC",X"A7",X"C0",X"32",
		X"C3",X"42",X"C3",X"74",X"08",X"3A",X"08",X"40",X"FE",X"07",X"30",X"03",X"3E",X"0A",X"C9",X"21",
		X"4F",X"1D",X"3A",X"85",X"42",X"BE",X"23",X"38",X"06",X"28",X"04",X"23",X"23",X"18",X"F6",X"5E",
		X"23",X"56",X"EB",X"3A",X"0D",X"43",X"A7",X"3A",X"0B",X"40",X"20",X"09",X"FE",X"10",X"38",X"05",
		X"3E",X"0C",X"32",X"0B",X"40",X"3D",X"BE",X"23",X"38",X"03",X"23",X"18",X"F9",X"7E",X"C9",X"04",
		X"5E",X"1D",X"08",X"72",X"1D",X"0C",X"82",X"1D",X"10",X"92",X"1D",X"FF",X"9E",X"1D",X"01",X"78",
		X"02",X"50",X"03",X"46",X"04",X"3C",X"05",X"37",X"06",X"32",X"07",X"50",X"08",X"2D",X"09",X"28",
		X"FF",X"23",X"01",X"64",X"02",X"3C",X"03",X"32",X"05",X"2D",X"06",X"28",X"07",X"3C",X"08",X"23",
		X"FF",X"1E",X"01",X"50",X"02",X"32",X"03",X"28",X"05",X"23",X"06",X"1E",X"07",X"32",X"08",X"1E",
		X"FF",X"19",X"01",X"50",X"02",X"28",X"06",X"1E",X"07",X"28",X"08",X"19",X"FF",X"14",X"01",X"3C",
		X"03",X"1E",X"05",X"19",X"06",X"14",X"07",X"1E",X"FF",X"14",X"21",X"8A",X"42",X"35",X"C0",X"36",
		X"1E",X"3A",X"08",X"40",X"A7",X"C8",X"3A",X"D0",X"42",X"3D",X"C0",X"3A",X"81",X"42",X"A7",X"C8",
		X"01",X"00",X"07",X"21",X"90",X"42",X"7E",X"2C",X"B6",X"28",X"01",X"0C",X"2C",X"10",X"F7",X"21",
		X"B0",X"1E",X"3A",X"08",X"40",X"3D",X"BE",X"23",X"38",X"04",X"23",X"23",X"18",X"F8",X"5E",X"23",
		X"56",X"EB",X"CD",X"33",X"1D",X"3D",X"B9",X"D8",X"CD",X"C8",X"1B",X"DD",X"21",X"00",X"40",X"DD",
		X"7E",X"00",X"DD",X"B6",X"02",X"DD",X"B6",X"04",X"DD",X"B6",X"06",X"A5",X"5F",X"DD",X"7E",X"01",
		X"DD",X"B6",X"03",X"DD",X"B6",X"05",X"DD",X"B6",X"07",X"A4",X"57",X"DD",X"21",X"8E",X"42",X"DD",
		X"23",X"DD",X"23",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"20",X"F4",X"7A",X"B3",X"CA",X"8C",X"1E",
		X"CD",X"E9",X"1F",X"21",X"09",X"40",X"87",X"38",X"01",X"2D",X"4F",X"07",X"07",X"07",X"3C",X"47",
		X"3E",X"80",X"07",X"10",X"FD",X"47",X"2D",X"2D",X"78",X"A6",X"28",X"FA",X"61",X"7D",X"D6",X"00",
		X"6F",X"E6",X"1E",X"0F",X"C6",X"C8",X"5F",X"7D",X"0F",X"CB",X"1C",X"87",X"87",X"87",X"87",X"C6",
		X"24",X"6F",X"16",X"42",X"1A",X"C6",X"07",X"84",X"67",X"DD",X"75",X"20",X"DD",X"74",X"21",X"3A",
		X"D3",X"42",X"C6",X"08",X"57",X"1E",X"C8",X"CD",X"E1",X"03",X"67",X"C6",X"40",X"FE",X"81",X"38",
		X"0B",X"FE",X"40",X"0E",X"6E",X"26",X"40",X"F2",X"7C",X"1E",X"26",X"C0",X"1E",X"1C",X"CD",X"97",
		X"03",X"DD",X"74",X"01",X"61",X"CD",X"97",X"03",X"DD",X"74",X"00",X"C9",X"06",X"07",X"FD",X"21",
		X"20",X"42",X"FD",X"7E",X"00",X"3D",X"20",X"07",X"FD",X"7E",X"50",X"FE",X"80",X"38",X"07",X"FD",
		X"23",X"FD",X"23",X"10",X"ED",X"C9",X"C6",X"0C",X"6F",X"FD",X"7E",X"51",X"C6",X"07",X"18",X"A8",
		X"06",X"BC",X"1E",X"12",X"C8",X"1E",X"1E",X"D4",X"1E",X"FF",X"DC",X"1E",X"01",X"03",X"02",X"04",
		X"06",X"05",X"07",X"04",X"0E",X"06",X"FF",X"07",X"01",X"02",X"02",X"03",X"06",X"04",X"07",X"03",
		X"0E",X"05",X"FF",X"06",X"02",X"02",X"07",X"03",X"0E",X"04",X"FF",X"05",X"07",X"02",X"0E",X"03",
		X"FF",X"04",X"21",X"88",X"42",X"35",X"C0",X"36",X"10",X"3A",X"D8",X"42",X"A7",X"C8",X"21",X"C4",
		X"42",X"7E",X"3C",X"FE",X"0C",X"38",X"01",X"AF",X"77",X"21",X"00",X"40",X"4E",X"06",X"08",X"CB",
		X"01",X"DC",X"0D",X"1F",X"10",X"F9",X"2C",X"7D",X"FE",X"08",X"38",X"F0",X"C9",X"E5",X"11",X"00",
		X"40",X"19",X"EB",X"CB",X"3B",X"78",X"30",X"02",X"C6",X"08",X"3D",X"6F",X"26",X"00",X"29",X"29",
		X"29",X"29",X"29",X"19",X"29",X"EB",X"FD",X"21",X"03",X"50",X"FD",X"19",X"3A",X"C5",X"42",X"A7",
		X"28",X"03",X"3A",X"C4",X"42",X"21",X"3E",X"1F",X"E7",X"CD",X"D7",X"19",X"E1",X"C9",X"B0",X"B4",
		X"B8",X"BC",X"B8",X"B4",X"B0",X"B4",X"B8",X"BC",X"B8",X"B4",X"01",X"00",X"07",X"11",X"20",X"42",
		X"1A",X"A7",X"20",X"01",X"0C",X"1C",X"1C",X"10",X"F7",X"79",X"FE",X"03",X"D8",X"3E",X"09",X"32",
		X"00",X"42",X"CD",X"C8",X"1B",X"11",X"00",X"40",X"01",X"10",X"00",X"1A",X"A5",X"C5",X"47",X"1C",
		X"1A",X"A4",X"B0",X"C1",X"28",X"02",X"04",X"37",X"CB",X"11",X"1C",X"30",X"EE",X"78",X"FE",X"03",
		X"D8",X"3E",X"FF",X"28",X"0C",X"3A",X"D7",X"42",X"E6",X"03",X"3C",X"47",X"3E",X"7F",X"07",X"10",
		X"FD",X"A1",X"06",X"04",X"05",X"0F",X"38",X"FC",X"78",X"32",X"01",X"42",X"87",X"C6",X"00",X"4F",
		X"06",X"04",X"21",X"00",X"40",X"79",X"BD",X"28",X"0B",X"C5",X"E5",X"CD",X"BF",X"1F",X"DD",X"36",
		X"00",X"05",X"E1",X"C1",X"2C",X"2C",X"10",X"ED",X"21",X"65",X"23",X"CD",X"1D",X"20",X"C9",X"E5",
		X"5E",X"2C",X"56",X"CD",X"E9",X"1F",X"E1",X"87",X"30",X"01",X"2C",X"07",X"07",X"07",X"4F",X"3C",
		X"47",X"3E",X"80",X"07",X"10",X"FD",X"AE",X"77",X"DD",X"21",X"20",X"42",X"DD",X"7E",X"00",X"A7",
		X"CA",X"6A",X"1C",X"DD",X"23",X"DD",X"23",X"18",X"F3",X"21",X"82",X"42",X"7E",X"07",X"07",X"86",
		X"3C",X"77",X"0F",X"0F",X"0F",X"0F",X"AE",X"E6",X"0F",X"3C",X"47",X"EB",X"AF",X"D6",X"10",X"29",
		X"30",X"FB",X"2C",X"10",X"F8",X"C9",X"A7",X"28",X"0C",X"47",X"3A",X"17",X"43",X"A7",X"C0",X"3A",
		X"0E",X"43",X"A7",X"C0",X"78",X"32",X"00",X"70",X"0F",X"32",X"02",X"70",X"C9",X"3A",X"17",X"43",
		X"A7",X"C0",X"3A",X"0E",X"43",X"A7",X"20",X"03",X"7E",X"87",X"D8",X"CD",X"5B",X"20",X"36",X"01",
		X"2C",X"36",X"00",X"C9",X"3A",X"17",X"43",X"A7",X"C0",X"3A",X"0E",X"43",X"A7",X"20",X"03",X"7E",
		X"87",X"D8",X"CD",X"5B",X"20",X"7E",X"A7",X"C0",X"34",X"2C",X"36",X"00",X"C9",X"CD",X"5B",X"20",
		X"36",X"00",X"3E",X"FF",X"32",X"28",X"43",X"32",X"00",X"78",X"C9",X"11",X"FB",X"20",X"1A",X"13",
		X"BD",X"20",X"04",X"1A",X"BC",X"28",X"03",X"13",X"18",X"F4",X"21",X"44",X"1F",X"19",X"C9",X"06",
		X"10",X"DD",X"21",X"40",X"40",X"C5",X"CD",X"93",X"20",X"C1",X"DD",X"23",X"DD",X"23",X"10",X"F5",
		X"3A",X"26",X"43",X"32",X"07",X"68",X"3A",X"27",X"43",X"32",X"06",X"68",X"3A",X"28",X"43",X"32",
		X"00",X"78",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"3E",X"10",X"90",X"87",X"21",X"FB",X"20",X"E7",
		X"5F",X"23",X"56",X"6B",X"62",X"DD",X"7E",X"00",X"E7",X"47",X"07",X"07",X"32",X"26",X"43",X"07",
		X"32",X"27",X"43",X"78",X"E6",X"1F",X"21",X"DB",X"20",X"E7",X"32",X"28",X"43",X"78",X"87",X"30",
		X"05",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"7E",X"01",X"D6",X"01",X"38",X"04",X"DD",X"77",X"01",
		X"C9",X"1A",X"E6",X"7F",X"DD",X"77",X"01",X"DD",X"34",X"00",X"C9",X"00",X"0E",X"1C",X"29",X"35",
		X"40",X"4B",X"55",X"5E",X"67",X"70",X"78",X"7F",X"87",X"8D",X"94",X"9A",X"9F",X"A5",X"AA",X"AF",
		X"B3",X"B7",X"BB",X"BF",X"C3",X"C6",X"C9",X"CC",X"CF",X"D2",X"FF",X"65",X"23",X"65",X"23",X"4B",
		X"22",X"4B",X"22",X"4B",X"22",X"4B",X"22",X"1D",X"21",X"93",X"22",X"1B",X"21",X"1B",X"21",X"1B",
		X"21",X"1B",X"21",X"85",X"22",X"07",X"22",X"75",X"22",X"6B",X"22",X"00",X"9F",X"80",X"11",X"13",
		X"11",X"13",X"11",X"13",X"11",X"13",X"1D",X"1C",X"1A",X"18",X"16",X"15",X"13",X"11",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"05",X"07",
		X"05",X"07",X"05",X"07",X"05",X"07",X"11",X"10",X"0E",X"0C",X"0A",X"09",X"07",X"05",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0C",X"0E",
		X"0C",X"0E",X"0C",X"0E",X"0C",X"0E",X"18",X"17",X"15",X"13",X"11",X"10",X"0E",X"0C",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"0C",X"0B",X"09",X"07",X"05",X"04",X"02",X"00",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"11",X"13",X"11",X"13",X"11",X"13",X"11",X"13",X"1D",X"1C",
		X"1A",X"18",X"16",X"15",X"13",X"11",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"05",X"07",X"05",X"07",X"05",X"07",X"05",X"07",X"11",X"10",
		X"0E",X"0C",X"0A",X"09",X"07",X"05",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0C",X"0E",X"0C",X"0E",X"0C",X"0E",X"0C",X"0E",X"18",X"17",
		X"15",X"13",X"11",X"10",X"0E",X"0C",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"0C",X"0B",
		X"09",X"07",X"05",X"04",X"02",X"00",X"9F",X"04",X"5A",X"5A",X"5A",X"1F",X"58",X"55",X"55",X"1F",
		X"53",X"5A",X"5A",X"1F",X"58",X"55",X"55",X"1F",X"53",X"5C",X"5A",X"58",X"57",X"55",X"53",X"52",
		X"50",X"4E",X"50",X"52",X"53",X"55",X"57",X"58",X"5A",X"5C",X"5A",X"5A",X"1F",X"58",X"55",X"55",
		X"1F",X"53",X"5A",X"5A",X"1F",X"58",X"55",X"55",X"1F",X"53",X"4E",X"50",X"4E",X"50",X"53",X"55",
		X"53",X"55",X"58",X"5A",X"58",X"5A",X"5C",X"5E",X"5C",X"5E",X"9F",X"00",X"00",X"11",X"02",X"13",
		X"05",X"18",X"0B",X"1D",X"0E",X"1E",X"00",X"1E",X"0E",X"00",X"1E",X"0E",X"1D",X"0C",X"1B",X"0A",
		X"10",X"08",X"17",X"05",X"14",X"03",X"12",X"02",X"11",X"01",X"9F",X"00",X"60",X"62",X"64",X"65",
		X"67",X"69",X"6B",X"6C",X"9F",X"04",X"7E",X"1F",X"7E",X"1F",X"7E",X"1F",X"7E",X"1F",X"7E",X"1F",
		X"7E",X"1F",X"7E",X"7E",X"9F",X"85",X"0C",X"0C",X"1F",X"07",X"09",X"1F",X"07",X"09",X"1F",X"0C",
		X"1F",X"0C",X"9F",X"80",X"00",X"02",X"03",X"04",X"05",X"04",X"03",X"02",X"01",X"03",X"04",X"05",
		X"06",X"05",X"04",X"03",X"02",X"04",X"05",X"06",X"07",X"06",X"05",X"04",X"03",X"05",X"06",X"07",
		X"08",X"07",X"06",X"05",X"04",X"06",X"07",X"08",X"09",X"08",X"07",X"06",X"05",X"07",X"08",X"09",
		X"0A",X"09",X"08",X"07",X"06",X"08",X"09",X"0A",X"0B",X"0A",X"09",X"08",X"07",X"09",X"0A",X"0B",
		X"0C",X"0B",X"0A",X"09",X"08",X"0A",X"0B",X"0C",X"0D",X"0C",X"0B",X"0A",X"09",X"0B",X"0C",X"0D",
		X"0E",X"0D",X"0C",X"0B",X"0A",X"0C",X"0D",X"0E",X"0F",X"0E",X"0D",X"0C",X"0B",X"0D",X"0E",X"0F",
		X"10",X"0F",X"0E",X"0D",X"0C",X"0E",X"0F",X"10",X"11",X"10",X"0F",X"0E",X"0D",X"0F",X"10",X"11",
		X"12",X"11",X"10",X"1F",X"0E",X"10",X"11",X"12",X"13",X"12",X"11",X"10",X"0F",X"11",X"12",X"13",
		X"14",X"13",X"12",X"11",X"10",X"12",X"13",X"14",X"15",X"14",X"13",X"12",X"11",X"13",X"14",X"15",
		X"16",X"15",X"14",X"13",X"12",X"14",X"15",X"16",X"17",X"16",X"15",X"14",X"13",X"15",X"16",X"17",
		X"18",X"17",X"16",X"15",X"14",X"16",X"17",X"18",X"19",X"18",X"17",X"16",X"15",X"17",X"18",X"19",
		X"1A",X"19",X"18",X"17",X"16",X"18",X"19",X"1A",X"1B",X"1A",X"19",X"18",X"17",X"19",X"1A",X"1B",
		X"1C",X"1B",X"1A",X"19",X"18",X"1A",X"1B",X"1C",X"1D",X"1C",X"1B",X"1A",X"19",X"1B",X"1C",X"1D",
		X"1E",X"1D",X"1C",X"1B",X"9F",X"00",X"10",X"0E",X"0D",X"0C",X"0B",X"0C",X"0D",X"0E",X"0F",X"0D",
		X"0C",X"0B",X"0A",X"0B",X"0C",X"0D",X"0E",X"0C",X"0B",X"0A",X"09",X"0A",X"0B",X"0C",X"0D",X"0B",
		X"0A",X"09",X"08",X"09",X"0A",X"0B",X"0C",X"0A",X"09",X"08",X"07",X"08",X"09",X"0A",X"0B",X"09",
		X"08",X"07",X"06",X"07",X"08",X"09",X"0A",X"08",X"07",X"06",X"05",X"06",X"07",X"08",X"09",X"08",
		X"07",X"06",X"05",X"04",X"05",X"06",X"07",X"08",X"06",X"05",X"04",X"03",X"04",X"05",X"06",X"07",
		X"05",X"04",X"03",X"02",X"03",X"04",X"05",X"06",X"05",X"04",X"03",X"02",X"01",X"02",X"03",X"04",
		X"05",X"03",X"02",X"01",X"00",X"01",X"02",X"03",X"9F",X"F5",X"23",X"48",X"24",X"00",X"40",X"0F",
		X"04",X"48",X"24",X"00",X"40",X"F0",X"04",X"CF",X"24",X"48",X"24",X"00",X"50",X"0F",X"04",X"48",
		X"24",X"00",X"50",X"F0",X"04",X"48",X"24",X"00",X"58",X"0F",X"01",X"48",X"24",X"00",X"58",X"F0",
		X"01",X"C6",X"24",X"E5",X"24",X"11",X"FC",X"26",X"21",X"00",X"00",X"01",X"00",X"10",X"3A",X"00",
		X"78",X"79",X"86",X"4F",X"2C",X"20",X"FA",X"24",X"10",X"F4",X"1A",X"B9",X"20",X"00",X"13",X"7B",
		X"FE",X"FE",X"38",X"E7",X"01",X"00",X"08",X"28",X"E5",X"3E",X"18",X"32",X"02",X"52",X"3E",X"14",
		X"18",X"03",X"7B",X"D6",X"FB",X"21",X"E2",X"51",X"77",X"06",X"18",X"21",X"A2",X"52",X"11",X"20",
		X"00",X"36",X"16",X"19",X"70",X"19",X"36",X"1B",X"FE",X"14",X"C8",X"3A",X"00",X"78",X"3A",X"00",
		X"60",X"CB",X"77",X"20",X"F6",X"C3",X"00",X"00",X"16",X"0F",X"E1",X"C1",X"5A",X"3A",X"00",X"78",
		X"7B",X"0F",X"0F",X"0F",X"0F",X"83",X"80",X"A1",X"77",X"7B",X"87",X"87",X"83",X"3C",X"5F",X"2C",
		X"20",X"EE",X"24",X"10",X"E8",X"3B",X"3B",X"3B",X"3B",X"E1",X"C1",X"5A",X"3A",X"00",X"78",X"7B",
		X"0F",X"0F",X"0F",X"0F",X"83",X"80",X"AE",X"A1",X"20",X"17",X"7B",X"87",X"87",X"83",X"3C",X"5F",
		X"2C",X"20",X"EC",X"24",X"10",X"E6",X"15",X"3B",X"3B",X"3B",X"3B",X"F2",X"4A",X"24",X"E1",X"C1",
		X"C9",X"79",X"E6",X"01",X"4F",X"7C",X"0F",X"0F",X"E6",X"06",X"20",X"02",X"3E",X"02",X"93",X"FE",
		X"03",X"38",X"17",X"4F",X"21",X"00",X"50",X"11",X"00",X"40",X"06",X"04",X"3A",X"00",X"78",X"1A",
		X"77",X"1C",X"2C",X"20",X"FA",X"14",X"24",X"10",X"F3",X"79",X"21",X"E4",X"51",X"77",X"06",X"0A",
		X"21",X"A4",X"52",X"C3",X"2E",X"24",X"3E",X"18",X"32",X"04",X"42",X"3E",X"14",X"18",X"D4",X"21",
		X"00",X"40",X"11",X"00",X"50",X"01",X"00",X"04",X"3A",X"00",X"78",X"1A",X"77",X"23",X"13",X"0B",
		X"79",X"B0",X"20",X"F4",X"C9",X"31",X"00",X"44",X"3A",X"00",X"78",X"21",X"00",X"58",X"01",X"00",
		X"80",X"71",X"2C",X"10",X"FC",X"01",X"05",X"20",X"21",X"01",X"58",X"71",X"2C",X"2C",X"10",X"FB",
		X"AF",X"32",X"04",X"70",X"01",X"00",X"28",X"3A",X"00",X"78",X"0D",X"20",X"FA",X"10",X"F8",X"3A",
		X"00",X"78",X"3A",X"00",X"68",X"CB",X"6F",X"20",X"00",X"3E",X"01",X"32",X"04",X"70",X"01",X"00",
		X"28",X"3A",X"00",X"78",X"0D",X"20",X"FA",X"10",X"F8",X"3A",X"00",X"78",X"3A",X"00",X"68",X"CB",
		X"6F",X"28",X"00",X"3A",X"00",X"78",X"3A",X"00",X"68",X"CB",X"6F",X"20",X"00",X"3E",X"01",X"32",
		X"00",X"60",X"32",X"01",X"60",X"32",X"02",X"60",X"32",X"04",X"43",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AF",X"00",X"00",X"32",X"01",X"70",X"32",X"04",X"43",X"3D",X"C3",X"82",X"25",X"21",
		X"00",X"50",X"01",X"00",X"04",X"36",X"F6",X"23",X"0B",X"79",X"B0",X"20",X"F8",X"01",X"00",X"00",
		X"3A",X"00",X"78",X"0D",X"20",X"FA",X"10",X"F8",X"3A",X"00",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"86",X"25",X"C9",X"25",X"13",X"E0",X"13",X"CD",X"93",X"13",X"CD",X"9F",X"25",
		X"CD",X"BF",X"25",X"CD",X"13",X"26",X"CD",X"45",X"26",X"CD",X"55",X"26",X"C3",X"1A",X"01",X"C9",
		X"01",X"B2",X"25",X"CF",X"21",X"10",X"43",X"C3",X"7A",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C9",X"3A",X"0B",X"43",X"21",X"14",X"43",X"34",X"96",X"C0",X"77",X"3C",X"C3",X"A0",X"02",
		X"3E",X"08",X"D7",X"7E",X"2F",X"E6",X"01",X"32",X"03",X"60",X"35",X"C2",X"85",X"02",X"C9",X"7D",
		X"FE",X"10",X"CA",X"C3",X"25",X"7E",X"2F",X"E6",X"01",X"32",X"04",X"68",X"35",X"C2",X"85",X"02",
		X"C9",X"24",X"32",X"08",X"52",X"28",X"02",X"3E",X"1C",X"32",X"28",X"52",X"3A",X"0C",X"43",X"32",
		X"E8",X"51",X"3D",X"3E",X"24",X"28",X"02",X"3E",X"1C",X"32",X"E8",X"50",X"F7",X"08",X"51",X"01",
		X"07",X"1D",X"12",X"0D",X"0E",X"1B",X"0C",X"24",X"F7",X"48",X"52",X"01",X"05",X"17",X"12",X"18",
		X"0C",X"24",X"C9",X"F7",X"2A",X"52",X"01",X"07",X"24",X"24",X"1C",X"1E",X"17",X"18",X"0B",X"3A",
		X"0A",X"43",X"3C",X"28",X"13",X"F7",X"4A",X"51",X"01",X"05",X"24",X"24",X"00",X"00",X"00",X"21",
		X"0A",X"52",X"11",X"0A",X"43",X"C3",X"BB",X"02",X"F7",X"4A",X"51",X"01",X"07",X"10",X"17",X"12",
		X"11",X"1D",X"18",X"17",X"C9",X"F7",X"8C",X"52",X"01",X"04",X"10",X"17",X"12",X"14",X"3A",X"09",
		X"43",X"32",X"EC",X"51",X"C9",X"3E",X"01",X"32",X"06",X"68",X"32",X"07",X"68",X"01",X"FF",X"0B",
		X"DD",X"21",X"CD",X"26",X"21",X"00",X"41",X"E5",X"DD",X"7E",X"00",X"E6",X"F8",X"57",X"1E",X"00",
		X"DD",X"7E",X"00",X"E6",X"07",X"3C",X"C5",X"47",X"1A",X"2F",X"0F",X"10",X"FD",X"C1",X"38",X"03",
		X"DD",X"4E",X"01",X"7E",X"17",X"77",X"E6",X"0F",X"FE",X"0C",X"CC",X"BF",X"26",X"E1",X"2C",X"DD",
		X"23",X"DD",X"23",X"10",X"D2",X"79",X"32",X"00",X"78",X"21",X"10",X"41",X"11",X"E3",X"26",X"06",
		X"10",X"1A",X"FE",X"FF",X"28",X"02",X"BE",X"C0",X"13",X"2C",X"10",X"F5",X"F7",X"78",X"51",X"01",
		X"0D",X"18",X"0C",X"16",X"0A",X"17",X"24",X"22",X"0B",X"24",X"0E",X"0D",X"0A",X"16",X"C9",X"C5",
		X"06",X"10",X"21",X"10",X"41",X"7E",X"71",X"2C",X"4F",X"10",X"FA",X"C1",X"C9",X"A2",X"00",X"A3",
		X"1C",X"A4",X"35",X"A8",X"40",X"A9",X"55",X"AA",X"67",X"AB",X"78",X"AC",X"7F",X"A7",X"8D",X"A0",
		X"9A",X"A1",X"9F",X"55",X"55",X"55",X"40",X"35",X"1C",X"00",X"1C",X"1C",X"40",X"35",X"35",X"55",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"B3",X"90",X"B1",
		X"00",X"03",X"06",X"09",X"0C",X"10",X"13",X"16",X"19",X"1C",X"1F",X"22",X"25",X"28",X"2B",X"2E",
		X"31",X"33",X"36",X"39",X"3C",X"3F",X"41",X"44",X"47",X"49",X"4C",X"4E",X"51",X"53",X"55",X"58",
		X"5A",X"5C",X"5E",X"60",X"62",X"64",X"66",X"68",X"6A",X"6B",X"6D",X"6F",X"70",X"71",X"73",X"74",
		X"75",X"76",X"78",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7C",X"7B",X"7A",X"7A",X"79",X"78",X"76",
		X"75",X"74",X"73",X"71",X"70",X"6F",X"6D",X"6B",X"6A",X"68",X"66",X"64",X"62",X"60",X"5E",X"5C",
		X"5A",X"58",X"55",X"53",X"51",X"4E",X"4C",X"49",X"47",X"44",X"41",X"3F",X"3C",X"39",X"36",X"33",
		X"31",X"2E",X"2B",X"28",X"25",X"22",X"1F",X"1C",X"19",X"16",X"13",X"10",X"0C",X"09",X"06",X"03",
		X"00",X"FD",X"FA",X"F7",X"F4",X"F0",X"ED",X"EA",X"E7",X"E4",X"E1",X"DE",X"DB",X"D8",X"D5",X"D2",
		X"CF",X"CD",X"CA",X"C7",X"C4",X"C1",X"BF",X"BC",X"B9",X"B7",X"B4",X"B2",X"AF",X"AD",X"AB",X"A8",
		X"A6",X"A4",X"A2",X"A0",X"9E",X"9C",X"9A",X"98",X"96",X"95",X"93",X"91",X"90",X"8F",X"8D",X"8C",
		X"8B",X"8A",X"88",X"87",X"86",X"86",X"85",X"84",X"83",X"83",X"82",X"82",X"82",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"84",X"85",X"86",X"86",X"87",X"88",X"8A",
		X"8B",X"8C",X"8D",X"8F",X"90",X"91",X"93",X"95",X"96",X"98",X"9A",X"9C",X"9E",X"A0",X"A2",X"A4",
		X"A6",X"A8",X"AB",X"AD",X"AF",X"B2",X"B4",X"B7",X"B9",X"BC",X"BF",X"C1",X"C4",X"C7",X"CA",X"CD",
		X"CF",X"D2",X"D5",X"D8",X"DB",X"DE",X"E1",X"E4",X"E7",X"EA",X"ED",X"F0",X"F4",X"F7",X"FA",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
