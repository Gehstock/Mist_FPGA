library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps26 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps26 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CD",X"C2",X"06",X"CD",X"99",X"50",X"01",X"00",X"51",X"CD",X"64",X"0A",X"21",X"1E",X"26",X"11",
		X"45",X"51",X"0E",X"19",X"CD",X"E6",X"02",X"21",X"1C",X"2A",X"11",X"60",X"51",X"0E",X"12",X"CD",
		X"E6",X"02",X"21",X"18",X"27",X"11",X"73",X"51",X"E5",X"00",X"1A",X"FE",X"FF",X"CA",X"3B",X"50",
		X"0E",X"03",X"CD",X"E6",X"02",X"E1",X"2D",X"2D",X"C3",X"28",X"50",X"E1",X"21",X"06",X"26",X"11",
		X"8F",X"51",X"0E",X"04",X"CD",X"E6",X"02",X"21",X"1A",X"2C",X"11",X"93",X"51",X"0E",X"10",X"CD",
		X"E6",X"02",X"21",X"18",X"2C",X"11",X"51",X"21",X"E5",X"D5",X"0E",X"02",X"1B",X"1A",X"13",X"FE",
		X"FF",X"CA",X"7B",X"50",X"1A",X"CD",X"30",X"03",X"1B",X"0D",X"C2",X"5C",X"50",X"3E",X"1C",X"CD",
		X"F2",X"02",X"D1",X"E1",X"13",X"13",X"2D",X"2D",X"C3",X"58",X"50",X"D1",X"E1",X"21",X"18",X"36",
		X"11",X"65",X"21",X"E5",X"1A",X"FE",X"FF",X"CA",X"95",X"50",X"0E",X"03",X"CD",X"54",X"03",X"E1",
		X"2D",X"2D",X"C3",X"83",X"50",X"E1",X"C3",X"73",X"03",X"21",X"14",X"23",X"11",X"50",X"21",X"06",
		X"02",X"CD",X"BB",X"04",X"C3",X"A0",X"04",X"CD",X"55",X"16",X"21",X"50",X"21",X"11",X"C0",X"50",
		X"06",X"34",X"CD",X"BB",X"04",X"21",X"50",X"22",X"11",X"C0",X"50",X"06",X"34",X"C3",X"F4",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"FF",X"CD",X"BB",X"04",X"3E",X"00",X"32",X"91",X"21",X"C9",X"00",X"00",X"00",
		X"1E",X"C6",X"01",X"30",X"06",X"1C",X"C6",X"01",X"30",X"02",X"1A",X"C6",X"01",X"30",X"03",X"18",
		X"C6",X"01",X"30",X"06",X"16",X"C6",X"01",X"30",X"02",X"14",X"C6",X"01",X"30",X"03",X"12",X"C6",
		X"01",X"30",X"05",X"10",X"C6",X"01",X"30",X"04",X"0E",X"C6",X"01",X"30",X"08",X"0C",X"C6",X"01",
		X"30",X"03",X"0A",X"C6",X"01",X"30",X"02",X"08",X"C6",X"01",X"30",X"04",X"06",X"C6",X"01",X"30",
		X"01",X"FF",X"00",X"00",X"00",X"29",X"1B",X"01",X"04",X"12",X"13",X"1B",X"12",X"02",X"0E",X"11",
		X"04",X"11",X"12",X"1B",X"0E",X"05",X"1B",X"13",X"0E",X"03",X"00",X"18",X"1B",X"29",X"00",X"00",
		X"29",X"1B",X"13",X"0E",X"0F",X"1B",X"1D",X"1C",X"1B",X"0F",X"0B",X"00",X"18",X"04",X"11",X"12",
		X"1B",X"29",X"00",X"1D",X"12",X"13",X"1E",X"0D",X"03",X"1F",X"11",X"03",X"20",X"13",X"07",X"21",
		X"13",X"07",X"22",X"13",X"07",X"23",X"13",X"07",X"24",X"13",X"07",X"25",X"13",X"07",X"FF",X"1D",
		X"1C",X"13",X"07",X"12",X"02",X"0E",X"11",X"04",X"1B",X"1B",X"1B",X"1B",X"08",X"0D",X"08",X"13",
		X"08",X"00",X"0B",X"00",X"00",X"00",X"00",X"3A",X"91",X"21",X"A7",X"CA",X"87",X"00",X"DB",X"01",
		X"E6",X"06",X"C4",X"D6",X"51",X"CD",X"05",X"04",X"E6",X"08",X"06",X"01",X"21",X"84",X"21",X"C2",
		X"CB",X"51",X"7E",X"A7",X"23",X"C2",X"CB",X"51",X"2B",X"06",X"00",X"70",X"2A",X"8E",X"21",X"23",
		X"22",X"8E",X"21",X"C3",X"87",X"00",X"3E",X"01",X"32",X"96",X"21",X"C9",X"3E",X"20",X"C3",X"78",
		X"03",X"3E",X"05",X"C3",X"78",X"03",X"01",X"50",X"06",X"CD",X"05",X"04",X"E6",X"50",X"CA",X"FA",
		X"51",X"0D",X"C2",X"E9",X"51",X"05",X"C2",X"E9",X"51",X"C9",X"E1",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"C5",X"E5",X"AF",X"77",X"23",X"77",X"23",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",X"C2",
		X"01",X"52",X"C9",X"FE",X"40",X"CC",X"39",X"54",X"C3",X"87",X"53",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"6E",X"03",X"21",X"84",X"21",X"11",X"84",X"56",X"06",X"14",X"CD",X"BB",X"04",X"00",X"00",
		X"CD",X"A0",X"04",X"01",X"00",X"56",X"CD",X"64",X"0A",X"21",X"19",X"26",X"11",X"33",X"56",X"0E",
		X"18",X"CD",X"E6",X"02",X"21",X"15",X"27",X"11",X"84",X"41",X"CD",X"40",X"53",X"21",X"13",X"27",
		X"CD",X"40",X"53",X"21",X"11",X"27",X"0E",X"05",X"CD",X"42",X"53",X"C3",X"52",X"53",X"00",X"00",
		X"0E",X"0B",X"06",X"05",X"CD",X"DB",X"03",X"C5",X"01",X"60",X"01",X"09",X"C1",X"0D",X"C2",X"42",
		X"53",X"C9",X"21",X"11",X"31",X"11",X"4B",X"56",X"06",X"28",X"CD",X"DB",X"03",X"21",X"0B",X"27",
		X"11",X"73",X"56",X"0E",X"0F",X"CD",X"E6",X"02",X"3A",X"91",X"21",X"A7",X"CA",X"32",X"55",X"3A",
		X"8F",X"21",X"FE",X"20",X"D2",X"32",X"55",X"CD",X"CA",X"53",X"CD",X"05",X"04",X"E6",X"50",X"FE",
		X"10",X"CC",X"E3",X"53",X"C3",X"13",X"52",X"3A",X"96",X"21",X"A7",X"C2",X"32",X"55",X"3A",X"85",
		X"21",X"A7",X"C2",X"83",X"54",X"01",X"30",X"01",X"CD",X"DA",X"53",X"00",X"00",X"00",X"3A",X"8F",
		X"21",X"FE",X"1D",X"C2",X"68",X"53",X"06",X"05",X"C5",X"21",X"0B",X"27",X"06",X"20",X"CD",X"01",
		X"52",X"CD",X"E1",X"51",X"11",X"73",X"56",X"21",X"0B",X"27",X"0E",X"07",X"CD",X"E6",X"02",X"CD",
		X"E1",X"51",X"C1",X"05",X"C2",X"A8",X"53",X"C3",X"68",X"53",X"2A",X"92",X"21",X"3E",X"2A",X"C3",
		X"F2",X"02",X"2A",X"92",X"21",X"3E",X"1B",X"C3",X"F2",X"02",X"0D",X"C2",X"DA",X"53",X"05",X"C2",
		X"DA",X"53",X"C9",X"CD",X"E6",X"51",X"CD",X"D2",X"53",X"2A",X"92",X"21",X"7D",X"FE",X"14",X"CA",
		X"14",X"54",X"FE",X"12",X"CA",X"1D",X"54",X"7C",X"FE",X"31",X"CA",X"28",X"54",X"24",X"24",X"7C",
		X"FE",X"33",X"D2",X"08",X"54",X"C3",X"0E",X"54",X"CD",X"D2",X"53",X"21",X"10",X"34",X"22",X"92",
		X"21",X"C3",X"CA",X"53",X"7C",X"FE",X"3B",X"D2",X"2D",X"54",X"C3",X"23",X"54",X"7C",X"FE",X"3B",
		X"D2",X"33",X"54",X"24",X"24",X"C3",X"0E",X"54",X"26",X"32",X"C3",X"FD",X"53",X"21",X"12",X"27",
		X"C3",X"0E",X"54",X"21",X"10",X"27",X"C3",X"0E",X"54",X"CD",X"E6",X"51",X"CD",X"D2",X"53",X"2A",
		X"92",X"21",X"7D",X"FE",X"14",X"CA",X"5D",X"54",X"FE",X"12",X"CA",X"6E",X"54",X"7C",X"FE",X"28",
		X"DA",X"77",X"54",X"FE",X"32",X"C2",X"63",X"54",X"26",X"31",X"C3",X"63",X"54",X"7C",X"FE",X"28",
		X"DA",X"68",X"54",X"25",X"25",X"C3",X"0E",X"54",X"21",X"14",X"27",X"C3",X"0E",X"54",X"7C",X"FE",
		X"28",X"DA",X"7D",X"54",X"C3",X"63",X"54",X"21",X"12",X"3B",X"C3",X"0E",X"54",X"21",X"14",X"3B",
		X"C3",X"0E",X"54",X"01",X"FF",X"20",X"CD",X"DA",X"53",X"3A",X"90",X"21",X"FE",X"03",X"D2",X"17",
		X"55",X"3A",X"92",X"21",X"FE",X"14",X"CA",X"B1",X"54",X"FE",X"12",X"CA",X"BA",X"54",X"3A",X"93",
		X"21",X"FE",X"30",X"D2",X"C2",X"54",X"CD",X"F5",X"54",X"C6",X"16",X"CD",X"FC",X"54",X"C3",X"68",
		X"53",X"CD",X"F5",X"54",X"CD",X"FC",X"54",X"C3",X"68",X"53",X"CD",X"F5",X"54",X"C6",X"0B",X"C3",
		X"B4",X"54",X"FE",X"33",X"D2",X"32",X"55",X"3A",X"90",X"21",X"A7",X"CA",X"E8",X"54",X"2A",X"94",
		X"21",X"25",X"22",X"94",X"21",X"3E",X"1B",X"CD",X"F2",X"02",X"21",X"90",X"21",X"35",X"21",X"88",
		X"21",X"3A",X"90",X"21",X"85",X"6F",X"36",X"1B",X"CD",X"EE",X"54",X"C3",X"68",X"53",X"21",X"00",
		X"00",X"22",X"84",X"21",X"C9",X"3A",X"93",X"21",X"D6",X"27",X"0F",X"C9",X"21",X"88",X"21",X"F5",
		X"3A",X"90",X"21",X"85",X"6F",X"F1",X"77",X"2A",X"94",X"21",X"CD",X"F2",X"02",X"22",X"94",X"21",
		X"21",X"90",X"21",X"34",X"C3",X"EE",X"54",X"3A",X"92",X"21",X"FE",X"10",X"C2",X"32",X"55",X"3A",
		X"93",X"21",X"FE",X"30",X"D2",X"2A",X"55",X"C3",X"32",X"55",X"FE",X"34",X"D2",X"32",X"55",X"C3",
		X"C7",X"54",X"AF",X"32",X"91",X"21",X"21",X"65",X"22",X"3A",X"98",X"21",X"3D",X"4F",X"81",X"81",
		X"4F",X"06",X"00",X"09",X"11",X"88",X"21",X"06",X"03",X"CD",X"BB",X"04",X"3A",X"98",X"21",X"FE",
		X"10",X"CA",X"6F",X"55",X"E5",X"21",X"65",X"21",X"3D",X"4F",X"81",X"81",X"4F",X"06",X"00",X"09",
		X"EB",X"E1",X"7E",X"FE",X"FF",X"CA",X"6F",X"55",X"1A",X"77",X"23",X"13",X"C3",X"62",X"55",X"21",
		X"65",X"21",X"11",X"65",X"22",X"06",X"1F",X"C3",X"BB",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"C7",X"01",X"2C",X"05",X"0B",X"C7",X"0B",X"30",X"04",X"11",X"D1",X"01",X"0C",X"06",X"0B",
		X"C7",X"01",X"16",X"06",X"0B",X"D5",X"01",X"02",X"06",X"14",X"C7",X"01",X"30",X"06",X"12",X"C7",
		X"01",X"30",X"06",X"10",X"C7",X"01",X"30",X"06",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"29",X"1B",X"08",X"0D",X"08",X"13",X"08",X"00",X"0B",X"1B",X"11",X"04",X"06",
		X"08",X"12",X"13",X"11",X"00",X"13",X"08",X"0E",X"0D",X"1B",X"29",X"00",X"1F",X"14",X"16",X"09",
		X"00",X"1E",X"01",X"01",X"1E",X"00",X"1F",X"15",X"15",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"15",X"15",X"11",X"00",X"1F",X"08",X"04",X"1F",X"00",X"1F",X"11",
		X"11",X"0E",X"00",X"08",X"0D",X"08",X"13",X"08",X"00",X"0B",X"1B",X"1B",X"1B",X"26",X"2A",X"2A",
		X"2A",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"00",X"00",
		X"00",X"01",X"14",X"27",X"0B",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"48",X"03",X"23",X"0E",X"00",X"11",X"51",X"22",X"E5",X"D5",X"CD",X"34",X"57",X"D1",X"E1",
		X"13",X"13",X"79",X"FE",X"0A",X"C2",X"09",X"57",X"21",X"50",X"21",X"11",X"50",X"22",X"06",X"02",
		X"CD",X"BB",X"04",X"21",X"14",X"23",X"11",X"50",X"21",X"06",X"02",X"CD",X"BB",X"04",X"C3",X"9A",
		X"04",X"00",X"00",X"00",X"0C",X"1A",X"BE",X"1B",X"2B",X"1A",X"CA",X"41",X"57",X"D0",X"C3",X"43",
		X"57",X"BE",X"D0",X"7E",X"12",X"13",X"23",X"7E",X"12",X"79",X"32",X"98",X"21",X"FE",X"0A",X"C2",
		X"63",X"57",X"21",X"50",X"21",X"11",X"50",X"22",X"06",X"14",X"CD",X"BB",X"04",X"D1",X"E1",X"E1",
		X"C3",X"85",X"57",X"21",X"50",X"21",X"CD",X"79",X"57",X"13",X"EB",X"7E",X"FE",X"FF",X"CA",X"52",
		X"57",X"1A",X"00",X"77",X"23",X"13",X"C3",X"6B",X"57",X"C5",X"3A",X"98",X"21",X"3D",X"87",X"4F",
		X"06",X"00",X"09",X"C1",X"C9",X"CD",X"00",X"53",X"C3",X"03",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
