library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_sound_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_sound_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"00",X"24",X"C3",X"72",X"00",X"FF",X"87",X"5F",X"16",X"00",X"19",X"D7",X"C9",X"FF",
		X"5E",X"23",X"56",X"23",X"EB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"D9",X"2A",X"E3",X"20",X"3A",X"00",X"30",
		X"77",X"23",X"22",X"E3",X"20",X"D9",X"08",X"FB",X"ED",X"4D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E5",X"21",X"E0",X"20",X"CB",X"C6",X"2A",X"00",X"40",X"E1",
		X"ED",X"45",X"ED",X"56",X"32",X"00",X"40",X"CD",X"2B",X"01",X"CD",X"EC",X"02",X"CD",X"99",X"00",
		X"21",X"E0",X"20",X"CB",X"4E",X"C4",X"53",X"01",X"CD",X"08",X"02",X"CD",X"B5",X"02",X"21",X"E0",
		X"20",X"CB",X"46",X"28",X"FC",X"CB",X"86",X"18",X"E1",X"2A",X"E3",X"20",X"11",X"E5",X"20",X"7B",
		X"BD",X"20",X"03",X"7A",X"BC",X"C8",X"F3",X"2A",X"E3",X"20",X"2B",X"22",X"E3",X"20",X"FB",X"7E",
		X"32",X"E1",X"20",X"E6",X"E0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",
		X"C4",X"00",X"CF",X"E9",X"05",X"01",X"D4",X"00",X"E2",X"00",X"23",X"01",X"DA",X"00",X"D9",X"00",
		X"D9",X"00",X"D9",X"00",X"21",X"E0",X"20",X"CB",X"CE",X"C9",X"01",X"05",X"00",X"21",X"6F",X"06",
		X"18",X"0E",X"3A",X"E1",X"20",X"E6",X"FF",X"FE",X"57",X"C8",X"01",X"05",X"00",X"21",X"2F",X"06",
		X"3A",X"E1",X"20",X"E6",X"1F",X"CF",X"7E",X"FE",X"FF",X"C8",X"E5",X"21",X"D3",X"05",X"CF",X"36",
		X"00",X"E1",X"09",X"18",X"F1",X"DD",X"21",X"00",X"20",X"11",X"20",X"00",X"06",X"06",X"DD",X"36",
		X"00",X"00",X"DD",X"36",X"04",X"00",X"DD",X"19",X"10",X"F4",X"F3",X"21",X"E5",X"20",X"22",X"E3",
		X"20",X"FB",X"C9",X"21",X"E0",X"20",X"CB",X"CE",X"CB",X"E6",X"C9",X"F3",X"FD",X"E1",X"21",X"00",
		X"20",X"06",X"04",X"36",X"00",X"2C",X"20",X"FB",X"24",X"10",X"F8",X"21",X"E5",X"20",X"22",X"E3",
		X"20",X"FB",X"3E",X"00",X"06",X"06",X"21",X"08",X"20",X"11",X"20",X"00",X"77",X"19",X"3C",X"10",
		X"FB",X"FD",X"E9",X"CB",X"8E",X"CB",X"66",X"21",X"2F",X"06",X"28",X"08",X"21",X"E0",X"20",X"CB",
		X"A6",X"21",X"6F",X"06",X"3A",X"E1",X"20",X"E6",X"1F",X"47",X"CF",X"7E",X"23",X"FE",X"FF",X"C8",
		X"E5",X"21",X"D3",X"05",X"CF",X"E5",X"DD",X"E1",X"E1",X"7E",X"23",X"FE",X"00",X"28",X"6A",X"DD",
		X"77",X"14",X"47",X"7E",X"23",X"DD",X"77",X"15",X"E5",X"78",X"21",X"94",X"01",X"3D",X"CF",X"11",
		X"C8",X"01",X"D5",X"E9",X"9A",X"01",X"B3",X"01",X"B3",X"01",X"DD",X"36",X"16",X"06",X"DD",X"36",
		X"17",X"00",X"DD",X"36",X"1A",X"06",X"DD",X"36",X"1B",X"00",X"DD",X"36",X"18",X"F0",X"DD",X"36",
		X"19",X"FF",X"C9",X"DD",X"36",X"16",X"10",X"DD",X"36",X"17",X"00",X"DD",X"36",X"18",X"0C",X"DD",
		X"36",X"19",X"FE",X"DD",X"36",X"1D",X"09",X"C9",X"E1",X"CD",X"D2",X"01",X"DD",X"36",X"00",X"02",
		X"18",X"23",X"D7",X"D5",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"D7",X"DD",X"75",X"12",X"DD",X"74",
		X"13",X"DD",X"73",X"10",X"DD",X"72",X"11",X"E1",X"C9",X"7E",X"23",X"DD",X"77",X"15",X"CD",X"D2",
		X"01",X"DD",X"36",X"00",X"01",X"DD",X"36",X"09",X"01",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"03",
		X"00",X"DD",X"36",X"1C",X"00",X"C3",X"6B",X"01",X"3E",X"00",X"32",X"C6",X"20",X"32",X"D6",X"20",
		X"32",X"CD",X"20",X"32",X"DD",X"20",X"3E",X"FF",X"32",X"C7",X"20",X"32",X"D7",X"20",X"FD",X"21",
		X"A0",X"20",X"06",X"06",X"C5",X"21",X"C7",X"20",X"FD",X"7E",X"08",X"FE",X"03",X"38",X"03",X"21",
		X"D7",X"20",X"FD",X"7E",X"00",X"B7",X"E5",X"28",X"64",X"CB",X"86",X"21",X"DF",X"05",X"FD",X"7E",
		X"08",X"CF",X"FD",X"7E",X"01",X"77",X"23",X"FD",X"7E",X"02",X"77",X"21",X"EB",X"05",X"FD",X"7E",
		X"08",X"CF",X"FD",X"7E",X"03",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"77",X"DD",X"21",
		X"C0",X"20",X"FD",X"7E",X"08",X"FE",X"03",X"38",X"04",X"DD",X"21",X"D0",X"20",X"CB",X"A6",X"FD",
		X"CB",X"05",X"7E",X"28",X"18",X"CB",X"E6",X"FD",X"7E",X"05",X"DD",X"77",X"0D",X"FD",X"CB",X"05",
		X"B6",X"FD",X"5E",X"06",X"FD",X"56",X"07",X"DD",X"73",X"0B",X"DD",X"72",X"0C",X"FD",X"CB",X"04",
		X"7E",X"28",X"0A",X"FD",X"7E",X"04",X"DD",X"77",X"06",X"E1",X"CB",X"9E",X"E5",X"11",X"E0",X"FF",
		X"FD",X"19",X"E1",X"C1",X"78",X"FE",X"04",X"28",X"07",X"FE",X"01",X"28",X"03",X"37",X"CB",X"16",
		X"05",X"C2",X"24",X"02",X"C9",X"DD",X"21",X"C0",X"20",X"0E",X"01",X"CD",X"C8",X"02",X"DD",X"21",
		X"D0",X"20",X"0E",X"81",X"CD",X"C8",X"02",X"C9",X"06",X"00",X"16",X"0D",X"DD",X"CB",X"0D",X"7E",
		X"28",X"08",X"DD",X"CB",X"0D",X"76",X"28",X"02",X"16",X"0F",X"78",X"ED",X"79",X"DD",X"7E",X"00",
		X"DD",X"23",X"0D",X"ED",X"79",X"0C",X"04",X"78",X"BA",X"20",X"EF",X"C9",X"06",X"06",X"DD",X"21",
		X"00",X"20",X"C5",X"DD",X"7E",X"00",X"FE",X"00",X"28",X"0C",X"FE",X"01",X"28",X"05",X"CD",X"0F",
		X"03",X"18",X"03",X"CD",X"C5",X"04",X"C1",X"11",X"20",X"00",X"DD",X"19",X"10",X"E4",X"C9",X"DD",
		X"6E",X"09",X"DD",X"66",X"0A",X"2B",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"7D",X"B4",X"CA",X"19",
		X"04",X"DD",X"CB",X"14",X"76",X"20",X"44",X"DD",X"CB",X"1C",X"46",X"20",X"63",X"DD",X"CB",X"14",
		X"66",X"28",X"1A",X"DD",X"7E",X"03",X"DD",X"86",X"18",X"38",X"07",X"DD",X"77",X"03",X"DD",X"BE",
		X"15",X"D8",X"DD",X"7E",X"15",X"DD",X"77",X"03",X"DD",X"CB",X"14",X"A6",X"C9",X"DD",X"CB",X"14",
		X"6E",X"CA",X"9D",X"03",X"DD",X"7E",X"14",X"E6",X"0F",X"FE",X"01",X"28",X"33",X"DD",X"7E",X"03",
		X"DD",X"86",X"19",X"FE",X"C0",X"20",X"32",X"3E",X"C0",X"18",X"2E",X"CD",X"EF",X"03",X"DD",X"34",
		X"1D",X"DD",X"7E",X"1D",X"FE",X"0C",X"C0",X"DD",X"7E",X"03",X"B7",X"C6",X"F0",X"FE",X"10",X"30",
		X"07",X"DD",X"36",X"03",X"00",X"C3",X"B0",X"04",X"DD",X"77",X"03",X"DD",X"36",X"1D",X"00",X"C9",
		X"DD",X"7E",X"03",X"FE",X"10",X"D8",X"DD",X"86",X"19",X"DD",X"77",X"03",X"C9",X"DD",X"7E",X"14",
		X"E6",X"0F",X"3D",X"21",X"13",X"04",X"CF",X"E9",X"DD",X"5E",X"09",X"DD",X"56",X"0A",X"DD",X"6E",
		X"16",X"DD",X"66",X"17",X"E5",X"EB",X"B7",X"ED",X"52",X"E1",X"38",X"16",X"2B",X"DD",X"75",X"16",
		X"DD",X"74",X"17",X"7D",X"B4",X"C0",X"DD",X"6E",X"1A",X"DD",X"66",X"1B",X"DD",X"75",X"16",X"DD",
		X"74",X"17",X"DD",X"CB",X"14",X"EE",X"C9",X"CD",X"EF",X"03",X"DD",X"6E",X"09",X"DD",X"66",X"0A",
		X"DD",X"5E",X"16",X"DD",X"56",X"17",X"B7",X"ED",X"52",X"D0",X"DD",X"CB",X"14",X"EE",X"C9",X"DD",
		X"7E",X"09",X"E6",X"0F",X"FE",X"01",X"C0",X"DD",X"CB",X"14",X"7E",X"20",X"0B",X"DD",X"34",X"01",
		X"DD",X"34",X"01",X"DD",X"CB",X"14",X"FE",X"C9",X"DD",X"35",X"01",X"DD",X"35",X"01",X"DD",X"CB",
		X"14",X"BE",X"C9",X"A8",X"03",X"DA",X"03",X"D7",X"03",X"DD",X"CB",X"1C",X"86",X"DD",X"6E",X"12",
		X"DD",X"66",X"13",X"7E",X"23",X"E5",X"FE",X"FF",X"28",X"44",X"FE",X"CC",X"20",X"06",X"DD",X"CB",
		X"1C",X"C6",X"18",X"26",X"47",X"E6",X"0F",X"21",X"F7",X"05",X"CF",X"CB",X"38",X"CB",X"38",X"CB",
		X"38",X"CB",X"38",X"04",X"18",X"04",X"CB",X"3C",X"CB",X"1D",X"10",X"FA",X"DD",X"75",X"01",X"DD",
		X"74",X"02",X"DD",X"CB",X"14",X"E6",X"DD",X"CB",X"14",X"AE",X"E1",X"7E",X"23",X"DD",X"75",X"12",
		X"DD",X"74",X"13",X"21",X"0F",X"06",X"CF",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"C9",X"DD",X"6E",
		X"10",X"DD",X"66",X"11",X"D7",X"7D",X"A4",X"FE",X"FF",X"28",X"21",X"FE",X"AA",X"28",X"0D",X"B4",
		X"FE",X"00",X"20",X"31",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"18",X"E8",X"DD",X"6E",X"0E",X"DD",
		X"66",X"0F",X"D7",X"EB",X"18",X"DE",X"7D",X"A4",X"FE",X"FF",X"20",X"19",X"DD",X"7E",X"14",X"E6",
		X"0F",X"FE",X"01",X"28",X"0A",X"DD",X"CB",X"14",X"F6",X"DD",X"36",X"09",X"FF",X"E1",X"C9",X"E1",
		X"DD",X"36",X"00",X"00",X"C9",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"73",X"10",X"DD",X"72",
		X"11",X"E1",X"C3",X"19",X"04",X"DD",X"35",X"09",X"28",X"39",X"DD",X"6E",X"01",X"DD",X"66",X"02",
		X"DD",X"5E",X"0B",X"DD",X"56",X"0C",X"19",X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"CB",X"05",
		X"7E",X"C0",X"DD",X"7E",X"03",X"DD",X"86",X"0D",X"DD",X"77",X"03",X"B7",X"DD",X"BE",X"15",X"D8",
		X"3E",X"80",X"DD",X"BE",X"15",X"38",X"07",X"DD",X"7E",X"15",X"DD",X"77",X"03",X"C9",X"DD",X"36",
		X"03",X"00",X"C9",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"FE",
		X"00",X"20",X"4D",X"DD",X"6E",X"10",X"DD",X"66",X"11",X"D7",X"7D",X"A4",X"FE",X"FF",X"28",X"18",
		X"7D",X"B4",X"FE",X"00",X"28",X"1B",X"FE",X"AA",X"28",X"2C",X"DD",X"75",X"12",X"DD",X"74",X"13",
		X"DD",X"73",X"10",X"DD",X"72",X"11",X"18",X"CB",X"DD",X"CB",X"04",X"BE",X"DD",X"36",X"00",X"00",
		X"C9",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"D7",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"73",
		X"10",X"DD",X"72",X"11",X"18",X"AD",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"D7",X"EB",X"18",X"E7",
		X"DD",X"77",X"09",X"DD",X"CB",X"05",X"BE",X"FD",X"CB",X"01",X"46",X"28",X"28",X"FD",X"7E",X"02",
		X"DD",X"BE",X"15",X"38",X"03",X"DD",X"7E",X"15",X"DD",X"77",X"03",X"DD",X"36",X"0D",X"00",X"FD",
		X"6E",X"03",X"FD",X"66",X"04",X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"36",X"0B",X"00",X"DD",
		X"36",X"0C",X"00",X"18",X"12",X"FD",X"7E",X"02",X"DD",X"77",X"0D",X"FD",X"6E",X"03",X"FD",X"66",
		X"04",X"DD",X"75",X"0B",X"DD",X"74",X"0C",X"DD",X"CB",X"04",X"BE",X"FD",X"CB",X"01",X"56",X"28",
		X"0A",X"FD",X"7E",X"07",X"DD",X"77",X"04",X"DD",X"CB",X"04",X"FE",X"11",X"05",X"00",X"FD",X"7E",
		X"01",X"FE",X"02",X"38",X"03",X"11",X"08",X"00",X"FD",X"E5",X"E1",X"19",X"DD",X"75",X"12",X"DD",
		X"74",X"13",X"C9",X"00",X"20",X"20",X"20",X"40",X"20",X"60",X"20",X"80",X"20",X"A0",X"20",X"C0",
		X"20",X"C2",X"20",X"C4",X"20",X"D0",X"20",X"D2",X"20",X"D4",X"20",X"C8",X"20",X"C9",X"20",X"CA",
		X"20",X"D8",X"20",X"D9",X"20",X"DA",X"20",X"EE",X"0E",X"17",X"0E",X"4D",X"0D",X"8E",X"0C",X"D9",
		X"0B",X"2F",X"0B",X"8E",X"0A",X"F7",X"09",X"67",X"09",X"E0",X"08",X"61",X"08",X"E8",X"07",X"02",
		X"00",X"04",X"00",X"08",X"00",X"0C",X"00",X"10",X"00",X"18",X"00",X"20",X"00",X"30",X"00",X"40",
		X"00",X"60",X"00",X"80",X"00",X"C0",X"00",X"50",X"00",X"68",X"00",X"28",X"00",X"00",X"01",X"23",
		X"0A",X"63",X"0A",X"48",X"0A",X"C2",X"09",X"5E",X"07",X"17",X"07",X"FE",X"07",X"D4",X"08",X"F9",
		X"08",X"11",X"09",X"51",X"08",X"5B",X"08",X"65",X"08",X"8F",X"06",X"26",X"0E",X"29",X"09",X"DD",
		X"09",X"F6",X"09",X"90",X"06",X"BB",X"06",X"E6",X"06",X"11",X"07",X"C4",X"07",X"28",X"08",X"B0",
		X"0A",X"9E",X"09",X"F7",X"0A",X"56",X"0B",X"8F",X"0B",X"A5",X"07",X"8F",X"06",X"8F",X"06",X"3D",
		X"0C",X"5D",X"0C",X"75",X"0C",X"99",X"0C",X"AA",X"0C",X"BD",X"0C",X"12",X"0D",X"3B",X"0D",X"46",
		X"0D",X"67",X"0D",X"B7",X"0D",X"D0",X"0D",X"01",X"0E",X"DC",X"0E",X"31",X"0F",X"5A",X"0F",X"FF",
		X"02",X"01",X"C0",X"96",X"06",X"FF",X"9A",X"06",X"00",X"00",X"40",X"08",X"40",X"08",X"37",X"08",
		X"40",X"06",X"3B",X"08",X"39",X"08",X"3B",X"06",X"40",X"06",X"3B",X"08",X"3B",X"08",X"37",X"08",
		X"3B",X"08",X"39",X"08",X"37",X"08",X"39",X"07",X"3B",X"04",X"FF",X"02",X"01",X"C0",X"C1",X"06",
		X"FF",X"C5",X"06",X"00",X"00",X"40",X"07",X"40",X"07",X"37",X"07",X"40",X"05",X"3B",X"07",X"39",
		X"07",X"3B",X"05",X"40",X"05",X"3B",X"07",X"3B",X"07",X"37",X"07",X"3B",X"07",X"39",X"07",X"37",
		X"07",X"39",X"07",X"3B",X"06",X"FF",X"02",X"01",X"C0",X"EC",X"06",X"FF",X"F0",X"06",X"00",X"00",
		X"40",X"06",X"40",X"06",X"37",X"06",X"40",X"04",X"3B",X"06",X"39",X"06",X"3B",X"04",X"40",X"04",
		X"3B",X"06",X"3B",X"06",X"37",X"06",X"3B",X"06",X"39",X"06",X"37",X"06",X"39",X"06",X"3B",X"04",
		X"FF",X"02",X"01",X"C0",X"EC",X"06",X"FF",X"00",X"00",X"FF",X"1D",X"07",X"FF",X"21",X"07",X"FF",
		X"FF",X"01",X"01",X"A0",X"34",X"01",X"14",X"00",X"08",X"EC",X"FF",X"1C",X"01",X"00",X"00",X"00",
		X"01",X"01",X"80",X"10",X"00",X"10",X"00",X"08",X"0A",X"00",X"1D",X"01",X"00",X"00",X"00",X"01",
		X"01",X"A0",X"32",X"01",X"14",X"00",X"08",X"EC",X"FF",X"1C",X"01",X"00",X"00",X"00",X"01",X"01",
		X"80",X"10",X"00",X"10",X"00",X"08",X"0E",X"00",X"1D",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"64",X"07",X"FF",X"68",X"07",X"FF",X"FF",X"01",X"01",X"A0",X"13",X"01",X"14",X"00",X"08",
		X"EF",X"FF",X"14",X"01",X"00",X"00",X"00",X"01",X"01",X"80",X"10",X"00",X"10",X"00",X"08",X"0A",
		X"00",X"18",X"01",X"00",X"00",X"00",X"01",X"01",X"A0",X"13",X"01",X"14",X"00",X"08",X"EF",X"FF",
		X"14",X"01",X"00",X"00",X"00",X"01",X"01",X"80",X"10",X"00",X"10",X"00",X"08",X"0A",X"00",X"18",
		X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"AB",X"07",X"FF",X"AF",X"07",X"FF",X"FF",X"01",
		X"01",X"80",X"A0",X"00",X"30",X"00",X"08",X"00",X"00",X"40",X"00",X"10",X"FF",X"FF",X"30",X"00",
		X"20",X"00",X"00",X"00",X"04",X"00",X"FF",X"CA",X"07",X"FF",X"CE",X"07",X"FF",X"FF",X"01",X"01",
		X"F0",X"FF",X"01",X"10",X"04",X"00",X"F0",X"FF",X"00",X"00",X"01",X"01",X"01",X"FE",X"60",X"00",
		X"10",X"04",X"FF",X"10",X"00",X"00",X"00",X"01",X"01",X"01",X"F0",X"60",X"01",X"20",X"04",X"00",
		X"FA",X"FF",X"00",X"00",X"01",X"40",X"04",X"FD",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"04",X"08",X"FF",X"08",X"08",X"FF",X"FF",X"01",X"01",X"DF",X"50",X"00",X"FF",X"02",X"0F",
		X"01",X"00",X"05",X"0F",X"00",X"70",X"01",X"00",X"70",X"00",X"01",X"01",X"E0",X"70",X"00",X"20",
		X"02",X"02",X"F9",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"DE",X"2E",X"08",X"FF",X"32",X"08",
		X"FF",X"FF",X"01",X"01",X"90",X"70",X"00",X"40",X"00",X"01",X"FF",X"FF",X"01",X"01",X"90",X"80",
		X"00",X"60",X"00",X"01",X"FF",X"FF",X"01",X"01",X"90",X"70",X"00",X"60",X"00",X"01",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"57",X"08",X"FF",X"6F",X"08",X"FF",X"FF",X"00",X"00",X"FF",X"61",X"08",
		X"FF",X"92",X"08",X"FF",X"FF",X"00",X"00",X"FF",X"6B",X"08",X"FF",X"B5",X"08",X"FF",X"FF",X"01",
		X"01",X"F0",X"30",X"01",X"10",X"00",X"00",X"F2",X"FF",X"10",X"01",X"00",X"00",X"00",X"01",X"01",
		X"B0",X"90",X"01",X"18",X"00",X"02",X"E3",X"FF",X"08",X"00",X"F0",X"2A",X"00",X"18",X"01",X"00",
		X"00",X"00",X"01",X"01",X"F0",X"1C",X"01",X"10",X"00",X"00",X"F2",X"FF",X"10",X"01",X"00",X"00",
		X"00",X"01",X"01",X"B0",X"80",X"01",X"18",X"00",X"02",X"E3",X"FF",X"08",X"00",X"F0",X"2A",X"00",
		X"18",X"01",X"00",X"00",X"00",X"01",X"01",X"F0",X"00",X"01",X"10",X"00",X"00",X"F2",X"FF",X"10",
		X"01",X"00",X"00",X"00",X"01",X"01",X"B0",X"70",X"01",X"18",X"00",X"02",X"E3",X"FF",X"08",X"00",
		X"F0",X"2A",X"00",X"00",X"00",X"00",X"FF",X"17",X"09",X"FF",X"DE",X"08",X"FF",X"FF",X"01",X"01",
		X"FE",X"10",X"03",X"10",X"02",X"00",X"E0",X"FF",X"60",X"00",X"00",X"01",X"01",X"FE",X"10",X"00",
		X"90",X"02",X"00",X"01",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"17",X"09",X"FF",X"03",
		X"09",X"FF",X"FF",X"01",X"01",X"FE",X"10",X"00",X"C8",X"02",X"00",X"02",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"17",X"09",X"FF",X"1B",X"09",X"FF",X"FF",X"01",X"01",X"FE",X"10",X"00",
		X"A0",X"02",X"00",X"03",X"00",X"60",X"00",X"00",X"00",X"01",X"01",X"E0",X"34",X"09",X"03",X"01",
		X"D0",X"38",X"09",X"FF",X"3C",X"09",X"FF",X"FF",X"6D",X"09",X"FF",X"FF",X"39",X"04",X"40",X"04",
		X"39",X"04",X"40",X"04",X"39",X"04",X"40",X"04",X"39",X"04",X"40",X"04",X"39",X"04",X"40",X"04",
		X"39",X"04",X"40",X"04",X"39",X"06",X"40",X"06",X"40",X"06",X"40",X"06",X"34",X"06",X"42",X"06",
		X"42",X"06",X"42",X"06",X"37",X"06",X"44",X"06",X"44",X"06",X"44",X"0F",X"FF",X"40",X"04",X"44",
		X"04",X"40",X"04",X"44",X"04",X"40",X"04",X"44",X"04",X"40",X"04",X"44",X"04",X"40",X"04",X"44",
		X"04",X"40",X"04",X"44",X"04",X"37",X"06",X"40",X"06",X"40",X"06",X"40",X"06",X"3B",X"06",X"44",
		X"06",X"44",X"06",X"44",X"06",X"42",X"06",X"47",X"06",X"47",X"06",X"47",X"0F",X"FF",X"03",X"01",
		X"E0",X"A4",X"09",X"FF",X"AC",X"09",X"AC",X"09",X"B7",X"09",X"FF",X"FF",X"50",X"03",X"52",X"03",
		X"54",X"03",X"55",X"03",X"57",X"08",X"FF",X"50",X"03",X"52",X"03",X"54",X"03",X"55",X"03",X"57",
		X"0F",X"FF",X"03",X"01",X"F0",X"C8",X"09",X"FF",X"CC",X"09",X"FF",X"FF",X"44",X"04",X"42",X"04",
		X"44",X"04",X"47",X"07",X"47",X"04",X"45",X"04",X"47",X"04",X"50",X"0F",X"FF",X"00",X"01",X"C0",
		X"E8",X"09",X"01",X"01",X"C0",X"EC",X"09",X"FF",X"F0",X"09",X"FF",X"FF",X"F3",X"09",X"FF",X"FF",
		X"47",X"0F",X"FF",X"44",X"0F",X"FF",X"03",X"01",X"D0",X"01",X"0A",X"01",X"01",X"D0",X"05",X"0A",
		X"FF",X"0B",X"0A",X"FF",X"FF",X"20",X"0A",X"0B",X"0A",X"FF",X"FF",X"47",X"0A",X"45",X"06",X"46",
		X"06",X"47",X"08",X"3A",X"06",X"3B",X"06",X"40",X"08",X"35",X"06",X"33",X"06",X"30",X"0F",X"FF",
		X"CC",X"03",X"FF",X"04",X"01",X"E0",X"2E",X"0A",X"05",X"01",X"E0",X"32",X"0A",X"FF",X"36",X"0A",
		X"FF",X"FF",X"3F",X"0A",X"FF",X"FF",X"44",X"04",X"42",X"04",X"44",X"04",X"47",X"0A",X"FF",X"47",
		X"04",X"45",X"04",X"47",X"04",X"50",X"0A",X"FF",X"01",X"01",X"D0",X"4E",X"0A",X"FF",X"52",X"0A",
		X"FF",X"FF",X"40",X"06",X"3B",X"06",X"39",X"06",X"3B",X"06",X"42",X"08",X"40",X"06",X"40",X"06",
		X"44",X"0F",X"FF",X"05",X"01",X"E0",X"6E",X"0A",X"02",X"01",X"D0",X"72",X"0A",X"FF",X"76",X"0A",
		X"FF",X"FF",X"93",X"0A",X"FF",X"FF",X"47",X"08",X"47",X"08",X"44",X"06",X"40",X"06",X"44",X"06",
		X"47",X"06",X"47",X"08",X"47",X"08",X"44",X"06",X"40",X"06",X"44",X"06",X"47",X"06",X"44",X"06",
		X"47",X"0F",X"FF",X"40",X"08",X"40",X"08",X"44",X"06",X"47",X"06",X"44",X"06",X"40",X"06",X"40",
		X"08",X"40",X"08",X"44",X"06",X"47",X"06",X"44",X"06",X"40",X"06",X"44",X"06",X"40",X"0F",X"FF",
		X"01",X"00",X"DF",X"B6",X"0A",X"FF",X"BA",X"0A",X"00",X"00",X"01",X"01",X"A0",X"A0",X"00",X"0C",
		X"00",X"04",X"00",X"00",X"0C",X"00",X"01",X"01",X"00",X"01",X"01",X"A0",X"90",X"00",X"0C",X"00",
		X"04",X"00",X"00",X"0C",X"00",X"01",X"01",X"00",X"01",X"01",X"DD",X"A0",X"00",X"0C",X"00",X"FF",
		X"00",X"00",X"0C",X"00",X"FF",X"FE",X"FF",X"01",X"01",X"DD",X"90",X"00",X"0C",X"00",X"FE",X"00",
		X"00",X"0C",X"00",X"FF",X"FE",X"FF",X"00",X"05",X"00",X"EF",X"FD",X"0A",X"FF",X"27",X"0B",X"45",
		X"0B",X"2D",X"0B",X"50",X"0B",X"33",X"0B",X"45",X"0B",X"39",X"0B",X"50",X"0B",X"3F",X"0B",X"45",
		X"0B",X"3F",X"0B",X"50",X"0B",X"39",X"0B",X"45",X"0B",X"33",X"0B",X"50",X"0B",X"2D",X"0B",X"45",
		X"0B",X"27",X"0B",X"50",X"0B",X"00",X"00",X"01",X"01",X"AA",X"8C",X"00",X"00",X"01",X"01",X"BB",
		X"70",X"00",X"00",X"01",X"01",X"AA",X"76",X"00",X"00",X"01",X"01",X"BB",X"60",X"00",X"00",X"01",
		X"01",X"AA",X"50",X"00",X"00",X"10",X"00",X"03",X"FF",X"FF",X"10",X"01",X"00",X"00",X"00",X"00",
		X"10",X"00",X"FE",X"FE",X"FF",X"00",X"05",X"01",X"E0",X"61",X"0B",X"04",X"01",X"D0",X"65",X"0B",
		X"FF",X"69",X"0B",X"FF",X"FF",X"7C",X"0B",X"FF",X"FF",X"47",X"03",X"45",X"02",X"47",X"03",X"44",
		X"02",X"47",X"03",X"45",X"02",X"47",X"03",X"49",X"02",X"50",X"0F",X"FF",X"44",X"03",X"42",X"02",
		X"44",X"03",X"40",X"02",X"44",X"03",X"42",X"02",X"44",X"03",X"47",X"02",X"49",X"0F",X"FF",X"00",
		X"01",X"C0",X"A4",X"0B",X"01",X"01",X"C0",X"A8",X"0B",X"02",X"01",X"C0",X"AC",X"0B",X"03",X"01",
		X"C0",X"B2",X"0B",X"FF",X"B8",X"0B",X"00",X"00",X"09",X"0C",X"00",X"00",X"3A",X"0C",X"B8",X"0B",
		X"AA",X"AA",X"3A",X"0C",X"09",X"0C",X"AA",X"AA",X"52",X"07",X"4B",X"05",X"47",X"09",X"4B",X"07",
		X"52",X"07",X"4B",X"07",X"47",X"05",X"44",X"09",X"47",X"07",X"4B",X"07",X"47",X"07",X"44",X"05",
		X"40",X"09",X"44",X"07",X"47",X"07",X"49",X"07",X"46",X"05",X"42",X"09",X"46",X"07",X"49",X"07",
		X"52",X"07",X"4B",X"05",X"47",X"09",X"4B",X"07",X"52",X"07",X"56",X"07",X"52",X"05",X"4B",X"09",
		X"52",X"07",X"56",X"07",X"57",X"07",X"54",X"05",X"50",X"09",X"54",X"07",X"57",X"07",X"59",X"07",
		X"56",X"05",X"52",X"09",X"56",X"07",X"59",X"07",X"FF",X"37",X"08",X"3B",X"09",X"42",X"09",X"34",
		X"08",X"37",X"09",X"3B",X"09",X"30",X"08",X"34",X"09",X"37",X"09",X"32",X"08",X"36",X"09",X"39",
		X"09",X"37",X"08",X"3B",X"09",X"42",X"09",X"3B",X"08",X"42",X"09",X"46",X"09",X"40",X"08",X"44",
		X"09",X"47",X"09",X"42",X"08",X"46",X"09",X"49",X"09",X"FF",X"CC",X"04",X"FF",X"00",X"01",X"C0",
		X"48",X"0C",X"FF",X"01",X"C0",X"48",X"0C",X"FF",X"4C",X"0C",X"00",X"00",X"47",X"05",X"44",X"05",
		X"47",X"05",X"44",X"05",X"45",X"05",X"42",X"05",X"45",X"05",X"42",X"05",X"FF",X"01",X"00",X"FF",
		X"63",X"0C",X"FF",X"67",X"0C",X"FF",X"FF",X"01",X"01",X"FD",X"00",X"03",X"20",X"04",X"00",X"E6",
		X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"7B",X"0C",X"FF",X"7F",X"0C",X"FF",X"FF",X"01",
		X"01",X"DA",X"80",X"00",X"14",X"00",X"01",X"02",X"00",X"10",X"01",X"00",X"A0",X"00",X"01",X"01",
		X"D0",X"A0",X"00",X"1A",X"00",X"01",X"FB",X"FF",X"00",X"02",X"01",X"E0",X"9F",X"0C",X"FF",X"A3",
		X"0C",X"FF",X"FF",X"54",X"02",X"50",X"02",X"57",X"02",X"FF",X"01",X"01",X"FF",X"B0",X"0C",X"FF",
		X"B4",X"0C",X"FF",X"FF",X"24",X"01",X"23",X"03",X"27",X"02",X"29",X"0F",X"FF",X"00",X"01",X"C0",
		X"C3",X"0C",X"FF",X"C7",X"0C",X"00",X"00",X"46",X"07",X"46",X"07",X"45",X"07",X"46",X"07",X"47",
		X"07",X"47",X"07",X"46",X"07",X"47",X"07",X"CC",X"07",X"49",X"07",X"49",X"07",X"49",X"07",X"46",
		X"07",X"46",X"07",X"48",X"07",X"4A",X"07",X"4B",X"09",X"4B",X"07",X"4B",X"07",X"49",X"07",X"49",
		X"07",X"4B",X"07",X"49",X"07",X"4B",X"09",X"4B",X"07",X"4B",X"07",X"49",X"07",X"49",X"07",X"4B",
		X"07",X"49",X"07",X"4A",X"09",X"4A",X"07",X"4A",X"07",X"4B",X"07",X"4B",X"07",X"4B",X"07",X"4B",
		X"07",X"FF",X"02",X"00",X"FF",X"18",X"0D",X"FF",X"1C",X"0D",X"FF",X"FF",X"01",X"01",X"F0",X"80",
		X"02",X"20",X"00",X"00",X"05",X"00",X"20",X"00",X"00",X"F8",X"FF",X"8C",X"01",X"00",X"00",X"00",
		X"01",X"01",X"FE",X"80",X"01",X"20",X"00",X"FE",X"F0",X"FF",X"00",X"04",X"01",X"C0",X"48",X"0C",
		X"FF",X"01",X"C0",X"48",X"0C",X"FF",X"01",X"00",X"FF",X"51",X"0D",X"05",X"00",X"FF",X"55",X"0D",
		X"FF",X"59",X"0D",X"FF",X"FF",X"59",X"0D",X"FF",X"FF",X"01",X"01",X"F6",X"07",X"00",X"18",X"04",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"00",X"FF",X"6D",X"0D",X"FF",X"7F",X"0D",X"9D",
		X"0D",X"85",X"0D",X"9D",X"0D",X"8B",X"0D",X"9D",X"0D",X"91",X"0D",X"9D",X"0D",X"FF",X"FF",X"01",
		X"01",X"F0",X"80",X"02",X"00",X"01",X"01",X"F0",X"60",X"02",X"00",X"01",X"01",X"F0",X"40",X"02",
		X"00",X"01",X"01",X"F0",X"20",X"02",X"00",X"01",X"01",X"F0",X"00",X"02",X"00",X"20",X"00",X"00",
		X"05",X"00",X"20",X"00",X"00",X"F8",X"FF",X"10",X"01",X"00",X"00",X"00",X"01",X"01",X"F0",X"80",
		X"01",X"20",X"00",X"FD",X"F0",X"FF",X"00",X"02",X"01",X"EF",X"BD",X"0D",X"FF",X"C1",X"0D",X"FF",
		X"FF",X"4B",X"01",X"47",X"01",X"44",X"01",X"40",X"01",X"44",X"01",X"47",X"01",X"49",X"01",X"FF",
		X"00",X"01",X"C0",X"D6",X"0D",X"FF",X"DA",X"0D",X"00",X"00",X"47",X"09",X"49",X"07",X"50",X"07",
		X"52",X"09",X"52",X"07",X"54",X"07",X"49",X"09",X"50",X"07",X"52",X"07",X"55",X"09",X"55",X"07",
		X"52",X"07",X"47",X"07",X"48",X"07",X"49",X"07",X"4B",X"07",X"50",X"09",X"50",X"07",X"49",X"07",
		X"FF",X"00",X"01",X"F0",X"0C",X"0E",X"05",X"03",X"B0",X"10",X"0E",X"FF",X"14",X"0E",X"FF",X"FF",
		X"25",X"0E",X"FF",X"FF",X"45",X"08",X"45",X"06",X"4A",X"09",X"51",X"06",X"51",X"06",X"51",X"06",
		X"4A",X"06",X"48",X"0F",X"FF",X"FF",X"00",X"00",X"FF",X"40",X"0E",X"01",X"00",X"FF",X"40",X"0E",
		X"02",X"00",X"FF",X"40",X"0E",X"03",X"00",X"FF",X"40",X"0E",X"04",X"00",X"FF",X"40",X"0E",X"FF",
		X"20",X"01",X"F0",X"7E",X"00",X"28",X"00",X"FE",X"00",X"00",X"12",X"01",X"F0",X"7E",X"00",X"06",
		X"00",X"F0",X"00",X"00",X"40",X"01",X"F0",X"7E",X"00",X"20",X"00",X"FF",X"00",X"00",X"30",X"01",
		X"F0",X"8E",X"00",X"00",X"20",X"01",X"F0",X"65",X"01",X"28",X"00",X"FE",X"00",X"00",X"18",X"01",
		X"F0",X"65",X"01",X"30",X"01",X"F0",X"2C",X"01",X"00",X"20",X"01",X"F0",X"FD",X"00",X"28",X"00",
		X"FE",X"00",X"00",X"12",X"01",X"F0",X"FD",X"00",X"06",X"00",X"F0",X"00",X"00",X"40",X"01",X"F0",
		X"FD",X"00",X"20",X"00",X"FF",X"00",X"00",X"30",X"01",X"F0",X"1C",X"01",X"00",X"20",X"01",X"F0",
		X"59",X"00",X"28",X"00",X"FE",X"00",X"00",X"18",X"01",X"F0",X"59",X"00",X"30",X"01",X"F0",X"4B",
		X"00",X"00",X"20",X"01",X"F0",X"3F",X"00",X"28",X"00",X"FE",X"00",X"00",X"12",X"01",X"F0",X"3F",
		X"00",X"06",X"00",X"F0",X"00",X"00",X"40",X"01",X"F0",X"3F",X"00",X"20",X"00",X"FF",X"00",X"00",
		X"30",X"01",X"F0",X"47",X"00",X"00",X"18",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"B0",X"E7",
		X"0E",X"FF",X"01",X"D0",X"EB",X"0E",X"FF",X"10",X"0F",X"00",X"00",X"10",X"0F",X"00",X"00",X"44",
		X"09",X"42",X"05",X"40",X"05",X"39",X"07",X"35",X"07",X"39",X"07",X"40",X"07",X"44",X"07",X"42",
		X"07",X"40",X"05",X"3B",X"05",X"37",X"07",X"34",X"07",X"37",X"07",X"3B",X"07",X"42",X"07",X"FF",
		X"52",X"09",X"50",X"05",X"4B",X"05",X"47",X"07",X"44",X"07",X"47",X"07",X"4B",X"07",X"52",X"07",
		X"50",X"09",X"4B",X"05",X"49",X"05",X"45",X"07",X"42",X"07",X"45",X"07",X"49",X"07",X"50",X"07",
		X"FF",X"01",X"00",X"FF",X"41",X"0F",X"00",X"01",X"B0",X"D6",X"0D",X"02",X"03",X"90",X"D6",X"0D",
		X"FF",X"45",X"0F",X"FF",X"FF",X"01",X"01",X"00",X"F6",X"01",X"50",X"00",X"24",X"00",X"00",X"30",
		X"00",X"18",X"01",X"00",X"20",X"00",X"10",X"01",X"00",X"00",X"02",X"00",X"FF",X"60",X"0F",X"FF",
		X"64",X"0F",X"FF",X"FF",X"01",X"01",X"00",X"10",X"00",X"50",X"04",X"03",X"01",X"00",X"00",X"00",
		X"00",X"30",X"04",X"00",X"01",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"01",X"00",X"00",X"00",
		X"00",X"40",X"04",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
