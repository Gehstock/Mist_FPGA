`define BUILD_DATE "210524"
`define BUILD_TIME "140250"
