library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg3_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg3_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"DC",X"EE",X"DC",X"FF",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"FF",X"FF",X"CC",X"CC",X"ED",X"DD",X"EE",X"EE",X"EF",X"CC",X"EE",X"CC",X"EE",X"EE",X"EE",X"EE",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",
		X"00",X"00",X"FF",X"00",X"CC",X"00",X"DC",X"FF",X"EE",X"CC",X"FF",X"CC",X"DC",X"DE",X"DC",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"00",X"CC",X"FF",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"EE",X"CC",X"FF",X"DC",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"FF",X"DC",X"FF",
		X"EE",X"FF",X"EE",X"CC",X"EE",X"DD",X"EE",X"EE",X"EE",X"FF",X"EE",X"CC",X"FF",X"DD",X"FF",X"EE",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"FF",X"DC",X"FF",X"11",X"11",X"44",X"44",
		X"FF",X"CC",X"DC",X"DD",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"23",X"33",X"32",X"33",X"33",X"32",X"33",X"23",X"33",X"23",X"33",X"32",X"32",X"33",X"23",X"33",
		X"EE",X"DD",X"CC",X"DE",X"DF",X"DE",X"FC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"11",X"11",X"77",X"77",X"99",X"99",X"11",X"11",X"16",X"66",X"16",X"AB",X"16",X"5A",X"17",X"AB",
		X"11",X"11",X"77",X"77",X"99",X"99",X"11",X"11",X"66",X"66",X"6B",X"AB",X"6A",X"BA",X"7B",X"AB",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"EF",X"18",X"EF",X"18",X"EF",X"17",X"EF",X"17",X"EF",X"1D",X"EE",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"EF",X"86",X"EF",X"8A",X"EF",X"7B",X"EF",X"7A",X"EF",X"7D",X"EE",
		X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",
		X"99",X"89",X"99",X"89",X"99",X"89",X"99",X"89",X"99",X"89",X"99",X"89",X"99",X"89",X"99",X"89",
		X"88",X"88",X"99",X"99",X"74",X"74",X"88",X"88",X"77",X"77",X"88",X"88",X"99",X"99",X"88",X"88",
		X"88",X"88",X"99",X"99",X"74",X"70",X"88",X"88",X"77",X"77",X"88",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"88",X"77",X"FF",X"77",X"CC",X"78",X"CC",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"88",X"88",X"77",X"77",X"99",X"99",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CD",X"CC",X"DD",
		X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"DD",X"DF",X"EF",X"F1",X"11",X"F1",X"DD",X"1D",X"CC",
		X"CC",X"FF",X"DD",X"11",X"FF",X"DD",X"11",X"CC",X"DD",X"EC",X"CC",X"1F",X"CC",X"C1",X"CC",X"CC",
		X"DD",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"1D",X"CC",X"1D",X"CC",
		X"11",X"11",X"BB",X"BB",X"22",X"22",X"00",X"64",X"11",X"11",X"BB",X"BB",X"22",X"22",X"00",X"64",
		X"11",X"11",X"BB",X"BB",X"22",X"22",X"12",X"63",X"11",X"11",X"BB",X"BB",X"22",X"22",X"12",X"63",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"33",X"00",X"70",X"00",
		X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",X"33",X"30",X"77",X"77",
		X"97",X"97",X"17",X"17",X"77",X"77",X"97",X"97",X"17",X"17",X"77",X"77",X"79",X"99",X"79",X"11",
		X"79",X"11",X"79",X"11",X"79",X"11",X"79",X"11",X"79",X"11",X"79",X"11",X"79",X"99",X"77",X"77",
		X"00",X"00",X"FF",X"00",X"CC",X"00",X"CC",X"FF",X"EE",X"CC",X"FE",X"CC",X"DC",X"DE",X"DC",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"F0",X"CC",X"CF",X"EE",X"CC",
		X"CC",X"FF",X"CC",X"CC",X"EE",X"CC",X"DC",X"DE",X"DC",X"FF",X"DC",X"FF",X"11",X"11",X"88",X"88",
		X"00",X"FF",X"F0",X"CE",X"CF",X"E0",X"CC",X"00",X"EC",X"E0",X"FE",X"CC",X"11",X"1E",X"88",X"00",
		X"77",X"77",X"91",X"91",X"77",X"77",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"11",X"11",X"77",X"77",X"88",X"80",X"88",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"77",X"CC",X"F7",X"CC",X"FF",X"CC",X"CF",X"FF",X"CC",X"EF",X"EC",X"FE",X"CD",X"FF",X"DE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"F7",X"77",X"FF",X"77",X"CF",X"77",X"CC",X"F7",
		X"99",X"EF",X"77",X"F9",X"11",X"99",X"FF",X"78",X"EE",X"17",X"EE",X"11",X"EE",X"FF",X"EE",X"EE",
		X"EC",X"FF",X"CD",X"CF",X"DE",X"CC",X"EF",X"EC",X"F9",X"CD",X"99",X"DE",X"78",X"EF",X"17",X"F9",
		X"97",X"97",X"17",X"17",X"87",X"87",X"97",X"97",X"17",X"17",X"87",X"87",X"97",X"97",X"17",X"17",
		X"77",X"77",X"17",X"77",X"11",X"77",X"99",X"77",X"17",X"17",X"87",X"11",X"97",X"91",X"17",X"17",
		X"87",X"87",X"97",X"97",X"17",X"17",X"87",X"87",X"97",X"97",X"17",X"17",X"87",X"DE",X"88",X"DE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"F7",X"77",X"CF",X"77",X"CC",X"77",X"EC",X"F7",X"CF",X"CF",
		X"DE",X"CC",X"EF",X"EC",X"F9",X"CD",X"99",X"DE",X"78",X"EF",X"17",X"F9",X"71",X"99",X"77",X"78",
		X"FF",X"FF",X"FC",X"CC",X"CF",X"CD",X"CC",X"DE",X"EC",X"FE",X"CD",X"CF",X"DE",X"CC",X"EF",X"EC",
		X"77",X"17",X"77",X"71",X"77",X"77",X"17",X"77",X"71",X"7D",X"79",X"77",X"79",X"DE",X"79",X"DE",
		X"F9",X"CD",X"99",X"DE",X"78",X"EF",X"17",X"F9",X"71",X"99",X"77",X"78",X"77",X"DE",X"77",X"DE",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"CD",X"EE",X"DE",X"FF",X"DE",X"DC",X"DE",X"DC",X"DE",X"FC",X"DE",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"CD",X"EE",X"DE",X"FF",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"CF",X"DE",X"CC",X"DE",X"CC",X"FF",X"FD",X"CC",X"EF",X"CC",X"F1",X"EE",X"99",X"CE",X"87",X"CE",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"FC",X"DE",X"CF",X"DE",X"CC",X"FE",X"EC",X"CF",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"DE",X"CC",X"E1",
		X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"ED",X"CC",X"ED",X"CC",
		X"CC",X"1D",X"CD",X"CC",X"DE",X"CC",X"E1",X"CC",X"1D",X"CC",X"DD",X"CC",X"DC",X"CC",X"CC",X"CC",
		X"EE",X"CC",X"1E",X"CC",X"1E",X"DD",X"D1",X"FF",X"DD",X"11",X"CD",X"DD",X"CD",X"DC",X"CD",X"DC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"CC",X"CD",X"DC",X"CD",X"DD",X"DE",X"FF",
		X"CD",X"DD",X"FF",X"FF",X"11",X"11",X"DD",X"DD",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"E1",X"11",X"1D",X"DD",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",
		X"CC",X"11",X"CC",X"C1",X"CC",X"C1",X"CC",X"DD",X"CC",X"DD",X"DD",X"DE",X"EE",X"EE",X"11",X"11",
		X"CC",X"CC",X"CC",X"CD",X"CC",X"D1",X"CC",X"D1",X"CD",X"D1",X"DD",X"E1",X"EE",X"E1",X"11",X"11",
		X"DC",X"DE",X"FF",X"DE",X"CC",X"DE",X"CC",X"FF",X"EE",X"CC",X"FE",X"CC",X"DC",X"DE",X"DC",X"DE",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"FF",X"DE",X"CC",X"FE",X"CC",X"CF",X"EE",X"CC",
		X"88",X"EE",X"88",X"DE",X"88",X"9D",X"88",X"88",X"88",X"88",X"81",X"11",X"17",X"17",X"17",X"17",
		X"71",X"87",X"77",X"98",X"77",X"19",X"77",X"71",X"77",X"77",X"97",X"77",X"11",X"77",X"17",X"77",
		X"87",X"87",X"97",X"97",X"17",X"17",X"17",X"17",X"87",X"87",X"17",X"97",X"17",X"DE",X"88",X"DE",
		X"87",X"17",X"97",X"91",X"17",X"17",X"17",X"17",X"87",X"87",X"97",X"97",X"17",X"DE",X"88",X"DE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"91",X"77",X"99",X"77",X"99",X"77",X"99",
		X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"11",X"11",X"11",X"11",X"18",X"AA",X"B8",X"11",X"18",
		X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"92",X"77",X"77",
		X"11",X"18",X"11",X"18",X"BB",X"B8",X"11",X"18",X"11",X"18",X"22",X"28",X"22",X"22",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"91",X"77",X"99",X"77",X"99",X"77",X"99",
		X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",
		X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"92",X"77",X"77",
		X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"22",X"77",X"22",X"77",X"77",X"77",
		X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"ED",X"FF",X"ED",X"FF",X"11",X"11",X"88",X"88",
		X"ED",X"CC",X"ED",X"CC",X"ED",X"DE",X"ED",X"DE",X"ED",X"FF",X"ED",X"FF",X"11",X"11",X"88",X"88",
		X"00",X"FF",X"FF",X"CC",X"CC",X"EE",X"CC",X"00",X"FF",X"CC",X"EF",X"FF",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"B3",X"BB",X"B3",X"BB",X"33",X"00",X"33",X"00",X"FF",X"00",X"EE",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"66",X"44",X"FF",X"77",X"CC",X"11",X"CC",
		X"77",X"77",X"77",X"77",X"77",X"77",X"F8",X"77",X"CF",X"66",X"CC",X"44",X"EC",X"F7",X"CF",X"CF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"27",X"77",X"27",X"77",X"27",X"77",X"27",X"77",X"27",X"77",X"27",X"77",X"27",X"77",X"27",X"77",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CD",X"CC",X"CD",X"CC",X"DE",X"CC",X"E1",X"DD",X"E1",
		X"1D",X"CC",X"1D",X"CC",X"DD",X"CC",X"DD",X"CC",X"DC",X"CC",X"CC",X"CC",X"DC",X"CC",X"ED",X"CC",
		X"FF",X"1D",X"11",X"ED",X"DD",X"1E",X"CC",X"C1",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"1E",X"CC",X"11",X"DD",X"D1",X"FF",X"FF",X"11",X"11",X"1D",X"CD",X"DD",X"1D",X"DC",X"C1",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"D1",X"DC",X"D1",X"ED",X"D1",X"ED",X"D1",X"1E",X"D1",X"D1",X"D1",X"D1",X"D1",X"DD",X"D1",X"FF",
		X"CC",X"CC",X"DD",X"DD",X"FF",X"FF",X"11",X"11",X"DD",X"DD",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"E1",X"11",X"11",X"DD",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"FF",X"CC",X"CC",X"CE",X"CC",X"DE",X"EE",X"DE",
		X"FF",X"CC",X"CC",X"CE",X"CC",X"DE",X"EE",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"33",X"11",X"11",X"11",X"55",X"55",X"66",X"66",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"11",X"55",X"55",X"66",X"66",
		X"77",X"77",X"91",X"91",X"77",X"77",X"98",X"98",X"98",X"98",X"99",X"99",X"89",X"89",X"88",X"88",
		X"99",X"99",X"99",X"99",X"99",X"19",X"99",X"19",X"88",X"18",X"88",X"18",X"77",X"17",X"77",X"97",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",X"FE",X"EF",X"FF",X"11",X"11",X"88",X"88",
		X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"FE",X"EF",X"FF",X"11",X"11",X"88",X"88",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DF",X"DC",X"FC",X"DF",X"CC",
		X"DC",X"DF",X"DC",X"FF",X"DC",X"CC",X"DF",X"CE",X"FC",X"EF",X"CC",X"F1",X"CE",X"DE",X"ED",X"CD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"CC",X"FC",X"CC",X"CC",X"DE",X"CE",X"DE",X"EE",X"DE",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"DE",X"DC",X"FF",X"FF",X"CC",X"CC",X"CC",
		X"DC",X"DE",X"DC",X"DE",X"DC",X"FF",X"DF",X"CC",X"FC",X"CC",X"CC",X"DE",X"CE",X"DE",X"EE",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"29",X"00",X"9A",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"28",X"02",X"A0",X"08",X"00",X"89",X"A0",X"AA",X"A2",X"A9",X"29",X"22",X"7A",X"99",X"A9",
		X"00",X"00",X"00",X"22",X"00",X"99",X"28",X"71",X"99",X"99",X"10",X"00",X"00",X"07",X"09",X"99",
		X"0A",X"99",X"AA",X"99",X"29",X"99",X"87",X"99",X"98",X"AA",X"99",X"77",X"99",X"A8",X"88",X"07",
		X"77",X"77",X"18",X"18",X"77",X"77",X"74",X"44",X"78",X"88",X"11",X"18",X"11",X"11",X"11",X"11",
		X"81",X"FE",X"74",X"FF",X"17",X"1F",X"71",X"81",X"87",X"78",X"88",X"74",X"88",X"17",X"11",X"71",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"77",X"77",X"77",X"77",
		X"11",X"87",X"91",X"88",X"99",X"18",X"99",X"91",X"99",X"99",X"88",X"99",X"88",X"88",X"77",X"88",
		X"44",X"44",X"47",X"77",X"47",X"11",X"47",X"99",X"47",X"79",X"47",X"99",X"47",X"66",X"47",X"67",
		X"44",X"44",X"77",X"77",X"11",X"11",X"66",X"66",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"66",X"66",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"99",X"91",X"66",X"91",X"76",X"91",X"77",X"91",X"77",X"91",
		X"11",X"11",X"91",X"11",X"99",X"11",X"99",X"11",X"99",X"11",X"99",X"11",X"99",X"22",X"92",X"22",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"0D",X"DD",X"DD",X"CC",X"0F",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"0D",X"EE",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"0D",X"EE",
		X"44",X"44",X"47",X"77",X"47",X"11",X"47",X"88",X"47",X"88",X"47",X"87",X"47",X"89",X"47",X"89",
		X"44",X"44",X"77",X"77",X"11",X"11",X"89",X"77",X"89",X"79",X"97",X"98",X"77",X"88",X"79",X"88",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CD",X"DD",X"DD",X"FF",X"FF",X"11",X"11",X"DD",X"DD",
		X"1D",X"CC",X"1D",X"CC",X"DD",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"DC",X"CC",X"ED",X"CC",
		X"CC",X"CD",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"ED",X"CC",X"1E",X"CC",X"1E",X"DD",X"D1",X"FF",X"DD",X"11",X"CD",X"DD",X"CD",X"DC",X"CC",X"DC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"DD",X"DD",X"FF",X"FF",X"11",X"11",X"DD",X"DD",
		X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1D",X"CC",X"1E",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"11",X"CC",X"D1",X"DD",X"D1",X"DD",X"DD",X"EE",X"CD",X"11",X"CC",X"DD",X"CC",X"DC",X"CC",X"DC",
		X"47",X"89",X"47",X"97",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"97",X"47",X"89",
		X"98",X"88",X"99",X"88",X"77",X"88",X"77",X"98",X"77",X"98",X"77",X"88",X"99",X"88",X"98",X"88",
		X"47",X"89",X"47",X"89",X"47",X"97",X"46",X"89",X"47",X"88",X"47",X"44",X"47",X"67",X"41",X"11",
		X"79",X"88",X"77",X"88",X"97",X"98",X"89",X"79",X"89",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"88",X"88",X"88",X"89",X"88",X"97",X"88",X"77",X"88",X"77",X"88",X"97",X"88",X"89",X"88",X"88",
		X"77",X"84",X"77",X"94",X"97",X"74",X"77",X"74",X"77",X"74",X"97",X"74",X"77",X"94",X"77",X"84",
		X"88",X"88",X"88",X"89",X"88",X"97",X"99",X"77",X"77",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"77",X"84",X"77",X"84",X"99",X"84",X"88",X"84",X"88",X"84",X"44",X"44",X"77",X"77",X"11",X"11",
		X"EE",X"EE",X"CC",X"CC",X"FF",X"FF",X"17",X"DF",X"17",X"DF",X"17",X"DF",X"17",X"DF",X"1E",X"DD",
		X"EE",X"EE",X"CC",X"CC",X"FF",X"FF",X"88",X"DF",X"88",X"DF",X"88",X"DF",X"88",X"DF",X"8E",X"DD",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"99",X"77",X"88",X"97",X"88",X"89",X"88",X"88",
		X"44",X"44",X"77",X"77",X"11",X"14",X"88",X"84",X"88",X"84",X"99",X"84",X"77",X"84",X"77",X"84",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"0D",X"EE",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"78",X"EF",X"78",X"EF",X"78",X"EF",X"78",X"EF",X"7D",X"EE",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"0D",X"EE",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"99",X"EF",X"99",X"EF",X"99",X"EF",X"99",X"EF",X"9D",X"EE",
		X"FF",X"77",X"CC",X"F7",X"CC",X"FF",X"EE",X"CF",X"FF",X"CC",X"11",X"EC",X"77",X"FE",X"77",X"1F",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"F7",X"77",X"FF",X"77",X"CF",X"77",X"CC",X"F7",
		X"88",X"71",X"77",X"77",X"11",X"87",X"FF",X"78",X"EE",X"17",X"EE",X"11",X"EE",X"FF",X"EE",X"EE",
		X"EC",X"FF",X"FE",X"CF",X"1F",X"CC",X"71",X"EC",X"77",X"FE",X"87",X"1F",X"78",X"71",X"17",X"77",
		X"97",X"97",X"17",X"17",X"97",X"97",X"97",X"97",X"17",X"17",X"97",X"97",X"97",X"97",X"17",X"17",
		X"77",X"77",X"17",X"77",X"11",X"77",X"99",X"77",X"17",X"17",X"97",X"11",X"97",X"91",X"17",X"17",
		X"97",X"97",X"97",X"97",X"17",X"17",X"97",X"97",X"97",X"97",X"17",X"17",X"97",X"DE",X"97",X"DE",
		X"77",X"77",X"97",X"77",X"99",X"77",X"F9",X"77",X"CF",X"97",X"CC",X"DD",X"EC",X"FE",X"FE",X"CF",
		X"44",X"44",X"18",X"88",X"17",X"77",X"17",X"99",X"17",X"48",X"17",X"48",X"17",X"84",X"17",X"84",
		X"44",X"44",X"18",X"88",X"77",X"77",X"99",X"99",X"48",X"49",X"48",X"49",X"84",X"89",X"84",X"89",
		X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",
		X"78",X"90",X"78",X"90",X"78",X"90",X"78",X"90",X"78",X"90",X"78",X"90",X"78",X"90",X"78",X"90",
		X"44",X"44",X"47",X"77",X"47",X"99",X"47",X"97",X"47",X"97",X"47",X"77",X"47",X"77",X"47",X"77",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"77",X"77",X"77",X"99",X"77",X"77",X"77",X"79",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"99",X"77",X"77",X"77",X"88",X"99",X"88",X"79",
		X"44",X"44",X"77",X"77",X"29",X"99",X"77",X"29",X"77",X"99",X"77",X"79",X"77",X"79",X"77",X"72",
		X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",
		X"79",X"79",X"79",X"87",X"97",X"88",X"97",X"88",X"97",X"99",X"97",X"99",X"79",X"97",X"79",X"78",
		X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"97",X"47",X"97",X"47",X"99",X"47",X"77",X"41",X"11",
		X"77",X"78",X"77",X"77",X"77",X"99",X"77",X"77",X"77",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"88",X"77",X"88",X"97",X"87",X"99",X"99",X"99",X"98",X"88",X"97",X"88",X"99",X"87",X"99",X"77",
		X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",
		X"99",X"79",X"99",X"99",X"77",X"77",X"99",X"77",X"77",X"77",X"44",X"44",X"77",X"77",X"11",X"11",
		X"77",X"72",X"77",X"79",X"77",X"79",X"77",X"99",X"77",X"29",X"29",X"99",X"77",X"77",X"11",X"11",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"0D",X"EE",
		X"DD",X"DD",X"CC",X"CC",X"FF",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"0D",X"EE",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"77",X"99",X"77",X"77",X"77",X"88",X"99",X"88",X"79",
		X"44",X"44",X"77",X"77",X"11",X"11",X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",X"77",X"74",
		X"00",X"27",X"02",X"98",X"00",X"A9",X"00",X"A9",X"00",X"98",X"02",X"89",X"00",X"87",X"0A",X"79",
		X"00",X"00",X"00",X"00",X"27",X"00",X"99",X"00",X"AA",X"70",X"00",X"80",X"00",X"80",X"20",X"00",
		X"0A",X"9A",X"0A",X"89",X"0A",X"88",X"0A",X"AA",X"00",X"A2",X"00",X"A2",X"02",X"A8",X"28",X"AA",
		X"00",X"00",X"98",X"00",X"99",X"92",X"A7",X"A9",X"99",X"99",X"90",X"00",X"AA",X"07",X"99",X"99",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"DD",X"EE",X"EE",X"FC",X"CF",X"0C",X"CF",X"0E",X"EF",X"0E",X"EF",
		X"FF",X"FF",X"CC",X"CC",X"CC",X"DD",X"CC",X"EE",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",
		X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",
		X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",
		X"77",X"77",X"11",X"27",X"98",X"79",X"79",X"91",X"87",X"18",X"27",X"98",X"79",X"98",X"91",X"79",
		X"77",X"77",X"11",X"27",X"98",X"79",X"79",X"91",X"87",X"18",X"27",X"98",X"79",X"98",X"91",X"79",
		X"18",X"87",X"98",X"27",X"98",X"79",X"79",X"91",X"87",X"18",X"27",X"98",X"77",X"78",X"99",X"99",
		X"18",X"87",X"98",X"27",X"98",X"79",X"79",X"91",X"87",X"18",X"97",X"98",X"77",X"78",X"99",X"99",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"64",X"77",X"64",X"77",X"64",X"77",X"64",X"77",X"64",X"77",X"64",X"77",X"64",X"77",X"64",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"66",X"44",X"44",X"77",X"77",X"11",X"11",
		X"77",X"94",X"77",X"94",X"76",X"94",X"66",X"94",X"99",X"94",X"44",X"44",X"77",X"77",X"11",X"11",
		X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",
		X"DC",X"CD",X"DC",X"CD",X"DC",X"CD",X"DC",X"CD",X"DC",X"CD",X"DC",X"CD",X"DC",X"CD",X"DC",X"CD",
		X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",
		X"EF",X"CE",X"EF",X"CE",X"EF",X"CE",X"EF",X"CE",X"EF",X"CE",X"EF",X"CE",X"EF",X"CE",X"EF",X"CE",
		X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",X"0F",X"FF",X"0C",X"CF",X"0D",X"DF",X"0E",X"EF",
		X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"CC",X"EF",X"FF",X"EF",X"FF",X"EF",X"FF",X"FF",
		X"00",X"00",X"00",X"EF",X"00",X"CC",X"00",X"EC",X"00",X"CE",X"0C",X"EE",X"0E",X"11",X"00",X"88",
		X"00",X"FC",X"FF",X"CC",X"CC",X"CE",X"CC",X"CE",X"EE",X"FE",X"FF",X"FF",X"11",X"11",X"88",X"88",
		X"02",X"27",X"00",X"19",X"00",X"72",X"00",X"81",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"91",X"91",X"77",X"77",X"18",X"18",X"18",X"18",X"11",X"11",X"11",X"11",X"11",X"11",
		X"EF",X"F1",X"EF",X"18",X"EF",X"84",X"EF",X"77",X"E1",X"71",X"18",X"17",X"84",X"78",X"77",X"88",
		X"77",X"77",X"71",X"81",X"17",X"77",X"78",X"44",X"88",X"88",X"88",X"11",X"11",X"11",X"11",X"11",
		X"71",X"81",X"17",X"11",X"78",X"19",X"88",X"99",X"88",X"99",X"99",X"98",X"98",X"88",X"88",X"88",
		X"11",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"77",X"77",X"77",
		X"88",X"88",X"09",X"99",X"00",X"47",X"00",X"88",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"77",X"00",X"DD",X"FF",X"EE",X"CC",X"DD",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CC",X"CC",X"DD",X"CD",X"EE",X"FF",X"FF",X"CC",X"EF",X"CC",X"FF",X"EF",X"CC",X"FF",
		X"FF",X"EF",X"CC",X"FF",X"CC",X"E1",X"EF",X"DE",X"FF",X"CF",X"E1",X"F8",X"DE",X"87",X"CF",X"11",
		X"CC",X"E1",X"EF",X"DE",X"EF",X"CF",X"DE",X"F8",X"CF",X"87",X"F7",X"11",X"88",X"DE",X"87",X"DE",
		X"F8",X"77",X"87",X"77",X"11",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"DE",X"77",X"DE",
		X"DE",X"91",X"CF",X"17",X"F8",X"77",X"99",X"77",X"11",X"77",X"77",X"77",X"77",X"71",X"7D",X"19",
		X"77",X"D9",X"77",X"98",X"77",X"88",X"79",X"88",X"98",X"11",X"81",X"19",X"11",X"19",X"19",X"19",
		X"77",X"99",X"77",X"19",X"11",X"19",X"19",X"19",X"89",X"99",X"19",X"19",X"19",X"DE",X"99",X"DE",
		X"99",X"99",X"19",X"19",X"19",X"19",X"19",X"19",X"99",X"99",X"19",X"19",X"19",X"DE",X"88",X"DE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"7F",X"77",X"FF",
		X"77",X"7F",X"77",X"FF",X"77",X"CC",X"7F",X"CC",X"FF",X"EE",X"CC",X"FF",X"CC",X"11",X"EE",X"77",
		X"77",X"CC",X"7F",X"CC",X"FF",X"EE",X"CC",X"FF",X"CC",X"11",X"EE",X"77",X"FF",X"77",X"11",X"88",
		X"FF",X"77",X"11",X"88",X"77",X"77",X"77",X"71",X"88",X"1F",X"77",X"FE",X"11",X"EE",X"FF",X"EE",
		X"88",X"88",X"77",X"77",X"17",X"97",X"17",X"17",X"17",X"17",X"87",X"87",X"87",X"87",X"17",X"17",
		X"88",X"88",X"77",X"77",X"97",X"99",X"17",X"18",X"17",X"18",X"87",X"88",X"87",X"88",X"17",X"18",
		X"88",X"88",X"87",X"77",X"87",X"97",X"87",X"17",X"87",X"17",X"87",X"87",X"87",X"87",X"87",X"17",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"17",X"87",X"17",X"87",X"77",X"87",X"97",X"87",X"17",X"87",X"17",X"87",X"17",X"87",X"17",
		X"17",X"17",X"17",X"17",X"77",X"77",X"97",X"97",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",
		X"87",X"77",X"87",X"97",X"87",X"17",X"87",X"17",X"87",X"17",X"87",X"87",X"87",X"77",X"89",X"99",
		X"77",X"77",X"97",X"97",X"17",X"17",X"17",X"17",X"17",X"17",X"87",X"87",X"77",X"77",X"99",X"99",
		X"17",X"18",X"17",X"18",X"77",X"77",X"97",X"98",X"17",X"18",X"17",X"18",X"17",X"18",X"17",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"97",X"98",X"17",X"18",X"17",X"18",X"17",X"18",X"87",X"88",X"77",X"77",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",X"47",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"47",X"67",X"47",X"66",X"47",X"99",X"47",X"79",X"47",X"99",X"47",X"44",X"47",X"77",X"11",X"11",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"66",X"44",X"44",X"77",X"77",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"EE",X"EE",X"CC",X"CC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"97",X"66",X"E9",X"EE",X"C9",X"CC",X"B9",X"EB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"66",X"87",X"EE",X"87",X"CC",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"BB",X"ED",X"BB",X"EE",X"BB",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"D7",X"DD",X"0D",X"BB",X"0D",X"BB",X"7D",X"BB",X"8D",X"BB",X"8D",X"BB",X"8D",X"BB",X"BD",
		X"DD",X"D8",X"DD",X"88",X"BB",X"88",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"BB",
		X"BD",X"DD",X"DD",X"DD",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"66",X"99",X"EE",X"99",X"DD",X"D9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"8B",X"66",X"BE",X"EE",X"BE",X"DD",X"BE",X"BB",X"ED",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"D9",X"D9",X"D9",X"DA",X"B9",X"BA",X"B9",X"BA",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"97",X"BB",X"97",X"BB",X"97",X"BB",X"97",X"7B",X"97",X"7B",X"97",X"7B",X"97",X"7B",X"97",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"7B",X"97",X"C7",X"C9",X"B7",X"79",X"B7",X"79",X"B7",X"79",X"B7",X"79",X"B7",X"79",X"87",X"79",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"EE",X"B7",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"88",X"BB",X"87",X"88",X"77",X"BB",X"87",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"BB",X"BD",X"BB",X"BD",X"BD",X"BD",X"BD",X"BD",X"DB",X"BD",X"DB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"D8",X"DD",X"88",X"BB",X"88",X"9B",X"B8",X"BD",X"B8",X"BB",X"B8",X"BB",X"B8",X"9B",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"BB",X"ED",X"BB",X"EE",X"BB",X"BE",X"BE",X"EB",X"BE",X"EB",X"BE",X"EB",X"BE",X"EB",X"BE",X"EB",
		X"DD",X"DE",X"DD",X"ED",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",
		X"BB",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"8D",X"D8",X"D8",X"88",X"B8",X"88",X"B8",X"B8",X"B8",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"8B",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"CB",X"BB",
		X"B9",X"9B",X"B9",X"9B",X"B9",X"9B",X"B9",X"9B",X"B9",X"9B",X"B9",X"9B",X"B9",X"9B",X"B9",X"9B",
		X"BB",X"ED",X"BB",X"EE",X"BB",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",
		X"DE",X"ED",X"DD",X"DD",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"BB",X"BB",
		X"EE",X"BE",X"EE",X"BE",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",X"EE",X"EB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"D9",X"D8",X"D9",X"88",X"BB",X"88",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"B8",X"BB",X"BB",
		X"9B",X"BE",X"9B",X"BE",X"B9",X"BE",X"B9",X"BE",X"B9",X"BE",X"B9",X"BE",X"B9",X"BE",X"B9",X"BE",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"22",X"66",X"2E",X"EE",X"EE",X"ED",X"EE",X"DB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"66",X"66",X"EE",X"EE",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"97",X"66",X"E9",X"EE",X"C9",X"CC",X"B9",X"EB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"66",X"87",X"EE",X"87",X"CC",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"EB",X"DB",X"EB",X"DB",X"EB",X"DB",X"EB",X"DB",X"EB",X"DB",X"EB",X"DB",X"EB",X"DB",X"EB",X"DB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"B9",X"EB",X"B9",X"EB",X"B9",X"EB",X"B9",X"EB",X"B9",X"EB",X"B9",X"EB",X"B9",X"EB",X"B9",X"EB",
		X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",
		X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",X"BB",X"EB",
		X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",
		X"BB",X"66",X"BE",X"EE",X"EE",X"ED",X"EE",X"DB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BD",X"97",X"DD",X"99",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"66",X"88",X"EE",X"88",X"DD",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"66",X"66",X"EE",X"E8",X"DD",X"88",X"BB",X"B8",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",X"BB",X"BE",
		X"BB",X"BB",X"66",X"66",X"EE",X"EE",X"DD",X"DD",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BE",X"BB",X"BE",X"BB",X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"BD",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"66",X"66",X"EE",X"EE",X"DD",X"D9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"66",X"99",X"EE",X"99",X"ED",X"98",X"BB",X"98",X"BB",X"98",X"BB",X"98",X"BB",X"98",X"BB",X"98",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"66",X"66",X"EE",X"EE",X"EE",X"ED",X"EE",X"DB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BD",X"97",X"DD",X"99",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"66",X"68",X"EE",X"88",X"DD",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"EE",X"9B",X"EE",X"99",X"DD",X"D9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"7B",X"EE",X"BE",X"EE",X"BE",X"DD",X"BE",X"BB",X"ED",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"BB",X"EE",X"BE",X"EE",X"EE",X"ED",X"EE",X"DB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BD",X"97",X"DD",X"99",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"EE",X"88",X"EE",X"88",X"DD",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"BB",X"EE",X"BB",X"EE",X"BE",X"ED",X"EE",X"DB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"EE",X"EE",X"EE",X"EE",X"CC",X"CC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"97",X"EE",X"E9",X"EE",X"C9",X"CC",X"B9",X"EB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"EE",X"88",X"EE",X"88",X"CC",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"ED",X"EE",X"DB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",X"EE",X"BB",
		X"BD",X"97",X"DD",X"99",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"EE",X"88",X"EE",X"88",X"DD",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",X"BB",X"87",
		X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",X"DB",X"88",
		X"66",X"9B",X"EE",X"99",X"DD",X"D9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"7B",X"66",X"BE",X"EE",X"BE",X"DD",X"BE",X"BB",X"ED",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",
		X"97",X"66",X"E9",X"EE",X"C9",X"CC",X"B9",X"EB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BD",X"D7",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",X"DD",X"77",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"EE",X"22",X"66",X"2E",X"66",X"C6",X"66",X"C6",X"CC",X"C6",X"EE",X"CC",X"EE",X"22",X"EE",
		X"2E",X"EE",X"66",X"66",X"DE",X"EE",X"EE",X"EE",X"DE",X"EE",X"DD",X"EE",X"ED",X"EE",X"EE",X"DE",
		X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",X"CE",X"22",X"CC",X"22",X"CC",X"22",X"BB",X"22",X"22",
		X"EE",X"DE",X"EE",X"DE",X"EE",X"DE",X"CC",X"CC",X"EC",X"BB",X"CB",X"B2",X"BB",X"22",X"22",X"22",
		X"22",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6D",X"66",X"DD",X"66",X"DD",
		X"26",X"66",X"66",X"6E",X"6E",X"66",X"66",X"66",X"66",X"CD",X"66",X"CD",X"66",X"CC",X"66",X"CC",
		X"66",X"66",X"DD",X"66",X"EE",X"DD",X"CC",X"EE",X"BB",X"CC",X"22",X"BC",X"22",X"BB",X"22",X"22",
		X"66",X"CC",X"66",X"EC",X"EE",X"CE",X"CC",X"BC",X"CB",X"2B",X"B2",X"22",X"22",X"22",X"22",X"22",
		X"22",X"66",X"66",X"6E",X"66",X"E6",X"66",X"66",X"66",X"EE",X"66",X"DE",X"66",X"DD",X"66",X"DD",
		X"66",X"66",X"EE",X"66",X"66",X"66",X"66",X"66",X"66",X"E6",X"66",X"E6",X"EE",X"66",X"DD",X"66",
		X"66",X"66",X"EE",X"66",X"DD",X"EE",X"CC",X"DD",X"BB",X"CD",X"22",X"BC",X"22",X"2B",X"22",X"22",
		X"DD",X"66",X"66",X"66",X"66",X"6E",X"66",X"EE",X"EE",X"DD",X"DD",X"CC",X"CC",X"BB",X"BB",X"22",
		X"00",X"66",X"66",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"60",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"66",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",X"00",X"00",X"00",X"00",
		X"40",X"14",X"04",X"10",X"10",X"24",X"14",X"20",X"10",X"41",X"14",X"0D",X"D0",X"24",X"2A",X"00",
		X"10",X"10",X"41",X"11",X"01",X"24",X"41",X"10",X"1D",X"4D",X"11",X"41",X"AD",X"01",X"41",X"DD",
		X"4D",X"4A",X"0A",X"0D",X"AE",X"4A",X"0A",X"AE",X"AE",X"AD",X"D0",X"EE",X"0E",X"EE",X"EE",X"EE",
		X"0A",X"4D",X"AA",X"0A",X"AA",X"A4",X"D0",X"00",X"0E",X"AA",X"EE",X"EA",X"EE",X"E0",X"EE",X"0E",
		X"41",X"01",X"14",X"10",X"20",X"4C",X"02",X"02",X"C4",X"C1",X"4C",X"40",X"10",X"0C",X"4C",X"C1",
		X"10",X"C1",X"12",X"14",X"01",X"0C",X"CC",X"14",X"24",X"02",X"4C",X"4C",X"2C",X"0C",X"0C",X"CB",
		X"0B",X"40",X"2B",X"B2",X"0B",X"40",X"B1",X"0B",X"B0",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"B4",X"1B",X"BC",X"B4",X"B4",X"1B",X"B0",X"04",X"BB",X"B0",X"BB",X"4B",X"BB",X"0B",X"BB",X"BB",
		X"00",X"14",X"0F",X"F0",X"10",X"24",X"C4",X"20",X"C0",X"FC",X"14",X"0C",X"B0",X"2F",X"2B",X"C0",
		X"10",X"F0",X"4C",X"C1",X"0C",X"C4",X"4F",X"10",X"CC",X"4C",X"C1",X"4F",X"BC",X"0C",X"B1",X"CB",
		X"4B",X"4B",X"0B",X"BF",X"BB",X"B0",X"4B",X"BF",X"0C",X"B0",X"BB",X"BB",X"BB",X"CB",X"BB",X"BB",
		X"BB",X"4C",X"BB",X"0B",X"BC",X"B4",X"BB",X"B0",X"BB",X"FB",X"BB",X"0B",X"CB",X"BB",X"BB",X"BB",
		X"F1",X"0F",X"14",X"10",X"2F",X"4F",X"02",X"02",X"A4",X"A1",X"4B",X"40",X"10",X"0B",X"4E",X"B1",
		X"10",X"A1",X"F2",X"F4",X"01",X"0B",X"AA",X"14",X"24",X"02",X"4B",X"4F",X"2B",X"0A",X"0B",X"AE",
		X"0F",X"40",X"2E",X"B2",X"0E",X"40",X"EF",X"0E",X"E0",X"BB",X"0E",X"EC",X"EE",X"EE",X"EE",X"EE",
		X"F4",X"FB",X"BB",X"A4",X"EF",X"1B",X"E0",X"0F",X"EE",X"BE",X"EE",X"F0",X"EE",X"0E",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"1A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"B2",X"22",X"21",X"21",X"18",X"11",X"11",X"11",X"22",X"82",X"22",X"22",X"20",X"20",X"00",X"00",
		X"22",X"22",X"21",X"21",X"11",X"11",X"11",X"81",X"22",X"22",X"21",X"22",X"20",X"20",X"00",X"00",
		X"0A",X"0A",X"AA",X"AA",X"AB",X"AB",X"BB",X"BB",X"BB",X"CB",X"EA",X"CC",X"EE",X"CC",X"EE",X"AC",
		X"0A",X"0A",X"AA",X"AA",X"AB",X"AB",X"BB",X"BC",X"BB",X"EC",X"BC",X"0A",X"CC",X"AC",X"DD",X"CC",
		X"22",X"13",X"22",X"21",X"26",X"22",X"11",X"26",X"31",X"13",X"11",X"11",X"01",X"11",X"00",X"00",
		X"21",X"21",X"21",X"22",X"02",X"22",X"12",X"22",X"31",X"01",X"11",X"11",X"00",X"11",X"00",X"00",
		X"A0",X"00",X"AA",X"DA",X"BA",X"DA",X"BB",X"DB",X"CC",X"DB",X"CC",X"DB",X"BC",X"DB",X"BB",X"DB",
		X"AA",X"00",X"AA",X"AA",X"BB",X"BB",X"BB",X"DB",X"BB",X"DB",X"AB",X"DB",X"AB",X"DD",X"AA",X"DD",
		X"81",X"58",X"05",X"50",X"10",X"01",X"52",X"11",X"08",X"22",X"25",X"52",X"20",X"02",X"0C",X"C0",
		X"18",X"15",X"50",X"50",X"01",X"05",X"11",X"10",X"25",X"11",X"50",X"05",X"0C",X"C0",X"BC",X"CC",
		X"CC",X"BC",X"CC",X"CC",X"CB",X"CC",X"CC",X"CC",X"CC",X"CB",X"BC",X"CC",X"CC",X"BB",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CB",X"CB",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CB",X"BB",X"CC",X"CC",X"CC",
		X"22",X"22",X"33",X"31",X"11",X"11",X"11",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"1A",X"10",
		X"21",X"22",X"12",X"33",X"12",X"11",X"11",X"00",X"01",X"00",X"01",X"AA",X"A1",X"AA",X"A1",X"AA",
		X"1A",X"10",X"1C",X"1A",X"0C",X"1C",X"0C",X"1C",X"AC",X"1D",X"AC",X"0D",X"CE",X"0D",X"CE",X"AD",
		X"B1",X"AA",X"B0",X"AA",X"BA",X"AA",X"BB",X"BA",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CA",X"CC",X"CA",X"CA",X"CB",X"CA",X"CC",X"CB",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"AC",X"CC",X"A0",X"CC",X"BC",X"CA",X"CC",X"CA",X"CC",X"CA",X"CC",X"CB",X"CC",X"CC",X"CC",
		X"BB",X"BB",X"BB",X"AB",X"BC",X"BA",X"BC",X"BA",X"BB",X"BC",X"BC",X"CB",X"CB",X"AB",X"CB",X"AB",
		X"CC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"CA",X"BB",X"BB",X"AB",X"BB",X"AB",X"BC",X"CC",X"CB",
		X"BC",X"BB",X"CB",X"BB",X"CB",X"CC",X"BB",X"BB",X"BB",X"AB",X"BC",X"BA",X"BC",X"BA",X"BB",X"BB",
		X"BB",X"CB",X"BB",X"BB",X"BB",X"BB",X"BB",X"AB",X"BC",X"BA",X"BC",X"BA",X"BB",X"BB",X"BB",X"BB",
		X"72",X"07",X"14",X"10",X"27",X"47",X"02",X"02",X"14",X"21",X"4D",X"40",X"10",X"0D",X"4D",X"E1",
		X"10",X"D1",X"71",X"74",X"01",X"01",X"12",X"14",X"24",X"02",X"12",X"47",X"2A",X"0B",X"0A",X"AB",
		X"07",X"40",X"2D",X"D2",X"0D",X"40",X"D7",X"0E",X"E0",X"EE",X"EE",X"EE",X"DE",X"EE",X"DE",X"EE",
		X"74",X"7A",X"BA",X"A4",X"B7",X"1A",X"B0",X"07",X"BB",X"A0",X"BB",X"7A",X"BB",X"0A",X"BB",X"BB",
		X"CD",X"ED",X"DD",X"ED",X"DD",X"ED",X"DE",X"ED",X"DE",X"ED",X"DE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"CC",X"EE",X"CC",X"EE",X"DC",X"ED",X"DC",X"ED",X"DC",X"ED",X"DC",X"EE",X"DC",X"EE",X"DC",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",
		X"DC",X"EE",X"DD",X"EE",X"DD",X"CE",X"DD",X"CD",X"DD",X"CD",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",
		X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"CC",X"DD",X"DC",X"DD",X"DC",X"DD",X"DE",X"DD",X"DE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"ED",X"EE",X"ED",X"EE",X"ED",X"EE",X"22",X"EE",
		X"DD",X"DE",X"DD",X"DE",X"DD",X"CE",X"DD",X"CE",X"DD",X"EE",X"DD",X"EE",X"DC",X"1E",X"11",X"12",
		X"AB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DB",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",
		X"AA",X"DD",X"AA",X"DD",X"AA",X"DB",X"AA",X"DB",X"AA",X"DB",X"AA",X"DD",X"BA",X"DD",X"BA",X"DD",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",X"BD",X"DB",
		X"BA",X"DD",X"BA",X"DD",X"BA",X"AD",X"BA",X"AB",X"BA",X"AB",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",
		X"BD",X"DB",X"AD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DB",X"DD",X"DD",X"DD",X"DD",
		X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"1D",X"DD",X"28",X"2D",
		X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"11",X"28",X"12",
		X"DE",X"CD",X"DD",X"CE",X"DD",X"CE",X"DD",X"EE",X"DD",X"EE",X"DD",X"DD",X"BD",X"EE",X"DD",X"EE",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BD",X"BB",X"AD",X"BA",X"BD",X"AB",X"BD",X"BB",X"BD",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"DD",X"DD",X"EE",X"DD",X"EE",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BA",X"DE",X"AB",X"DE",
		X"DD",X"DE",X"BD",X"DE",X"BD",X"DE",X"BD",X"DE",X"BD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DD",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BA",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"11",X"11",X"12",X"11",X"22",X"22",
		X"AB",X"DD",X"BD",X"DD",X"BD",X"DD",X"BD",X"DB",X"B1",X"EB",X"B1",X"E1",X"21",X"12",X"22",X"22",
		X"BB",X"DE",X"AB",X"DE",X"EA",X"DE",X"EA",X"DE",X"EA",X"DE",X"AA",X"EE",X"A0",X"EE",X"C0",X"EB",
		X"EB",X"CB",X"EB",X"BB",X"BB",X"AA",X"BB",X"0A",X"BB",X"0D",X"BB",X"BD",X"BA",X"BC",X"BA",X"B0",
		X"AA",X"AB",X"AC",X"AC",X"AA",X"AE",X"A0",X"EE",X"AA",X"EE",X"CB",X"EE",X"BD",X"EE",X"11",X"EE",
		X"BB",X"B0",X"BB",X"BB",X"AC",X"BB",X"AA",X"BB",X"AA",X"AB",X"AE",X"AA",X"1E",X"AA",X"11",X"A1",
		X"BB",X"DE",X"AB",X"DE",X"EA",X"DE",X"EA",X"DE",X"EA",X"DE",X"AA",X"EE",X"A0",X"EE",X"C0",X"EB",
		X"EB",X"CB",X"EB",X"BB",X"BB",X"AA",X"BB",X"0A",X"BB",X"0D",X"BB",X"BD",X"BA",X"BC",X"BA",X"B0",
		X"AA",X"AB",X"AC",X"AC",X"AA",X"AE",X"A0",X"EE",X"AA",X"EE",X"CB",X"EE",X"BD",X"EE",X"BD",X"EE",
		X"BB",X"B0",X"BB",X"BB",X"AC",X"BB",X"AA",X"BB",X"AA",X"AB",X"AE",X"AA",X"AE",X"AA",X"AE",X"EA",
		X"BB",X"BD",X"BC",X"DD",X"CA",X"DD",X"AA",X"AD",X"AA",X"AC",X"AE",X"AC",X"EE",X"AA",X"DE",X"AA",
		X"EA",X"CC",X"EE",X"BC",X"EA",X"BC",X"AA",X"BC",X"A0",X"BC",X"BB",X"BC",X"BC",X"BB",X"CC",X"AB",
		X"BD",X"A0",X"DD",X"0B",X"DD",X"BB",X"DD",X"BC",X"DD",X"CC",X"DD",X"CC",X"DB",X"CD",X"DB",X"DD",
		X"CD",X"AA",X"DD",X"AA",X"DD",X"AA",X"DD",X"DA",X"DD",X"D0",X"BB",X"0D",X"AA",X"DD",X"AA",X"CD",
		X"DD",X"DE",X"BD",X"DE",X"BD",X"DE",X"BD",X"DE",X"BD",X"DE",X"DD",X"DE",X"DD",X"DE",X"DD",X"DD",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BA",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AB",X"DD",X"BD",X"DD",X"BD",X"DD",X"BD",X"DB",X"B1",X"EB",X"B1",X"E1",X"11",X"11",X"11",X"11",
		X"DB",X"DB",X"BD",X"BD",X"CB",X"DB",X"DC",X"CC",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"CC",X"DD",
		X"DB",X"DB",X"BD",X"CC",X"CC",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"CC",X"CC",X"DE",
		X"CC",X"CC",X"DE",X"DE",X"ED",X"ED",X"DE",X"DE",X"ED",X"ED",X"CC",X"DE",X"DD",X"CC",X"BD",X"BD",
		X"ED",X"ED",X"DE",X"DE",X"ED",X"ED",X"DE",X"DE",X"ED",X"CC",X"CC",X"BD",X"DB",X"DB",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"06",X"00",X"00",X"06",X"00",X"60",X"00",X"60",X"00",X"06",X"06",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
