`define BUILD_DATE "180607"
`define BUILD_TIME "201354"
