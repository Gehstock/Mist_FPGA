-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity INVADERS_ROM_H is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of INVADERS_ROM_H is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"00",x"00",x"C3",x"D4",x"18",x"00",x"00", -- 0x0000
    x"F5",x"C5",x"D5",x"E5",x"C3",x"8C",x"00",x"00", -- 0x0008
    x"F5",x"C5",x"D5",x"E5",x"3E",x"80",x"32",x"72", -- 0x0010
    x"20",x"21",x"C0",x"20",x"35",x"CD",x"CD",x"17", -- 0x0018
    x"DB",x"01",x"0F",x"DA",x"67",x"00",x"3A",x"EA", -- 0x0020
    x"20",x"A7",x"CA",x"42",x"00",x"3A",x"EB",x"20", -- 0x0028
    x"FE",x"99",x"CA",x"3E",x"00",x"C6",x"01",x"27", -- 0x0030
    x"32",x"EB",x"20",x"CD",x"47",x"19",x"AF",x"32", -- 0x0038
    x"EA",x"20",x"3A",x"E9",x"20",x"A7",x"CA",x"82", -- 0x0040
    x"00",x"3A",x"EF",x"20",x"A7",x"C2",x"6F",x"00", -- 0x0048
    x"3A",x"EB",x"20",x"A7",x"C2",x"5D",x"00",x"CD", -- 0x0050
    x"BF",x"0A",x"C3",x"82",x"00",x"3A",x"93",x"20", -- 0x0058
    x"A7",x"C2",x"82",x"00",x"C3",x"65",x"07",x"3E", -- 0x0060
    x"01",x"32",x"EA",x"20",x"C3",x"3F",x"00",x"CD", -- 0x0068
    x"40",x"17",x"3A",x"32",x"20",x"32",x"80",x"20", -- 0x0070
    x"CD",x"00",x"01",x"CD",x"48",x"02",x"CD",x"13", -- 0x0078
    x"09",x"00",x"E1",x"D1",x"C1",x"F1",x"FB",x"C9", -- 0x0080
    x"00",x"00",x"00",x"00",x"AF",x"32",x"72",x"20", -- 0x0088
    x"3A",x"E9",x"20",x"A7",x"CA",x"82",x"00",x"3A", -- 0x0090
    x"EF",x"20",x"A7",x"C2",x"A5",x"00",x"3A",x"C1", -- 0x0098
    x"20",x"0F",x"D2",x"82",x"00",x"21",x"20",x"20", -- 0x00A0
    x"CD",x"4B",x"02",x"CD",x"41",x"01",x"C3",x"82", -- 0x00A8
    x"00",x"CD",x"86",x"08",x"E5",x"7E",x"23",x"66", -- 0x00B0
    x"6F",x"22",x"09",x"20",x"22",x"0B",x"20",x"E1", -- 0x00B8
    x"2B",x"7E",x"FE",x"03",x"C2",x"C8",x"00",x"3D", -- 0x00C0
    x"32",x"08",x"20",x"FE",x"FE",x"3E",x"00",x"C2", -- 0x00C8
    x"D3",x"00",x"3C",x"32",x"0D",x"20",x"C9",x"3E", -- 0x00D0
    x"02",x"32",x"FB",x"21",x"32",x"FB",x"22",x"C3", -- 0x00D8
    x"E4",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"21",x"02",x"20",x"7E",x"A7",x"C2",x"38",x"15", -- 0x0100
    x"E5",x"3A",x"06",x"20",x"6F",x"3A",x"67",x"20", -- 0x0108
    x"67",x"7E",x"A7",x"E1",x"CA",x"36",x"01",x"23", -- 0x0110
    x"23",x"7E",x"23",x"46",x"E6",x"FE",x"07",x"07", -- 0x0118
    x"07",x"5F",x"16",x"00",x"21",x"00",x"1C",x"19", -- 0x0120
    x"EB",x"78",x"A7",x"C4",x"3B",x"01",x"2A",x"0B", -- 0x0128
    x"20",x"06",x"10",x"CD",x"D3",x"15",x"AF",x"32", -- 0x0130
    x"00",x"20",x"C9",x"21",x"30",x"00",x"19",x"EB", -- 0x0138
    x"C9",x"3A",x"68",x"20",x"A7",x"C8",x"3A",x"00", -- 0x0140
    x"20",x"A7",x"C0",x"3A",x"67",x"20",x"67",x"3A", -- 0x0148
    x"06",x"20",x"16",x"02",x"3C",x"FE",x"37",x"CC", -- 0x0150
    x"A1",x"01",x"6F",x"46",x"05",x"C2",x"54",x"01", -- 0x0158
    x"32",x"06",x"20",x"CD",x"7A",x"01",x"61",x"22", -- 0x0160
    x"0B",x"20",x"7D",x"FE",x"28",x"DA",x"71",x"19", -- 0x0168
    x"7A",x"32",x"04",x"20",x"3E",x"01",x"32",x"00", -- 0x0170
    x"20",x"C9",x"16",x"00",x"7D",x"21",x"09",x"20", -- 0x0178
    x"46",x"23",x"4E",x"FE",x"0B",x"FA",x"94",x"01", -- 0x0180
    x"DE",x"0B",x"5F",x"78",x"C6",x"10",x"47",x"7B", -- 0x0188
    x"14",x"C3",x"83",x"01",x"68",x"A7",x"C8",x"5F", -- 0x0190
    x"79",x"C6",x"10",x"4F",x"7B",x"3D",x"C3",x"95", -- 0x0198
    x"01",x"15",x"CA",x"CD",x"01",x"21",x"06",x"20", -- 0x01A0
    x"36",x"00",x"23",x"4E",x"36",x"00",x"CD",x"D9", -- 0x01A8
    x"01",x"21",x"05",x"20",x"7E",x"3C",x"E6",x"01", -- 0x01B0
    x"77",x"AF",x"21",x"67",x"20",x"66",x"C9",x"00", -- 0x01B8
    x"21",x"00",x"21",x"06",x"37",x"36",x"01",x"23", -- 0x01C0
    x"05",x"C2",x"C5",x"01",x"C9",x"E1",x"C9",x"3E", -- 0x01C8
    x"01",x"06",x"E0",x"21",x"02",x"24",x"C3",x"CC", -- 0x01D0
    x"14",x"23",x"46",x"23",x"79",x"86",x"77",x"23", -- 0x01D8
    x"78",x"86",x"77",x"C9",x"06",x"C0",x"11",x"00", -- 0x01E0
    x"1B",x"21",x"00",x"20",x"C3",x"32",x"1A",x"21", -- 0x01E8
    x"42",x"21",x"C3",x"F8",x"01",x"21",x"42",x"22", -- 0x01F0
    x"0E",x"04",x"11",x"20",x"1D",x"D5",x"06",x"2C", -- 0x01F8
    x"CD",x"32",x"1A",x"D1",x"0D",x"C2",x"FD",x"01", -- 0x0200
    x"C9",x"3E",x"01",x"C3",x"1B",x"02",x"3E",x"01", -- 0x0208
    x"C3",x"14",x"02",x"AF",x"11",x"42",x"22",x"C3", -- 0x0210
    x"1E",x"02",x"AF",x"11",x"42",x"21",x"32",x"81", -- 0x0218
    x"20",x"01",x"02",x"16",x"21",x"06",x"28",x"3E", -- 0x0220
    x"04",x"F5",x"C5",x"3A",x"81",x"20",x"A7",x"C2", -- 0x0228
    x"42",x"02",x"CD",x"69",x"1A",x"C1",x"F1",x"3D", -- 0x0230
    x"C8",x"D5",x"11",x"E0",x"02",x"19",x"D1",x"C3", -- 0x0238
    x"29",x"02",x"CD",x"7C",x"14",x"C3",x"35",x"02", -- 0x0240
    x"21",x"10",x"20",x"7E",x"FE",x"FF",x"C8",x"FE", -- 0x0248
    x"FE",x"CA",x"81",x"02",x"23",x"46",x"4F",x"B0", -- 0x0250
    x"79",x"C2",x"77",x"02",x"23",x"7E",x"A7",x"C2", -- 0x0258
    x"88",x"02",x"23",x"5E",x"23",x"56",x"E5",x"EB", -- 0x0260
    x"E5",x"21",x"6F",x"02",x"E3",x"D5",x"E9",x"E1", -- 0x0268
    x"11",x"0C",x"00",x"19",x"C3",x"4B",x"02",x"05", -- 0x0270
    x"04",x"C2",x"7D",x"02",x"3D",x"05",x"70",x"2B", -- 0x0278
    x"77",x"11",x"10",x"00",x"19",x"C3",x"4B",x"02", -- 0x0280
    x"35",x"2B",x"2B",x"C3",x"81",x"02",x"E1",x"23", -- 0x0288
    x"7E",x"FE",x"FF",x"CA",x"3B",x"03",x"23",x"35", -- 0x0290
    x"C0",x"47",x"AF",x"32",x"68",x"20",x"32",x"69", -- 0x0298
    x"20",x"3E",x"30",x"32",x"6A",x"20",x"78",x"36", -- 0x02A0
    x"05",x"23",x"35",x"C2",x"9B",x"03",x"2A",x"1A", -- 0x02A8
    x"20",x"06",x"10",x"CD",x"24",x"14",x"21",x"10", -- 0x02B0
    x"20",x"11",x"10",x"1B",x"06",x"10",x"CD",x"32", -- 0x02B8
    x"1A",x"06",x"00",x"CD",x"DC",x"19",x"3A",x"6D", -- 0x02C0
    x"20",x"A7",x"C0",x"3A",x"EF",x"20",x"A7",x"C8", -- 0x02C8
    x"31",x"00",x"24",x"FB",x"CD",x"D7",x"19",x"CD", -- 0x02D0
    x"2E",x"09",x"A7",x"CA",x"6D",x"16",x"CD",x"E7", -- 0x02D8
    x"18",x"7E",x"A7",x"CA",x"2C",x"03",x"3A",x"CE", -- 0x02E0
    x"20",x"A7",x"CA",x"2C",x"03",x"3A",x"67",x"20", -- 0x02E8
    x"F5",x"0F",x"DA",x"32",x"03",x"CD",x"0E",x"02", -- 0x02F0
    x"CD",x"78",x"08",x"73",x"23",x"72",x"2B",x"2B", -- 0x02F8
    x"70",x"00",x"CD",x"E4",x"01",x"F1",x"0F",x"3E", -- 0x0300
    x"21",x"06",x"00",x"D2",x"12",x"03",x"06",x"20", -- 0x0308
    x"3E",x"22",x"32",x"67",x"20",x"CD",x"B6",x"0A", -- 0x0310
    x"AF",x"32",x"11",x"20",x"78",x"D3",x"05",x"3C", -- 0x0318
    x"32",x"98",x"20",x"CD",x"D6",x"09",x"CD",x"7F", -- 0x0320
    x"1A",x"C3",x"F9",x"07",x"CD",x"7F",x"1A",x"C3", -- 0x0328
    x"17",x"08",x"CD",x"09",x"02",x"C3",x"F8",x"02", -- 0x0330
    x"00",x"00",x"00",x"21",x"68",x"20",x"36",x"01", -- 0x0338
    x"23",x"7E",x"A7",x"C3",x"B0",x"03",x"00",x"2B", -- 0x0340
    x"36",x"01",x"3A",x"1B",x"20",x"47",x"3A",x"EF", -- 0x0348
    x"20",x"A7",x"C2",x"63",x"03",x"3A",x"1D",x"20", -- 0x0350
    x"0F",x"DA",x"81",x"03",x"0F",x"DA",x"8E",x"03", -- 0x0358
    x"C3",x"6F",x"03",x"CD",x"C0",x"17",x"07",x"07", -- 0x0360
    x"DA",x"81",x"03",x"07",x"DA",x"8E",x"03",x"21", -- 0x0368
    x"18",x"20",x"CD",x"3B",x"1A",x"CD",x"47",x"1A", -- 0x0370
    x"CD",x"39",x"14",x"3E",x"00",x"32",x"12",x"20", -- 0x0378
    x"C9",x"78",x"FE",x"D9",x"CA",x"6F",x"03",x"3C", -- 0x0380
    x"32",x"1B",x"20",x"C3",x"6F",x"03",x"78",x"FE", -- 0x0388
    x"30",x"CA",x"6F",x"03",x"3D",x"32",x"1B",x"20", -- 0x0390
    x"C3",x"6F",x"03",x"3C",x"E6",x"01",x"32",x"15", -- 0x0398
    x"20",x"07",x"07",x"07",x"07",x"21",x"70",x"1C", -- 0x03A0
    x"85",x"6F",x"22",x"18",x"20",x"C3",x"6F",x"03", -- 0x03A8
    x"C2",x"4A",x"03",x"23",x"35",x"C2",x"4A",x"03", -- 0x03B0
    x"C3",x"46",x"03",x"11",x"2A",x"20",x"CD",x"06", -- 0x03B8
    x"1A",x"E1",x"D0",x"23",x"7E",x"A7",x"C8",x"FE", -- 0x03C0
    x"01",x"CA",x"FA",x"03",x"FE",x"02",x"CA",x"0A", -- 0x03C8
    x"04",x"23",x"FE",x"03",x"C2",x"2A",x"04",x"35", -- 0x03D0
    x"CA",x"36",x"04",x"7E",x"FE",x"0F",x"C0",x"E5", -- 0x03D8
    x"CD",x"30",x"04",x"CD",x"52",x"14",x"E1",x"23", -- 0x03E0
    x"34",x"23",x"23",x"35",x"35",x"23",x"35",x"35", -- 0x03E8
    x"35",x"23",x"36",x"08",x"CD",x"30",x"04",x"C3", -- 0x03F0
    x"00",x"14",x"3C",x"77",x"3A",x"1B",x"20",x"C6", -- 0x03F8
    x"08",x"32",x"2A",x"20",x"CD",x"30",x"04",x"C3", -- 0x0400
    x"00",x"14",x"CD",x"30",x"04",x"D5",x"E5",x"C5", -- 0x0408
    x"CD",x"52",x"14",x"C1",x"E1",x"D1",x"3A",x"2C", -- 0x0410
    x"20",x"85",x"6F",x"32",x"29",x"20",x"CD",x"91", -- 0x0418
    x"14",x"3A",x"61",x"20",x"A7",x"C8",x"32",x"02", -- 0x0420
    x"20",x"C9",x"FE",x"05",x"C8",x"C3",x"36",x"04", -- 0x0428
    x"21",x"27",x"20",x"C3",x"3B",x"1A",x"CD",x"30", -- 0x0430
    x"04",x"CD",x"52",x"14",x"21",x"25",x"20",x"11", -- 0x0438
    x"25",x"1B",x"06",x"07",x"CD",x"32",x"1A",x"2A", -- 0x0440
    x"8D",x"20",x"2C",x"7D",x"FE",x"63",x"DA",x"53", -- 0x0448
    x"04",x"2E",x"54",x"22",x"8D",x"20",x"2A",x"8F", -- 0x0450
    x"20",x"2C",x"22",x"8F",x"20",x"3A",x"84",x"20", -- 0x0458
    x"A7",x"C0",x"7E",x"E6",x"01",x"01",x"29",x"02", -- 0x0460
    x"C2",x"6E",x"04",x"01",x"E0",x"FE",x"21",x"8A", -- 0x0468
    x"20",x"71",x"23",x"23",x"70",x"C9",x"E1",x"3A", -- 0x0470
    x"32",x"1B",x"32",x"32",x"20",x"2A",x"38",x"20", -- 0x0478
    x"7D",x"B4",x"C2",x"8A",x"04",x"2B",x"22",x"38", -- 0x0480
    x"20",x"C9",x"11",x"35",x"20",x"3E",x"F9",x"CD", -- 0x0488
    x"50",x"05",x"3A",x"46",x"20",x"32",x"70",x"20", -- 0x0490
    x"3A",x"56",x"20",x"32",x"71",x"20",x"CD",x"63", -- 0x0498
    x"05",x"3A",x"78",x"20",x"A7",x"21",x"35",x"20", -- 0x04A0
    x"C2",x"5B",x"05",x"11",x"30",x"1B",x"21",x"30", -- 0x04A8
    x"20",x"06",x"10",x"C3",x"32",x"1A",x"E1",x"3A", -- 0x04B0
    x"6E",x"20",x"A7",x"C0",x"3A",x"80",x"20",x"FE", -- 0x04B8
    x"01",x"C0",x"11",x"45",x"20",x"3E",x"ED",x"CD", -- 0x04C0
    x"50",x"05",x"3A",x"36",x"20",x"32",x"70",x"20", -- 0x04C8
    x"3A",x"56",x"20",x"32",x"71",x"20",x"CD",x"63", -- 0x04D0
    x"05",x"3A",x"76",x"20",x"FE",x"10",x"DA",x"E7", -- 0x04D8
    x"04",x"3A",x"48",x"1B",x"32",x"76",x"20",x"3A", -- 0x04E0
    x"78",x"20",x"A7",x"21",x"45",x"20",x"C2",x"5B", -- 0x04E8
    x"05",x"11",x"40",x"1B",x"21",x"40",x"20",x"06", -- 0x04F0
    x"10",x"CD",x"32",x"1A",x"3A",x"82",x"20",x"3D", -- 0x04F8
    x"C2",x"08",x"05",x"3E",x"01",x"32",x"6E",x"20", -- 0x0500
    x"2A",x"76",x"20",x"C3",x"7E",x"06",x"E1",x"11", -- 0x0508
    x"55",x"20",x"3E",x"DB",x"CD",x"50",x"05",x"3A", -- 0x0510
    x"46",x"20",x"32",x"70",x"20",x"3A",x"36",x"20", -- 0x0518
    x"32",x"71",x"20",x"CD",x"63",x"05",x"3A",x"76", -- 0x0520
    x"20",x"FE",x"15",x"DA",x"34",x"05",x"3A",x"58", -- 0x0528
    x"1B",x"32",x"76",x"20",x"3A",x"78",x"20",x"A7", -- 0x0530
    x"21",x"55",x"20",x"C2",x"5B",x"05",x"11",x"50", -- 0x0538
    x"1B",x"21",x"50",x"20",x"06",x"10",x"CD",x"32", -- 0x0540
    x"1A",x"2A",x"76",x"20",x"22",x"58",x"20",x"C9", -- 0x0548
    x"32",x"7F",x"20",x"21",x"73",x"20",x"06",x"0B", -- 0x0550
    x"C3",x"32",x"1A",x"11",x"73",x"20",x"06",x"0B", -- 0x0558
    x"C3",x"32",x"1A",x"21",x"73",x"20",x"7E",x"E6", -- 0x0560
    x"80",x"C2",x"C1",x"05",x"3A",x"C1",x"20",x"FE", -- 0x0568
    x"04",x"3A",x"69",x"20",x"CA",x"B7",x"05",x"A7", -- 0x0570
    x"C8",x"23",x"36",x"00",x"3A",x"70",x"20",x"A7", -- 0x0578
    x"CA",x"89",x"05",x"47",x"3A",x"CF",x"20",x"B8", -- 0x0580
    x"D0",x"3A",x"71",x"20",x"A7",x"CA",x"96",x"05", -- 0x0588
    x"47",x"3A",x"CF",x"20",x"B8",x"D0",x"23",x"7E", -- 0x0590
    x"A7",x"CA",x"1B",x"06",x"2A",x"76",x"20",x"4E", -- 0x0598
    x"23",x"00",x"22",x"76",x"20",x"CD",x"2F",x"06", -- 0x05A0
    x"D0",x"CD",x"7A",x"01",x"79",x"C6",x"07",x"67", -- 0x05A8
    x"7D",x"D6",x"0A",x"6F",x"22",x"7B",x"20",x"21", -- 0x05B0
    x"73",x"20",x"7E",x"F6",x"80",x"77",x"23",x"34", -- 0x05B8
    x"C9",x"11",x"7C",x"20",x"CD",x"06",x"1A",x"D0", -- 0x05C0
    x"23",x"7E",x"E6",x"01",x"C2",x"44",x"06",x"23", -- 0x05C8
    x"34",x"CD",x"75",x"06",x"3A",x"79",x"20",x"C6", -- 0x05D0
    x"03",x"21",x"7F",x"20",x"BE",x"DA",x"E2",x"05", -- 0x05D8
    x"D6",x"0C",x"32",x"79",x"20",x"3A",x"7B",x"20", -- 0x05E0
    x"47",x"3A",x"7E",x"20",x"80",x"32",x"7B",x"20", -- 0x05E8
    x"CD",x"6C",x"06",x"3A",x"7B",x"20",x"FE",x"15", -- 0x05F0
    x"DA",x"12",x"06",x"3A",x"61",x"20",x"A7",x"C8", -- 0x05F8
    x"3A",x"7B",x"20",x"FE",x"1E",x"DA",x"12",x"06", -- 0x0600
    x"FE",x"27",x"00",x"D2",x"12",x"06",x"97",x"32", -- 0x0608
    x"15",x"20",x"3A",x"73",x"20",x"F6",x"01",x"32", -- 0x0610
    x"73",x"20",x"C9",x"3A",x"1B",x"20",x"C6",x"08", -- 0x0618
    x"67",x"CD",x"6F",x"15",x"79",x"FE",x"0C",x"DA", -- 0x0620
    x"A5",x"05",x"0E",x"0B",x"C3",x"A5",x"05",x"0D", -- 0x0628
    x"3A",x"67",x"20",x"67",x"69",x"16",x"05",x"7E", -- 0x0630
    x"A7",x"37",x"C0",x"7D",x"C6",x"0B",x"6F",x"15", -- 0x0638
    x"C2",x"37",x"06",x"C9",x"21",x"78",x"20",x"35", -- 0x0640
    x"7E",x"FE",x"03",x"C2",x"67",x"06",x"CD",x"75", -- 0x0648
    x"06",x"21",x"DC",x"1C",x"22",x"79",x"20",x"21", -- 0x0650
    x"7C",x"20",x"35",x"35",x"2B",x"35",x"35",x"3E", -- 0x0658
    x"06",x"32",x"7D",x"20",x"C3",x"6C",x"06",x"A7", -- 0x0660
    x"C0",x"C3",x"75",x"06",x"21",x"79",x"20",x"CD", -- 0x0668
    x"3B",x"1A",x"C3",x"91",x"14",x"21",x"79",x"20", -- 0x0670
    x"CD",x"3B",x"1A",x"C3",x"52",x"14",x"22",x"48", -- 0x0678
    x"20",x"C9",x"E1",x"3A",x"80",x"20",x"FE",x"02", -- 0x0680
    x"C0",x"21",x"83",x"20",x"7E",x"A7",x"CA",x"0F", -- 0x0688
    x"05",x"3A",x"56",x"20",x"A7",x"C2",x"0F",x"05", -- 0x0690
    x"23",x"7E",x"A7",x"C2",x"AB",x"06",x"3A",x"82", -- 0x0698
    x"20",x"FE",x"08",x"DA",x"0F",x"05",x"36",x"01", -- 0x06A0
    x"CD",x"3C",x"07",x"11",x"8A",x"20",x"CD",x"06", -- 0x06A8
    x"1A",x"D0",x"21",x"85",x"20",x"7E",x"A7",x"C2", -- 0x06B0
    x"D6",x"06",x"21",x"8A",x"20",x"7E",x"23",x"23", -- 0x06B8
    x"86",x"32",x"8A",x"20",x"CD",x"3C",x"07",x"21", -- 0x06C0
    x"8A",x"20",x"7E",x"FE",x"28",x"DA",x"F9",x"06", -- 0x06C8
    x"FE",x"E1",x"D2",x"F9",x"06",x"C9",x"06",x"FE", -- 0x06D0
    x"CD",x"DC",x"19",x"23",x"35",x"7E",x"FE",x"1F", -- 0x06D8
    x"CA",x"4B",x"07",x"FE",x"18",x"CA",x"0C",x"07", -- 0x06E0
    x"A7",x"C0",x"06",x"EF",x"21",x"98",x"20",x"7E", -- 0x06E8
    x"A0",x"77",x"E6",x"20",x"D3",x"05",x"00",x"00", -- 0x06F0
    x"00",x"CD",x"42",x"07",x"CD",x"CB",x"14",x"21", -- 0x06F8
    x"83",x"20",x"06",x"0A",x"CD",x"5F",x"07",x"06", -- 0x0700
    x"FE",x"C3",x"DC",x"19",x"3E",x"01",x"32",x"F1", -- 0x0708
    x"20",x"2A",x"8D",x"20",x"46",x"0E",x"04",x"21", -- 0x0710
    x"50",x"1D",x"11",x"4C",x"1D",x"1A",x"B8",x"CA", -- 0x0718
    x"28",x"07",x"23",x"13",x"0D",x"C2",x"1D",x"07", -- 0x0720
    x"7E",x"32",x"87",x"20",x"26",x"00",x"68",x"29", -- 0x0728
    x"29",x"29",x"29",x"22",x"F2",x"20",x"CD",x"42", -- 0x0730
    x"07",x"C3",x"F1",x"08",x"CD",x"42",x"07",x"C3", -- 0x0738
    x"39",x"14",x"21",x"87",x"20",x"CD",x"3B",x"1A", -- 0x0740
    x"C3",x"47",x"1A",x"06",x"10",x"21",x"98",x"20", -- 0x0748
    x"7E",x"B0",x"77",x"CD",x"70",x"17",x"21",x"7C", -- 0x0750
    x"1D",x"22",x"87",x"20",x"C3",x"3C",x"07",x"11", -- 0x0758
    x"83",x"1B",x"C3",x"32",x"1A",x"3E",x"01",x"32", -- 0x0760
    x"93",x"20",x"31",x"00",x"24",x"FB",x"CD",x"79", -- 0x0768
    x"19",x"CD",x"D6",x"09",x"21",x"13",x"30",x"11", -- 0x0770
    x"F3",x"1F",x"0E",x"04",x"CD",x"F3",x"08",x"3A", -- 0x0778
    x"EB",x"20",x"3D",x"21",x"10",x"28",x"0E",x"14", -- 0x0780
    x"C2",x"57",x"08",x"11",x"CF",x"1A",x"CD",x"F3", -- 0x0788
    x"08",x"DB",x"01",x"E6",x"04",x"CA",x"7F",x"07", -- 0x0790
    x"06",x"99",x"AF",x"32",x"CE",x"20",x"3A",x"EB", -- 0x0798
    x"20",x"80",x"27",x"32",x"EB",x"20",x"CD",x"47", -- 0x07A0
    x"19",x"21",x"00",x"00",x"22",x"F8",x"20",x"22", -- 0x07A8
    x"FC",x"20",x"CD",x"25",x"19",x"CD",x"2B",x"19", -- 0x07B0
    x"CD",x"D7",x"19",x"21",x"01",x"01",x"7C",x"32", -- 0x07B8
    x"EF",x"20",x"22",x"E7",x"20",x"22",x"E5",x"20", -- 0x07C0
    x"CD",x"56",x"19",x"CD",x"EF",x"01",x"CD",x"F5", -- 0x07C8
    x"01",x"CD",x"D1",x"08",x"32",x"FF",x"21",x"32", -- 0x07D0
    x"FF",x"22",x"CD",x"D7",x"00",x"AF",x"32",x"FE", -- 0x07D8
    x"21",x"32",x"FE",x"22",x"CD",x"C0",x"01",x"CD", -- 0x07E0
    x"04",x"19",x"21",x"78",x"38",x"22",x"FC",x"21", -- 0x07E8
    x"22",x"FC",x"22",x"CD",x"E4",x"01",x"CD",x"7F", -- 0x07F0
    x"1A",x"CD",x"8D",x"08",x"CD",x"D6",x"09",x"00"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
