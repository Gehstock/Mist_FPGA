library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"C6",X"C6",X"82",X"C6",X"C6",X"7C",X"00",X"00",X"00",X"FE",X"FE",X"8E",X"00",X"00",
		X"00",X"66",X"F2",X"BA",X"9E",X"8E",X"C6",X"62",X"00",X"FE",X"FE",X"92",X"92",X"82",X"C6",X"C6",
		X"00",X"18",X"FE",X"1E",X"1A",X"D8",X"F8",X"F8",X"00",X"9C",X"BE",X"B2",X"B2",X"B2",X"F6",X"F6",
		X"00",X"4C",X"DE",X"92",X"92",X"92",X"FE",X"7C",X"00",X"E0",X"F0",X"98",X"8E",X"86",X"C2",X"E0",
		X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"7C",X"FE",X"92",X"92",X"92",X"F6",X"64",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"24",X"24",X"18",X"00",X"00",
		X"3E",X"7F",X"F8",X"F8",X"F8",X"C0",X"C1",X"43",X"00",X"00",X"04",X"18",X"18",X"00",X"80",X"C0",
		X"03",X"01",X"00",X"18",X"18",X"20",X"00",X"00",X"C0",X"80",X"00",X"18",X"18",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"D6",X"D0",X"D0",X"D0",X"D6",X"7E",
		X"00",X"44",X"EE",X"BA",X"92",X"82",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"7C",X"FE",X"82",X"82",X"BA",X"FE",X"FE",X"00",X"C6",X"C6",X"92",X"92",X"92",X"FE",X"FE",
		X"00",X"C0",X"C0",X"90",X"92",X"96",X"FE",X"FE",X"00",X"6C",X"EE",X"8A",X"8A",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"D0",X"10",X"16",X"FE",X"FE",X"00",X"00",X"C6",X"FE",X"FE",X"FE",X"C6",X"00",
		X"00",X"FC",X"FE",X"C2",X"06",X"0E",X"0C",X"08",X"00",X"82",X"C6",X"EE",X"38",X"92",X"FE",X"FE",
		X"00",X"1E",X"0E",X"06",X"02",X"E2",X"FE",X"FE",X"00",X"FE",X"C6",X"60",X"30",X"60",X"C6",X"FE",
		X"00",X"FE",X"CE",X"9C",X"38",X"72",X"E6",X"FE",X"00",X"7C",X"EE",X"C6",X"C6",X"C6",X"EE",X"7C",
		X"00",X"60",X"F0",X"90",X"90",X"92",X"FE",X"FE",X"00",X"06",X"7E",X"F6",X"CE",X"C6",X"DE",X"7C",
		X"00",X"62",X"F6",X"9E",X"90",X"96",X"FE",X"FE",X"00",X"C4",X"8E",X"9A",X"9A",X"B2",X"F2",X"66",
		X"00",X"F0",X"C2",X"FE",X"FE",X"FE",X"C2",X"F0",X"00",X"FC",X"FE",X"FA",X"02",X"02",X"FE",X"FC",
		X"00",X"C0",X"F8",X"FC",X"0E",X"FC",X"F8",X"C0",X"00",X"FE",X"C6",X"0C",X"18",X"0C",X"C6",X"FE",
		X"00",X"C6",X"C6",X"28",X"10",X"28",X"C6",X"C6",X"00",X"FE",X"FE",X"D2",X"12",X"16",X"F6",X"F6",
		X"00",X"CE",X"E2",X"F2",X"BA",X"9E",X"8E",X"E6",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"06",X"0B",X"3F",X"3F",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"00",X"00",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"04",X"0C",X"00",X"00",
		X"00",X"00",X"18",X"24",X"28",X"18",X"00",X"00",X"00",X"00",X"18",X"0A",X"36",X"08",X"0C",X"00",
		X"00",X"78",X"C8",X"8C",X"A4",X"C8",X"38",X"00",X"38",X"04",X"BC",X"78",X"86",X"64",X"38",X"00",
		X"00",X"A8",X"86",X"02",X"44",X"10",X"14",X"10",X"04",X"10",X"20",X"00",X"00",X"00",X"02",X"0C",
		X"02",X"08",X"10",X"00",X"00",X"00",X"01",X"06",X"05",X"08",X"00",X"00",X"00",X"01",X"00",X"02",
		X"06",X"0E",X"1E",X"1E",X"1E",X"1E",X"0E",X"06",X"18",X"38",X"78",X"78",X"78",X"78",X"38",X"18",
		X"30",X"70",X"90",X"F0",X"F0",X"90",X"70",X"30",X"18",X"38",X"48",X"78",X"78",X"48",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F1",
		X"00",X"00",X"00",X"00",X"F1",X"11",X"1F",X"11",X"00",X"00",X"1F",X"11",X"F1",X"11",X"1F",X"11",
		X"F1",X"11",X"1F",X"11",X"F1",X"11",X"1F",X"11",X"F1",X"11",X"1F",X"11",X"F1",X"11",X"00",X"00",
		X"F1",X"11",X"1F",X"11",X"00",X"00",X"00",X"00",X"F1",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"38",X"54",X"7C",X"54",X"38",X"81",X"83",X"F0",X"08",X"E4",X"12",X"C9",X"25",X"95",X"D5",
		X"AB",X"A9",X"A4",X"93",X"48",X"27",X"10",X"0F",X"D5",X"95",X"25",X"C9",X"12",X"E4",X"08",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"03",X"01",X"06",X"0E",X"13",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"09",X"11",X"05",X"01",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"3C",X"04",X"00",X"00",X"00",X"00",
		X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"C4",X"64",X"34",X"18",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"04",X"00",X"00",X"00",X"00",
		X"11",X"30",X"04",X"0C",X"18",X"30",X"60",X"00",X"84",X"04",X"04",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"04",X"00",X"00",X"00",X"80",
		X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"04",X"04",X"88",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"01",X"03",X"03",X"02",X"10",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"40",X"81",X"05",X"0A",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"22",X"02",X"06",X"04",X"82",X"81",X"00",
		X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"01",X"01",X"0B",X"02",X"20",X"42",X"44",X"00",
		X"20",X"98",X"8B",X"7C",X"18",X"2E",X"42",X"44",X"30",X"88",X"48",X"66",X"01",X"34",X"44",X"43",
		X"30",X"08",X"08",X"7E",X"99",X"A5",X"14",X"23",X"83",X"4C",X"69",X"06",X"00",X"24",X"42",X"C1",
		X"02",X"02",X"00",X"00",X"08",X"18",X"00",X"00",X"20",X"41",X"11",X"22",X"20",X"00",X"00",X"00",
		X"00",X"00",X"20",X"40",X"02",X"04",X"00",X"00",X"01",X"03",X"41",X"50",X"2C",X"02",X"C0",X"80",
		X"08",X"09",X"05",X"00",X"00",X"30",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"85",X"08",X"02",X"03",X"00",X"00",X"00",X"0C",X"40",X"A0",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"13",X"01",X"08",X"12",X"20",X"00",X"40",X"80",X"00",X"00",X"40",X"80",X"00",
		X"00",X"40",X"01",X"02",X"0F",X"10",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"4E",X"A4",X"96",X"64",X"0E",X"1C",X"00",X"3C",X"4E",X"84",X"86",X"94",X"6E",X"1C",X"00",
		X"3C",X"4C",X"86",X"84",X"86",X"8C",X"9C",X"58",X"3C",X"4C",X"86",X"84",X"96",X"6C",X"1C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FE",
		X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F3",X"1F",X"0F",X"03",X"06",X"00",X"00",X"00",X"06",X"F8",X"E0",X"E0",X"18",
		X"06",X"03",X"0F",X"1F",X"F3",X"00",X"00",X"00",X"18",X"E0",X"E0",X"F8",X"06",X"00",X"00",X"00",
		X"80",X"63",X"37",X"1F",X"0F",X"02",X"03",X"06",X"02",X"0C",X"B8",X"F0",X"E0",X"00",X"E0",X"18",
		X"06",X"03",X"02",X"0F",X"1F",X"37",X"63",X"80",X"18",X"E0",X"00",X"E0",X"F0",X"B8",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"81",X"E1",X"81",X"E1",X"81",X"E1",X"7E",X"3C",X"42",X"72",X"42",X"72",X"42",X"72",X"3C",
		X"18",X"24",X"3C",X"24",X"3C",X"24",X"3C",X"18",X"3C",X"42",X"72",X"42",X"72",X"42",X"72",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"92",X"FF",
		X"FF",X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"B6",X"04",X"04",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"B6",X"04",X"0A",X"11",X"00",X"00",X"00",
		X"01",X"03",X"03",X"01",X"03",X"03",X"01",X"03",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"03",X"01",X"03",X"13",X"09",X"06",X"0B",X"11",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"01",X"03",X"03",X"01",X"03",X"03",X"01",X"03",X"00",X"80",X"C0",X"80",X"80",X"C0",X"80",X"80",
		X"03",X"01",X"03",X"03",X"11",X"0F",X"12",X"01",X"C0",X"80",X"80",X"C0",X"80",X"80",X"C0",X"80",
		X"00",X"1F",X"20",X"5C",X"BC",X"B0",X"B0",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"84",X"24",
		X"80",X"BC",X"B0",X"B0",X"5C",X"20",X"1F",X"00",X"84",X"24",X"04",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"5C",X"B0",X"B8",X"BC",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"84",X"24",
		X"80",X"B0",X"B8",X"BC",X"5C",X"20",X"1F",X"00",X"04",X"84",X"24",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"5C",X"A4",X"AC",X"BC",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"04",X"04",
		X"80",X"A4",X"AC",X"BC",X"5C",X"20",X"1F",X"00",X"04",X"04",X"04",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"5C",X"BC",X"AC",X"A4",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"04",X"04",
		X"80",X"BC",X"AC",X"A4",X"5C",X"20",X"1F",X"00",X"04",X"04",X"04",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"03",X"06",X"0E",X"1E",X"1E",X"3E",X"3F",X"00",X"C0",X"60",X"70",X"78",X"78",X"7C",X"FC",
		X"3F",X"3E",X"1E",X"1E",X"0E",X"06",X"03",X"00",X"FC",X"7C",X"78",X"78",X"70",X"60",X"C0",X"00",
		X"00",X"03",X"06",X"0C",X"1C",X"1C",X"3C",X"3D",X"00",X"C0",X"60",X"30",X"38",X"38",X"3C",X"BC",
		X"3D",X"3C",X"1C",X"1C",X"0C",X"06",X"03",X"00",X"BC",X"3C",X"38",X"38",X"30",X"60",X"C0",X"00",
		X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"31",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"8C",
		X"31",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"8C",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"1E",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"78",
		X"1E",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"78",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"20",X"F0",X"E0",X"60",
		X"06",X"07",X"0F",X"04",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"06",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"60",
		X"06",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"60",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"60",
		X"06",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"60",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0F",X"08",X"1A",X"18",X"1F",X"00",X"00",X"0E",X"10",X"A0",X"C0",X"C0",X"C0",
		X"18",X"1A",X"08",X"0F",X"06",X"00",X"00",X"00",X"C0",X"C0",X"A0",X"10",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"30",X"78",X"44",X"E7",X"F7",X"FF",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"C7",X"E7",X"74",X"78",X"30",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"20",X"30",X"E8",X"F6",X"78",X"38",X"18",X"F8",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"78",X"38",X"18",X"F6",X"E8",X"30",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"22",X"02",X"02",X"02",X"00",X"00",
		X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"20",X"40",X"00",X"00",X"20",X"20",
		X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"0C",X"24",X"24",
		X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"20",X"40",X"00",X"00",X"04",X"04",
		X"20",X"60",X"00",X"00",X"01",X"00",X"00",X"00",X"04",X"04",X"08",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"08",X"08",X"08",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"04",X"04",X"04",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"10",X"00",X"00",X"00",X"40",X"44",X"04",X"04",X"04",X"00",
		X"00",X"10",X"18",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"10",X"08",X"08",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"10",X"00",X"00",X"20",X"20",X"04",X"04",X"04",X"04",X"00",
		X"00",X"10",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"10",X"01",X"00",X"00",X"04",X"04",X"04",X"C4",X"40",X"FE",
		X"01",X"10",X"18",X"00",X"00",X"00",X"00",X"00",X"FE",X"40",X"C4",X"04",X"04",X"04",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
