library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity c1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of c1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CD",X"1F",X"48",X"CD",X"5C",X"48",X"CD",X"FF",X"49",X"C9",X"C3",X"58",X"49",X"C3",X"69",X"4C",
		X"C3",X"57",X"4C",X"00",X"00",X"00",X"C3",X"4C",X"4E",X"C3",X"A9",X"4A",X"C3",X"BA",X"4F",X"3A",
		X"12",X"20",X"E6",X"01",X"C8",X"CD",X"98",X"4E",X"3A",X"22",X"20",X"B7",X"C8",X"21",X"C4",X"21",
		X"AF",X"BE",X"C2",X"53",X"48",X"3A",X"F6",X"22",X"21",X"CF",X"22",X"B6",X"C0",X"2B",X"DB",X"00",
		X"E6",X"40",X"CA",X"4A",X"48",X"7E",X"B7",X"C8",X"35",X"C9",X"7E",X"B7",X"C0",X"36",X"01",X"CD",
		X"DE",X"4B",X"C9",X"23",X"23",X"BE",X"C8",X"77",X"CD",X"DE",X"4B",X"C9",X"3A",X"CF",X"22",X"B7",
		X"C8",X"21",X"0E",X"22",X"22",X"00",X"23",X"2A",X"02",X"22",X"11",X"10",X"22",X"CD",X"AA",X"49",
		X"DA",X"67",X"4B",X"21",X"2E",X"22",X"22",X"00",X"23",X"2A",X"22",X"22",X"11",X"30",X"22",X"CD",
		X"AA",X"49",X"DA",X"67",X"4B",X"21",X"4E",X"22",X"22",X"00",X"23",X"2A",X"42",X"22",X"11",X"50",
		X"22",X"CD",X"AA",X"49",X"DA",X"67",X"4B",X"21",X"6E",X"22",X"22",X"00",X"23",X"2A",X"62",X"22",
		X"11",X"70",X"22",X"CD",X"AA",X"49",X"DA",X"67",X"4B",X"21",X"D2",X"22",X"22",X"00",X"23",X"2A",
		X"D2",X"22",X"11",X"DF",X"22",X"CD",X"C2",X"49",X"DA",X"D3",X"49",X"21",X"E2",X"22",X"22",X"00",
		X"23",X"2A",X"E2",X"22",X"11",X"EF",X"22",X"CD",X"C2",X"49",X"DA",X"D3",X"49",X"21",X"8E",X"22",
		X"22",X"00",X"23",X"2A",X"82",X"22",X"11",X"90",X"22",X"CD",X"95",X"49",X"DA",X"F6",X"4A",X"21",
		X"AE",X"22",X"22",X"00",X"23",X"2A",X"A2",X"22",X"11",X"B0",X"22",X"CD",X"95",X"49",X"DA",X"F6",
		X"4A",X"CD",X"F8",X"48",X"DA",X"28",X"49",X"C9",X"3A",X"E3",X"21",X"FE",X"03",X"CA",X"07",X"49",
		X"FE",X"04",X"CA",X"07",X"49",X"B7",X"C9",X"21",X"C3",X"22",X"3A",X"E5",X"21",X"57",X"47",X"FE",
		X"0A",X"DA",X"16",X"49",X"16",X"0A",X"3A",X"0A",X"20",X"C6",X"11",X"90",X"82",X"42",X"57",X"1E",
		X"80",X"0E",X"0F",X"C3",X"B8",X"49",X"00",X"10",X"21",X"00",X"00",X"22",X"C2",X"22",X"CD",X"3C",
		X"49",X"3E",X"05",X"32",X"E3",X"21",X"21",X"E6",X"21",X"36",X"20",X"C9",X"3A",X"54",X"23",X"C6",
		X"07",X"D6",X"82",X"0F",X"0F",X"0F",X"E6",X"0F",X"67",X"2E",X"00",X"22",X"86",X"21",X"21",X"86",
		X"21",X"22",X"00",X"23",X"CD",X"39",X"4C",X"C9",X"3A",X"22",X"20",X"B7",X"C8",X"3A",X"6B",X"20",
		X"FE",X"C8",X"D0",X"D6",X"60",X"D2",X"6A",X"49",X"3E",X"00",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"21",X"8D",X"49",X"85",X"D2",X"78",X"49",X"24",X"6F",X"7E",X"21",X"34",X"20",X"86",X"77",X"D0",
		X"11",X"2E",X"20",X"21",X"8A",X"49",X"CD",X"10",X"48",X"C9",X"01",X"00",X"00",X"80",X"40",X"20",
		X"14",X"0C",X"08",X"06",X"04",X"1A",X"B7",X"C8",X"13",X"1A",X"B7",X"C0",X"11",X"0E",X"08",X"19",
		X"EB",X"21",X"C3",X"22",X"01",X"12",X"10",X"C3",X"B8",X"49",X"1A",X"B7",X"C8",X"11",X"07",X"0D",
		X"19",X"EB",X"21",X"C3",X"22",X"01",X"0B",X"10",X"7A",X"96",X"B8",X"D0",X"7B",X"2B",X"96",X"B9",
		X"D0",X"C9",X"1A",X"B7",X"C8",X"11",X"03",X"05",X"19",X"EB",X"21",X"C3",X"22",X"01",X"04",X"0A",
		X"C3",X"B8",X"49",X"2A",X"00",X"23",X"AF",X"77",X"23",X"77",X"21",X"00",X"00",X"22",X"C2",X"22",
		X"C9",X"1A",X"B7",X"C8",X"13",X"1A",X"B7",X"C0",X"11",X"0E",X"08",X"19",X"EB",X"21",X"6B",X"20",
		X"01",X"1E",X"18",X"C3",X"B8",X"49",X"2A",X"00",X"23",X"36",X"E8",X"CD",X"19",X"48",X"C9",X"3A",
		X"22",X"20",X"B7",X"C8",X"3A",X"4E",X"20",X"B7",X"C0",X"21",X"D3",X"22",X"22",X"00",X"23",X"2A",
		X"D2",X"22",X"11",X"DF",X"22",X"CD",X"4B",X"4B",X"DA",X"5C",X"4B",X"21",X"E3",X"22",X"22",X"00",
		X"23",X"2A",X"E2",X"22",X"11",X"EF",X"22",X"CD",X"4B",X"4B",X"DA",X"5C",X"4B",X"21",X"03",X"22",
		X"22",X"00",X"23",X"2A",X"02",X"22",X"11",X"10",X"22",X"CD",X"3A",X"4B",X"DA",X"9A",X"4A",X"21",
		X"23",X"22",X"22",X"00",X"23",X"2A",X"22",X"22",X"11",X"30",X"22",X"CD",X"3A",X"4B",X"DA",X"9A",
		X"4A",X"21",X"43",X"22",X"22",X"00",X"23",X"2A",X"42",X"22",X"11",X"50",X"22",X"CD",X"3A",X"4B",
		X"DA",X"9A",X"4A",X"21",X"63",X"22",X"22",X"00",X"23",X"2A",X"62",X"22",X"11",X"70",X"22",X"CD",
		X"3A",X"4B",X"DA",X"9A",X"4A",X"21",X"83",X"22",X"22",X"00",X"23",X"2A",X"82",X"22",X"11",X"90",
		X"22",X"CD",X"E1",X"49",X"DA",X"F6",X"49",X"21",X"A3",X"22",X"22",X"00",X"23",X"2A",X"A2",X"22",
		X"11",X"B0",X"22",X"CD",X"E1",X"49",X"DA",X"F6",X"49",X"C9",X"2A",X"00",X"23",X"36",X"E8",X"7D",
		X"C6",X"0E",X"6F",X"36",X"FF",X"CD",X"19",X"48",X"C9",X"AF",X"32",X"22",X"20",X"32",X"D9",X"20",
		X"21",X"E3",X"21",X"7E",X"FE",X"02",X"DA",X"BB",X"4A",X"36",X"07",X"3E",X"FF",X"32",X"D7",X"20",
		X"32",X"62",X"20",X"21",X"00",X"00",X"22",X"C2",X"22",X"22",X"D2",X"22",X"22",X"E2",X"22",X"3E",
		X"10",X"32",X"C2",X"21",X"11",X"C0",X"21",X"21",X"71",X"20",X"36",X"FE",X"3A",X"6A",X"20",X"21",
		X"6E",X"20",X"FE",X"78",X"DA",X"EF",X"4A",X"36",X"FE",X"3E",X"FF",X"12",X"1B",X"12",X"C9",X"36",
		X"02",X"AF",X"12",X"1B",X"12",X"C9",X"21",X"00",X"00",X"22",X"C2",X"22",X"CD",X"39",X"4C",X"2A",
		X"00",X"23",X"E5",X"23",X"23",X"23",X"36",X"FF",X"E1",X"2B",X"E5",X"CD",X"29",X"4B",X"E1",X"11",
		X"40",X"12",X"72",X"2B",X"73",X"2B",X"2B",X"2B",X"36",X"00",X"2B",X"2B",X"2B",X"36",X"00",X"7D",
		X"C6",X"10",X"6F",X"36",X"10",X"CD",X"C0",X"4B",X"C9",X"46",X"2B",X"4E",X"7D",X"C6",X"07",X"6F",
		X"3E",X"FF",X"BE",X"C8",X"77",X"23",X"71",X"23",X"70",X"C9",X"1A",X"B7",X"C8",X"11",X"06",X"0D",
		X"19",X"EB",X"21",X"6B",X"20",X"01",X"16",X"1D",X"C3",X"B8",X"49",X"1A",X"B7",X"C8",X"11",X"03",
		X"05",X"19",X"EB",X"21",X"6B",X"20",X"01",X"13",X"15",X"C3",X"B8",X"49",X"2A",X"00",X"23",X"AF",
		X"77",X"2B",X"77",X"CD",X"19",X"48",X"C9",X"21",X"00",X"00",X"22",X"C2",X"22",X"CD",X"39",X"4C",
		X"2A",X"00",X"23",X"23",X"23",X"23",X"3E",X"FF",X"BE",X"CA",X"B3",X"4B",X"77",X"2B",X"2B",X"2B",
		X"2B",X"E5",X"CD",X"29",X"4B",X"E1",X"11",X"00",X"40",X"72",X"2B",X"73",X"2B",X"00",X"00",X"2B",
		X"36",X"E0",X"2B",X"36",X"FC",X"2B",X"36",X"01",X"2B",X"36",X"01",X"2B",X"7E",X"FE",X"80",X"D2",
		X"AE",X"4B",X"36",X"04",X"2B",X"36",X"01",X"2B",X"36",X"01",X"CD",X"C0",X"4B",X"C9",X"36",X"FC",
		X"C3",X"A4",X"4B",X"7D",X"D6",X"0E",X"6F",X"36",X"D0",X"2B",X"36",X"00",X"CD",X"C0",X"4B",X"C9",
		X"21",X"A6",X"21",X"36",X"FF",X"23",X"7E",X"B7",X"C2",X"D1",X"4B",X"36",X"01",X"23",X"36",X"01",
		X"C9",X"36",X"08",X"23",X"36",X"04",X"3A",X"A1",X"21",X"7E",X"E6",X"EF",X"77",X"C9",X"2A",X"6A",
		X"20",X"01",X"06",X"02",X"11",X"C0",X"22",X"CD",X"20",X"4C",X"7E",X"32",X"C4",X"22",X"23",X"7E",
		X"32",X"C6",X"22",X"21",X"C9",X"22",X"36",X"FC",X"21",X"CF",X"22",X"36",X"FF",X"3A",X"6B",X"20",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"21",X"1C",X"4E",X"85",X"D2",X"0E",X"4C",X"24",X"6F",X"7E",
		X"32",X"CB",X"22",X"21",X"A1",X"21",X"7E",X"F6",X"20",X"77",X"21",X"A3",X"21",X"36",X"01",X"C9",
		X"09",X"EB",X"73",X"23",X"72",X"23",X"73",X"23",X"72",X"2B",X"7E",X"EB",X"CD",X"A7",X"4D",X"21",
		X"2C",X"4E",X"85",X"D2",X"37",X"4C",X"24",X"6F",X"C9",X"3A",X"01",X"20",X"B7",X"C0",X"2A",X"00",
		X"23",X"11",X"86",X"21",X"7E",X"12",X"23",X"13",X"7E",X"12",X"AF",X"13",X"12",X"21",X"86",X"21",
		X"11",X"28",X"20",X"CD",X"10",X"48",X"C9",X"B7",X"1A",X"86",X"27",X"12",X"13",X"23",X"1A",X"8E",
		X"27",X"12",X"13",X"23",X"1A",X"8E",X"27",X"12",X"C9",X"3A",X"22",X"20",X"B7",X"C8",X"3A",X"12",
		X"20",X"E6",X"01",X"CA",X"92",X"4C",X"C3",X"79",X"4C",X"21",X"F2",X"22",X"7E",X"B7",X"CA",X"70",
		X"4D",X"3A",X"12",X"20",X"E6",X"06",X"C0",X"EB",X"21",X"EE",X"22",X"7E",X"23",X"B6",X"C0",X"EB",
		X"EF",X"C9",X"21",X"F1",X"22",X"7E",X"B7",X"CA",X"CA",X"4C",X"3A",X"12",X"20",X"E6",X"06",X"C0",
		X"EB",X"21",X"DE",X"22",X"7E",X"23",X"B6",X"C0",X"EB",X"EF",X"C9",X"01",X"16",X"4E",X"3A",X"39",
		X"20",X"FE",X"AA",X"CC",X"C7",X"4C",X"FE",X"00",X"CC",X"C7",X"4C",X"3A",X"8C",X"21",X"81",X"D2",
		X"C3",X"4C",X"04",X"4F",X"0A",X"77",X"C9",X"03",X"03",X"C9",X"22",X"F1",X"21",X"3A",X"F3",X"22",
		X"B7",X"CD",X"8B",X"4D",X"11",X"D2",X"22",X"21",X"30",X"22",X"7E",X"B7",X"CA",X"97",X"4D",X"2F",
		X"23",X"B6",X"C0",X"21",X"23",X"22",X"3A",X"6B",X"20",X"D6",X"20",X"96",X"D8",X"D6",X"0A",X"47",
		X"2B",X"7E",X"FE",X"78",X"DA",X"5D",X"4D",X"CD",X"D2",X"4D",X"86",X"D8",X"4F",X"3A",X"6A",X"20",
		X"C6",X"10",X"91",X"D8",X"FE",X"10",X"D0",X"7E",X"C6",X"03",X"4F",X"12",X"1B",X"1B",X"12",X"23",
		X"13",X"7E",X"C6",X"0A",X"12",X"13",X"13",X"12",X"79",X"CD",X"BC",X"4D",X"21",X"F6",X"4D",X"85",
		X"D2",X"24",X"4D",X"24",X"6F",X"13",X"7E",X"12",X"13",X"13",X"26",X"01",X"79",X"FE",X"80",X"D2",
		X"34",X"4D",X"26",X"FF",X"3A",X"F5",X"22",X"B7",X"7C",X"CA",X"3D",X"4D",X"84",X"12",X"7B",X"C6",
		X"09",X"5F",X"3E",X"FF",X"12",X"2A",X"F1",X"21",X"CD",X"AB",X"4C",X"3E",X"10",X"32",X"A4",X"21",
		X"21",X"A2",X"21",X"7E",X"E6",X"FD",X"77",X"21",X"A5",X"21",X"36",X"00",X"C9",X"CD",X"D2",X"4D",
		X"4F",X"7E",X"91",X"D8",X"4F",X"3A",X"6A",X"20",X"91",X"D0",X"FE",X"F0",X"D8",X"C3",X"07",X"4D",
		X"22",X"F1",X"21",X"3A",X"F4",X"22",X"B7",X"CD",X"8B",X"4D",X"21",X"50",X"22",X"7E",X"2F",X"23",
		X"B6",X"C0",X"21",X"43",X"22",X"11",X"E2",X"22",X"C3",X"E6",X"4C",X"3E",X"FF",X"32",X"F5",X"22",
		X"C0",X"3E",X"00",X"32",X"F5",X"22",X"C9",X"3A",X"B0",X"22",X"B7",X"C8",X"C3",X"DF",X"4F",X"3A",
		X"6B",X"20",X"D6",X"10",X"C3",X"EB",X"4C",X"FE",X"38",X"D2",X"AE",X"4D",X"3E",X"38",X"FE",X"B7",
		X"DA",X"B5",X"4D",X"3E",X"B7",X"D6",X"38",X"0F",X"0F",X"E6",X"1E",X"C9",X"FE",X"40",X"D2",X"C3",
		X"4D",X"3E",X"40",X"FE",X"BF",X"DA",X"CA",X"4D",X"3E",X"BF",X"D6",X"40",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"C9",X"D5",X"7E",X"C6",X"03",X"CD",X"BC",X"4D",X"11",X"06",X"4E",X"83",X"D2",X"E1",X"4D",
		X"14",X"5F",X"1A",X"57",X"78",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"0E",X"04",X"AF",X"92",X"82",
		X"0D",X"C2",X"EF",X"4D",X"D1",X"C9",X"01",X"01",X"01",X"01",X"02",X"03",X"04",X"08",X"08",X"04",
		X"03",X"02",X"01",X"01",X"01",X"01",X"10",X"10",X"10",X"08",X"06",X"04",X"02",X"02",X"04",X"05",
		X"06",X"07",X"08",X"40",X"40",X"40",X"08",X"04",X"02",X"01",X"01",X"01",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"38",X"40",X"48",X"50",X"58",X"60",X"68",X"70",X"78",X"01",X"02",X"03",X"05",
		X"02",X"03",X"03",X"04",X"01",X"01",X"02",X"01",X"04",X"01",X"08",X"01",X"08",X"FF",X"04",X"FF",
		X"02",X"FF",X"01",X"FF",X"03",X"FC",X"02",X"FD",X"03",X"FB",X"01",X"FE",X"CD",X"71",X"4E",X"CD",
		X"A6",X"4E",X"CD",X"91",X"4F",X"3A",X"12",X"20",X"07",X"E6",X"06",X"21",X"69",X"4E",X"85",X"D2",
		X"63",X"4E",X"24",X"6F",X"5E",X"23",X"56",X"EB",X"E9",X"F5",X"4E",X"4D",X"4F",X"67",X"4F",X"90",
		X"4F",X"3A",X"12",X"20",X"E6",X"07",X"C0",X"3A",X"6B",X"20",X"FE",X"CF",X"DA",X"81",X"4E",X"3E",
		X"CF",X"D6",X"50",X"D2",X"88",X"4E",X"3E",X"00",X"0F",X"0F",X"0F",X"2F",X"E6",X"0F",X"47",X"21",
		X"A1",X"21",X"7E",X"E6",X"F0",X"B0",X"77",X"C9",X"21",X"A3",X"21",X"EF",X"C0",X"3A",X"A1",X"21",
		X"E6",X"DF",X"32",X"A1",X"21",X"C9",X"3A",X"12",X"20",X"E6",X"01",X"C0",X"3A",X"DF",X"22",X"21",
		X"EF",X"22",X"B6",X"CA",X"D6",X"4E",X"21",X"A4",X"21",X"7E",X"B7",X"C8",X"23",X"EF",X"C0",X"2B",
		X"35",X"7E",X"11",X"E5",X"4E",X"83",X"D2",X"CA",X"4E",X"14",X"5F",X"1A",X"23",X"77",X"21",X"A2",
		X"21",X"7E",X"EE",X"02",X"77",X"C9",X"AF",X"32",X"A4",X"21",X"32",X"A5",X"21",X"21",X"A2",X"21",
		X"7E",X"E6",X"FD",X"77",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",
		X"05",X"00",X"03",X"00",X"02",X"11",X"A1",X"21",X"01",X"A2",X"21",X"21",X"A6",X"21",X"7E",X"B7",
		X"C8",X"23",X"EF",X"D2",X"19",X"4F",X"0A",X"E6",X"0C",X"C2",X"15",X"4F",X"0A",X"F6",X"0C",X"02",
		X"36",X"08",X"C3",X"19",X"4F",X"0A",X"E6",X"F3",X"02",X"23",X"EF",X"DA",X"26",X"4F",X"C0",X"2B",
		X"B6",X"C0",X"2B",X"36",X"00",X"C9",X"1A",X"E6",X"10",X"C2",X"3B",X"4F",X"1A",X"F6",X"10",X"12",
		X"3A",X"A0",X"21",X"F6",X"04",X"32",X"A0",X"21",X"36",X"04",X"C9",X"1A",X"E6",X"EF",X"12",X"3A",
		X"22",X"20",X"B7",X"C8",X"3A",X"A0",X"21",X"E6",X"FB",X"32",X"A0",X"21",X"C9",X"21",X"A0",X"21",
		X"3A",X"22",X"20",X"B7",X"CA",X"62",X"4F",X"3A",X"A1",X"21",X"E6",X"10",X"C0",X"7E",X"E6",X"FB",
		X"77",X"C9",X"7E",X"F6",X"04",X"77",X"C9",X"21",X"AD",X"21",X"3A",X"43",X"20",X"E6",X"08",X"C2",
		X"81",X"4F",X"36",X"02",X"21",X"A0",X"21",X"7E",X"F6",X"04",X"77",X"23",X"7E",X"F6",X"1F",X"77",
		X"C9",X"EF",X"D0",X"21",X"A0",X"21",X"7E",X"E6",X"FB",X"77",X"23",X"7E",X"E6",X"E0",X"77",X"C9",
		X"C9",X"11",X"A2",X"21",X"1A",X"E6",X"DF",X"12",X"CD",X"A1",X"4F",X"C8",X"1A",X"F6",X"20",X"12",
		X"C9",X"3A",X"EC",X"21",X"FE",X"FF",X"C0",X"3A",X"E3",X"21",X"FE",X"01",X"C8",X"FE",X"02",X"C8",
		X"FE",X"03",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"3A",X"12",X"20",X"E6",X"03",X"C0",
		X"01",X"A2",X"21",X"21",X"A7",X"21",X"EF",X"7E",X"FE",X"08",X"D0",X"0A",X"E6",X"08",X"C2",X"D8",
		X"4F",X"0A",X"F6",X"08",X"02",X"36",X"10",X"C9",X"0A",X"E6",X"F7",X"02",X"36",X"35",X"C9",X"3A",
		X"B1",X"22",X"B7",X"C0",X"21",X"A3",X"22",X"C3",X"9F",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
