library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_sound is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7E",X"F0",X"32",X"7E",X"F0",X"11",X"7E",X"F0",X"09",X"7C",X"00",X"8F",X"86",X"00",X"97",X"BF",
		X"3B",X"B7",X"90",X"00",X"86",X"0D",X"97",X"03",X"C6",X"0E",X"D7",X"02",X"C6",X"0C",X"4F",X"97",
		X"03",X"97",X"00",X"D7",X"03",X"96",X"02",X"5F",X"D7",X"03",X"5A",X"D7",X"00",X"84",X"1F",X"97",
		X"90",X"3B",X"8E",X"00",X"FF",X"0F",X"CE",X"FF",X"FF",X"FF",X"00",X"00",X"BD",X"F0",X"42",X"7E",
		X"F0",X"7A",X"CC",X"00",X"20",X"BD",X"F0",X"4C",X"5A",X"2A",X"FA",X"39",X"37",X"36",X"C1",X"10",
		X"2A",X"19",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"08",X"D7",X"03",X"5C",X"32",X"97",X"02",
		X"A5",X"00",X"A5",X"00",X"D7",X"03",X"5A",X"D7",X"03",X"33",X"39",X"86",X"15",X"97",X"03",X"C4",
		X"0F",X"D7",X"02",X"C6",X"10",X"20",X"E3",X"7E",X"F1",X"20",X"CE",X"00",X"80",X"CC",X"00",X"60",
		X"A7",X"00",X"08",X"5A",X"2A",X"FA",X"86",X"BF",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"0E",
		X"96",X"90",X"27",X"E3",X"C6",X"00",X"D7",X"90",X"81",X"01",X"26",X"05",X"BD",X"F2",X"06",X"20",
		X"D6",X"81",X"05",X"26",X"05",X"BD",X"F2",X"88",X"20",X"CD",X"81",X"02",X"26",X"05",X"BD",X"F5",
		X"16",X"20",X"C4",X"81",X"07",X"27",X"04",X"81",X"04",X"26",X"05",X"BD",X"F3",X"83",X"20",X"B7",
		X"81",X"0B",X"27",X"EA",X"81",X"08",X"26",X"05",X"BD",X"F4",X"04",X"20",X"53",X"81",X"09",X"26",
		X"05",X"BD",X"F4",X"8D",X"20",X"4A",X"81",X"03",X"26",X"05",X"BD",X"F3",X"02",X"20",X"41",X"81",
		X"06",X"26",X"05",X"BD",X"F5",X"97",X"20",X"38",X"81",X"10",X"26",X"17",X"96",X"C9",X"81",X"00",
		X"26",X"11",X"86",X"01",X"97",X"C9",X"86",X"FC",X"97",X"C2",X"BD",X"F5",X"D1",X"BD",X"F8",X"4D",
		X"7E",X"F1",X"20",X"81",X"11",X"26",X"16",X"CC",X"00",X"18",X"BD",X"F0",X"4C",X"CC",X"00",X"19",
		X"BD",X"F0",X"4C",X"CC",X"00",X"1A",X"BD",X"F0",X"4C",X"86",X"00",X"97",X"C9",X"BD",X"F8",X"C0",
		X"96",X"BF",X"26",X"1D",X"0F",X"BD",X"F1",X"BD",X"BD",X"F2",X"40",X"BD",X"F2",X"B6",X"BD",X"F3",
		X"3C",X"BD",X"F3",X"BD",X"BD",X"F4",X"3E",X"BD",X"F4",X"C7",X"BD",X"F5",X"50",X"7C",X"00",X"BF",
		X"0E",X"96",X"8F",X"8B",X"FC",X"24",X"37",X"86",X"00",X"B7",X"00",X"8F",X"0F",X"BD",X"F6",X"08",
		X"BD",X"F8",X"4A",X"0E",X"7E",X"F0",X"90",X"BD",X"F2",X"06",X"96",X"81",X"26",X"FC",X"BD",X"F1",
		X"81",X"BD",X"F2",X"88",X"96",X"87",X"26",X"FC",X"BD",X"F1",X"81",X"BD",X"F2",X"AE",X"96",X"87",
		X"26",X"FC",X"BD",X"F1",X"81",X"7E",X"F0",X"90",X"BD",X"F2",X"06",X"7E",X"F1",X"5A",X"7E",X"F0",
		X"90",X"CC",X"20",X"00",X"5A",X"26",X"FD",X"4A",X"26",X"FA",X"39",X"D6",X"8B",X"5C",X"86",X"F0",
		X"DD",X"8D",X"DE",X"8D",X"A6",X"00",X"9B",X"8C",X"97",X"8C",X"9B",X"8B",X"97",X"8B",X"39",X"0F",
		X"0F",X"0E",X"0E",X"0D",X"0D",X"0C",X"0C",X"0B",X"0B",X"0A",X"0A",X"09",X"09",X"08",X"08",X"07",
		X"07",X"06",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"96",X"81",X"26",
		X"01",X"39",X"7A",X"00",X"84",X"27",X"01",X"39",X"86",X"02",X"97",X"84",X"DC",X"82",X"C3",X"00",
		X"03",X"DD",X"82",X"96",X"83",X"C6",X"00",X"96",X"83",X"BD",X"F0",X"4C",X"C6",X"01",X"96",X"82",
		X"BD",X"F0",X"4C",X"7A",X"00",X"85",X"26",X"DF",X"86",X"00",X"97",X"81",X"97",X"82",X"97",X"83",
		X"97",X"84",X"97",X"85",X"96",X"80",X"8A",X"01",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",
		X"00",X"08",X"BD",X"F0",X"4C",X"39",X"CC",X"00",X"08",X"BD",X"F0",X"4C",X"86",X"01",X"97",X"81",
		X"CC",X"00",X"10",X"DD",X"82",X"86",X"04",X"97",X"84",X"86",X"00",X"97",X"85",X"96",X"80",X"84",
		X"FE",X"8A",X"08",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"C6",X"00",X"96",X"83",X"BD",X"F0",
		X"4C",X"C6",X"01",X"96",X"82",X"BD",X"F0",X"4C",X"C6",X"08",X"86",X"0F",X"BD",X"F0",X"4C",X"39",
		X"96",X"87",X"26",X"01",X"39",X"7A",X"00",X"8A",X"26",X"FA",X"86",X"80",X"97",X"8A",X"7C",X"00",
		X"89",X"96",X"89",X"81",X"20",X"26",X"1C",X"86",X"00",X"97",X"87",X"97",X"88",X"97",X"89",X"97",
		X"8A",X"96",X"80",X"8A",X"12",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"86",X"00",X"C6",X"09",
		X"7E",X"F0",X"4C",X"96",X"89",X"C6",X"06",X"BD",X"F8",X"80",X"D6",X"89",X"CE",X"F1",X"9F",X"3A",
		X"A6",X"00",X"C6",X"09",X"BD",X"F0",X"4C",X"39",X"CC",X"00",X"06",X"BD",X"F0",X"4C",X"96",X"80",
		X"84",X"EF",X"8A",X"02",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",X"0F",X"09",X"BD",X"F0",
		X"4C",X"86",X"01",X"97",X"87",X"86",X"00",X"97",X"89",X"86",X"20",X"97",X"8A",X"39",X"BD",X"F2",
		X"88",X"86",X"08",X"97",X"89",X"39",X"96",X"91",X"26",X"01",X"39",X"7A",X"00",X"94",X"27",X"01",
		X"39",X"86",X"05",X"97",X"94",X"DC",X"92",X"83",X"00",X"01",X"DD",X"92",X"BD",X"F1",X"8B",X"84",
		X"3F",X"9B",X"93",X"C6",X"04",X"BD",X"F0",X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",X"4C",X"7A",
		X"00",X"95",X"26",X"DC",X"86",X"00",X"97",X"91",X"97",X"92",X"97",X"93",X"97",X"94",X"97",X"95",
		X"96",X"80",X"8A",X"04",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",X"00",X"0A",X"BD",X"F0",
		X"4C",X"39",X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"86",X"01",X"97",X"91",X"CC",X"01",X"00",X"DD",
		X"92",X"86",X"04",X"97",X"94",X"86",X"D0",X"97",X"95",X"96",X"80",X"84",X"FB",X"8A",X"20",X"97",
		X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"C6",X"04",X"96",X"93",X"BD",X"F0",X"4C",X"C6",X"05",X"96",
		X"92",X"BD",X"F0",X"4C",X"C6",X"0A",X"86",X"0F",X"BD",X"F0",X"4C",X"39",X"96",X"96",X"26",X"01",
		X"39",X"7A",X"00",X"94",X"27",X"01",X"39",X"86",X"10",X"97",X"94",X"DC",X"92",X"83",X"00",X"04",
		X"DD",X"92",X"96",X"93",X"C6",X"04",X"BD",X"F0",X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",X"4C",
		X"7A",X"00",X"95",X"26",X"E1",X"86",X"00",X"97",X"96",X"97",X"92",X"97",X"93",X"97",X"94",X"97",
		X"95",X"96",X"80",X"8A",X"04",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",X"00",X"0A",X"BD",
		X"F0",X"4C",X"39",X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"86",X"01",X"97",X"96",X"CC",X"01",X"80",
		X"DD",X"92",X"86",X"04",X"97",X"94",X"86",X"80",X"97",X"95",X"96",X"80",X"84",X"FB",X"8A",X"20",
		X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"C6",X"04",X"96",X"93",X"BD",X"F0",X"4C",X"C6",X"05",
		X"96",X"92",X"BD",X"F0",X"4C",X"C6",X"0A",X"86",X"0F",X"BD",X"F0",X"4C",X"39",X"96",X"97",X"26",
		X"01",X"39",X"7A",X"00",X"94",X"27",X"01",X"39",X"86",X"02",X"97",X"94",X"DC",X"92",X"C3",X"00",
		X"08",X"DD",X"92",X"96",X"93",X"C6",X"04",X"BD",X"F0",X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",
		X"4C",X"7A",X"00",X"95",X"26",X"E1",X"86",X"00",X"97",X"97",X"97",X"92",X"97",X"93",X"97",X"94",
		X"97",X"95",X"96",X"80",X"8A",X"04",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",X"00",X"0A",
		X"BD",X"F0",X"4C",X"39",X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"86",X"01",X"97",X"97",X"CC",X"00",
		X"01",X"DD",X"92",X"86",X"04",X"97",X"94",X"86",X"00",X"97",X"95",X"96",X"80",X"84",X"FB",X"8A",
		X"20",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"C6",X"04",X"96",X"93",X"BD",X"F0",X"4C",X"C6",
		X"05",X"96",X"92",X"BD",X"F0",X"4C",X"C6",X"0A",X"86",X"0F",X"BD",X"F0",X"4C",X"39",X"96",X"98",
		X"26",X"01",X"39",X"7A",X"00",X"94",X"27",X"01",X"39",X"86",X"08",X"97",X"94",X"DC",X"92",X"C3",
		X"00",X"08",X"DD",X"92",X"96",X"93",X"D6",X"95",X"C4",X"08",X"27",X"02",X"88",X"FF",X"C6",X"04",
		X"BD",X"F0",X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",X"4C",X"7A",X"00",X"95",X"26",X"D9",X"86",
		X"00",X"97",X"98",X"97",X"92",X"97",X"93",X"97",X"94",X"97",X"95",X"96",X"80",X"8A",X"04",X"97",
		X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"39",X"CC",X"00",X"0A",
		X"BD",X"F0",X"4C",X"86",X"01",X"97",X"98",X"CC",X"00",X"01",X"DD",X"92",X"86",X"04",X"97",X"94",
		X"86",X"80",X"97",X"95",X"96",X"80",X"84",X"FB",X"8A",X"20",X"97",X"80",X"C6",X"07",X"BD",X"F0",
		X"4C",X"C6",X"04",X"96",X"93",X"BD",X"F0",X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",X"4C",X"C6",
		X"0A",X"86",X"0F",X"BD",X"F0",X"4C",X"39",X"96",X"99",X"26",X"01",X"39",X"7A",X"00",X"94",X"27",
		X"01",X"39",X"86",X"0B",X"97",X"94",X"DC",X"92",X"83",X"00",X"01",X"DD",X"92",X"96",X"93",X"D6",
		X"95",X"C4",X"08",X"26",X"02",X"88",X"FF",X"C6",X"04",X"BD",X"F0",X"4C",X"C6",X"05",X"96",X"92",
		X"BD",X"F0",X"4C",X"7A",X"00",X"95",X"26",X"D9",X"86",X"00",X"97",X"99",X"97",X"92",X"97",X"93",
		X"97",X"94",X"97",X"95",X"96",X"80",X"8A",X"04",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"CC",
		X"00",X"0A",X"BD",X"F0",X"4C",X"39",X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"86",X"01",X"97",X"99",
		X"CC",X"01",X"00",X"DD",X"92",X"86",X"04",X"97",X"94",X"86",X"58",X"97",X"95",X"96",X"80",X"84",
		X"FB",X"8A",X"20",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"C6",X"04",X"96",X"93",X"BD",X"F0",
		X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",X"4C",X"C6",X"0A",X"86",X"0F",X"BD",X"F0",X"4C",X"39",
		X"96",X"9A",X"26",X"01",X"39",X"7A",X"00",X"94",X"27",X"01",X"39",X"86",X"10",X"97",X"94",X"DC",
		X"92",X"C3",X"00",X"04",X"DD",X"92",X"96",X"93",X"C6",X"04",X"BD",X"F0",X"4C",X"C6",X"05",X"96",
		X"92",X"BD",X"F0",X"4C",X"7A",X"00",X"95",X"26",X"E1",X"86",X"00",X"97",X"9A",X"97",X"92",X"97",
		X"93",X"97",X"94",X"97",X"95",X"96",X"80",X"8A",X"04",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",
		X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"39",X"CC",X"00",X"0A",X"BD",X"F0",X"4C",X"86",X"01",X"97",
		X"9A",X"CC",X"01",X"00",X"DD",X"92",X"86",X"04",X"97",X"94",X"86",X"50",X"97",X"95",X"96",X"80",
		X"84",X"FB",X"8A",X"20",X"97",X"80",X"C6",X"07",X"BD",X"F0",X"4C",X"C6",X"04",X"96",X"93",X"BD",
		X"F0",X"4C",X"C6",X"05",X"96",X"92",X"BD",X"F0",X"4C",X"C6",X"0A",X"86",X"0F",X"BD",X"F0",X"4C",
		X"39",X"CC",X"FC",X"17",X"BD",X"F0",X"4C",X"86",X"00",X"97",X"A0",X"97",X"A1",X"97",X"A2",X"97",
		X"A3",X"97",X"A4",X"97",X"A6",X"CE",X"00",X"A0",X"86",X"FD",X"97",X"C2",X"BD",X"F6",X"A5",X"86",
		X"00",X"97",X"A8",X"97",X"A9",X"97",X"AA",X"97",X"AB",X"97",X"AC",X"97",X"AD",X"CE",X"00",X"A8",
		X"86",X"FC",X"97",X"C2",X"BD",X"F6",X"A5",X"39",X"7A",X"00",X"CC",X"26",X"0B",X"86",X"08",X"97",
		X"CC",X"BD",X"F8",X"0E",X"96",X"C9",X"26",X"01",X"39",X"CE",X"00",X"A0",X"86",X"FD",X"97",X"C2",
		X"BD",X"F6",X"9C",X"CE",X"00",X"A8",X"86",X"FC",X"97",X"C2",X"BD",X"F6",X"9C",X"7A",X"00",X"CC",
		X"26",X"05",X"86",X"01",X"B7",X"00",X"CC",X"7A",X"00",X"CB",X"26",X"04",X"86",X"01",X"97",X"CB",
		X"D6",X"CC",X"86",X"00",X"C3",X"F6",X"80",X"DD",X"C0",X"DE",X"C0",X"A6",X"00",X"C6",X"18",X"BD",
		X"F0",X"4C",X"D6",X"CB",X"86",X"00",X"C3",X"F6",X"65",X"DD",X"C0",X"DE",X"C0",X"A6",X"00",X"C6",
		X"19",X"BD",X"F0",X"4C",X"39",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"0A",X"0C",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"01",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"6A",X"01",X"27",X"01",
		X"39",X"BD",X"F6",X"A5",X"39",X"DF",X"C0",X"E6",X"00",X"C4",X"7F",X"96",X"C2",X"DD",X"C3",X"DE",
		X"C3",X"A6",X"00",X"97",X"C5",X"A6",X"80",X"97",X"C6",X"DE",X"C0",X"6C",X"00",X"96",X"C5",X"81",
		X"C7",X"26",X"0F",X"86",X"00",X"A7",X"00",X"A7",X"01",X"A7",X"02",X"A7",X"03",X"A7",X"04",X"7E",
		X"F6",X"A5",X"81",X"C2",X"26",X"07",X"A6",X"00",X"A7",X"04",X"7E",X"F6",X"A5",X"81",X"C0",X"26",
		X"18",X"A6",X"03",X"27",X"05",X"6A",X"03",X"7E",X"F6",X"A5",X"A6",X"04",X"84",X"7F",X"A7",X"00",
		X"6C",X"02",X"A6",X"02",X"A7",X"03",X"7E",X"F6",X"A5",X"96",X"C6",X"84",X"01",X"27",X"0A",X"BD",
		X"F7",X"5D",X"96",X"C6",X"84",X"FE",X"A7",X"01",X"39",X"96",X"C6",X"A7",X"01",X"C6",X"60",X"D0",
		X"C5",X"86",X"00",X"58",X"49",X"C3",X"FE",X"00",X"DD",X"C3",X"DE",X"C3",X"EC",X"00",X"DD",X"C7",
		X"96",X"C1",X"81",X"A0",X"26",X"1A",X"96",X"C8",X"C6",X"10",X"BD",X"F0",X"4C",X"96",X"C7",X"C6",
		X"11",X"BD",X"F0",X"4C",X"86",X"0F",X"C6",X"18",X"BD",X"F0",X"4C",X"86",X"14",X"97",X"CC",X"39",
		X"96",X"C8",X"C6",X"12",X"BD",X"F0",X"4C",X"96",X"C7",X"C6",X"13",X"BD",X"F0",X"4C",X"86",X"0F",
		X"C6",X"19",X"BD",X"F0",X"4C",X"86",X"14",X"97",X"CB",X"39",X"7E",X"F6",X"A5",X"96",X"C1",X"81",
		X"A0",X"26",X"07",X"86",X"00",X"C6",X"18",X"7E",X"F0",X"4C",X"86",X"00",X"C6",X"19",X"7E",X"F0",
		X"4C",X"39",X"B2",X"81",X"02",X"26",X"31",X"7A",X"00",X"B1",X"96",X"B1",X"26",X"2A",X"86",X"02",
		X"97",X"B1",X"DC",X"B7",X"C3",X"00",X"09",X"DD",X"B7",X"36",X"17",X"C6",X"14",X"BD",X"F0",X"4C",
		X"32",X"C6",X"15",X"BD",X"F0",X"4C",X"7A",X"00",X"B6",X"96",X"B6",X"26",X"0B",X"86",X"00",X"97",
		X"B2",X"86",X"00",X"C6",X"1A",X"BD",X"F0",X"4C",X"39",X"39",X"01",X"00",X"DD",X"B7",X"C6",X"14",
		X"86",X"00",X"BD",X"F0",X"4C",X"C6",X"15",X"86",X"02",X"BD",X"F0",X"4C",X"86",X"F8",X"C6",X"17",
		X"BD",X"F0",X"4C",X"86",X"0E",X"C6",X"1A",X"BD",X"F0",X"4C",X"86",X"08",X"C6",X"1C",X"BD",X"F0",
		X"4C",X"86",X"00",X"C6",X"1D",X"BD",X"F0",X"4C",X"86",X"02",X"97",X"B2",X"86",X"40",X"97",X"B6",
		X"86",X"02",X"97",X"B1",X"39",X"39",X"01",X"97",X"B2",X"86",X"17",X"C6",X"16",X"BD",X"F0",X"4C",
		X"86",X"10",X"C6",X"1A",X"BD",X"F0",X"4C",X"86",X"00",X"C6",X"1D",X"BD",X"F0",X"4C",X"86",X"08",
		X"C6",X"1C",X"BD",X"F0",X"4C",X"86",X"DC",X"C6",X"17",X"BD",X"F0",X"4C",X"39",X"39",X"96",X"C9",
		X"81",X"01",X"20",X"F9",X"7A",X"00",X"B3",X"26",X"F4",X"86",X"20",X"97",X"B3",X"86",X"00",X"C6",
		X"1A",X"BD",X"F0",X"4C",X"86",X"00",X"97",X"B2",X"96",X"B4",X"49",X"24",X"02",X"8A",X"01",X"97",
		X"B4",X"84",X"01",X"27",X"04",X"BD",X"F7",X"E5",X"39",X"39",X"B5",X"49",X"24",X"02",X"8A",X"01",
		X"97",X"B5",X"84",X"01",X"27",X"03",X"BD",X"F7",X"A9",X"39",X"7E",X"F7",X"71",X"86",X"00",X"97",
		X"B4",X"86",X"02",X"97",X"B5",X"86",X"01",X"97",X"B3",X"86",X"00",X"97",X"B2",X"39",X"B2",X"39",
		X"CE",X"00",X"80",X"CC",X"00",X"60",X"A7",X"00",X"08",X"5A",X"2A",X"FA",X"86",X"BF",X"97",X"80",
		X"86",X"07",X"BD",X"FC",X"00",X"CE",X"F0",X"00",X"86",X"01",X"97",X"81",X"7E",X"FC",X"E3",X"FF",
		X"8B",X"9A",X"3C",X"DE",X"D8",X"3C",X"37",X"16",X"86",X"F8",X"DD",X"D8",X"DE",X"D8",X"A6",X"00",
		X"33",X"38",X"DF",X"D8",X"38",X"C6",X"06",X"7E",X"F0",X"4C",X"1F",X"1F",X"1F",X"0E",X"10",X"12",
		X"14",X"16",X"18",X"1A",X"1C",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"18",X"10",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"0A",X"26",X"03",X"7E",X"FC",X"E0",X"96",X"BF",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"8E",X"00",X"FF",X"CE",X"FF",X"FF",X"DF",X"00",X"86",X"3F",X"C6",X"17",X"BD",X"FC",X"00",
		X"BD",X"F9",X"00",X"BD",X"F0",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"C6",X"1F",
		X"BD",X"FC",X"80",X"84",X"0F",X"81",X"01",X"26",X"07",X"BD",X"F8",X"28",X"20",X"F0",X"01",X"01",
		X"81",X"02",X"26",X"08",X"BD",X"F8",X"38",X"20",X"E5",X"01",X"01",X"01",X"81",X"03",X"26",X"08",
		X"BD",X"F8",X"50",X"20",X"D9",X"01",X"01",X"01",X"81",X"04",X"26",X"D2",X"BD",X"F8",X"80",X"20",
		X"CD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DE",X"57",X"49",X"4E",X"44",X"53",X"4F",X"52",X"20",X"41",X"4E",X"44",X"20",X"48",X"4F",X"44",
		X"47",X"45",X"54",X"54",X"53",X"20",X"44",X"4F",X"20",X"49",X"54",X"20",X"41",X"47",X"41",X"49",
		X"4E",X"20",X"53",X"55",X"4E",X"20",X"31",X"30",X"54",X"48",X"20",X"41",X"50",X"52",X"49",X"4C",
		X"20",X"31",X"39",X"38",X"38",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C2",X"28",X"28",X"1C",X"21",X"1A",X"1C",X"1F",X"1A",X"1C",X"21",X"1A",X"1C",X"26",X"1A",X"1C",
		X"28",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C2",X"1F",X"2B",X"1F",X"26",X"1D",X"1F",X"26",
		X"1D",X"1F",X"2B",X"1D",X"1F",X"2B",X"1D",X"1F",X"2B",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C2",X"21",X"2D",X"21",X"26",X"1F",X"21",X"28",X"1F",X"21",X"2B",X"1F",X"21",
		X"2D",X"1F",X"21",X"2D",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"20",X"40",X"20",X"20",X"40",X"20",X"20",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"C7",X"C7",X"C7",X"C7",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CE",X"FA",X"00",X"B6",X"B0",X"00",X"01",X"AD",X"00",X"86",X"05",X"CE",X"00",X"00",X"09",X"26",
		X"FD",X"4A",X"26",X"FA",X"20",X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"E0",
		X"C2",X"2F",X"2F",X"28",X"1C",X"28",X"1C",X"26",X"28",X"1C",X"2B",X"2D",X"21",X"2F",X"1F",X"2B",
		X"28",X"26",X"23",X"26",X"1A",X"28",X"1C",X"2B",X"1F",X"28",X"1C",X"26",X"23",X"28",X"1C",X"2D",
		X"21",X"2B",X"1F",X"28",X"26",X"28",X"1C",X"26",X"1A",X"28",X"26",X"2B",X"28",X"2D",X"2B",X"2F",
		X"23",X"C7",X"C7",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"20",X"20",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0F",X"00",X"10",
		X"00",X"11",X"00",X"12",X"00",X"13",X"00",X"14",X"00",X"15",X"00",X"16",X"00",X"18",X"00",X"19",
		X"00",X"1B",X"00",X"1C",X"00",X"1E",X"00",X"20",X"00",X"22",X"00",X"24",X"00",X"26",X"00",X"28",
		X"00",X"2A",X"00",X"2D",X"00",X"30",X"00",X"32",X"00",X"35",X"00",X"39",X"00",X"3C",X"00",X"3F",
		X"00",X"43",X"00",X"47",X"00",X"4B",X"00",X"50",X"00",X"55",X"00",X"5A",X"00",X"5F",X"00",X"65",
		X"00",X"6B",X"00",X"71",X"00",X"78",X"00",X"7F",X"00",X"87",X"00",X"8F",X"00",X"97",X"00",X"A0",
		X"00",X"A9",X"00",X"B4",X"00",X"BE",X"00",X"CA",X"00",X"D6",X"00",X"E2",X"00",X"F0",X"00",X"FE",
		X"01",X"0D",X"01",X"1D",X"01",X"2E",X"01",X"40",X"01",X"53",X"01",X"67",X"01",X"7C",X"01",X"93",
		X"01",X"AB",X"01",X"C4",X"01",X"DF",X"01",X"FC",X"02",X"1A",X"02",X"3A",X"02",X"5C",X"02",X"80",
		X"02",X"A6",X"02",X"CE",X"02",X"F9",X"03",X"26",X"03",X"56",X"03",X"89",X"03",X"BF",X"03",X"F8",
		X"04",X"34",X"04",X"74",X"04",X"B8",X"05",X"00",X"05",X"4C",X"05",X"9D",X"05",X"F2",X"06",X"4C",
		X"06",X"AC",X"07",X"12",X"07",X"7E",X"07",X"F0",X"08",X"68",X"08",X"E8",X"09",X"70",X"0A",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"03",X"F0",X"00",X"F0",X"09",X"F0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
