library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_P1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_P1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"20",X"75",X"28",X"A5",X"80",X"6A",X"90",X"03",X"4C",X"91",X"28",X"A9",X"3E",X"8D",X"21",X"0B",
		X"8D",X"3D",X"0B",X"A9",X"3F",X"8D",X"42",X"0B",X"8D",X"5E",X"0B",X"A6",X"89",X"E8",X"86",X"89",
		X"E0",X"0F",X"D0",X"10",X"A2",X"00",X"86",X"89",X"E6",X"88",X"A5",X"88",X"C9",X"04",X"D0",X"04",
		X"A9",X"00",X"85",X"88",X"20",X"38",X"28",X"60",X"A9",X"00",X"85",X"8E",X"A4",X"88",X"98",X"0A",
		X"0A",X"18",X"65",X"8E",X"AA",X"BD",X"46",X"29",X"85",X"8C",X"A9",X"0B",X"85",X"8D",X"A5",X"89",
		X"0A",X"0A",X"65",X"8E",X"AA",X"BD",X"56",X"29",X"C9",X"00",X"F0",X"08",X"88",X"30",X"05",X"18",
		X"69",X"25",X"90",X"F8",X"A0",X"00",X"91",X"8C",X"A0",X"1C",X"91",X"8C",X"E6",X"8E",X"A5",X"8E",
		X"C9",X"04",X"D0",X"C8",X"60",X"A5",X"88",X"48",X"A5",X"89",X"48",X"A9",X"0F",X"85",X"89",X"A2",
		X"03",X"86",X"88",X"20",X"38",X"28",X"C6",X"88",X"10",X"F9",X"68",X"85",X"89",X"68",X"85",X"88",
		X"60",X"A0",X"1C",X"98",X"4A",X"29",X"02",X"AA",X"A5",X"CF",X"10",X"21",X"A5",X"E4",X"F0",X"1D",
		X"AD",X"60",X"08",X"38",X"E9",X"04",X"10",X"02",X"A9",X"3F",X"8D",X"60",X"08",X"29",X"30",X"F0",
		X"06",X"85",X"65",X"85",X"67",X"D0",X"1D",X"85",X"64",X"85",X"66",X"F0",X"17",X"BD",X"60",X"08",
		X"D0",X"04",X"95",X"64",X"F0",X"0E",X"DE",X"60",X"08",X"A5",X"63",X"6A",X"90",X"04",X"A5",X"CF",
		X"10",X"02",X"95",X"65",X"B5",X"98",X"4A",X"4A",X"29",X"38",X"85",X"8C",X"B5",X"90",X"2A",X"2A",
		X"2A",X"2A",X"29",X"07",X"05",X"8C",X"AA",X"86",X"8E",X"A5",X"88",X"0A",X"0A",X"0A",X"0A",X"05",
		X"89",X"DD",X"06",X"2A",X"F0",X"19",X"98",X"4A",X"29",X"02",X"AA",X"D6",X"85",X"10",X"3D",X"F6",
		X"84",X"84",X"8C",X"B4",X"84",X"B9",X"3E",X"2A",X"95",X"85",X"A4",X"8C",X"4C",X"2B",X"29",X"98",
		X"4A",X"29",X"02",X"AA",X"24",X"CF",X"10",X"04",X"A5",X"E4",X"D0",X"05",X"A9",X"30",X"9D",X"60",
		X"08",X"A9",X"00",X"95",X"85",X"95",X"84",X"A5",X"8E",X"95",X"C9",X"B5",X"C9",X"AA",X"BD",X"96",
		X"29",X"85",X"8C",X"A9",X"0B",X"85",X"8D",X"BD",X"CE",X"29",X"91",X"8C",X"C0",X"00",X"F0",X"05",
		X"A0",X"00",X"4C",X"93",X"28",X"60",X"02",X"03",X"22",X"23",X"43",X"63",X"42",X"62",X"61",X"60",
		X"41",X"40",X"20",X"00",X"21",X"01",X"44",X"41",X"43",X"42",X"46",X"41",X"45",X"42",X"48",X"41",
		X"47",X"42",X"4A",X"41",X"49",X"42",X"4C",X"41",X"4B",X"42",X"4E",X"41",X"4D",X"42",X"50",X"51",
		X"4F",X"42",X"53",X"54",X"52",X"42",X"40",X"57",X"55",X"56",X"40",X"5A",X"58",X"59",X"40",X"41",
		X"5B",X"5C",X"40",X"41",X"5D",X"5E",X"40",X"41",X"5F",X"60",X"40",X"41",X"61",X"62",X"40",X"41",
		X"63",X"64",X"40",X"41",X"00",X"42",X"00",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"00",X"00",
		X"01",X"01",X"02",X"02",X"03",X"03",X"20",X"20",X"20",X"21",X"22",X"22",X"23",X"23",X"20",X"20",
		X"21",X"21",X"22",X"22",X"23",X"23",X"40",X"40",X"41",X"41",X"42",X"42",X"43",X"43",X"40",X"40",
		X"41",X"41",X"42",X"42",X"43",X"43",X"60",X"60",X"61",X"61",X"62",X"62",X"63",X"63",X"EC",X"EC",
		X"ED",X"EF",X"D4",X"D6",X"D7",X"D7",X"EC",X"EC",X"ED",X"EE",X"D5",X"D6",X"D7",X"D7",X"EB",X"EB",
		X"EB",X"F8",X"F0",X"F8",X"D8",X"D8",X"EA",X"EA",X"F2",X"FA",X"F2",X"FA",X"D9",X"DA",X"E8",X"E8",
		X"F1",X"F9",X"F1",X"F9",X"DB",X"DC",X"E6",X"E6",X"F3",X"FB",X"F3",X"FB",X"DD",X"DD",X"E5",X"E5",
		X"E4",X"E3",X"E1",X"DF",X"DE",X"DE",X"38",X"38",X"3A",X"3D",X"01",X"05",X"08",X"08",X"38",X"38",
		X"3A",X"3D",X"02",X"05",X"08",X"08",X"36",X"36",X"36",X"3A",X"01",X"06",X"0A",X"0A",X"31",X"31",
		X"33",X"37",X"01",X"0B",X"0D",X"0E",X"2E",X"2E",X"2A",X"24",X"1C",X"15",X"12",X"11",X"2A",X"2A",
		X"27",X"22",X"1E",X"19",X"15",X"15",X"28",X"28",X"26",X"21",X"1E",X"1A",X"18",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"40",
		X"A2",X"02",X"BD",X"20",X"00",X"0A",X"B5",X"DF",X"29",X"1F",X"90",X"37",X"F0",X"10",X"C9",X"1B",
		X"B0",X"0A",X"A8",X"A5",X"CD",X"29",X"07",X"C9",X"07",X"98",X"90",X"02",X"E9",X"01",X"95",X"DF",
		X"AD",X"02",X"00",X"29",X"80",X"D0",X"04",X"A9",X"F0",X"85",X"E2",X"A5",X"E2",X"F0",X"08",X"C6",
		X"E2",X"A9",X"00",X"95",X"DF",X"95",X"DE",X"18",X"B5",X"DE",X"F0",X"23",X"D6",X"DE",X"D0",X"1F",
		X"38",X"B0",X"1C",X"C9",X"1B",X"B0",X"09",X"B5",X"DF",X"69",X"20",X"90",X"D1",X"F0",X"01",X"18",
		X"A9",X"1F",X"B0",X"CA",X"95",X"DF",X"B5",X"DE",X"F0",X"01",X"38",X"A9",X"78",X"95",X"DE",X"90",
		X"04",X"E6",X"97",X"E6",X"E3",X"CA",X"CA",X"10",X"99",X"E6",X"CD",X"A5",X"CD",X"4A",X"A5",X"E3",
		X"B0",X"0C",X"F0",X"0A",X"C9",X"10",X"B0",X"02",X"69",X"FF",X"69",X"EF",X"85",X"E3",X"0A",X"60",
		X"A4",X"00",X"00",X"00",X"00",X"00",X"24",X"CF",X"50",X"26",X"A5",X"CF",X"29",X"BF",X"85",X"CF",
		X"A9",X"FF",X"85",X"E4",X"A5",X"63",X"29",X"02",X"F0",X"08",X"A5",X"61",X"6A",X"B0",X"03",X"20",
		X"70",X"2D",X"20",X"3E",X"31",X"A9",X"00",X"85",X"C5",X"85",X"C7",X"85",X"00",X"20",X"6F",X"31",
		X"20",X"10",X"31",X"E6",X"80",X"20",X"CD",X"31",X"A5",X"E4",X"F0",X"02",X"C6",X"E4",X"A2",X"02",
		X"36",X"91",X"18",X"76",X"91",X"95",X"6D",X"B5",X"A1",X"D0",X"03",X"4C",X"3E",X"2B",X"D6",X"A1",
		X"F0",X"16",X"36",X"91",X"38",X"76",X"91",X"A0",X"C0",X"A5",X"80",X"29",X"02",X"F0",X"04",X"B4",
		X"C4",X"95",X"6C",X"94",X"99",X"4C",X"5E",X"2B",X"20",X"87",X"30",X"4C",X"5E",X"2B",X"B5",X"A0",
		X"29",X"0A",X"F0",X"0F",X"A5",X"80",X"29",X"04",X"F0",X"09",X"A5",X"CF",X"F0",X"05",X"36",X"91",
		X"38",X"76",X"91",X"B5",X"C4",X"95",X"99",X"A5",X"E4",X"D0",X"03",X"20",X"A9",X"2E",X"CA",X"CA",
		X"30",X"03",X"4C",X"10",X"2B",X"20",X"00",X"28",X"20",X"2A",X"36",X"20",X"BA",X"32",X"20",X"87",
		X"32",X"A2",X"0A",X"A0",X"00",X"8A",X"6A",X"6A",X"90",X"02",X"A0",X"02",X"B9",X"25",X"00",X"10",
		X"08",X"B9",X"A0",X"00",X"29",X"EF",X"99",X"A0",X"00",X"B5",X"A0",X"30",X"03",X"4C",X"B6",X"2B",
		X"B5",X"A1",X"D0",X"06",X"20",X"A9",X"2E",X"4C",X"41",X"2C",X"D6",X"A1",X"F0",X"0F",X"A0",X"C1",
		X"A5",X"80",X"29",X"02",X"F0",X"02",X"A0",X"C9",X"94",X"C4",X"4C",X"41",X"2C",X"B5",X"A0",X"29",
		X"7F",X"95",X"A0",X"4C",X"DC",X"2B",X"B9",X"A1",X"00",X"D0",X"21",X"C0",X"00",X"F0",X"04",X"A5",
		X"A1",X"10",X"02",X"A5",X"A3",X"D0",X"15",X"A5",X"E4",X"D0",X"11",X"B9",X"A0",X"00",X"10",X"4C",
		X"B9",X"25",X"00",X"30",X"07",X"B9",X"A0",X"00",X"29",X"10",X"F0",X"07",X"A9",X"F9",X"95",X"C4",
		X"4C",X"41",X"2C",X"B9",X"A0",X"00",X"09",X"10",X"99",X"A0",X"00",X"B9",X"99",X"00",X"09",X"01",
		X"95",X"C4",X"B9",X"B8",X"00",X"95",X"B8",X"99",X"D5",X"00",X"B9",X"B9",X"00",X"95",X"B9",X"99",
		X"D6",X"00",X"A9",X"3F",X"99",X"61",X"08",X"A5",X"CF",X"10",X"06",X"A5",X"95",X"09",X"0F",X"85",
		X"95",X"A9",X"80",X"95",X"A0",X"A9",X"00",X"95",X"A1",X"4C",X"41",X"2C",X"B9",X"40",X"08",X"F0",
		X"0A",X"B9",X"41",X"08",X"D0",X"B6",X"20",X"C6",X"35",X"90",X"B1",X"86",X"8C",X"20",X"9A",X"35",
		X"BD",X"F4",X"3B",X"99",X"40",X"08",X"BD",X"00",X"3C",X"99",X"41",X"08",X"A6",X"8C",X"4C",X"E3",
		X"2B",X"CA",X"CA",X"E0",X"02",X"F0",X"0A",X"4C",X"73",X"2B",X"B4",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A5",X"97",X"F0",X"10",X"A5",X"61",X"6A",X"B0",X"06",X"A5",X"63",X"29",X"02",X"D0",X"05",
		X"C6",X"97",X"20",X"70",X"2D",X"24",X"CF",X"10",X"43",X"70",X"70",X"A5",X"E4",X"D0",X"6C",X"F8",
		X"A5",X"81",X"D0",X"22",X"A5",X"82",X"D0",X"11",X"A5",X"83",X"F0",X"27",X"A9",X"59",X"85",X"82",
		X"A5",X"83",X"38",X"E9",X"01",X"85",X"83",X"10",X"07",X"A5",X"82",X"38",X"E9",X"01",X"85",X"82",
		X"A9",X"59",X"85",X"81",X"10",X"07",X"A5",X"81",X"38",X"E9",X"01",X"85",X"81",X"A5",X"CF",X"09",
		X"80",X"30",X"36",X"A9",X"FF",X"85",X"E4",X"A9",X"03",X"8D",X"82",X"08",X"A5",X"61",X"6A",X"90",
		X"11",X"A5",X"E4",X"D0",X"0D",X"20",X"AB",X"38",X"BD",X"0C",X"3C",X"85",X"82",X"BD",X"0D",X"3C",
		X"85",X"83",X"A5",X"26",X"30",X"03",X"4C",X"1C",X"3C",X"A5",X"A0",X"29",X"7F",X"85",X"A0",X"A5",
		X"A2",X"29",X"7F",X"85",X"A2",X"A5",X"CF",X"29",X"7F",X"85",X"CF",X"D8",X"A5",X"83",X"C9",X"A0",
		X"90",X"03",X"4C",X"1C",X"3C",X"20",X"8C",X"34",X"4C",X"D6",X"2A",X"48",X"8A",X"48",X"98",X"48",
		X"D8",X"A5",X"8A",X"C9",X"55",X"D0",X"0E",X"A5",X"8B",X"C9",X"AA",X"D0",X"08",X"BA",X"BD",X"06",
		X"01",X"C9",X"40",X"90",X"03",X"4C",X"1C",X"3C",X"A2",X"02",X"A5",X"E4",X"D0",X"50",X"B5",X"A0",
		X"30",X"03",X"4C",X"8D",X"2D",X"B5",X"05",X"10",X"14",X"B5",X"04",X"10",X"08",X"A9",X"60",X"15",
		X"A0",X"95",X"A0",X"D0",X"08",X"A9",X"40",X"15",X"A0",X"29",X"DF",X"95",X"A0",X"2C",X"24",X"00",
		X"30",X"2C",X"B5",X"A0",X"0A",X"10",X"27",X"0A",X"30",X"11",X"A9",X"FE",X"18",X"75",X"C4",X"95",
		X"C4",X"29",X"F8",X"C9",X"F8",X"D0",X"11",X"A9",X"B8",X"30",X"0B",X"A9",X"02",X"18",X"75",X"C4",
		X"C9",X"C0",X"90",X"02",X"A9",X"00",X"95",X"C4",X"A9",X"BF",X"35",X"A0",X"95",X"A0",X"CA",X"CA",
		X"30",X"03",X"4C",X"0A",X"2D",X"85",X"20",X"20",X"50",X"2A",X"68",X"A8",X"68",X"AA",X"68",X"40",
		X"F8",X"20",X"AB",X"38",X"BD",X"0C",X"3C",X"18",X"65",X"82",X"C9",X"60",X"90",X"02",X"E9",X"60",
		X"85",X"82",X"BD",X"0D",X"3C",X"65",X"83",X"B0",X"02",X"85",X"83",X"D8",X"60",X"B5",X"A0",X"29",
		X"08",X"F0",X"0A",X"A5",X"80",X"10",X"03",X"4C",X"25",X"2D",X"4C",X"1D",X"2D",X"2C",X"24",X"00",
		X"10",X"03",X"4C",X"2D",X"2D",X"86",X"D9",X"8A",X"A8",X"20",X"9A",X"35",X"86",X"DA",X"BD",X"06",
		X"3C",X"A6",X"D9",X"25",X"80",X"F0",X"03",X"4C",X"2D",X"2D",X"A0",X"00",X"E0",X"00",X"D0",X"02",
		X"A0",X"02",X"A5",X"DA",X"C9",X"05",X"90",X"0F",X"B9",X"98",X"00",X"99",X"D6",X"00",X"B9",X"90",
		X"00",X"99",X"D5",X"00",X"4C",X"F9",X"2D",X"B9",X"61",X"08",X"D0",X"1D",X"B9",X"85",X"00",X"F0",
		X"03",X"4C",X"2D",X"2D",X"B9",X"C9",X"00",X"48",X"0A",X"0A",X"29",X"E0",X"99",X"D6",X"00",X"68",
		X"6A",X"6A",X"6A",X"6A",X"29",X"E0",X"99",X"D5",X"00",X"A9",X"00",X"85",X"D9",X"B5",X"B8",X"38",
		X"F9",X"D5",X"00",X"85",X"DA",X"26",X"D9",X"A5",X"D9",X"4A",X"B0",X"07",X"A9",X"00",X"38",X"E5",
		X"DA",X"85",X"DA",X"B5",X"B9",X"38",X"F9",X"D6",X"00",X"85",X"DB",X"26",X"D9",X"A5",X"D9",X"4A",
		X"B0",X"07",X"A9",X"00",X"38",X"E5",X"DB",X"85",X"DB",X"A5",X"DB",X"85",X"DC",X"F0",X"20",X"A9",
		X"FF",X"85",X"DC",X"A4",X"DA",X"F0",X"18",X"A9",X"00",X"85",X"DC",X"A0",X"0C",X"06",X"DC",X"26",
		X"DA",X"2A",X"B0",X"04",X"C5",X"DB",X"90",X"04",X"E5",X"DB",X"E6",X"DC",X"88",X"D0",X"EE",X"A0",
		X"06",X"A5",X"DA",X"D0",X"1A",X"88",X"F0",X"17",X"B9",X"9E",X"2E",X"C5",X"DC",X"90",X"F6",X"38",
		X"E5",X"DC",X"85",X"DD",X"B9",X"9F",X"2E",X"38",X"E5",X"DC",X"C5",X"DD",X"B0",X"01",X"C8",X"84",
		X"DA",X"A4",X"D9",X"B9",X"A5",X"2E",X"18",X"65",X"DA",X"85",X"DA",X"B5",X"99",X"4A",X"4A",X"4A",
		X"C9",X"18",X"B0",X"05",X"38",X"E5",X"DA",X"D0",X"03",X"4C",X"2D",X"2D",X"90",X"06",X"C9",X"0C",
		X"90",X"06",X"B0",X"07",X"C9",X"F4",X"B0",X"03",X"4C",X"25",X"2D",X"4C",X"1D",X"2D",X"FF",X"3C",
		X"1C",X"10",X"09",X"04",X"00",X"06",X"00",X"0C",X"12",X"B5",X"A0",X"29",X"F7",X"95",X"A0",X"86",
		X"8C",X"A9",X"0C",X"E0",X"03",X"90",X"03",X"18",X"69",X"10",X"85",X"8E",X"B5",X"C4",X"4A",X"4A",
		X"4A",X"85",X"8D",X"AA",X"18",X"BD",X"F1",X"39",X"F0",X"0F",X"AA",X"20",X"E4",X"2F",X"A6",X"8C",
		X"A5",X"D2",X"18",X"75",X"AC",X"95",X"AC",X"A5",X"D3",X"A6",X"8C",X"75",X"B8",X"85",X"D0",X"A6",
		X"8D",X"18",X"BD",X"EB",X"39",X"F0",X"0F",X"AA",X"20",X"E4",X"2F",X"A6",X"8C",X"A5",X"D2",X"18",
		X"75",X"AD",X"95",X"AD",X"A5",X"D3",X"A6",X"8C",X"75",X"B9",X"85",X"D1",X"A6",X"8D",X"A4",X"8C",
		X"C0",X"03",X"90",X"06",X"BD",X"3D",X"34",X"4C",X"0D",X"2F",X"BD",X"21",X"3A",X"18",X"65",X"D0",
		X"85",X"8E",X"C0",X"03",X"90",X"06",X"BD",X"25",X"34",X"4C",X"1F",X"2F",X"BD",X"09",X"3A",X"18",
		X"65",X"D1",X"85",X"8F",X"20",X"16",X"30",X"B0",X"0D",X"A5",X"D0",X"99",X"B8",X"00",X"A5",X"D1",
		X"99",X"B9",X"00",X"4C",X"92",X"2F",X"C0",X"03",X"B0",X"09",X"A5",X"CF",X"09",X"01",X"85",X"CF",
		X"4C",X"4D",X"2F",X"A9",X"3F",X"8D",X"81",X"08",X"A9",X"20",X"99",X"A1",X"00",X"B9",X"A0",X"00",
		X"09",X"08",X"99",X"A0",X"00",X"A6",X"8D",X"BD",X"21",X"3A",X"18",X"65",X"D0",X"85",X"8E",X"BD",
		X"09",X"3A",X"18",X"79",X"B9",X"00",X"85",X"8F",X"20",X"16",X"30",X"B0",X"08",X"A5",X"D0",X"99",
		X"B8",X"00",X"4C",X"92",X"2F",X"A6",X"8D",X"BD",X"21",X"3A",X"18",X"79",X"B8",X"00",X"85",X"8E",
		X"BD",X"09",X"3A",X"18",X"65",X"D1",X"85",X"8F",X"20",X"16",X"30",X"B0",X"05",X"A5",X"D1",X"99",
		X"B9",X"00",X"A6",X"8D",X"C0",X"03",X"90",X"06",X"BD",X"3D",X"34",X"4C",X"A1",X"2F",X"BD",X"21",
		X"3A",X"49",X"FF",X"38",X"79",X"B8",X"00",X"85",X"8E",X"C0",X"03",X"90",X"06",X"BD",X"25",X"34",
		X"4C",X"B6",X"2F",X"BD",X"09",X"3A",X"49",X"FF",X"38",X"79",X"B9",X"00",X"85",X"8F",X"20",X"16",
		X"30",X"90",X"1E",X"C0",X"03",X"B0",X"08",X"A5",X"CF",X"09",X"01",X"85",X"CF",X"D0",X"0A",X"A9",
		X"3F",X"8D",X"81",X"08",X"A9",X"20",X"99",X"A1",X"00",X"B9",X"A0",X"00",X"09",X"08",X"99",X"A0",
		X"00",X"A6",X"8C",X"60",X"86",X"8F",X"8A",X"10",X"04",X"49",X"FF",X"AA",X"E8",X"A9",X"00",X"85",
		X"D2",X"85",X"D3",X"A5",X"D2",X"18",X"65",X"8E",X"85",X"D2",X"90",X"02",X"E6",X"D3",X"CA",X"D0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
