library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"DC",X"01",X"E9",X"02",X"CC",X"02",X"CC",X"02",X"CC",X"02",X"CC",X"01",X"E9",X"01",X"E4",
		X"01",X"E6",X"01",X"E1",X"01",X"E4",X"02",X"E6",X"01",X"D9",X"01",X"D9",X"01",X"DB",X"01",X"DC",
		X"01",X"D9",X"01",X"DB",X"02",X"E1",X"01",X"E9",X"01",X"E1",X"01",X"D9",X"02",X"DB",X"02",X"D9",
		X"01",X"80",X"01",X"D9",X"02",X"BC",X"02",X"BC",X"02",X"BC",X"02",X"BC",X"01",X"D9",X"01",X"D4",
		X"01",X"D6",X"01",X"D1",X"01",X"D4",X"02",X"D6",X"01",X"C9",X"01",X"C9",X"01",X"CB",X"01",X"CC",
		X"01",X"C9",X"01",X"CB",X"02",X"D1",X"01",X"C9",X"01",X"D1",X"01",X"C9",X"02",X"CB",X"02",X"C9",
		X"02",X"80",X"02",X"B9",X"02",X"C1",X"02",X"C1",X"02",X"B9",X"02",X"BB",X"02",X"C2",X"02",X"C2",
		X"02",X"B4",X"02",X"B9",X"02",X"C1",X"02",X"C1",X"02",X"B9",X"02",X"BB",X"02",X"C2",X"02",X"C2",
		X"02",X"B4",X"04",X"B5",X"02",X"B4",X"02",X"B4",X"04",X"B5",X"02",X"B4",X"02",X"80",X"02",X"99",
		X"02",X"80",X"02",X"A9",X"02",X"80",X"02",X"B9",X"02",X"80",X"02",X"C9",X"02",X"80",X"02",X"C9",
		X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"D1",X"02",X"D1",X"02",X"D1",X"02",X"D1",X"02",X"CC",
		X"02",X"CC",X"02",X"D1",X"02",X"D1",X"02",X"D1",X"02",X"D2",X"02",X"D1",X"02",X"80",X"02",X"B9",
		X"02",X"B9",X"02",X"B9",X"02",X"B9",X"02",X"C1",X"02",X"C1",X"02",X"C1",X"02",X"C1",X"02",X"BC",
		X"02",X"BC",X"02",X"C1",X"02",X"C1",X"02",X"C1",X"02",X"C2",X"02",X"C1",X"02",X"80",X"02",X"A9",
		X"02",X"B9",X"02",X"B9",X"02",X"A9",X"02",X"AB",X"02",X"B8",X"02",X"B8",X"02",X"A4",X"02",X"A9",
		X"02",X"B9",X"02",X"B9",X"02",X"A9",X"02",X"AB",X"02",X"B8",X"02",X"B8",X"02",X"A4",X"04",X"A5",
		X"02",X"A4",X"02",X"A4",X"04",X"A5",X"02",X"A4",X"02",X"80",X"02",X"99",X"02",X"80",X"02",X"A9",
		X"02",X"80",X"02",X"B9",X"02",X"80",X"02",X"C9",X"02",X"80",X"02",X"C6",X"02",X"C6",X"02",X"C6",
		X"02",X"C6",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",
		X"02",X"C9",X"02",X"C9",X"02",X"C8",X"02",X"C9",X"02",X"80",X"02",X"B6",X"02",X"B6",X"02",X"B6",
		X"02",X"B6",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",
		X"02",X"C9",X"02",X"B9",X"02",X"B8",X"02",X"B9",X"02",X"A0",X"02",X"80",X"02",X"B4",X"02",X"B4",
		X"02",X"80",X"02",X"80",X"02",X"B4",X"02",X"B4",X"02",X"80",X"02",X"80",X"02",X"B4",X"02",X"B4",
		X"02",X"80",X"02",X"80",X"02",X"B4",X"02",X"B4",X"02",X"80",X"08",X"80",X"08",X"80",X"08",X"80",
		X"08",X"80",X"02",X"C3",X"02",X"C3",X"02",X"C3",X"02",X"C3",X"02",X"C4",X"02",X"C4",X"02",X"C4",
		X"02",X"C4",X"02",X"C5",X"02",X"C5",X"02",X"C4",X"02",X"C4",X"02",X"C4",X"02",X"C4",X"04",X"80",
		X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B4",X"02",X"B4",X"02",X"B4",X"02",X"B4",
		X"02",X"B5",X"02",X"B5",X"02",X"B4",X"02",X"B4",X"02",X"B4",X"02",X"B4",X"04",X"80",X"18",X"03",
		X"03",X"03",X"03",X"03",X"03",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",X"FF",
		X"0F",X"FF",X"0F",X"22",X"D7",X"09",X"10",X"10",X"6C",X"0E",X"0A",X"1B",X"0A",X"27",X"0A",X"33",
		X"0A",X"3F",X"0A",X"41",X"0A",X"08",X"18",X"03",X"03",X"03",X"03",X"03",X"03",X"19",X"FF",X"0F",
		X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"22",X"FF",X"09",X"10",X"10",
		X"6C",X"0E",X"0A",X"1B",X"0A",X"27",X"0A",X"33",X"0A",X"3F",X"0A",X"41",X"0A",X"03",X"02",X"B1",
		X"02",X"B5",X"02",X"B8",X"04",X"C1",X"02",X"B8",X"04",X"C1",X"00",X"02",X"B8",X"02",X"C1",X"02",
		X"C5",X"04",X"C8",X"02",X"C5",X"04",X"C8",X"02",X"B5",X"02",X"B8",X"02",X"C1",X"04",X"C5",X"02",
		X"C1",X"04",X"C5",X"02",X"C8",X"02",X"D1",X"02",X"D5",X"04",X"D8",X"02",X"D5",X"04",X"D8",X"10",
		X"80",X"10",X"80",X"19",X"A0",X"00",X"F0",X"00",X"40",X"01",X"1D",X"07",X"09",X"07",X"1E",X"00",
		X"00",X"00",X"07",X"0F",X"00",X"05",X"81",X"13",X"05",X"81",X"10",X"19",X"A0",X"00",X"F0",X"00",
		X"40",X"01",X"1D",X"03",X"04",X"03",X"1E",X"00",X"00",X"00",X"07",X"0F",X"00",X"05",X"81",X"13",
		X"05",X"81",X"10",X"19",X"12",X"00",X"15",X"00",X"20",X"00",X"1D",X"0D",X"0F",X"0D",X"1E",X"00",
		X"00",X"00",X"07",X"05",X"00",X"05",X"81",X"13",X"05",X"81",X"10",X"18",X"03",X"03",X"03",X"03",
		X"03",X"03",X"06",X"00",X"00",X"81",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",
		X"FF",X"0F",X"FF",X"0F",X"22",X"A8",X"0A",X"10",X"08",X"55",X"E3",X"0A",X"EE",X"0A",X"F2",X"0A",
		X"F6",X"0A",X"FA",X"0A",X"FE",X"0A",X"0A",X"18",X"03",X"03",X"03",X"03",X"03",X"03",X"06",X"00",
		X"00",X"81",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",
		X"22",X"D4",X"0A",X"10",X"08",X"55",X"E3",X"0A",X"EE",X"0A",X"F2",X"0A",X"F6",X"0A",X"FA",X"0A",
		X"FE",X"0A",X"04",X"02",X"C1",X"04",X"C3",X"02",X"BC",X"02",X"C1",X"06",X"C3",X"00",X"08",X"80",
		X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",
		X"08",X"80",X"18",X"03",X"03",X"03",X"03",X"03",X"03",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",
		X"1A",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"22",X"1C",X"0B",X"02",X"FB",X"48",X"1E",X"54",X"0B",
		X"E1",X"0C",X"1B",X"0E",X"54",X"0B",X"E1",X"0C",X"1B",X"0E",X"07",X"18",X"03",X"03",X"03",X"03",
		X"03",X"03",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",
		X"22",X"45",X"0B",X"02",X"FB",X"48",X"1E",X"54",X"0B",X"E1",X"0C",X"1B",X"0E",X"54",X"0B",X"E1",
		X"0C",X"1B",X"0E",X"03",X"06",X"D1",X"06",X"C8",X"06",X"D4",X"06",X"D4",X"06",X"D1",X"06",X"D8",
		X"12",X"D8",X"12",X"C8",X"06",X"D1",X"06",X"D3",X"06",X"D4",X"06",X"D6",X"06",X"D8",X"06",X"D9",
		X"06",X"CC",X"06",X"D9",X"06",X"D8",X"06",X"D6",X"06",X"D4",X"06",X"D3",X"12",X"D4",X"18",X"D1",
		X"06",X"CC",X"06",X"D1",X"06",X"D3",X"06",X"D4",X"06",X"D6",X"06",X"D4",X"06",X"D6",X"06",X"D4",
		X"06",X"D3",X"06",X"D4",X"06",X"D1",X"24",X"D8",X"0C",X"80",X"06",X"D8",X"0C",X"D1",X"06",X"D4",
		X"0C",X"C6",X"18",X"80",X"0C",X"80",X"06",X"D6",X"0C",X"CB",X"06",X"D3",X"0C",X"C4",X"18",X"80",
		X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",
		X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",
		X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",
		X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",
		X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",X"02",X"D4",X"02",X"D6",
		X"02",X"D4",X"02",X"D6",X"06",X"D6",X"18",X"D3",X"03",X"D8",X"03",X"D6",X"03",X"D4",X"03",X"D3",
		X"03",X"D1",X"03",X"D3",X"03",X"D1",X"03",X"CB",X"03",X"CA",X"03",X"C8",X"06",X"C7",X"03",X"DA",
		X"03",X"D8",X"03",X"D7",X"03",X"D5",X"03",X"D3",X"03",X"D4",X"03",X"D3",X"03",X"D1",X"03",X"CB",
		X"03",X"CA",X"24",X"CB",X"12",X"CA",X"12",X"D7",X"12",X"D8",X"12",X"80",X"24",X"80",X"06",X"C8",
		X"06",X"C3",X"06",X"CB",X"06",X"CB",X"06",X"C8",X"06",X"D3",X"12",X"D3",X"12",X"C3",X"06",X"C8",
		X"06",X"CA",X"06",X"CB",X"06",X"D1",X"06",X"D3",X"06",X"D4",X"06",X"C7",X"06",X"D4",X"06",X"D3",
		X"06",X"D1",X"06",X"CB",X"06",X"CA",X"0C",X"CB",X"18",X"80",X"03",X"80",X"03",X"C8",X"03",X"CA",
		X"03",X"CB",X"03",X"D1",X"03",X"D3",X"03",X"D4",X"03",X"D6",X"03",X"D4",X"03",X"D3",X"03",X"D1",
		X"03",X"CB",X"0C",X"CA",X"18",X"80",X"03",X"80",X"03",X"C6",X"03",X"C8",X"03",X"CA",X"03",X"CB",
		X"03",X"D1",X"03",X"D3",X"03",X"D4",X"03",X"D3",X"03",X"D1",X"03",X"CB",X"03",X"CA",X"0C",X"C8",
		X"12",X"80",X"06",X"C8",X"0C",X"C6",X"12",X"80",X"06",X"C8",X"0C",X"C4",X"12",X"80",X"06",X"C6",
		X"0C",X"C3",X"06",X"D3",X"1E",X"CB",X"06",X"D4",X"12",X"D1",X"12",X"80",X"18",X"CB",X"06",X"CA",
		X"06",X"C8",X"12",X"C7",X"06",X"C8",X"06",X"C3",X"06",X"CB",X"06",X"CB",X"06",X"C8",X"06",X"D2",
		X"24",X"D2",X"06",X"80",X"06",X"CB",X"06",X"D5",X"06",X"D5",X"06",X"D1",X"06",X"D8",X"24",X"D9",
		X"00",X"48",X"80",X"48",X"80",X"06",X"C1",X"06",X"B8",X"06",X"C4",X"06",X"C4",X"06",X"C1",X"06",
		X"C8",X"12",X"C8",X"12",X"B8",X"06",X"C1",X"06",X"C3",X"06",X"C4",X"06",X"C6",X"06",X"C8",X"06",
		X"C9",X"06",X"BC",X"06",X"C9",X"06",X"C8",X"06",X"C6",X"06",X"C4",X"06",X"C3",X"0C",X"C4",X"1B",
		X"80",X"03",X"C1",X"03",X"C3",X"03",X"C4",X"03",X"C6",X"03",X"C8",X"03",X"C9",X"03",X"CB",X"03",
		X"C9",X"03",X"C8",X"03",X"C6",X"03",X"C4",X"0C",X"C3",X"1B",X"80",X"03",X"BB",X"03",X"C1",X"03",
		X"C3",X"03",X"C4",X"03",X"C6",X"03",X"C8",X"03",X"C9",X"03",X"C8",X"03",X"C6",X"03",X"C4",X"03",
		X"C3",X"0C",X"C1",X"12",X"80",X"06",X"D1",X"1E",X"CB",X"06",X"D1",X"1E",X"C9",X"06",X"CB",X"0C",
		X"C8",X"18",X"80",X"48",X"80",X"06",X"C7",X"06",X"C5",X"06",X"C3",X"06",X"D1",X"06",X"CB",X"06",
		X"CA",X"06",X"CB",X"06",X"D1",X"06",X"CB",X"06",X"CA",X"06",X"CB",X"06",X"C8",X"06",X"D3",X"06",
		X"D1",X"06",X"CB",X"06",X"CA",X"06",X"C8",X"06",X"C7",X"0C",X"C8",X"06",X"80",X"0C",X"C3",X"06",
		X"80",X"0C",X"CA",X"06",X"80",X"0C",X"C7",X"06",X"80",X"0C",X"C8",X"18",X"80",X"2A",X"80",X"06",
		X"C3",X"06",X"CB",X"06",X"CB",X"06",X"C8",X"06",X"D3",X"0C",X"C4",X"18",X"80",X"06",X"C6",X"06",
		X"C1",X"06",X"CA",X"06",X"CA",X"06",X"C6",X"06",X"D1",X"0C",X"C3",X"18",X"80",X"06",X"C4",X"06",
		X"BB",X"06",X"C8",X"06",X"C8",X"06",X"C4",X"06",X"CB",X"06",X"C3",X"06",X"BB",X"06",X"C6",X"06",
		X"C6",X"06",X"C3",X"06",X"CB",X"06",X"C1",X"06",X"C3",X"06",X"C4",X"06",X"C6",X"06",X"C8",X"06",
		X"CA",X"0C",X"BB",X"12",X"80",X"06",X"C8",X"1E",X"C4",X"06",X"CA",X"06",X"C7",X"03",X"D3",X"03",
		X"D1",X"03",X"CB",X"03",X"CA",X"03",X"C8",X"03",X"CA",X"03",X"C8",X"03",X"C6",X"03",X"C4",X"03",
		X"C3",X"18",X"C4",X"06",X"BA",X"06",X"C1",X"0C",X"BB",X"24",X"80",X"06",X"CB",X"0C",X"C8",X"06",
		X"CB",X"0C",X"C5",X"1B",X"80",X"03",X"D6",X"03",X"D4",X"03",X"D2",X"03",X"D1",X"03",X"CB",X"03",
		X"C9",X"03",X"CB",X"03",X"C9",X"03",X"C8",X"03",X"C6",X"03",X"C4",X"12",X"B1",X"12",X"C1",X"06",
		X"BC",X"06",X"BA",X"06",X"B8",X"06",X"C6",X"06",X"C4",X"06",X"C3",X"0C",X"C4",X"06",X"C1",X"0C",
		X"B9",X"06",X"B6",X"0C",X"B8",X"06",X"BA",X"0C",X"BC",X"06",X"B8",X"0C",X"C1",X"3C",X"80",X"48",
		X"80",X"06",X"C1",X"06",X"B8",X"06",X"C4",X"06",X"C4",X"06",X"C1",X"06",X"C8",X"0C",X"B9",X"18",
		X"80",X"06",X"BB",X"06",X"B6",X"06",X"C3",X"06",X"C3",X"06",X"BB",X"06",X"C6",X"0C",X"B8",X"18",
		X"80",X"06",X"B9",X"06",X"B4",X"06",X"C1",X"06",X"C1",X"06",X"B9",X"06",X"C4",X"06",X"B8",X"06",
		X"B4",X"06",X"BB",X"06",X"BB",X"06",X"B8",X"06",X"C4",X"06",X"B6",X"06",X"B8",X"06",X"B9",X"06",
		X"BB",X"06",X"C1",X"06",X"C3",X"12",X"B4",X"12",X"C4",X"12",X"C3",X"12",X"B7",X"06",X"B8",X"06",
		X"B3",X"06",X"BB",X"06",X"BB",X"06",X"B8",X"06",X"C3",X"12",X"C3",X"12",X"B3",X"06",X"B8",X"06",
		X"BA",X"06",X"BB",X"06",X"C1",X"06",X"C3",X"06",X"C4",X"06",X"B7",X"06",X"C4",X"06",X"C3",X"06",
		X"C1",X"06",X"BB",X"06",X"BA",X"12",X"BB",X"12",X"B8",X"06",X"80",X"06",X"B7",X"06",X"B8",X"06",
		X"BA",X"06",X"BB",X"06",X"C1",X"06",X"BB",X"06",X"C1",X"06",X"BB",X"06",X"BA",X"06",X"BB",X"06",
		X"B8",X"06",X"C3",X"06",X"C1",X"06",X"BB",X"06",X"BA",X"06",X"B8",X"06",X"B7",X"0C",X"B8",X"06",
		X"C3",X"0C",X"B8",X"06",X"BB",X"0C",X"B1",X"24",X"80",X"06",X"C1",X"0C",X"B6",X"06",X"BA",X"0C",
		X"AB",X"18",X"80",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",
		X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",
		X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",
		X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",
		X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",
		X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"02",X"B1",X"02",X"AB",X"12",X"AA",X"06",
		X"80",X"03",X"B3",X"03",X"B1",X"03",X"AB",X"03",X"AA",X"03",X"A8",X"03",X"AA",X"03",X"A8",X"03",
		X"A6",X"03",X"A4",X"03",X"A3",X"06",X"A1",X"03",X"B4",X"03",X"B3",X"03",X"B1",X"03",X"AB",X"03",
		X"AA",X"03",X"AB",X"03",X"AA",X"03",X"A8",X"03",X"A7",X"03",X"A5",X"12",X"A3",X"09",X"80",X"03",
		X"A8",X"03",X"AA",X"03",X"AB",X"03",X"B1",X"03",X"AB",X"03",X"B1",X"03",X"B3",X"03",X"B4",X"03",
		X"B1",X"03",X"B3",X"03",X"B4",X"03",X"B3",X"03",X"B1",X"03",X"AB",X"03",X"AA",X"0C",X"A8",X"1E",
		X"80",X"03",X"BB",X"03",X"B9",X"03",X"B8",X"03",X"B6",X"03",X"B5",X"03",X"B6",X"03",X"B5",X"03",
		X"B3",X"03",X"B1",X"03",X"AB",X"03",X"A9",X"03",X"B6",X"03",X"B5",X"03",X"B3",X"03",X"B1",X"03",
		X"AB",X"03",X"A9",X"03",X"AB",X"03",X"A9",X"03",X"A8",X"03",X"A6",X"03",X"A5",X"0C",X"A6",X"18",
		X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
