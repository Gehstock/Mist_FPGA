library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"11",X"3F",X"FC",X"BF",X"81",X"11",X"3F",X"25",X"C6",X"81",X"11",X"3F",X"2A",X"D5",X"81",X"0E",
		X"03",X"C0",X"81",X"04",X"04",X"0B",X"0E",X"03",X"CF",X"81",X"0F",X"0F",X"0F",X"0F",X"02",X"B8",
		X"81",X"5D",X"0D",X"AE",X"06",X"06",X"08",X"98",X"81",X"14",X"C4",X"0A",X"0A",X"01",X"C0",X"81",
		X"0A",X"01",X"C1",X"81",X"03",X"98",X"81",X"F1",X"14",X"E8",X"0A",X"11",X"00",X"F8",X"CE",X"81",
		X"0F",X"03",X"B8",X"81",X"AE",X"06",X"4D",X"05",X"75",X"04",X"0F",X"03",X"C7",X"81",X"3B",X"02",
		X"AC",X"01",X"53",X"01",X"14",X"C4",X"0A",X"07",X"68",X"01",X"CB",X"81",X"07",X"CF",X"02",X"BA",
		X"81",X"14",X"D6",X"0A",X"14",X"D6",X"0A",X"14",X"21",X"0B",X"11",X"00",X"FC",X"BF",X"81",X"07",
		X"5D",X"0D",X"B8",X"81",X"14",X"E8",X"0A",X"11",X"00",X"F8",X"BF",X"81",X"11",X"00",X"F8",X"CE",
		X"81",X"0E",X"03",X"CF",X"81",X"0E",X"0F",X"0F",X"0F",X"03",X"B8",X"81",X"AE",X"06",X"9E",X"05",
		X"75",X"04",X"0F",X"03",X"C7",X"81",X"AC",X"01",X"68",X"01",X"1D",X"01",X"14",X"C4",X"0A",X"0F",
		X"02",X"C7",X"81",X"D6",X"00",X"53",X"01",X"07",X"4D",X"05",X"BA",X"81",X"14",X"D6",X"0A",X"14",
		X"D6",X"0A",X"14",X"21",X"0B",X"11",X"00",X"FC",X"BF",X"81",X"07",X"5D",X"0D",X"B8",X"81",X"14",
		X"E8",X"0A",X"14",X"D6",X"0A",X"11",X"3F",X"F8",X"BF",X"81",X"11",X"3F",X"F8",X"CE",X"81",X"0E",
		X"03",X"CF",X"81",X"0F",X"0F",X"0F",X"0F",X"03",X"B8",X"81",X"AE",X"06",X"4D",X"05",X"75",X"04",
		X"0F",X"03",X"C7",X"81",X"3B",X"02",X"53",X"01",X"AC",X"01",X"14",X"C4",X"0A",X"0F",X"02",X"C7",
		X"81",X"40",X"01",X"FE",X"00",X"0F",X"02",X"BA",X"81",X"01",X"05",X"F9",X"03",X"14",X"D6",X"0A",
		X"12",X"3C",X"CE",X"81",X"0F",X"03",X"B8",X"81",X"01",X"05",X"F9",X"03",X"57",X"03",X"0F",X"02",
		X"C7",X"81",X"81",X"02",X"FC",X"01",X"14",X"CD",X"0A",X"0F",X"02",X"C7",X"81",X"3B",X"02",X"C5",
		X"01",X"14",X"CD",X"0A",X"0F",X"02",X"C7",X"81",X"FC",X"01",X"AC",X"01",X"14",X"C4",X"0A",X"14",
		X"D6",X"0A",X"0E",X"03",X"C0",X"81",X"0D",X"0D",X"0D",X"0E",X"03",X"CF",X"81",X"0F",X"0F",X"0F",
		X"11",X"00",X"F8",X"BF",X"81",X"11",X"00",X"F8",X"CE",X"81",X"0F",X"03",X"B8",X"81",X"F4",X"05",
		X"01",X"05",X"57",X"03",X"0F",X"03",X"C7",X"81",X"1B",X"02",X"AC",X"01",X"7D",X"01",X"14",X"DF",
		X"0A",X"12",X"FC",X"BF",X"81",X"0F",X"02",X"B8",X"81",X"EB",X"08",X"4D",X"05",X"0F",X"03",X"C7",
		X"81",X"3B",X"02",X"AC",X"01",X"53",X"01",X"14",X"C4",X"0A",X"12",X"FC",X"CE",X"81",X"0F",X"02",
		X"B8",X"81",X"EB",X"08",X"01",X"05",X"0F",X"02",X"C7",X"81",X"7D",X"01",X"40",X"01",X"14",X"C4",
		X"0A",X"11",X"00",X"F8",X"BF",X"81",X"11",X"00",X"F8",X"CE",X"81",X"0F",X"03",X"B8",X"81",X"EB",
		X"08",X"AE",X"06",X"4D",X"05",X"0F",X"03",X"C7",X"81",X"AC",X"01",X"53",X"01",X"1D",X"01",X"14",
		X"DF",X"0A",X"0E",X"03",X"C0",X"81",X"0D",X"0D",X"0D",X"0E",X"03",X"CF",X"81",X"0D",X"0D",X"0D",
		X"12",X"FE",X"BF",X"81",X"07",X"57",X"03",X"B8",X"81",X"14",X"C4",X"0A",X"07",X"75",X"04",X"B8",
		X"81",X"14",X"C4",X"0A",X"07",X"4D",X"05",X"B8",X"81",X"14",X"C4",X"0A",X"07",X"AE",X"06",X"B8",
		X"81",X"0E",X"03",X"C0",X"81",X"0C",X"0C",X"0C",X"0E",X"03",X"CF",X"81",X"0F",X"0F",X"0F",X"12",
		X"FC",X"BF",X"81",X"0F",X"02",X"C7",X"81",X"AC",X"01",X"53",X"01",X"14",X"CD",X"0A",X"0F",X"02",
		X"C7",X"81",X"7D",X"01",X"40",X"01",X"14",X"CD",X"0A",X"0F",X"03",X"C7",X"81",X"AC",X"01",X"53",
		X"01",X"1D",X"01",X"0F",X"03",X"B8",X"81",X"AE",X"06",X"4D",X"05",X"75",X"04",X"11",X"00",X"F8",
		X"BF",X"81",X"11",X"00",X"F8",X"CE",X"81",X"14",X"D6",X"0A",X"0E",X"03",X"C0",X"81",X"0B",X"0B",
		X"0C",X"0E",X"03",X"CF",X"81",X"0F",X"0F",X"0F",X"0F",X"03",X"B8",X"81",X"AE",X"06",X"4D",X"05",
		X"F9",X"03",X"0F",X"03",X"C7",X"81",X"AC",X"01",X"53",X"01",X"FE",X"00",X"14",X"DF",X"0A",X"0F",
		X"03",X"B8",X"81",X"F4",X"05",X"75",X"04",X"8A",X"03",X"0F",X"03",X"C7",X"81",X"7D",X"01",X"1D",
		X"01",X"E2",X"00",X"14",X"DF",X"0A",X"0F",X"03",X"B8",X"81",X"AE",X"06",X"4D",X"05",X"75",X"04",
		X"0F",X"03",X"C7",X"81",X"53",X"01",X"1D",X"01",X"D6",X"00",X"14",X"D6",X"0A",X"14",X"D6",X"0A",
		X"14",X"DF",X"0A",X"12",X"3E",X"BF",X"81",X"12",X"3F",X"CE",X"81",X"06",X"08",X"C0",X"81",X"07",
		X"AE",X"06",X"B8",X"81",X"14",X"D6",X"0A",X"14",X"D6",X"0A",X"12",X"3F",X"BF",X"81",X"01",X"10",
		X"07",X"AE",X"06",X"BA",X"81",X"14",X"C4",X"0A",X"03",X"98",X"81",X"F4",X"15",X"06",X"00",X"C5",
		X"81",X"01",X"06",X"03",X"C5",X"81",X"07",X"00",X"0D",X"C3",X"81",X"07",X"64",X"00",X"A8",X"81",
		X"13",X"A8",X"81",X"15",X"07",X"96",X"00",X"A8",X"81",X"13",X"A8",X"81",X"15",X"07",X"4B",X"00",
		X"A8",X"81",X"13",X"A8",X"81",X"15",X"07",X"58",X"02",X"A8",X"81",X"13",X"A8",X"81",X"15",X"07",
		X"2C",X"01",X"A8",X"81",X"13",X"A8",X"81",X"15",X"11",X"00",X"F8",X"BF",X"81",X"0E",X"03",X"C0",
		X"81",X"0B",X"0B",X"0F",X"07",X"57",X"03",X"BC",X"81",X"06",X"04",X"98",X"81",X"14",X"A0",X"0A",
		X"07",X"3B",X"02",X"BC",X"81",X"06",X"04",X"98",X"81",X"14",X"A0",X"0A",X"07",X"AC",X"01",X"BC",
		X"81",X"06",X"07",X"98",X"81",X"14",X"A0",X"0A",X"07",X"C2",X"01",X"A8",X"81",X"13",X"A8",X"81",
		X"15",X"0E",X"03",X"C0",X"81",X"10",X"00",X"00",X"11",X"00",X"FE",X"BF",X"81",X"11",X"03",X"3E",
		X"C6",X"81",X"07",X"AE",X"06",X"B8",X"81",X"14",X"AD",X"0A",X"0E",X"03",X"CF",X"81",X"00",X"00",
		X"00",X"07",X"EB",X"08",X"B8",X"81",X"14",X"AD",X"0A",X"06",X"05",X"98",X"81",X"07",X"AE",X"06",
		X"B8",X"81",X"14",X"AD",X"0A",X"07",X"EB",X"08",X"B8",X"81",X"14",X"AD",X"0A",X"03",X"98",X"81",
		X"EC",X"06",X"0C",X"C0",X"81",X"11",X"03",X"3D",X"C6",X"81",X"15",X"07",X"00",X"00",X"49",X"81",
		X"07",X"00",X"00",X"6F",X"81",X"07",X"00",X"00",X"95",X"81",X"12",X"3F",X"CE",X"81",X"11",X"3F",
		X"FC",X"BF",X"81",X"11",X"3F",X"25",X"C6",X"81",X"11",X"3F",X"2A",X"D5",X"81",X"0E",X"03",X"C0",
		X"81",X"04",X"04",X"0B",X"0E",X"03",X"CF",X"81",X"0F",X"0F",X"0F",X"0F",X"02",X"B8",X"81",X"5D",
		X"0D",X"AE",X"06",X"06",X"08",X"98",X"81",X"14",X"C4",X"0A",X"0A",X"01",X"C0",X"81",X"0A",X"01",
		X"C1",X"81",X"03",X"98",X"81",X"F1",X"14",X"E8",X"0A",X"11",X"00",X"F8",X"CE",X"81",X"0F",X"03",
		X"B8",X"81",X"AE",X"06",X"4D",X"05",X"75",X"04",X"0F",X"03",X"C7",X"81",X"3B",X"02",X"AC",X"01",
		X"53",X"01",X"14",X"C4",X"0A",X"07",X"68",X"01",X"CB",X"81",X"07",X"CF",X"02",X"BA",X"81",X"14",
		X"D6",X"0A",X"14",X"D6",X"0A",X"12",X"3F",X"BF",X"81",X"12",X"3F",X"CE",X"81",X"00",X"0E",X"03",
		X"C3",X"81",X"00",X"00",X"00",X"01",X"07",X"60",X"03",X"BC",X"81",X"07",X"00",X"13",X"C3",X"81",
		X"06",X"03",X"C5",X"81",X"11",X"24",X"FB",X"BF",X"81",X"11",X"30",X"1F",X"C6",X"81",X"06",X"10",
		X"C2",X"81",X"07",X"F4",X"01",X"98",X"81",X"13",X"98",X"81",X"06",X"00",X"C2",X"81",X"12",X"24",
		X"BF",X"81",X"00",X"10",X"0E",X"03",X"C0",X"81",X"0D",X"0C",X"0B",X"11",X"3F",X"F8",X"BF",X"81",
		X"11",X"3F",X"2A",X"C6",X"81",X"0F",X"03",X"B8",X"81",X"6B",X"00",X"55",X"00",X"47",X"00",X"06",
		X"14",X"A6",X"81",X"06",X"0C",X"A4",X"81",X"01",X"0B",X"1A",X"00",X"B8",X"81",X"0B",X"16",X"00",
		X"BA",X"81",X"0B",X"10",X"00",X"BC",X"81",X"03",X"A4",X"81",X"EC",X"06",X"0C",X"A4",X"81",X"01",
		X"0B",X"E6",X"FF",X"B8",X"81",X"0B",X"EA",X"FF",X"BA",X"81",X"0B",X"F0",X"FF",X"BC",X"81",X"03",
		X"A4",X"81",X"EC",X"03",X"A6",X"81",X"CC",X"12",X"3F",X"BF",X"81",X"00",X"0E",X"02",X"C0",X"81",
		X"09",X"09",X"0F",X"02",X"B8",X"81",X"AC",X"01",X"53",X"01",X"0F",X"02",X"98",X"81",X"14",X"00",
		X"14",X"00",X"14",X"B2",X"0C",X"02",X"F3",X"0E",X"02",X"C0",X"81",X"07",X"07",X"0F",X"02",X"B8",
		X"81",X"3B",X"02",X"AC",X"01",X"0F",X"02",X"98",X"81",X"38",X"00",X"38",X"00",X"14",X"B2",X"0C",
		X"02",X"F3",X"11",X"1B",X"FC",X"BF",X"81",X"11",X"3F",X"2A",X"C6",X"81",X"01",X"0B",X"10",X"00",
		X"B8",X"81",X"0B",X"0C",X"00",X"BA",X"81",X"03",X"98",X"81",X"F1",X"01",X"0B",X"F0",X"FF",X"B8",
		X"81",X"0B",X"F4",X"FF",X"BA",X"81",X"03",X"9A",X"81",X"F1",X"15",X"11",X"3F",X"FF",X"BF",X"81",
		X"0E",X"03",X"C3",X"81",X"00",X"00",X"00",X"01",X"11",X"1B",X"FC",X"BF",X"81",X"11",X"0F",X"3F",
		X"C6",X"81",X"0E",X"03",X"C0",X"81",X"10",X"10",X"00",X"0F",X"02",X"B8",X"81",X"80",X"00",X"00",
		X"00",X"07",X"00",X"0C",X"C3",X"81",X"07",X"03",X"00",X"C5",X"81",X"06",X"02",X"98",X"81",X"06",
		X"6E",X"9A",X"81",X"01",X"0B",X"03",X"00",X"B8",X"81",X"0B",X"04",X"00",X"BA",X"81",X"03",X"9A",
		X"81",X"F1",X"16",X"03",X"98",X"81",X"E8",X"12",X"1B",X"BF",X"81",X"00",X"11",X"3F",X"FF",X"CE",
		X"81",X"0E",X"03",X"D2",X"81",X"00",X"00",X"00",X"01",X"11",X"09",X"FE",X"CE",X"81",X"11",X"03",
		X"3D",X"D5",X"81",X"06",X"10",X"CF",X"81",X"07",X"48",X"00",X"C7",X"81",X"07",X"04",X"18",X"D2",
		X"81",X"07",X"03",X"00",X"D4",X"81",X"06",X"50",X"A8",X"81",X"06",X"06",X"AA",X"81",X"13",X"AA",
		X"81",X"0B",X"04",X"00",X"C7",X"81",X"03",X"A8",X"81",X"F0",X"12",X"1B",X"CE",X"81",X"00",X"11",
		X"24",X"FB",X"BF",X"81",X"11",X"30",X"2F",X"C6",X"81",X"06",X"0F",X"C2",X"81",X"07",X"48",X"00",
		X"BC",X"81",X"06",X"20",X"A2",X"81",X"06",X"20",X"A0",X"81",X"01",X"0A",X"08",X"BC",X"81",X"03",
		X"A0",X"81",X"F7",X"06",X"10",X"A0",X"81",X"01",X"0A",X"F7",X"BC",X"81",X"03",X"A0",X"81",X"F7",
		X"03",X"A2",X"81",X"E2",X"12",X"24",X"BF",X"81",X"00",X"11",X"3F",X"F8",X"CE",X"81",X"11",X"3F",
		X"2A",X"D5",X"81",X"0E",X"03",X"CF",X"81",X"0B",X"0C",X"0C",X"0F",X"03",X"C7",X"81",X"32",X"00",
		X"32",X"00",X"32",X"00",X"06",X"02",X"B6",X"81",X"06",X"20",X"B4",X"81",X"07",X"32",X"00",X"C7",
		X"81",X"01",X"0B",X"0F",X"00",X"C7",X"81",X"0B",X"11",X"00",X"C9",X"81",X"0B",X"10",X"00",X"CB",
		X"81",X"03",X"B4",X"81",X"EC",X"03",X"B6",X"81",X"DF",X"06",X"A4",X"B4",X"81",X"01",X"0B",X"0A",
		X"00",X"C7",X"81",X"0B",X"0D",X"00",X"C9",X"81",X"0B",X"0F",X"00",X"CB",X"81",X"03",X"B4",X"81",
		X"EC",X"12",X"3F",X"CE",X"81",X"00",X"0E",X"03",X"CF",X"81",X"0F",X"0F",X"0F",X"11",X"3F",X"F8",
		X"CE",X"81",X"11",X"3F",X"2A",X"D5",X"81",X"0F",X"03",X"C7",X"81",X"C8",X"00",X"3C",X"00",X"28",
		X"00",X"06",X"14",X"B0",X"81",X"06",X"14",X"B2",X"81",X"01",X"0B",X"14",X"00",X"C7",X"81",X"0B",
		X"06",X"00",X"C9",X"81",X"0B",X"04",X"00",X"CB",X"81",X"03",X"B2",X"81",X"EC",X"06",X"14",X"B2",
		X"81",X"01",X"0B",X"EC",X"FF",X"C7",X"81",X"0B",X"FA",X"FF",X"C9",X"81",X"0B",X"FC",X"FF",X"CB",
		X"81",X"03",X"B2",X"81",X"EC",X"03",X"B0",X"81",X"CC",X"12",X"3F",X"CE",X"81",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
