library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity crater_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of crater_bg_bits_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"6A",X"AA",X"95",X"55",
		X"55",X"55",X"55",X"61",X"55",X"55",X"66",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"56",X"AA",
		X"55",X"55",X"54",X"85",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"58",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"68",X"A6",X"15",X"55",X"55",X"55",
		X"55",X"55",X"60",X"AA",X"85",X"55",X"55",X"55",X"55",X"55",X"2A",X"AA",X"85",X"55",X"55",X"55",
		X"55",X"55",X"8A",X"AA",X"85",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A1",X"55",X"55",X"55",
		X"55",X"54",X"AA",X"AA",X"A1",X"55",X"55",X"50",X"55",X"9A",X"AA",X"AA",X"25",X"55",X"55",X"55",
		X"54",X"9A",X"AA",X"AA",X"A9",X"55",X"55",X"45",X"5A",X"AA",X"AA",X"AA",X"29",X"55",X"55",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"5A",X"AA",X"55",X"55",X"5A",X"AA",X"A5",X"55",
		X"56",X"95",X"56",X"A9",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"6A",X"A5",X"55",X"55",X"55",
		X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"45",X"55",X"55",X"55",X"56",X"55",X"55",X"51",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"51",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"55",X"95",X"55",
		X"54",X"2A",X"A5",X"56",X"66",X"AA",X"55",X"55",X"55",X"55",X"6A",X"A5",X"55",X"95",X"55",X"95",
		X"55",X"55",X"55",X"AA",X"65",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"95",X"55",X"56",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"59",
		X"55",X"55",X"55",X"55",X"55",X"55",X"48",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"A1",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A2",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"86",X"55",
		X"95",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"69",X"64",X"55",X"55",X"55",
		X"56",X"A5",X"5A",X"95",X"A4",X"55",X"55",X"55",X"55",X"42",X"AA",X"82",X"55",X"00",X"00",X"05",
		X"55",X"AA",X"A5",X"96",X"95",X"55",X"40",X"45",X"55",X"45",X"15",X"56",X"55",X"55",X"55",X"50",
		X"55",X"65",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"05",X"55",X"6A",X"95",X"55",X"55",X"55",X"55",X"99",X"55",X"29",X"55",X"55",X"55",X"55",
		X"55",X"25",X"55",X"95",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"96",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"96",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A6",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"92",X"45",X"95",X"55",X"55",X"55",
		X"51",X"50",X"25",X"54",X"4A",X"85",X"55",X"55",X"52",X"55",X"55",X"55",X"55",X"50",X"15",X"69",
		X"40",X"50",X"55",X"55",X"55",X"5A",X"A6",X"99",X"05",X"55",X"55",X"55",X"55",X"19",X"69",X"95",
		X"55",X"55",X"55",X"54",X"41",X"55",X"59",X"A5",X"55",X"55",X"55",X"55",X"54",X"55",X"59",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"99",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"54",X"55",X"5A",X"AA",X"58",
		X"55",X"40",X"21",X"A9",X"45",X"A8",X"51",X"55",X"55",X"55",X"52",X"05",X"55",X"AA",X"55",X"44",
		X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"46",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"05",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"21",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"09",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"A1",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"81",X"55",X"55",X"55",X"55",X"55",X"55",
		X"52",X"99",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",
		X"52",X"A1",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"86",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"2A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"0A",X"55",X"55",X"55",X"55",X"55",X"55",X"58",X"AA",
		X"55",X"55",X"6A",X"55",X"55",X"55",X"5A",X"AA",X"55",X"55",X"68",X"55",X"55",X"55",X"4A",X"88",
		X"55",X"55",X"8A",X"65",X"55",X"55",X"68",X"AA",X"55",X"56",X"AA",X"85",X"55",X"55",X"28",X"8A",
		X"AA",X"4A",X"AA",X"AA",X"95",X"55",X"55",X"55",X"AA",X"8A",X"AA",X"AA",X"55",X"55",X"51",X"45",
		X"AA",X"2A",X"AA",X"A9",X"55",X"55",X"55",X"95",X"A8",X"AA",X"AA",X"A9",X"55",X"55",X"54",X"A5",
		X"9A",X"AA",X"AA",X"A1",X"55",X"55",X"55",X"59",X"A6",X"AA",X"AA",X"A5",X"59",X"55",X"55",X"65",
		X"AA",X"AA",X"AA",X"85",X"61",X"55",X"55",X"65",X"AA",X"AA",X"AA",X"85",X"69",X"65",X"55",X"55",
		X"AA",X"A9",X"8A",X"86",X"A9",X"85",X"55",X"59",X"A4",X"A6",X"2A",X"96",X"28",X"AA",X"95",X"55",
		X"A2",X"92",X"AA",X"9A",X"A9",X"A6",X"55",X"55",X"2A",X"52",X"AA",X"9A",X"AA",X"A9",X"55",X"55",
		X"89",X"5A",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"A5",X"5A",X"AA",X"AA",X"AA",X"81",X"55",X"55",
		X"A5",X"4A",X"AA",X"6A",X"AA",X"A5",X"55",X"55",X"95",X"2A",X"AA",X"A6",X"A2",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"8A",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"8A",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"2A",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"66",X"55",
		X"55",X"55",X"55",X"55",X"55",X"62",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A9",X"55",
		X"55",X"55",X"55",X"55",X"55",X"6A",X"A9",X"59",X"55",X"55",X"55",X"55",X"55",X"AA",X"A5",X"65",
		X"55",X"55",X"55",X"55",X"55",X"A9",X"A5",X"A5",X"55",X"55",X"55",X"55",X"55",X"AA",X"A6",X"55",
		X"55",X"55",X"55",X"55",X"55",X"AA",X"95",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"99",X"95",
		X"55",X"55",X"55",X"55",X"66",X"A9",X"56",X"15",X"55",X"55",X"55",X"55",X"AA",X"AA",X"5A",X"95",
		X"55",X"55",X"55",X"55",X"8A",X"AA",X"68",X"55",X"55",X"55",X"55",X"56",X"A2",X"AA",X"A9",X"55",
		X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"A5",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"55",
		X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",
		X"58",X"88",X"55",X"55",X"55",X"55",X"55",X"55",X"52",X"A1",X"55",X"55",X"55",X"55",X"55",X"55",
		X"52",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"A9",X"85",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"A9",X"A5",X"55",X"55",X"55",X"55",X"95",X"5A",X"A9",X"A5",X"55",X"55",X"55",X"55",X"95",
		X"5A",X"A5",X"65",X"55",X"55",X"55",X"55",X"95",X"5A",X"A6",X"A5",X"55",X"55",X"55",X"AA",X"95",
		X"5A",X"A5",X"29",X"55",X"55",X"55",X"AA",X"59",X"6A",X"A6",X"29",X"55",X"55",X"6A",X"95",X"55",
		X"62",X"AA",X"09",X"55",X"55",X"69",X"55",X"55",X"42",X"AA",X"29",X"95",X"55",X"55",X"65",X"55",
		X"8A",X"A6",X"29",X"95",X"55",X"55",X"55",X"55",X"5A",X"AA",X"2A",X"95",X"55",X"55",X"55",X"55",
		X"4A",X"A6",X"29",X"95",X"55",X"55",X"55",X"59",X"2A",X"AA",X"22",X"95",X"55",X"55",X"55",X"65",
		X"55",X"56",X"9A",X"95",X"55",X"56",X"6A",X"AA",X"55",X"5A",X"66",X"85",X"55",X"69",X"AA",X"69",
		X"55",X"52",X"56",X"25",X"15",X"9A",X"66",X"A5",X"55",X"4A",X"95",X"85",X"95",X"69",X"A9",X"55",
		X"55",X"28",X"56",X"26",X"15",X"6A",X"65",X"55",X"54",X"29",X"56",X"8A",X"59",X"56",X"6A",X"59",
		X"54",X"A5",X"9A",X"22",X"95",X"55",X"55",X"59",X"54",X"95",X"A8",X"88",X"A9",X"55",X"55",X"55",
		X"5A",X"95",X"A5",X"4A",X"22",X"A5",X"55",X"59",X"52",X"56",X"56",X"AA",X"A9",X"15",X"55",X"55",
		X"4A",X"55",X"69",X"5A",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"45",X"56",X"15",X"55",
		X"55",X"AA",X"8A",X"95",X"8A",X"55",X"55",X"55",X"55",X"AA",X"6A",X"99",X"AA",X"55",X"55",X"55",
		X"55",X"A4",X"6A",X"6A",X"A9",X"55",X"55",X"55",X"5A",X"59",X"A9",X"AA",X"A9",X"A1",X"55",X"55",
		X"AA",X"5A",X"A5",X"AA",X"6A",X"99",X"55",X"55",X"A5",X"56",X"A9",X"AA",X"AA",X"68",X"55",X"55",
		X"59",X"5A",X"AA",X"AA",X"AA",X"9A",X"95",X"55",X"55",X"5A",X"A9",X"5A",X"AA",X"AA",X"A5",X"55",
		X"55",X"66",X"A5",X"6A",X"AA",X"AA",X"65",X"55",X"55",X"AA",X"A5",X"95",X"AA",X"AA",X"95",X"55",
		X"55",X"55",X"65",X"55",X"AA",X"AA",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"AA",X"99",X"55",
		X"55",X"55",X"55",X"55",X"55",X"6A",X"A8",X"81",X"55",X"96",X"55",X"59",X"55",X"55",X"6A",X"A1",
		X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"89",X"55",X"55",X"56",X"55",X"55",X"55",X"56",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"55",X"56",X"86",X"AA",X"A2",X"55",
		X"55",X"55",X"55",X"99",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"16",X"2A",X"AA",X"A9",X"55",
		X"55",X"55",X"54",X"99",X"A6",X"AA",X"A9",X"55",X"55",X"55",X"56",X"96",X"AA",X"AA",X"85",X"55",
		X"55",X"55",X"56",X"56",X"9A",X"AA",X"95",X"55",X"55",X"55",X"52",X"56",X"AA",X"AA",X"95",X"55",
		X"55",X"55",X"52",X"56",X"6A",X"AA",X"55",X"55",X"55",X"55",X"5A",X"55",X"AA",X"A9",X"95",X"55",
		X"55",X"55",X"59",X"56",X"AA",X"AA",X"55",X"55",X"55",X"55",X"19",X"56",X"AA",X"A9",X"55",X"65",
		X"55",X"54",X"29",X"56",X"AA",X"6A",X"56",X"65",X"55",X"56",X"A5",X"5A",X"AA",X"AA",X"59",X"55",
		X"55",X"42",X"29",X"6A",X"AA",X"AA",X"55",X"65",X"55",X"28",X"A5",X"5A",X"AA",X"A9",X"65",X"5A",
		X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"61",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"65",X"85",X"55",X"55",X"55",X"55",X"55",X"55",X"A6",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"A1",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"99",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"99",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"46",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"49",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",
		X"29",X"A6",X"2A",X"95",X"55",X"55",X"56",X"A5",X"28",X"AA",X"8A",X"95",X"55",X"55",X"55",X"55",
		X"88",X"6A",X"6A",X"95",X"55",X"55",X"69",X"55",X"0A",X"16",X"5A",X"95",X"55",X"55",X"55",X"55",
		X"42",X"5A",X"AA",X"05",X"55",X"55",X"55",X"55",X"65",X"5A",X"68",X"85",X"55",X"55",X"55",X"55",
		X"85",X"6A",X"9A",X"85",X"55",X"55",X"55",X"55",X"2A",X"9A",X"AA",X"85",X"55",X"55",X"55",X"55",
		X"9A",X"69",X"66",X"85",X"55",X"55",X"55",X"55",X"6A",X"6A",X"52",X"05",X"55",X"55",X"55",X"55",
		X"A6",X"9A",X"4A",X"15",X"55",X"55",X"55",X"55",X"96",X"A6",X"26",X"95",X"55",X"55",X"55",X"55",
		X"9A",X"96",X"26",X"15",X"55",X"55",X"55",X"55",X"99",X"9A",X"06",X"95",X"55",X"55",X"55",X"55",
		X"99",X"AA",X"8A",X"A5",X"55",X"55",X"55",X"55",X"AA",X"69",X"8A",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"59",X"59",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"56",X"55",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"58",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"2A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"A6",X"95",X"2A",X"55",X"6A",
		X"55",X"55",X"55",X"54",X"58",X"99",X"99",X"55",X"55",X"55",X"55",X"69",X"A6",X"A9",X"A5",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"59",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A0",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"24",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"98",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"A0",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"8A",X"65",X"55",X"55",X"A9",X"55",X"55",X"55",X"22",X"95",X"55",X"56",X"24",X"95",X"55",X"55",
		X"48",X"55",X"59",X"92",X"82",X"55",X"55",X"55",X"52",X"95",X"56",X"28",X"2A",X"A5",X"55",X"55",
		X"56",X"55",X"55",X"41",X"4A",X"95",X"55",X"55",X"55",X"55",X"55",X"41",X"16",X"95",X"55",X"55",
		X"55",X"55",X"55",X"26",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"A5",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"52",X"95",X"2A",X"AA",X"A5",X"AA",X"6A",X"55",X"49",X"98",X"8A",X"6A",X"69",X"AA",X"6A",
		X"55",X"AA",X"8A",X"AA",X"AA",X"A6",X"AA",X"A9",X"55",X"56",X"AA",X"AA",X"A6",X"AA",X"AA",X"A5",
		X"55",X"68",X"22",X"29",X"AA",X"AA",X"AA",X"85",X"55",X"4A",X"2A",X"AA",X"AA",X"9A",X"AA",X"A5",
		X"55",X"92",X"2A",X"AA",X"6A",X"AA",X"AA",X"25",X"55",X"68",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",
		X"56",X"82",X"AA",X"AA",X"9A",X"AA",X"99",X"95",X"55",X"2A",X"AA",X"AA",X"A6",X"AA",X"A2",X"55",
		X"56",X"8A",X"66",X"AA",X"9A",X"AA",X"99",X"55",X"5A",X"A9",X"9A",X"A9",X"5A",X"AA",X"69",X"55",
		X"59",X"69",X"55",X"59",X"6A",X"AA",X"95",X"56",X"55",X"65",X"55",X"55",X"56",X"A6",X"95",X"55",
		X"99",X"55",X"69",X"55",X"59",X"AA",X"55",X"5A",X"55",X"55",X"69",X"55",X"55",X"56",X"55",X"55",
		X"AA",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"5A",X"95",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"59",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"A6",X"9A",X"55",X"55",X"55",X"55",X"55",X"5A",X"5A",X"AA",X"55",X"55",X"55",X"55",X"55",
		X"69",X"9A",X"AA",X"95",X"55",X"55",X"55",X"55",X"59",X"5A",X"A8",X"A5",X"55",X"55",X"55",X"55",
		X"59",X"5A",X"A8",X"A5",X"55",X"55",X"55",X"55",X"59",X"AA",X"A8",X"A5",X"55",X"55",X"55",X"55",
		X"65",X"6A",X"AA",X"25",X"55",X"55",X"55",X"55",X"95",X"AA",X"AA",X"29",X"55",X"55",X"55",X"55",
		X"56",X"5A",X"AA",X"29",X"55",X"55",X"55",X"55",X"55",X"A9",X"AA",X"A9",X"55",X"55",X"55",X"55",
		X"96",X"AA",X"A8",X"A9",X"55",X"55",X"55",X"55",X"69",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",
		X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"25",X"55",X"55",
		X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"42",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"45",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"4A",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"48",
		X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"8A",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"8A",
		X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"AA",
		X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"AA",X"55",X"55",X"55",X"66",X"54",X"55",X"55",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"55",X"55",X"55",X"A6",X"55",X"55",X"59",X"AA",
		X"55",X"55",X"56",X"95",X"55",X"55",X"56",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"66",X"A9",
		X"A9",X"A6",X"AA",X"65",X"55",X"55",X"55",X"55",X"A5",X"A9",X"21",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"29",X"55",X"55",X"55",X"55",X"55",X"A5",X"AA",X"85",X"55",X"55",X"55",X"55",X"55",
		X"A9",X"AA",X"A9",X"55",X"55",X"55",X"55",X"55",X"A9",X"AA",X"15",X"55",X"55",X"55",X"55",X"55",
		X"9A",X"AA",X"16",X"55",X"55",X"55",X"55",X"55",X"AA",X"A8",X"99",X"55",X"55",X"55",X"55",X"55",
		X"A9",X"A8",X"99",X"55",X"55",X"55",X"55",X"55",X"A9",X"A0",X"95",X"65",X"55",X"55",X"55",X"55",
		X"A6",X"A0",X"59",X"65",X"55",X"55",X"55",X"55",X"6A",X"21",X"56",X"55",X"55",X"55",X"55",X"55",
		X"66",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"09",X"56",X"55",X"55",X"55",X"55",X"55",
		X"69",X"A9",X"55",X"65",X"55",X"55",X"55",X"55",X"9A",X"69",X"95",X"65",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"52",X"9A",
		X"55",X"41",X"59",X"55",X"55",X"55",X"56",X"25",X"55",X"15",X"56",X"6A",X"55",X"55",X"5A",X"55",
		X"55",X"45",X"55",X"A5",X"65",X"55",X"51",X"65",X"55",X"55",X"55",X"95",X"55",X"55",X"6A",X"55",
		X"55",X"55",X"55",X"A5",X"55",X"55",X"65",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"5A",X"55",
		X"55",X"55",X"56",X"55",X"56",X"55",X"66",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"59",X"55",
		X"55",X"59",X"55",X"55",X"55",X"55",X"66",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"66",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"59",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"99",X"A5",X"55",X"55",
		X"55",X"55",X"59",X"55",X"96",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"65",
		X"55",X"55",X"56",X"55",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A6",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"99",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"A5",X"A8",X"89",X"55",X"55",X"55",X"55",X"55",X"55",X"62",X"A9",X"55",X"55",X"55",X"55",
		X"59",X"55",X"6A",X"85",X"55",X"55",X"55",X"55",X"55",X"65",X"59",X"85",X"55",X"55",X"55",X"55",
		X"55",X"65",X"56",X"A5",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A6",X"55",X"55",X"55",X"55",X"15",X"55",X"9A",X"A9",
		X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"95",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"58",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"66",X"A5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"AA",X"2A",X"55",X"55",X"55",X"55",X"55",X"55",X"9A",X"A5",X"55",X"58",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"A9",X"55",X"69",X"55",X"55",X"55",X"55",X"59",X"A9",X"96",X"56",X"15",X"55",X"55",X"55",
		X"55",X"A9",X"55",X"68",X"95",X"55",X"55",X"55",X"99",X"65",X"59",X"6A",X"95",X"55",X"55",X"55",
		X"55",X"65",X"56",X"6A",X"15",X"55",X"55",X"55",X"59",X"69",X"56",X"9A",X"15",X"55",X"55",X"55",
		X"55",X"65",X"69",X"69",X"A5",X"55",X"55",X"55",X"55",X"69",X"55",X"59",X"A5",X"55",X"55",X"55",
		X"55",X"65",X"55",X"56",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"59",X"55",X"55",
		X"55",X"5A",X"55",X"55",X"55",X"65",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"66",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"95",X"51",X"55",X"55",X"55",X"55",
		X"55",X"59",X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"45",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"66",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"96",X"55",X"55",X"55",
		X"6A",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"A6",X"55",X"55",X"55",X"96",X"55",X"55",X"95",
		X"5A",X"55",X"55",X"55",X"95",X"55",X"56",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"56",X"A5",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"95",X"55",
		X"55",X"59",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"55",
		X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"15",
		X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"69",X"56",X"95",
		X"55",X"55",X"54",X"95",X"56",X"29",X"54",X"15",X"55",X"51",X"58",X"A5",X"54",X"AA",X"58",X"15",
		X"55",X"52",X"61",X"A9",X"5A",X"A5",X"62",X"55",X"55",X"42",X"A5",X"56",X"6A",X"55",X"6A",X"55",
		X"55",X"49",X"AA",X"55",X"55",X"55",X"A1",X"55",X"50",X"AA",X"55",X"59",X"55",X"55",X"AA",X"95",
		X"58",X"A9",X"56",X"55",X"55",X"56",X"69",X"95",X"20",X"56",X"A5",X"55",X"55",X"5A",X"AA",X"A5",
		X"56",X"A9",X"55",X"55",X"55",X"6A",X"99",X"65",X"5A",X"55",X"55",X"55",X"55",X"55",X"59",X"59",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"51",X"55",
		X"55",X"55",X"59",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A4",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"15",X"55",X"55",X"55",
		X"55",X"5A",X"95",X"55",X"15",X"55",X"55",X"55",X"55",X"88",X"6A",X"55",X"15",X"55",X"55",X"55",
		X"55",X"A5",X"55",X"96",X"95",X"55",X"55",X"55",X"54",X"99",X"55",X"56",X"25",X"55",X"55",X"55",
		X"5A",X"A5",X"55",X"56",X"85",X"55",X"55",X"55",X"59",X"95",X"55",X"56",X"A5",X"55",X"55",X"55",
		X"55",X"95",X"55",X"5A",X"85",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"25",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5A",X"A5",X"55",X"55",X"55",X"55",X"55",X"15",X"69",X"85",X"55",X"55",X"55",
		X"55",X"56",X"55",X"89",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"95",X"55",X"55",X"55",
		X"AA",X"EA",X"B5",X"7A",X"B7",X"AA",X"FA",X"9D",X"AA",X"EA",X"D5",X"7A",X"B7",X"AA",X"FA",X"9D",
		X"AA",X"6A",X"D5",X"7A",X"B7",X"AA",X"FA",X"9F",X"AA",X"6A",X"D5",X"7A",X"B7",X"A9",X"FA",X"AB",
		X"AA",X"6A",X"D5",X"7A",X"B7",X"A9",X"FA",X"AA",X"AA",X"6A",X"D5",X"7E",X"B7",X"A9",X"FA",X"AA",
		X"6A",X"6A",X"D5",X"5E",X"B7",X"A9",X"FA",X"AA",X"62",X"48",X"D5",X"5C",X"B7",X"21",X"F8",X"88",
		X"40",X"40",X"F5",X"5C",X"37",X"01",X"C0",X"15",X"40",X"40",X"F5",X"5C",X"37",X"01",X"C0",X"15",
		X"40",X"40",X"35",X"5C",X"37",X"01",X"C0",X"1F",X"40",X"40",X"0F",X"FC",X"37",X"01",X"C0",X"1D",
		X"40",X"10",X"00",X"00",X"37",X"01",X"C0",X"75",X"40",X"14",X"00",X"00",X"0C",X"01",X"C0",X"75",
		X"00",X"35",X"00",X"00",X"0C",X"00",X"C0",X"75",X"00",X"35",X"55",X"55",X"5F",X"55",X"C0",X"75",
		X"00",X"3D",X"55",X"55",X"5F",X"55",X"D5",X"75",X"05",X"5F",X"FF",X"FF",X"FF",X"D5",X"55",X"75",
		X"57",X"FD",X"55",X"55",X"55",X"7F",X"FF",X"F5",X"FD",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"48",X"00",X"00",X"45",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"15",X"55",
		X"55",X"00",X"55",X"55",X"55",X"54",X"01",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"40",X"55",
		X"51",X"55",X"55",X"55",X"55",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",
		X"55",X"55",X"55",X"95",X"55",X"55",X"5A",X"66",X"55",X"59",X"56",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"59",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"59",X"56",X"59",X"55",X"A6",X"59",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"56",X"65",X"65",X"65",X"59",X"95",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"56",X"55",X"95",X"56",X"55",X"65",X"55",X"65",X"55",X"59",X"55",X"55",X"55",X"5A",
		X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"59",X"65",X"55",X"65",X"59",
		X"55",X"55",X"55",X"55",X"56",X"56",X"55",X"55",X"55",X"55",X"5A",X"56",X"65",X"65",X"95",X"55",
		X"55",X"55",X"55",X"65",X"95",X"55",X"95",X"55",X"55",X"55",X"95",X"55",X"56",X"55",X"55",X"55",
		X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"65",X"56",X"95",X"55",X"55",X"55",X"55",
		X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"A9",X"95",X"55",X"55",X"55",X"54",X"95",X"56",X"A6",X"95",X"56",X"55",X"55",
		X"59",X"55",X"5A",X"AA",X"55",X"52",X"55",X"55",X"55",X"55",X"56",X"68",X"95",X"55",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"A2",X"55",X"55",X"55",X"55",
		X"55",X"55",X"64",X"AA",X"95",X"55",X"55",X"55",X"55",X"55",X"A6",X"62",X"95",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"66",X"95",X"55",X"55",X"55",X"55",X"56",X"A2",X"AA",X"65",X"55",X"55",X"55",
		X"55",X"5A",X"A9",X"99",X"99",X"55",X"55",X"55",X"55",X"55",X"99",X"A9",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"69",X"55",X"55",X"55",X"55",X"55",X"56",X"59",X"55",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"95",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"41",X"55",X"55",X"55",X"FC",X"15",X"55",X"54",X"15",X"55",X"55",X"55",X"57",X"C1",X"55",
		X"51",X"55",X"5A",X"AA",X"AA",X"55",X"7C",X"55",X"45",X"56",X"AA",X"AA",X"AA",X"A9",X"57",X"15",
		X"15",X"6A",X"AA",X"AA",X"AA",X"AA",X"A5",X"C5",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"71",
		X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"71",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9C",
		X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9C",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9D",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AC",X"3A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"90",
		X"0E",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"41",X"40",X"EA",X"AA",X"AA",X"AA",X"AA",X"A8",X"05",
		X"50",X"0E",X"AA",X"AA",X"AA",X"AB",X"00",X"15",X"55",X"00",X"3E",X"AA",X"AB",X"C0",X"01",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"44",X"00",X"00",X"45",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"15",X"55",
		X"55",X"00",X"55",X"55",X"55",X"54",X"01",X"55",X"50",X"15",X"55",X"55",X"55",X"55",X"40",X"15",
		X"41",X"55",X"55",X"55",X"55",X"55",X"54",X"05",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"01",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",
		X"55",X"55",X"55",X"55",X"59",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"96",X"59",X"99",X"56",
		X"55",X"55",X"55",X"55",X"55",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"55",X"9A",X"55",X"55",X"95",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"15",X"55",
		X"55",X"59",X"55",X"55",X"55",X"55",X"51",X"55",X"59",X"65",X"95",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"66",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"55",X"40",
		X"55",X"55",X"54",X"15",X"55",X"55",X"54",X"15",X"55",X"55",X"41",X"55",X"55",X"55",X"41",X"54",
		X"55",X"54",X"15",X"55",X"55",X"F4",X"15",X"57",X"55",X"41",X"55",X"55",X"57",X"D1",X"53",X"55",
		X"54",X"15",X"55",X"55",X"5F",X"45",X"5D",X"55",X"41",X"55",X"55",X"55",X"7D",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"00",X"00",X"15",
		X"45",X"55",X"55",X"00",X"55",X"55",X"55",X"55",X"51",X"55",X"50",X"05",X"55",X"55",X"55",X"55",
		X"54",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"07",X"55",X"55",X"55",X"5D",X"05",X"55",
		X"05",X"41",X"FF",X"FF",X"FF",X"F4",X"15",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",
		X"55",X"54",X"3F",X"FF",X"FF",X"C1",X"55",X"55",X"D5",X"55",X"10",X"00",X"00",X"45",X"55",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",
		X"55",X"55",X"70",X"00",X"00",X"D5",X"55",X"05",X"55",X"5C",X"05",X"55",X"55",X"03",X"55",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"15",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"54",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"55",X"40",X"55",X"55",
		X"55",X"54",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"4A",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"62",X"95",X"55",X"65",X"55",X"55",
		X"55",X"55",X"2A",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"99",X"85",X"55",X"55",X"55",X"55",
		X"55",X"6A",X"99",X"89",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"21",X"55",X"55",X"55",X"55",
		X"55",X"59",X"9A",X"A9",X"55",X"55",X"55",X"55",X"55",X"6A",X"A6",X"9A",X"55",X"55",X"55",X"55",
		X"55",X"56",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"65",X"55",X"55",X"55",X"55",
		X"55",X"5A",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"9A",X"95",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"66",X"5A",X"15",X"55",X"55",X"55",X"55",X"55",
		X"59",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"A2",X"95",X"A5",X"55",X"55",X"55",
		X"55",X"56",X"16",X"A5",X"5A",X"95",X"55",X"55",X"55",X"58",X"55",X"59",X"56",X"55",X"55",X"55",
		X"55",X"52",X"95",X"55",X"85",X"55",X"55",X"55",X"55",X"66",X"55",X"58",X"99",X"55",X"55",X"55",
		X"55",X"5A",X"55",X"54",X"15",X"96",X"55",X"55",X"55",X"6A",X"55",X"50",X"55",X"55",X"A6",X"A5",
		X"55",X"19",X"55",X"69",X"55",X"55",X"59",X"55",X"55",X"A9",X"55",X"68",X"55",X"55",X"55",X"95",
		X"55",X"89",X"55",X"61",X"55",X"51",X"59",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"51",X"86",X"9A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"05",X"55",X"55",X"65",X"65",X"56",
		X"55",X"55",X"15",X"55",X"55",X"55",X"5A",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",
		X"51",X"55",X"55",X"59",X"56",X"6A",X"55",X"55",X"45",X"55",X"66",X"56",X"AA",X"95",X"65",X"55",
		X"55",X"55",X"55",X"5A",X"55",X"55",X"65",X"55",X"55",X"55",X"AA",X"A5",X"55",X"55",X"65",X"55",
		X"55",X"6A",X"55",X"55",X"55",X"55",X"59",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"65",X"55",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"41",X"55",X"55",X"55",X"59",X"5A",X"A5",
		X"55",X"45",X"55",X"5A",X"AA",X"AA",X"A6",X"A5",X"65",X"55",X"55",X"55",X"AA",X"55",X"55",X"55",
		X"56",X"5A",X"AA",X"95",X"55",X"55",X"55",X"55",X"AA",X"A9",X"55",X"59",X"55",X"55",X"55",X"55",
		X"95",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"54",
		X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"7C",X"01",X"55",X"55",X"F5",X"55",X"55",X"55",X"5F",X"FC",X"00",X"15",X"C0",X"05",X"55",X"55",
		X"55",X"5F",X"FF",X"C7",X"D5",X"50",X"01",X"55",X"55",X"55",X"55",X"FF",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"7F",X"F5",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"10",X"55",X"55",X"50",
		X"55",X"55",X"55",X"55",X"15",X"01",X"55",X"50",X"55",X"55",X"00",X"1D",X"10",X"55",X"55",X"50",
		X"00",X"00",X"15",X"5D",X"15",X"55",X"55",X"54",X"15",X"55",X"55",X"5D",X"15",X"5F",X"C1",X"54",
		X"15",X"55",X"55",X"5F",X"57",X"FC",X"15",X"55",X"C5",X"55",X"55",X"57",X"7F",X"01",X"55",X"55",
		X"71",X"55",X"55",X"57",X"C0",X"55",X"55",X"55",X"5C",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",
		X"55",X"41",X"55",X"55",X"55",X"54",X"15",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"41",X"55",
		X"51",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"15",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"74",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"35",X"55",X"55",X"55",X"55",X"55",X"55",X"41",
		X"0D",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"40",X"D5",X"55",X"55",X"55",X"55",X"50",X"15",
		X"50",X"0D",X"55",X"55",X"55",X"57",X"00",X"55",X"55",X"00",X"1D",X"55",X"57",X"40",X"05",X"55",
		X"15",X"55",X"55",X"54",X"55",X"54",X"01",X"55",X"45",X"55",X"00",X"54",X"00",X"01",X"55",X"55",
		X"54",X"00",X"55",X"54",X"15",X"55",X"55",X"55",X"55",X"55",X"7F",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"FF",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"44",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"01",X"55",X"05",X"55",X"55",X"45",X"55",X"55",X"55",
		X"55",X"F0",X"55",X"55",X"45",X"55",X"55",X"55",X"54",X"5F",X"01",X"55",X"45",X"55",X"55",X"55",
		X"51",X"55",X"FC",X"05",X"45",X"55",X"55",X"55",X"45",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"59",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"69",X"9A",X"55",X"55",X"55",X"55",X"55",X"65",X"A5",X"A6",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"96",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"A6",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"55",
		X"55",X"55",X"56",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"65",X"55",X"A5",X"55",X"48",X"24",X"14",X"56",X"65",X"55",X"65",X"55",X"48",X"54",X"90",
		X"56",X"95",X"56",X"95",X"55",X"54",X"56",X"55",X"56",X"95",X"56",X"95",X"55",X"54",X"1A",X"55",
		X"56",X"55",X"56",X"55",X"55",X"54",X"99",X"55",X"56",X"55",X"5A",X"55",X"55",X"50",X"59",X"05",
		X"55",X"55",X"59",X"56",X"55",X"42",X"69",X"55",X"55",X"55",X"59",X"58",X"55",X"21",X"45",X"45",
		X"55",X"55",X"69",X"61",X"55",X"01",X"95",X"05",X"55",X"55",X"AA",X"61",X"54",X"45",X"15",X"41",
		X"55",X"56",X"9A",X"A5",X"55",X"46",X"16",X"95",X"55",X"55",X"AA",X"65",X"54",X"14",X"56",X"55",
		X"55",X"55",X"A6",X"95",X"54",X"52",X"55",X"55",X"55",X"55",X"96",X"55",X"54",X"52",X"55",X"56",
		X"55",X"56",X"AA",X"55",X"54",X"5A",X"55",X"55",X"55",X"56",X"A5",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"59",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",
		X"55",X"56",X"AA",X"95",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"69",
		X"55",X"55",X"55",X"5A",X"A5",X"55",X"5A",X"95",X"55",X"55",X"55",X"55",X"55",X"AA",X"55",X"55",
		X"5C",X"55",X"55",X"55",X"75",X"55",X"F5",X"55",X"57",X"15",X"55",X"40",X"FC",X"15",X"D5",X"55",
		X"55",X"C5",X"54",X"3F",X"57",X"C5",X"55",X"55",X"55",X"71",X"43",X"D5",X"55",X"F1",X"55",X"F5",
		X"55",X"5C",X"3D",X"55",X"55",X"7C",X"55",X"D5",X"55",X"57",X"D5",X"55",X"55",X"5F",X"05",X"55",
		X"55",X"55",X"55",X"55",X"55",X"57",X"F0",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"51",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"5F",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"50",X"05",X"00",X"01",X"00",X"55",X"55",X"55",X"55",X"50",X"05",X"00",X"55",X"55",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"50",X"55",
		X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"15",X"55",X"44",X"00",X"01",X"15",X"55",X"45",
		X"55",X"55",X"15",X"55",X"55",X"45",X"55",X"51",X"55",X"54",X"57",X"FF",X"FD",X"51",X"55",X"54",
		X"5D",X"51",X"55",X"55",X"55",X"54",X"57",X"55",X"D5",X"45",X"55",X"55",X"55",X"55",X"15",X"55",
		X"70",X"17",X"FF",X"FF",X"FF",X"FD",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"15",X"75",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"54",X"05",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"FF",X"FF",X"FF",X"FF",X"F5",
		X"55",X"55",X"7E",X"AA",X"AA",X"AA",X"A5",X"D5",X"F5",X"55",X"7A",X"AA",X"AA",X"AA",X"A5",X"D5",
		X"BD",X"55",X"7A",X"AA",X"AA",X"AA",X"97",X"55",X"AD",X"55",X"7A",X"AA",X"AA",X"AA",X"97",X"55",
		X"AB",X"55",X"7A",X"AA",X"AA",X"AA",X"97",X"55",X"69",X"D5",X"7A",X"AA",X"55",X"6A",X"5D",X"55",
		X"A9",X"D5",X"7E",X"AA",X"7F",X"EA",X"5D",X"55",X"A9",X"F5",X"5E",X"AA",X"75",X"EA",X"5D",X"55",
		X"E9",X"B5",X"5F",X"AA",X"9D",X"EA",X"75",X"55",X"A9",X"9D",X"57",X"AA",X"9D",X"EA",X"75",X"55",
		X"56",X"9D",X"55",X"EA",X"A5",X"AA",X"75",X"55",X"7A",X"97",X"55",X"EA",X"A5",X"AA",X"75",X"55",
		X"7A",X"A7",X"55",X"7A",X"A9",X"AA",X"75",X"55",X"5E",X"A7",X"55",X"7A",X"A9",X"AA",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"BF",X"FF",X"FD",
		X"FF",X"D5",X"55",X"7F",X"AF",X"AA",X"9E",X"AF",X"AB",X"55",X"55",X"FA",X"AF",X"AA",X"9E",X"AA",
		X"AB",X"55",X"57",X"EA",X"B7",X"AA",X"BE",X"AA",X"AD",X"55",X"5E",X"AA",X"B5",X"AA",X"76",X"AA",
		X"AA",X"6A",X"A6",X"AA",X"B6",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"AA",X"BA",X"AA",X"AA",X"55",
		X"56",X"55",X"69",X"6A",X"69",X"A9",X"56",X"6A",X"AA",X"6A",X"AA",X"69",X"A5",X"AA",X"AA",X"66",
		X"56",X"55",X"6A",X"69",X"AA",X"A9",X"56",X"67",X"A6",X"6A",X"AA",X"6A",X"95",X"AA",X"DE",X"6A",
		X"A5",X"F5",X"56",X"59",X"75",X"56",X"DE",X"65",X"AA",X"EA",X"AF",X"7A",X"B7",X"AA",X"DE",X"A7",
		X"AA",X"EA",X"AD",X"7A",X"B7",X"AA",X"FA",X"A7",X"AA",X"EA",X"B5",X"7A",X"B7",X"AA",X"FA",X"9D",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"7E",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",
		X"55",X"FA",X"AA",X"AA",X"AA",X"B6",X"AA",X"AA",X"57",X"6A",X"AA",X"AA",X"AA",X"B6",X"AA",X"AA",
		X"5D",X"6A",X"AA",X"AA",X"AA",X"B6",X"AA",X"5A",X"5D",X"6A",X"AA",X"AA",X"AA",X"B5",X"AA",X"5A",
		X"5D",X"6A",X"AA",X"AA",X"AA",X"B5",X"55",X"59",X"5D",X"6A",X"A9",X"55",X"6A",X"BD",X"FF",X"5A",
		X"5D",X"5A",X"AB",X"FF",X"5A",X"AD",X"AA",X"99",X"5D",X"5A",X"AA",X"B5",X"DA",X"AD",X"A9",X"6A",
		X"57",X"56",X"AA",X"B5",X"DA",X"AD",X"A9",X"56",X"55",X"D5",X"AA",X"AF",X"DA",X"AD",X"6A",X"AA",
		X"55",X"75",X"6A",X"AA",X"D6",X"AD",X"6A",X"AA",X"55",X"5D",X"5A",X"AA",X"D6",X"AF",X"6A",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"49",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"56",X"95",X"25",X"55",X"55",X"55",X"55",X"A9",X"5A",X"96",X"45",X"55",X"55",X"55",X"55",
		X"A9",X"6A",X"55",X"85",X"55",X"55",X"55",X"55",X"99",X"5A",X"56",X"25",X"55",X"55",X"55",X"55",
		X"99",X"5A",X"96",X"85",X"55",X"55",X"55",X"55",X"A9",X"9A",X"9A",X"A9",X"55",X"55",X"55",X"55",
		X"A6",X"95",X"96",X"21",X"55",X"55",X"55",X"55",X"66",X"55",X"90",X"A8",X"55",X"55",X"55",X"55",
		X"6A",X"55",X"58",X"8A",X"55",X"55",X"55",X"55",X"65",X"95",X"52",X"19",X"55",X"55",X"55",X"55",
		X"55",X"55",X"40",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"48",X"AA",X"55",X"55",X"55",X"55",
		X"55",X"55",X"62",X"86",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"26",X"95",X"55",X"55",X"55",
		X"55",X"55",X"6A",X"1A",X"95",X"55",X"55",X"55",X"55",X"55",X"AA",X"9A",X"A5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"58",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"05",X"55",X"55",
		X"55",X"55",X"55",X"55",X"66",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"85",X"55",X"55",
		X"55",X"55",X"55",X"55",X"6A",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"45",X"55",X"55",
		X"55",X"55",X"55",X"56",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"69",X"9A",X"45",X"55",
		X"55",X"55",X"55",X"55",X"6A",X"6A",X"62",X"55",X"55",X"55",X"55",X"55",X"95",X"5A",X"9A",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",
		X"55",X"55",X"55",X"55",X"56",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"56",X"AA",X"96",X"AB",X"55",X"55",X"55",X"55",X"D5",X"AA",X"A6",X"AB",X"7F",X"FD",
		X"55",X"55",X"75",X"6A",X"AA",X"AB",X"55",X"5D",X"55",X"55",X"5D",X"56",X"AA",X"AB",X"55",X"5D",
		X"55",X"55",X"57",X"56",X"AA",X"AB",X"55",X"5D",X"55",X"55",X"55",X"D6",X"AA",X"AB",X"55",X"5D",
		X"55",X"55",X"55",X"DA",X"AA",X"AB",X"55",X"57",X"55",X"55",X"55",X"D2",X"22",X"22",X"D5",X"57",
		X"55",X"55",X"55",X"D0",X"00",X"00",X"D5",X"57",X"55",X"55",X"55",X"D0",X"01",X"40",X"D5",X"57",
		X"55",X"55",X"57",X"40",X"05",X"40",X"D5",X"57",X"55",X"55",X"57",X"40",X"0F",X"40",X"D5",X"57",
		X"55",X"55",X"57",X"40",X"37",X"40",X"D5",X"57",X"55",X"55",X"57",X"40",X"37",X"40",X"3F",X"FF",
		X"55",X"55",X"57",X"40",X"D7",X"50",X"30",X"00",X"55",X"55",X"57",X"40",X"D5",X"D0",X"30",X"00",
		X"5E",X"A7",X"55",X"5E",X"A5",X"A9",X"75",X"55",X"5E",X"A7",X"55",X"7E",X"AA",X"A9",X"75",X"55",
		X"5E",X"A7",X"55",X"FA",X"AA",X"A9",X"75",X"55",X"FE",X"A7",X"55",X"EA",X"AA",X"A9",X"75",X"55",
		X"AA",X"A7",X"57",X"EA",X"AA",X"A9",X"D5",X"55",X"AA",X"A7",X"57",X"AA",X"AA",X"A9",X"D5",X"55",
		X"AA",X"9D",X"5F",X"AA",X"AA",X"A5",X"D5",X"55",X"22",X"1D",X"5E",X"22",X"58",X"85",X"D5",X"55",
		X"00",X"1D",X"7C",X"01",X"50",X"05",X"D5",X"55",X"50",X"1D",X"70",X"05",X"70",X"05",X"D5",X"55",
		X"F0",X"1D",X"F0",X"15",X"F0",X"05",X"D5",X"55",X"70",X"1D",X"C0",X"57",X"70",X"05",X"D5",X"55",
		X"70",X"1F",X"C1",X"5D",X"70",X"05",X"D5",X"55",X"70",X"1F",X"05",X"75",X"C0",X"07",X"55",X"55",
		X"C0",X"1C",X"15",X"D5",X"C0",X"17",X"55",X"55",X"C0",X"50",X"17",X"55",X"C0",X"17",X"55",X"55",
		X"55",X"55",X"A8",X"94",X"65",X"55",X"55",X"55",X"55",X"55",X"6A",X"54",X"95",X"55",X"55",X"55",
		X"55",X"55",X"68",X"54",X"95",X"55",X"55",X"55",X"55",X"55",X"26",X"55",X"95",X"55",X"55",X"55",
		X"55",X"55",X"99",X"52",X"55",X"55",X"55",X"55",X"55",X"56",X"A5",X"99",X"55",X"55",X"55",X"55",
		X"55",X"55",X"A2",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"89",X"96",X"95",X"55",X"55",X"55",
		X"55",X"54",X"89",X"95",X"65",X"55",X"55",X"55",X"55",X"5A",X"2A",X"95",X"55",X"55",X"55",X"55",
		X"55",X"59",X"A9",X"95",X"55",X"55",X"55",X"55",X"55",X"6A",X"95",X"65",X"55",X"55",X"55",X"55",
		X"55",X"A9",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"54",X"55",X"55",X"55",X"55",X"56",X"95",
		X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"69",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"55",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"95",X"59",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"59",X"56",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"95",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"65",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"65",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"56",X"55",X"55",X"55",X"55",
		X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"56",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"69",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"56",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",
		X"55",X"55",X"55",X"55",X"55",X"66",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"95",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"40",X"5D",X"55",X"C0",X"17",X"55",X"55",X"55",X"41",X"5D",X"55",X"C0",X"17",X"55",X"55",
		X"F5",X"05",X"75",X"57",X"00",X"17",X"55",X"55",X"5F",X"05",X"D5",X"57",X"00",X"17",X"55",X"55",
		X"55",X"05",X"D5",X"57",X"00",X"17",X"55",X"55",X"55",X"17",X"55",X"57",X"00",X"17",X"55",X"55",
		X"55",X"17",X"55",X"5D",X"00",X"17",X"55",X"55",X"55",X"F7",X"55",X"5D",X"40",X"17",X"55",X"55",
		X"57",X"FD",X"55",X"57",X"D5",X"07",X"55",X"55",X"57",X"F5",X"55",X"55",X"F5",X"57",X"55",X"55",
		X"57",X"F5",X"55",X"55",X"5F",X"57",X"55",X"55",X"57",X"D5",X"55",X"55",X"55",X"FF",X"D5",X"55",
		X"55",X"D5",X"55",X"55",X"55",X"57",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"59",X"55",X"99",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"59",X"55",X"55",X"55",X"55",X"54",X"55",
		X"55",X"55",X"59",X"55",X"55",X"56",X"55",X"55",X"65",X"65",X"65",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"55",X"55",X"56",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"59",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"59",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"59",X"55",X"55",X"55",X"55",X"65",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"99",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"56",X"D9",X"55",X"55",X"55",
		X"55",X"65",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"55",X"65",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"65",X"65",X"55",X"55",X"55",X"59",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"95",X"65",X"59",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"69",X"55",X"55",X"55",X"55",X"55",
		X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"66",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"5D",X"03",X"55",X"D0",X"30",X"00",X"55",X"55",X"5D",X"03",X"55",X"D0",X"00",X"00",
		X"55",X"55",X"5D",X"03",X"55",X"D4",X"04",X"15",X"55",X"55",X"5D",X"0D",X"55",X"74",X"15",X"55",
		X"55",X"55",X"5D",X"0D",X"55",X"75",X"55",X"7F",X"55",X"55",X"5D",X"0D",X"55",X"75",X"5F",X"D5",
		X"55",X"55",X"5D",X"0D",X"55",X"75",X"F5",X"55",X"55",X"55",X"5D",X"35",X"55",X"FF",X"55",X"55",
		X"55",X"55",X"5D",X"35",X"55",X"D5",X"55",X"55",X"55",X"55",X"5F",X"35",X"55",X"55",X"55",X"55",
		X"55",X"55",X"5F",X"35",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"58",X"99",X"55",X"55",X"55",X"55",X"55",X"65",X"96",X"55",X"55",X"55",
		X"55",X"55",X"55",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"99",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"59",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"55",X"55",X"95",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"65",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"56",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"59",X"55",
		X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",
		X"55",X"65",X"96",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",
		X"65",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"55",X"95",X"55",X"55",X"55",X"55",X"59",X"55",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"59",
		X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"59",X"55",
		X"56",X"55",X"55",X"95",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"95",X"56",X"55",X"55",X"55",X"55",
		X"55",X"A1",X"56",X"55",X"55",X"55",X"55",X"55",X"59",X"85",X"65",X"55",X"55",X"55",X"55",X"55",
		X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"65",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"95",X"55",X"55",
		X"65",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"65",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"95",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"65",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"44",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"59",X"95",X"55",X"55",
		X"55",X"55",X"65",X"55",X"56",X"56",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"95",X"55",X"55",X"55",X"55",X"55",X"56",X"56",X"A5",X"55",X"55",X"55",X"55",X"55",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"D5",X"7D",X"5F",X"F5",X"55",X"55",X"55",X"5D",X"75",X"D7",X"55",X"D5",X"55",
		X"56",X"55",X"5D",X"75",X"D7",X"57",X"55",X"55",X"5A",X"55",X"5D",X"75",X"D7",X"5F",X"55",X"55",
		X"5A",X"95",X"5D",X"75",X"D7",X"5C",X"75",X"56",X"56",X"A5",X"57",X"D5",X"7D",X"57",X"D5",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"D5",X"7D",X"57",X"F5",X"55",X"55",X"55",X"5D",X"75",X"D7",X"5D",X"55",X"55",
		X"56",X"55",X"5D",X"75",X"D7",X"5D",X"55",X"55",X"5A",X"55",X"5D",X"75",X"D7",X"57",X"D5",X"55",
		X"5A",X"95",X"5D",X"75",X"D7",X"5D",X"55",X"56",X"56",X"A5",X"57",X"D5",X"7D",X"5F",X"F5",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"D5",X"7D",X"5D",X"55",X"55",X"55",X"55",X"5D",X"75",X"D7",X"5D",X"55",X"55",
		X"56",X"55",X"5D",X"75",X"D7",X"5F",X"F5",X"55",X"5A",X"55",X"5D",X"75",X"D7",X"5D",X"D5",X"55",
		X"5A",X"95",X"5D",X"75",X"D7",X"5F",X"55",X"56",X"56",X"A5",X"57",X"D5",X"7D",X"5D",X"55",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"D5",X"7D",X"57",X"D5",X"55",X"55",X"55",X"5D",X"75",X"D7",X"5D",X"75",X"55",
		X"56",X"55",X"5D",X"75",X"D7",X"5D",X"75",X"55",X"5A",X"55",X"5D",X"75",X"D7",X"57",X"F5",X"55",
		X"5A",X"95",X"5D",X"75",X"D7",X"55",X"75",X"56",X"56",X"A5",X"57",X"D5",X"7D",X"5F",X"D5",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"D5",X"7D",X"57",X"D5",X"55",X"55",X"55",X"5D",X"75",X"D7",X"5D",X"75",X"55",
		X"56",X"55",X"5D",X"75",X"D7",X"5D",X"75",X"55",X"5A",X"55",X"5D",X"75",X"D7",X"57",X"D5",X"55",
		X"5A",X"95",X"5D",X"75",X"D7",X"5D",X"75",X"56",X"56",X"A5",X"57",X"D5",X"7D",X"57",X"D5",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"7D",X"57",X"D5",X"FF",X"5D",X"55",X"55",X"55",X"D7",X"5D",X"75",X"5D",X"5D",X"55",
		X"56",X"55",X"D7",X"5D",X"75",X"75",X"5D",X"55",X"5A",X"55",X"D7",X"5D",X"75",X"F5",X"5F",X"55",
		X"5A",X"95",X"D7",X"5D",X"75",X"D7",X"5D",X"56",X"56",X"A5",X"7D",X"57",X"D5",X"7D",X"5D",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"7D",X"57",X"D5",X"7D",X"5D",X"55",X"55",X"55",X"D7",X"5D",X"75",X"D7",X"5D",X"55",
		X"56",X"55",X"D7",X"5D",X"75",X"D7",X"5D",X"55",X"5A",X"55",X"D7",X"5D",X"75",X"7F",X"5F",X"55",
		X"5A",X"95",X"D7",X"5D",X"75",X"57",X"5D",X"56",X"56",X"A5",X"7D",X"57",X"D5",X"FD",X"5D",X"5A",
		X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"A9",X"55",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",X"55",X"55",X"56",X"6A",X"AA",X"A6",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
