library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog_rom_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog_rom_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"02",X"85",X"06",X"98",X"7D",X"8C",X"02",X"C9",X"18",X"90",X"08",X"F0",X"04",X"A9",X"17",X"D0",
		X"02",X"A9",X"00",X"9D",X"8C",X"02",X"85",X"07",X"BD",X"00",X"02",X"A0",X"E0",X"4A",X"B0",X"07",
		X"A0",X"F0",X"4A",X"B0",X"02",X"A0",X"00",X"20",X"FE",X"72",X"4C",X"5E",X"6F",X"AD",X"F8",X"02",
		X"8D",X"F7",X"02",X"A9",X"00",X"8D",X"1C",X"02",X"8D",X"3F",X"02",X"8D",X"62",X"02",X"60",X"A5",
		X"1C",X"F0",X"42",X"AD",X"1B",X"02",X"30",X"3D",X"AD",X"FA",X"02",X"F0",X"39",X"CE",X"FA",X"02",
		X"D0",X"33",X"A4",X"59",X"30",X"19",X"D0",X"10",X"20",X"39",X"71",X"D0",X"24",X"AC",X"1C",X"02",
		X"F0",X"06",X"A0",X"02",X"8C",X"FA",X"02",X"60",X"A9",X"01",X"8D",X"1B",X"02",X"D0",X"12",X"A9",
		X"A0",X"8D",X"1B",X"02",X"A2",X"3E",X"86",X"69",X"A6",X"18",X"D6",X"57",X"A9",X"81",X"8D",X"FA",
		X"02",X"A9",X"00",X"85",X"59",X"60",X"AD",X"07",X"24",X"10",X"04",X"A9",X"03",X"D0",X"07",X"AD",
		X"06",X"24",X"10",X"07",X"A9",X"FD",X"18",X"65",X"61",X"85",X"61",X"A5",X"5C",X"4A",X"B0",X"E5",
		X"AD",X"05",X"24",X"10",X"3C",X"A9",X"80",X"8D",X"03",X"3C",X"A0",X"00",X"A5",X"61",X"20",X"D2",
		X"77",X"10",X"01",X"88",X"0A",X"18",X"65",X"64",X"AA",X"98",X"6D",X"3E",X"02",X"20",X"25",X"71",
		X"8D",X"3E",X"02",X"86",X"64",X"A0",X"00",X"A5",X"61",X"20",X"D5",X"77",X"10",X"01",X"88",X"0A",
		X"18",X"65",X"65",X"AA",X"98",X"6D",X"61",X"02",X"20",X"25",X"71",X"8D",X"61",X"02",X"86",X"65",
		X"60",X"A9",X"00",X"8D",X"03",X"3C",X"AD",X"3E",X"02",X"05",X"64",X"F0",X"18",X"AD",X"3E",X"02",
		X"0A",X"A2",X"FF",X"18",X"49",X"FF",X"30",X"02",X"E8",X"38",X"65",X"64",X"85",X"64",X"8A",X"6D",
		X"3E",X"02",X"8D",X"3E",X"02",X"A5",X"65",X"0D",X"61",X"02",X"F0",X"18",X"AD",X"61",X"02",X"0A",
		X"A2",X"FF",X"18",X"49",X"FF",X"30",X"02",X"38",X"E8",X"65",X"65",X"85",X"65",X"8A",X"6D",X"61",
		X"02",X"8D",X"61",X"02",X"60",X"30",X"09",X"C9",X"40",X"90",X"0D",X"A2",X"FF",X"A9",X"3F",X"60",
		X"C9",X"C0",X"B0",X"04",X"A2",X"01",X"A9",X"C0",X"60",X"A2",X"1C",X"BD",X"00",X"02",X"F0",X"1E",
		X"BD",X"69",X"02",X"38",X"ED",X"84",X"02",X"C9",X"04",X"90",X"04",X"C9",X"FC",X"90",X"0F",X"BD",
		X"8C",X"02",X"38",X"ED",X"A7",X"02",X"C9",X"04",X"90",X"09",X"C9",X"FC",X"B0",X"05",X"CA",X"10",
		X"DA",X"E8",X"60",X"EE",X"FA",X"02",X"60",X"90",X"A2",X"1A",X"AD",X"FB",X"02",X"D0",X"70",X"AD",
		X"1C",X"02",X"D0",X"73",X"8D",X"3F",X"02",X"8D",X"62",X"02",X"EE",X"FD",X"02",X"AD",X"FD",X"02",
		X"C9",X"0B",X"90",X"03",X"CE",X"FD",X"02",X"AD",X"F5",X"02",X"18",X"69",X"02",X"C9",X"0B",X"90",
		X"02",X"A9",X"0B",X"8D",X"F6",X"02",X"8D",X"F5",X"02",X"85",X"08",X"A0",X"1C",X"20",X"B5",X"77",
		X"29",X"18",X"09",X"04",X"9D",X"00",X"02",X"20",X"03",X"72",X"20",X"B5",X"77",X"4A",X"29",X"1F",
		X"90",X"13",X"C9",X"18",X"90",X"02",X"29",X"17",X"9D",X"8C",X"02",X"A9",X"00",X"9D",X"69",X"02",
		X"9D",X"AF",X"02",X"F0",X"0B",X"9D",X"69",X"02",X"A9",X"00",X"9D",X"8C",X"02",X"9D",X"D2",X"02",
		X"CA",X"C6",X"08",X"D0",X"C8",X"A9",X"7F",X"8D",X"F7",X"02",X"A9",X"30",X"8D",X"FC",X"02",X"A9",
		X"00",X"9D",X"00",X"02",X"CA",X"10",X"FA",X"60",X"A9",X"60",X"8D",X"CA",X"02",X"8D",X"ED",X"02",
		X"A9",X"00",X"8D",X"3E",X"02",X"8D",X"61",X"02",X"A9",X"10",X"8D",X"84",X"02",X"A9",X"0C",X"8D",
		X"A7",X"02",X"60",X"20",X"B5",X"77",X"29",X"8F",X"10",X"02",X"09",X"F0",X"18",X"79",X"23",X"02",
		X"20",X"33",X"72",X"9D",X"23",X"02",X"20",X"B5",X"77",X"20",X"B5",X"77",X"20",X"B5",X"77",X"20",
		X"B5",X"77",X"29",X"8F",X"10",X"02",X"09",X"F0",X"18",X"79",X"46",X"02",X"20",X"33",X"72",X"9D",
		X"46",X"02",X"60",X"10",X"0D",X"C9",X"E1",X"B0",X"02",X"A9",X"E1",X"C9",X"FB",X"90",X"0F",X"A9",
		X"FA",X"60",X"C9",X"06",X"B0",X"02",X"A9",X"06",X"C9",X"20",X"90",X"02",X"A9",X"1F",X"60",X"A9",
		X"10",X"85",X"00",X"A9",X"50",X"A2",X"A4",X"20",X"FC",X"7B",X"A9",X"19",X"A2",X"DB",X"20",X"03",
		X"7C",X"A9",X"70",X"20",X"DE",X"7C",X"A2",X"00",X"A5",X"1C",X"C9",X"02",X"D0",X"18",X"A5",X"18",
		X"D0",X"14",X"A2",X"20",X"AD",X"1B",X"02",X"05",X"59",X"D0",X"0B",X"AD",X"FA",X"02",X"30",X"06",
		X"A5",X"5C",X"29",X"10",X"F0",X"0D",X"A9",X"52",X"A0",X"02",X"38",X"20",X"3F",X"77",X"A9",X"00",
		X"20",X"8B",X"77",X"A9",X"28",X"A4",X"57",X"20",X"3E",X"6F",X"A9",X"00",X"85",X"00",X"A9",X"78",
		X"A2",X"DB",X"20",X"03",X"7C",X"A9",X"50",X"20",X"DE",X"7C",X"A9",X"1D",X"A0",X"02",X"38",X"20",
		X"3F",X"77",X"A9",X"00",X"20",X"D1",X"7B",X"A9",X"10",X"85",X"00",X"A9",X"C0",X"A2",X"DB",X"20",
		X"03",X"7C",X"A9",X"50",X"20",X"DE",X"7C",X"A2",X"00",X"A5",X"1C",X"C9",X"01",X"F0",X"2E",X"90",
		X"18",X"A5",X"18",X"F0",X"14",X"A2",X"20",X"AD",X"1B",X"02",X"05",X"59",X"D0",X"0B",X"AD",X"FA",
		X"02",X"30",X"06",X"A5",X"5C",X"29",X"10",X"F0",X"0D",X"A9",X"54",X"A0",X"02",X"38",X"20",X"3F",
		X"77",X"A9",X"00",X"20",X"8B",X"77",X"A9",X"CF",X"A4",X"58",X"4C",X"3E",X"6F",X"60",X"84",X"00",
		X"86",X"0D",X"A5",X"05",X"4A",X"66",X"04",X"4A",X"66",X"04",X"4A",X"66",X"04",X"85",X"05",X"A5",
		X"07",X"18",X"69",X"04",X"4A",X"66",X"06",X"4A",X"66",X"06",X"4A",X"66",X"06",X"85",X"07",X"A2",
		X"04",X"20",X"1C",X"7C",X"A9",X"70",X"38",X"E5",X"00",X"C9",X"A0",X"90",X"0E",X"48",X"A9",X"90",
		X"20",X"DE",X"7C",X"68",X"38",X"E9",X"10",X"C9",X"A0",X"B0",X"F2",X"20",X"DE",X"7C",X"A6",X"0D",
		X"BD",X"00",X"02",X"10",X"16",X"E0",X"1B",X"F0",X"0C",X"29",X"0C",X"4A",X"A8",X"B9",X"F8",X"50",
		X"BE",X"F9",X"50",X"D0",X"1B",X"20",X"65",X"74",X"A6",X"0D",X"60",X"E0",X"1B",X"F0",X"17",X"E0",
		X"1C",X"F0",X"19",X"B0",X"1F",X"29",X"18",X"4A",X"4A",X"A8",X"B9",X"DE",X"51",X"BE",X"DF",X"51",
		X"20",X"45",X"7D",X"A6",X"0D",X"60",X"20",X"0B",X"75",X"A6",X"0D",X"60",X"AD",X"50",X"52",X"AE",
		X"51",X"52",X"D0",X"EC",X"A9",X"70",X"A2",X"F0",X"20",X"E0",X"7C",X"A6",X"0D",X"A5",X"5C",X"29",
		X"03",X"D0",X"03",X"DE",X"00",X"02",X"60",X"F8",X"75",X"52",X"95",X"52",X"90",X"12",X"B5",X"53",
		X"69",X"00",X"95",X"53",X"29",X"0F",X"D0",X"08",X"A9",X"B0",X"85",X"68",X"A6",X"18",X"F6",X"57",
		X"D8",X"60",X"A5",X"18",X"0A",X"0A",X"85",X"08",X"A5",X"6F",X"29",X"FB",X"05",X"08",X"85",X"6F",
		X"8D",X"00",X"32",X"60",X"A5",X"1C",X"F0",X"02",X"18",X"60",X"A5",X"5D",X"29",X"04",X"D0",X"F8",
		X"A5",X"1D",X"05",X"1E",X"F0",X"F2",X"A0",X"00",X"20",X"F6",X"77",X"A2",X"00",X"86",X"10",X"A9",
		X"01",X"85",X"00",X"A9",X"A7",X"85",X"0E",X"A9",X"10",X"85",X"00",X"B5",X"1D",X"15",X"1E",X"F0",
		X"67",X"86",X"0F",X"A9",X"5F",X"A6",X"0E",X"20",X"03",X"7C",X"A9",X"40",X"20",X"DE",X"7C",X"A5",
		X"0F",X"4A",X"F8",X"69",X"01",X"D8",X"85",X"0D",X"A9",X"0D",X"38",X"A0",X"01",X"A2",X"00",X"20",
		X"3F",X"77",X"A9",X"40",X"AA",X"20",X"E0",X"7C",X"A0",X"00",X"20",X"35",X"6F",X"A5",X"0F",X"18",
		X"69",X"1D",X"A0",X"02",X"38",X"A2",X"00",X"20",X"3F",X"77",X"A9",X"00",X"20",X"D1",X"7B",X"A0",
		X"00",X"20",X"35",X"6F",X"A4",X"10",X"20",X"1A",X"6F",X"E6",X"10",X"A4",X"10",X"20",X"1A",X"6F",
		X"E6",X"10",X"A4",X"10",X"20",X"1A",X"6F",X"E6",X"10",X"A5",X"0E",X"38",X"E9",X"08",X"85",X"0E",
		X"A6",X"0F",X"E8",X"E8",X"E0",X"14",X"90",X"93",X"38",X"60",X"A2",X"1A",X"BD",X"00",X"02",X"F0",
		X"03",X"CA",X"10",X"F8",X"60",X"AD",X"1B",X"02",X"C9",X"A2",X"B0",X"22",X"A2",X"0A",X"BD",X"EC",
		X"50",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"F8",X"49",X"F8",X"95",X"7E",X"BD",X"ED",X"50",X"4A",
		X"4A",X"4A",X"4A",X"18",X"69",X"F8",X"49",X"F8",X"95",X"8A",X"CA",X"CA",X"10",X"E0",X"AD",X"1B",
		X"02",X"49",X"FF",X"29",X"70",X"4A",X"4A",X"4A",X"AA",X"86",X"09",X"A0",X"00",X"BD",X"EC",X"50",
		X"10",X"01",X"88",X"18",X"75",X"7D",X"95",X"7D",X"98",X"75",X"7E",X"95",X"7E",X"85",X"04",X"84",
		X"05",X"A0",X"00",X"BD",X"ED",X"50",X"10",X"01",X"88",X"18",X"75",X"89",X"95",X"89",X"98",X"75",
		X"8A",X"95",X"8A",X"85",X"06",X"84",X"07",X"A5",X"02",X"85",X"0B",X"A5",X"03",X"85",X"0C",X"20",
		X"49",X"7C",X"A4",X"09",X"B9",X"E0",X"50",X"BE",X"E1",X"50",X"20",X"45",X"7D",X"A4",X"09",X"B9",
		X"E1",X"50",X"49",X"04",X"AA",X"B9",X"E0",X"50",X"29",X"0F",X"49",X"04",X"20",X"45",X"7D",X"A0",
		X"FF",X"C8",X"B1",X"0B",X"91",X"02",X"C8",X"B1",X"0B",X"49",X"04",X"91",X"02",X"C0",X"03",X"90",
		X"F0",X"20",X"39",X"7C",X"A6",X"09",X"CA",X"CA",X"10",X"8F",X"60",X"A2",X"00",X"86",X"17",X"A0",
		X"00",X"A5",X"61",X"10",X"06",X"A0",X"04",X"8A",X"38",X"E5",X"61",X"85",X"08",X"24",X"08",X"30",
		X"02",X"50",X"07",X"A2",X"04",X"A9",X"80",X"38",X"E5",X"08",X"86",X"08",X"84",X"09",X"4A",X"29",
		X"FE",X"A8",X"B9",X"6E",X"52",X"BE",X"6F",X"52",X"20",X"D3",X"6A",X"AD",X"05",X"24",X"10",X"14",
		X"A5",X"5C",X"29",X"04",X"F0",X"0E",X"C8",X"C8",X"38",X"A6",X"0C",X"98",X"65",X"0B",X"90",X"01",
		X"E8",X"20",X"D3",X"6A",X"60",X"A5",X"1C",X"D0",X"01",X"60",X"A2",X"00",X"AD",X"1C",X"02",X"30",
		X"0A",X"F0",X"08",X"6A",X"6A",X"6A",X"8D",X"02",X"3C",X"A2",X"80",X"8E",X"00",X"3C",X"A2",X"01",
		X"20",X"CD",X"75",X"8D",X"01",X"3C",X"CA",X"20",X"CD",X"75",X"8D",X"04",X"3C",X"AD",X"1B",X"02",
		X"C9",X"01",X"F0",X"04",X"8A",X"8D",X"03",X"3C",X"AD",X"F6",X"02",X"F0",X"11",X"AD",X"1B",X"02",
		X"30",X"0C",X"05",X"59",X"F0",X"08",X"A5",X"6D",X"F0",X"14",X"C6",X"6D",X"D0",X"21",X"A5",X"6C",
		X"29",X"0F",X"85",X"6C",X"8D",X"00",X"3A",X"AD",X"FC",X"02",X"85",X"6E",X"10",X"11",X"C6",X"6E",
		X"D0",X"0D",X"A9",X"04",X"85",X"6D",X"A5",X"6C",X"49",X"14",X"85",X"6C",X"8D",X"00",X"3A",X"A5",
		X"69",X"AA",X"29",X"3F",X"F0",X"01",X"CA",X"86",X"69",X"8E",X"00",X"36",X"60",X"B5",X"6A",X"30",
		X"0C",X"B5",X"66",X"10",X"12",X"A9",X"10",X"95",X"66",X"A9",X"80",X"30",X"0C",X"B5",X"66",X"F0",
		X"06",X"30",X"04",X"D6",X"66",X"D0",X"F2",X"A9",X"00",X"95",X"6A",X"60",X"86",X"0D",X"A9",X"50",
		X"8D",X"F9",X"02",X"B9",X"00",X"02",X"29",X"78",X"85",X"0E",X"B9",X"00",X"02",X"29",X"07",X"4A",
		X"AA",X"F0",X"02",X"05",X"0E",X"99",X"00",X"02",X"A5",X"1C",X"F0",X"11",X"A5",X"0D",X"F0",X"04",
		X"C9",X"04",X"90",X"09",X"BD",X"59",X"76",X"A6",X"19",X"18",X"20",X"97",X"73",X"BE",X"00",X"02",
		X"F0",X"34",X"20",X"5A",X"74",X"30",X"2F",X"EE",X"F6",X"02",X"20",X"9D",X"6A",X"20",X"03",X"72",
		X"BD",X"23",X"02",X"29",X"1F",X"0A",X"5D",X"AF",X"02",X"9D",X"AF",X"02",X"20",X"5C",X"74",X"30",
		X"15",X"EE",X"F6",X"02",X"20",X"9D",X"6A",X"20",X"03",X"72",X"BD",X"46",X"02",X"29",X"1F",X"0A",
		X"5D",X"D2",X"02",X"9D",X"D2",X"02",X"A6",X"0D",X"60",X"10",X"05",X"02",X"A5",X"1C",X"10",X"38",
		X"A2",X"02",X"85",X"5D",X"85",X"32",X"85",X"33",X"A0",X"00",X"B9",X"1D",X"00",X"D5",X"52",X"B9",
		X"1E",X"00",X"F5",X"53",X"90",X"23",X"C8",X"C8",X"C0",X"14",X"90",X"EE",X"CA",X"CA",X"10",X"E8",
		X"A5",X"33",X"30",X"0E",X"C5",X"32",X"90",X"0A",X"69",X"02",X"C9",X"1E",X"90",X"02",X"A9",X"FF",
		X"85",X"33",X"A9",X"00",X"85",X"1C",X"85",X"31",X"60",X"86",X"0B",X"84",X"0C",X"8A",X"4A",X"AA",
		X"98",X"4A",X"65",X"0C",X"85",X"0D",X"95",X"32",X"A2",X"1B",X"A0",X"12",X"E4",X"0D",X"F0",X"1F",
		X"B5",X"31",X"95",X"34",X"B5",X"32",X"95",X"35",X"B5",X"33",X"95",X"36",X"B9",X"1B",X"00",X"99",
		X"1D",X"00",X"B9",X"1C",X"00",X"99",X"1E",X"00",X"88",X"88",X"CA",X"CA",X"CA",X"D0",X"DD",X"A9",
		X"0B",X"95",X"34",X"A9",X"00",X"95",X"35",X"95",X"36",X"A9",X"F0",X"85",X"5D",X"A6",X"0B",X"A4",
		X"0C",X"B5",X"53",X"99",X"1E",X"00",X"B5",X"52",X"99",X"1D",X"00",X"A0",X"00",X"F0",X"8D",X"6E",
		X"98",X"10",X"09",X"20",X"08",X"77",X"20",X"FC",X"76",X"4C",X"08",X"77",X"A8",X"8A",X"10",X"0E",
		X"20",X"08",X"77",X"20",X"0E",X"77",X"49",X"80",X"49",X"FF",X"18",X"69",X"01",X"60",X"85",X"0C",
		X"98",X"C5",X"0C",X"F0",X"10",X"90",X"11",X"A4",X"0C",X"85",X"0C",X"98",X"20",X"28",X"77",X"38",
		X"E9",X"40",X"4C",X"08",X"77",X"A9",X"20",X"60",X"20",X"6C",X"77",X"BD",X"2F",X"77",X"60",X"00",
		X"02",X"05",X"07",X"0A",X"0C",X"0F",X"11",X"13",X"15",X"17",X"19",X"1A",X"1C",X"1D",X"1F",X"08",
		X"86",X"17",X"88",X"84",X"16",X"18",X"65",X"16",X"85",X"15",X"28",X"AA",X"08",X"B5",X"00",X"4A",
		X"4A",X"4A",X"4A",X"28",X"20",X"85",X"77",X"A5",X"16",X"D0",X"01",X"18",X"A6",X"15",X"B5",X"00",
		X"20",X"85",X"77",X"C6",X"15",X"A6",X"15",X"C6",X"16",X"10",X"E1",X"60",X"A0",X"00",X"84",X"0B",
		X"A0",X"04",X"26",X"0B",X"2A",X"C5",X"0C",X"90",X"02",X"E5",X"0C",X"88",X"D0",X"F4",X"A5",X"0B",
		X"2A",X"29",X"0F",X"AA",X"60",X"90",X"04",X"29",X"0F",X"F0",X"27",X"A6",X"17",X"F0",X"23",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A8",X"B9",X"D4",X"56",X"0A",X"85",X"0B",X"B9",X"D5",X"56",
		X"2A",X"29",X"1F",X"09",X"40",X"85",X"0C",X"A9",X"00",X"85",X"08",X"85",X"09",X"20",X"D7",X"6A",
		X"28",X"60",X"4C",X"CB",X"7B",X"06",X"5F",X"26",X"60",X"10",X"02",X"E6",X"5F",X"A5",X"5F",X"2C",
		X"D1",X"77",X"F0",X"04",X"49",X"01",X"85",X"5F",X"05",X"60",X"D0",X"02",X"E6",X"5F",X"A5",X"5F",
		X"60",X"02",X"18",X"69",X"40",X"10",X"08",X"29",X"7F",X"20",X"DF",X"77",X"4C",X"08",X"77",X"C9",
		X"41",X"90",X"04",X"49",X"7F",X"69",X"00",X"AA",X"BD",X"B9",X"57",X"60",X"06",X"0B",X"2A",X"06",
		X"0B",X"2A",X"38",X"E5",X"0C",X"60",X"AD",X"03",X"28",X"29",X"03",X"0A",X"AA",X"A9",X"10",X"85");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
