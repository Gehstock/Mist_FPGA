library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity chargen is
    generic(
        AddrWidth   : integer := 11
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end chargen;

architecture rtl of chargen is
    signal romAddr : integer range 0 to 2**AddrWidth-1;
    type rom2048x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom2048x8 := (
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0000
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0008
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0010
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0018
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0020
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0028
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0030
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0038
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0040
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0048
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0050
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0058
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0060
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0068
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0070
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0078
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0080
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0088
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0090
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0098
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0100
         x"10",  x"10",  x"10",  x"10",  x"00",  x"00",  x"10",  x"00", -- 0108
         x"28",  x"28",  x"28",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0110
         x"28",  x"28",  x"7c",  x"28",  x"7c",  x"28",  x"28",  x"00", -- 0118
         x"10",  x"3c",  x"50",  x"38",  x"14",  x"78",  x"10",  x"00", -- 0120
         x"60",  x"64",  x"08",  x"10",  x"20",  x"4c",  x"0c",  x"00", -- 0128
         x"10",  x"28",  x"28",  x"30",  x"54",  x"48",  x"34",  x"00", -- 0130
         x"04",  x"10",  x"20",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"08",  x"10",  x"20",  x"20",  x"20",  x"10",  x"08",  x"00", -- 0140
         x"20",  x"10",  x"08",  x"08",  x"08",  x"10",  x"20",  x"00", -- 0148
         x"00",  x"10",  x"54",  x"38",  x"54",  x"10",  x"00",  x"00", -- 0150
         x"00",  x"10",  x"10",  x"7c",  x"10",  x"10",  x"00",  x"00", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"10",  x"10",  x"20",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"7c",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"30",  x"30",  x"00", -- 0170
         x"00",  x"04",  x"08",  x"10",  x"20",  x"40",  x"00",  x"00", -- 0178
         x"38",  x"44",  x"4c",  x"54",  x"64",  x"44",  x"38",  x"00", -- 0180
         x"10",  x"30",  x"10",  x"10",  x"10",  x"10",  x"38",  x"00", -- 0188
         x"38",  x"44",  x"04",  x"08",  x"10",  x"20",  x"7c",  x"00", -- 0190
         x"7c",  x"08",  x"10",  x"08",  x"04",  x"44",  x"38",  x"00", -- 0198
         x"08",  x"18",  x"28",  x"48",  x"7c",  x"08",  x"08",  x"00", -- 01A0
         x"7c",  x"40",  x"78",  x"04",  x"04",  x"44",  x"38",  x"00", -- 01A8
         x"18",  x"20",  x"40",  x"78",  x"44",  x"44",  x"38",  x"00", -- 01B0
         x"7c",  x"04",  x"08",  x"10",  x"20",  x"20",  x"20",  x"00", -- 01B8
         x"38",  x"44",  x"44",  x"38",  x"44",  x"44",  x"38",  x"00", -- 01C0
         x"38",  x"44",  x"44",  x"3c",  x"04",  x"08",  x"30",  x"00", -- 01C8
         x"00",  x"30",  x"30",  x"00",  x"30",  x"30",  x"00",  x"00", -- 01D0
         x"00",  x"00",  x"10",  x"00",  x"10",  x"10",  x"20",  x"00", -- 01D8
         x"08",  x"10",  x"20",  x"40",  x"20",  x"10",  x"08",  x"00", -- 01E0
         x"00",  x"00",  x"7c",  x"00",  x"7c",  x"00",  x"00",  x"00", -- 01E8
         x"20",  x"10",  x"08",  x"04",  x"08",  x"10",  x"20",  x"00", -- 01F0
         x"38",  x"44",  x"04",  x"08",  x"10",  x"10",  x"10",  x"00", -- 01F8
         x"38",  x"44",  x"5c",  x"54",  x"5c",  x"40",  x"3c",  x"00", -- 0200
         x"38",  x"44",  x"44",  x"7c",  x"44",  x"44",  x"44",  x"00", -- 0208
         x"78",  x"44",  x"44",  x"78",  x"44",  x"44",  x"78",  x"00", -- 0210
         x"38",  x"44",  x"40",  x"40",  x"40",  x"44",  x"38",  x"00", -- 0218
         x"78",  x"24",  x"24",  x"24",  x"24",  x"24",  x"78",  x"00", -- 0220
         x"7c",  x"40",  x"40",  x"78",  x"40",  x"40",  x"7c",  x"00", -- 0228
         x"7c",  x"40",  x"40",  x"78",  x"40",  x"40",  x"40",  x"00", -- 0230
         x"38",  x"44",  x"40",  x"40",  x"4c",  x"44",  x"3c",  x"00", -- 0238
         x"44",  x"44",  x"44",  x"7c",  x"44",  x"44",  x"44",  x"00", -- 0240
         x"38",  x"10",  x"10",  x"10",  x"10",  x"10",  x"38",  x"00", -- 0248
         x"1c",  x"08",  x"08",  x"08",  x"08",  x"48",  x"30",  x"00", -- 0250
         x"44",  x"48",  x"50",  x"60",  x"50",  x"48",  x"44",  x"00", -- 0258
         x"40",  x"40",  x"40",  x"40",  x"40",  x"40",  x"7c",  x"00", -- 0260
         x"44",  x"6c",  x"54",  x"54",  x"44",  x"44",  x"44",  x"00", -- 0268
         x"44",  x"44",  x"64",  x"54",  x"4c",  x"44",  x"44",  x"00", -- 0270
         x"38",  x"44",  x"44",  x"44",  x"44",  x"44",  x"38",  x"00", -- 0278
         x"78",  x"44",  x"44",  x"78",  x"40",  x"40",  x"40",  x"00", -- 0280
         x"38",  x"44",  x"44",  x"44",  x"54",  x"48",  x"34",  x"00", -- 0288
         x"78",  x"44",  x"44",  x"78",  x"50",  x"48",  x"44",  x"00", -- 0290
         x"3c",  x"40",  x"40",  x"38",  x"04",  x"04",  x"78",  x"00", -- 0298
         x"7c",  x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"00", -- 02A0
         x"44",  x"44",  x"44",  x"44",  x"44",  x"44",  x"38",  x"00", -- 02A8
         x"44",  x"44",  x"44",  x"44",  x"44",  x"28",  x"10",  x"00", -- 02B0
         x"44",  x"44",  x"44",  x"54",  x"54",  x"6c",  x"44",  x"00", -- 02B8
         x"44",  x"44",  x"28",  x"10",  x"28",  x"44",  x"44",  x"00", -- 02C0
         x"44",  x"44",  x"44",  x"28",  x"10",  x"10",  x"10",  x"00", -- 02C8
         x"7c",  x"04",  x"08",  x"10",  x"20",  x"40",  x"7c",  x"00", -- 02D0
         x"38",  x"20",  x"20",  x"20",  x"20",  x"20",  x"38",  x"00", -- 02D8
         x"00",  x"40",  x"20",  x"10",  x"08",  x"04",  x"00",  x"00", -- 02E0
         x"38",  x"08",  x"08",  x"08",  x"08",  x"08",  x"38",  x"00", -- 02E8
         x"10",  x"10",  x"10",  x"28",  x"28",  x"44",  x"44",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"7c",  x"00",  x"00", -- 02F8
         x"00",  x"20",  x"10",  x"08",  x"00",  x"00",  x"00",  x"00", -- 0300
         x"00",  x"00",  x"34",  x"4c",  x"44",  x"44",  x"3a",  x"00", -- 0308
         x"40",  x"40",  x"58",  x"64",  x"44",  x"44",  x"78",  x"00", -- 0310
         x"00",  x"00",  x"38",  x"44",  x"40",  x"44",  x"38",  x"00", -- 0318
         x"04",  x"04",  x"34",  x"4c",  x"44",  x"44",  x"3a",  x"00", -- 0320
         x"00",  x"00",  x"38",  x"4c",  x"7c",  x"40",  x"38",  x"00", -- 0328
         x"08",  x"10",  x"38",  x"10",  x"10",  x"10",  x"10",  x"00", -- 0330
         x"00",  x"00",  x"34",  x"4c",  x"44",  x"3c",  x"04",  x"38", -- 0338
         x"40",  x"40",  x"58",  x"64",  x"44",  x"44",  x"44",  x"00", -- 0340
         x"10",  x"00",  x"10",  x"10",  x"10",  x"10",  x"08",  x"00", -- 0348
         x"10",  x"00",  x"10",  x"10",  x"10",  x"10",  x"10",  x"20", -- 0350
         x"40",  x"40",  x"48",  x"50",  x"70",  x"48",  x"44",  x"00", -- 0358
         x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"08",  x"00", -- 0360
         x"00",  x"00",  x"68",  x"54",  x"54",  x"54",  x"54",  x"00", -- 0368
         x"00",  x"00",  x"58",  x"64",  x"44",  x"44",  x"44",  x"00", -- 0370
         x"00",  x"00",  x"38",  x"44",  x"44",  x"44",  x"38",  x"00", -- 0378
         x"00",  x"00",  x"58",  x"64",  x"44",  x"78",  x"40",  x"40", -- 0380
         x"00",  x"00",  x"34",  x"4c",  x"44",  x"3c",  x"04",  x"04", -- 0388
         x"00",  x"00",  x"58",  x"64",  x"40",  x"40",  x"40",  x"00", -- 0390
         x"00",  x"00",  x"38",  x"40",  x"38",  x"04",  x"78",  x"00", -- 0398
         x"10",  x"10",  x"38",  x"10",  x"10",  x"10",  x"08",  x"00", -- 03A0
         x"00",  x"00",  x"44",  x"44",  x"44",  x"4c",  x"34",  x"00", -- 03A8
         x"00",  x"00",  x"44",  x"44",  x"44",  x"28",  x"10",  x"00", -- 03B0
         x"00",  x"00",  x"54",  x"54",  x"54",  x"54",  x"28",  x"00", -- 03B8
         x"00",  x"00",  x"44",  x"28",  x"10",  x"28",  x"44",  x"00", -- 03C0
         x"00",  x"00",  x"44",  x"44",  x"44",  x"3c",  x"04",  x"38", -- 03C8
         x"00",  x"00",  x"7c",  x"08",  x"10",  x"20",  x"7c",  x"00", -- 03D0
         x"08",  x"10",  x"10",  x"20",  x"10",  x"10",  x"08",  x"00", -- 03D8
         x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"00", -- 03E0
         x"20",  x"10",  x"10",  x"08",  x"10",  x"10",  x"20",  x"00", -- 03E8
         x"00",  x"00",  x"00",  x"32",  x"4c",  x"00",  x"00",  x"00", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F8
         x"c0",  x"20",  x"10",  x"10",  x"10",  x"10",  x"20",  x"c0", -- 0400
         x"03",  x"04",  x"08",  x"08",  x"08",  x"08",  x"04",  x"03", -- 0408
         x"81",  x"81",  x"42",  x"3c",  x"00",  x"00",  x"00",  x"00", -- 0410
         x"00",  x"00",  x"00",  x"00",  x"3c",  x"42",  x"81",  x"81", -- 0418
         x"10",  x"10",  x"20",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 0420
         x"08",  x"08",  x"04",  x"03",  x"00",  x"00",  x"00",  x"00", -- 0428
         x"00",  x"00",  x"00",  x"00",  x"03",  x"04",  x"08",  x"08", -- 0430
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"20",  x"10",  x"10", -- 0438
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"ff", -- 0440
         x"ff",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01", -- 0448
         x"00",  x"10",  x"28",  x"44",  x"82",  x"44",  x"28",  x"10", -- 0450
         x"ff",  x"ef",  x"c7",  x"83",  x"01",  x"83",  x"c7",  x"ef", -- 0458
         x"3c",  x"42",  x"81",  x"81",  x"81",  x"81",  x"42",  x"3c", -- 0460
         x"c3",  x"81",  x"00",  x"00",  x"00",  x"00",  x"81",  x"c3", -- 0468
         x"ff",  x"fe",  x"fc",  x"f8",  x"f0",  x"e0",  x"c0",  x"80", -- 0470
         x"80",  x"c0",  x"e0",  x"f0",  x"f8",  x"fc",  x"fe",  x"ff", -- 0478
         x"01",  x"02",  x"04",  x"08",  x"10",  x"20",  x"40",  x"80", -- 0480
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"01", -- 0488
         x"00",  x"00",  x"00",  x"00",  x"03",  x"0c",  x"30",  x"c0", -- 0490
         x"03",  x"0c",  x"30",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 0498
         x"03",  x"0c",  x"30",  x"c0",  x"c0",  x"30",  x"0c",  x"03", -- 04A0
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"30",  x"0c",  x"03", -- 04A8
         x"c0",  x"30",  x"0c",  x"03",  x"00",  x"00",  x"00",  x"00", -- 04B0
         x"c0",  x"30",  x"0c",  x"03",  x"03",  x"0c",  x"30",  x"c0", -- 04B8
         x"10",  x"10",  x"20",  x"20",  x"40",  x"40",  x"80",  x"80", -- 04C0
         x"01",  x"01",  x"02",  x"02",  x"04",  x"04",  x"08",  x"08", -- 04C8
         x"81",  x"81",  x"42",  x"42",  x"24",  x"24",  x"18",  x"18", -- 04D0
         x"80",  x"80",  x"40",  x"40",  x"20",  x"20",  x"10",  x"10", -- 04D8
         x"08",  x"08",  x"04",  x"04",  x"02",  x"02",  x"01",  x"01", -- 04E0
         x"18",  x"18",  x"24",  x"24",  x"42",  x"42",  x"81",  x"81", -- 04E8
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 04F0
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80", -- 04F8
         x"00",  x"00",  x"00",  x"ff",  x"ff",  x"00",  x"00",  x"00", -- 0500
         x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18", -- 0508
         x"18",  x"18",  x"18",  x"ff",  x"ff",  x"00",  x"00",  x"00", -- 0510
         x"18",  x"18",  x"18",  x"1f",  x"1f",  x"18",  x"18",  x"18", -- 0518
         x"00",  x"00",  x"00",  x"ff",  x"ff",  x"18",  x"18",  x"18", -- 0520
         x"18",  x"18",  x"18",  x"f8",  x"f8",  x"18",  x"18",  x"18", -- 0528
         x"18",  x"18",  x"18",  x"ff",  x"ff",  x"18",  x"18",  x"18", -- 0530
         x"18",  x"18",  x"18",  x"1f",  x"1f",  x"00",  x"00",  x"00", -- 0538
         x"00",  x"00",  x"00",  x"1f",  x"1f",  x"18",  x"18",  x"18", -- 0540
         x"00",  x"00",  x"00",  x"f8",  x"f8",  x"18",  x"18",  x"18", -- 0548
         x"18",  x"18",  x"18",  x"f8",  x"f8",  x"00",  x"00",  x"00", -- 0550
         x"80",  x"80",  x"80",  x"40",  x"40",  x"20",  x"18",  x"07", -- 0558
         x"01",  x"01",  x"01",  x"02",  x"02",  x"04",  x"18",  x"e0", -- 0560
         x"e0",  x"18",  x"04",  x"02",  x"02",  x"01",  x"01",  x"01", -- 0568
         x"07",  x"18",  x"20",  x"40",  x"40",  x"80",  x"80",  x"80", -- 0570
         x"81",  x"42",  x"24",  x"18",  x"18",  x"24",  x"42",  x"81", -- 0578
         x"f0",  x"f0",  x"f0",  x"f0",  x"00",  x"00",  x"00",  x"00", -- 0580
         x"0f",  x"0f",  x"0f",  x"0f",  x"00",  x"00",  x"00",  x"00", -- 0588
         x"00",  x"00",  x"00",  x"00",  x"0f",  x"0f",  x"0f",  x"0f", -- 0590
         x"00",  x"00",  x"00",  x"00",  x"f0",  x"f0",  x"f0",  x"f0", -- 0598
         x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0", -- 05A0
         x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f", -- 05A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 05B0
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff", -- 05B8
         x"f0",  x"f0",  x"f0",  x"f0",  x"0f",  x"0f",  x"0f",  x"0f", -- 05C0
         x"0f",  x"0f",  x"0f",  x"0f",  x"f0",  x"f0",  x"f0",  x"f0", -- 05C8
         x"0f",  x"0f",  x"0f",  x"0f",  x"ff",  x"ff",  x"ff",  x"ff", -- 05D0
         x"f0",  x"f0",  x"f0",  x"f0",  x"ff",  x"ff",  x"ff",  x"ff", -- 05D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"f0",  x"f0",  x"f0",  x"f0", -- 05E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"0f",  x"0f",  x"0f",  x"0f", -- 05E8
         x"01",  x"03",  x"07",  x"0f",  x"1f",  x"3f",  x"7f",  x"ff", -- 05F0
         x"ff",  x"7f",  x"3f",  x"1f",  x"0f",  x"07",  x"03",  x"01", -- 05F8
         x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01", -- 0600
         x"ff",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80", -- 0608
         x"ff",  x"80",  x"80",  x"9c",  x"9c",  x"9c",  x"80",  x"80", -- 0610
         x"ff",  x"ff",  x"ff",  x"e3",  x"e3",  x"e3",  x"ff",  x"ff", -- 0618
         x"18",  x"3c",  x"7e",  x"3c",  x"18",  x"3c",  x"7e",  x"ff", -- 0620
         x"ff",  x"00",  x"ff",  x"00",  x"ff",  x"00",  x"ff",  x"00", -- 0628
         x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa", -- 0630
         x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa", -- 0638
         x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"ff", -- 0640
         x"00",  x"10",  x"38",  x"7c",  x"fe",  x"7c",  x"38",  x"10", -- 0648
         x"38",  x"10",  x"92",  x"fe",  x"92",  x"10",  x"38",  x"7c", -- 0650
         x"00",  x"6c",  x"fe",  x"fe",  x"fe",  x"7c",  x"38",  x"10", -- 0658
         x"10",  x"38",  x"7c",  x"fe",  x"fe",  x"7c",  x"10",  x"7c", -- 0660
         x"e7",  x"e7",  x"42",  x"ff",  x"ff",  x"42",  x"e7",  x"e7", -- 0668
         x"db",  x"ff",  x"db",  x"18",  x"18",  x"db",  x"ff",  x"db", -- 0670
         x"3c",  x"7e",  x"ff",  x"ff",  x"ff",  x"ff",  x"7e",  x"3c", -- 0678
         x"c0",  x"c0",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0680
         x"30",  x"30",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0688
         x"0c",  x"0c",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0690
         x"03",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0698
         x"00",  x"00",  x"c0",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 06A0
         x"00",  x"00",  x"30",  x"30",  x"00",  x"00",  x"00",  x"00", -- 06A8
         x"00",  x"00",  x"0c",  x"0c",  x"00",  x"00",  x"00",  x"00", -- 06B0
         x"00",  x"00",  x"03",  x"03",  x"00",  x"00",  x"00",  x"00", -- 06B8
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"c0",  x"00",  x"00", -- 06C0
         x"00",  x"00",  x"00",  x"00",  x"30",  x"30",  x"00",  x"00", -- 06C8
         x"00",  x"00",  x"00",  x"00",  x"0c",  x"0c",  x"00",  x"00", -- 06D0
         x"00",  x"00",  x"00",  x"00",  x"03",  x"03",  x"00",  x"00", -- 06D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"c0", -- 06E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"30",  x"30", -- 06E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"0c",  x"0c", -- 06F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"03", -- 06F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"0f",  x"0f", -- 0700
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"3f",  x"3f", -- 0708
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 0710
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"fc",  x"fc", -- 0718
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"f0",  x"f0", -- 0720
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"c0", -- 0728
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"c0",  x"c0",  x"c0", -- 0730
         x"00",  x"00",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0", -- 0738
         x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0", -- 0740
         x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"00",  x"00", -- 0748
         x"c0",  x"c0",  x"c0",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 0750
         x"c0",  x"c0",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0758
         x"f0",  x"f0",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0760
         x"fc",  x"fc",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0768
         x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0770
         x"3f",  x"3f",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0778
         x"0f",  x"0f",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0780
         x"03",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0788
         x"03",  x"03",  x"03",  x"03",  x"00",  x"00",  x"00",  x"00", -- 0790
         x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"00",  x"00", -- 0798
         x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03", -- 07A0
         x"00",  x"00",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03", -- 07A8
         x"00",  x"00",  x"00",  x"00",  x"03",  x"03",  x"03",  x"03", -- 07B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"03", -- 07B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 07C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 07C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff", -- 07D0
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff", -- 07D8
         x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07E0
         x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07E8
         x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 07F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
