library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx4 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"CC",X"0B",X"CC",X"BB",X"CF",X"BB",X"CC",X"CB",X"BB",
		X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"CC",X"4C",X"CC",X"44",X"CF",X"44",X"BC",X"44",X"BB",X"44",
		X"0C",X"BB",X"00",X"CC",X"0B",X"BF",X"0B",X"BF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"BB",X"BF",
		X"BB",X"CC",X"CC",X"00",X"FF",X"44",X"FF",X"44",X"FF",X"C0",X"FF",X"4C",X"FF",X"4C",X"FF",X"44",
		X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"CB",X"00",X"CB",X"00",X"BC",X"00",X"CC",X"0B",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"C4",X"BB",X"C4",X"BC",X"44",X"BC",X"C4",X"BC",X"C4",
		X"0B",X"CC",X"0C",X"BB",X"00",X"BB",X"00",X"CC",X"0B",X"BB",X"00",X"BB",X"00",X"BF",X"00",X"FF",
		X"BB",X"C4",X"BB",X"44",X"CB",X"4C",X"BC",X"C4",X"BB",X"44",X"FF",X"4C",X"FF",X"44",X"FF",X"F4",
		X"00",X"BC",X"00",X"CB",X"00",X"CB",X"00",X"BC",X"00",X"CC",X"0B",X"CC",X"0B",X"CC",X"0C",X"BB",
		X"00",X"BC",X"00",X"C4",X"BB",X"C4",X"BC",X"44",X"BC",X"C4",X"BC",X"C4",X"BB",X"C4",X"BB",X"44",
		X"00",X"BB",X"00",X"CC",X"00",X"BB",X"00",X"CB",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"00",X"BB",
		X"CB",X"4C",X"FC",X"C0",X"FF",X"44",X"FF",X"C4",X"FF",X"4C",X"FF",X"F4",X"FF",X"44",X"FF",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"BB",X"0B",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"BB",X"4C",X"CC",X"44",
		X"BB",X"CC",X"BB",X"CF",X"CB",X"CC",X"0C",X"BB",X"00",X"CC",X"0B",X"BF",X"0B",X"CF",X"0C",X"CF",
		X"CC",X"44",X"CF",X"44",X"BC",X"44",X"BB",X"CC",X"CC",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"CC",X"0B",X"CC",X"BB",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"CC",X"4C",X"CC",X"44",X"CF",X"44",
		X"BC",X"CC",X"CB",X"BB",X"0B",X"BB",X"0B",X"CC",X"0B",X"BB",X"0C",X"BF",X"00",X"FF",X"00",X"FF",
		X"BC",X"44",X"BB",X"44",X"BB",X"CC",X"CC",X"44",X"BB",X"44",X"FF",X"CC",X"FF",X"4C",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"BC",X"0B",X"CC",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"BC",X"4C",X"BC",X"C4",X"BC",X"C4",
		X"BB",X"CC",X"CB",X"BB",X"0C",X"BC",X"0B",X"CC",X"0B",X"BB",X"0C",X"BF",X"00",X"FF",X"00",X"FF",
		X"BB",X"C4",X"BB",X"44",X"CB",X"CC",X"BC",X"44",X"BB",X"44",X"FF",X"CC",X"FF",X"4C",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"00",X"4B",X"00",X"BB",X"0B",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"BB",X"4C",X"BB",X"4C",X"BC",X"44",
		X"BB",X"CC",X"BB",X"CC",X"CB",X"CC",X"0C",X"BB",X"00",X"CC",X"0B",X"CF",X"0C",X"BC",X"00",X"BB",
		X"BC",X"C4",X"BC",X"C4",X"BB",X"C4",X"CB",X"CC",X"FC",X"44",X"FF",X"44",X"FF",X"CC",X"FF",X"4C",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"CF",X"00",X"CC",X"0B",X"BB",X"BB",X"BC",X"BB",X"BB",X"CB",X"BF",
		X"00",X"00",X"00",X"00",X"CF",X"00",X"BC",X"4C",X"BB",X"44",X"CC",X"44",X"CB",X"44",X"FF",X"44",
		X"0B",X"FF",X"0C",X"FF",X"0B",X"FF",X"44",X"FF",X"44",X"FF",X"C4",X"FF",X"04",X"4F",X"0C",X"44",
		X"FF",X"44",X"FF",X"4C",X"FF",X"F4",X"FF",X"F4",X"FF",X"F4",X"FF",X"44",X"FF",X"44",X"44",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CB",X"0B",X"BB",X"0B",X"BF",X"0B",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"4C",X"CB",X"44",X"FF",X"44",X"FF",X"44",
		X"0C",X"FF",X"0B",X"FF",X"44",X"FF",X"44",X"FF",X"C4",X"FF",X"04",X"4F",X"0C",X"44",X"00",X"CC",
		X"FF",X"4C",X"FF",X"F4",X"FF",X"F4",X"FF",X"F4",X"FF",X"44",X"FF",X"44",X"44",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CB",X"0B",X"BF",X"0B",X"FF",X"0B",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"4C",X"FB",X"44",X"FF",X"44",X"FF",X"44",
		X"0C",X"FF",X"BB",X"FF",X"44",X"FF",X"CC",X"FF",X"44",X"FF",X"44",X"4F",X"C4",X"44",X"0C",X"CC",
		X"FF",X"FC",X"FF",X"F4",X"FF",X"F4",X"FF",X"FC",X"FF",X"C4",X"FF",X"44",X"44",X"44",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"00",X"BB",X"0B",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"BB",X"4C",X"BB",X"4C",X"CC",X"44",
		X"BB",X"CC",X"BB",X"CF",X"CB",X"CC",X"0C",X"CB",X"0B",X"CC",X"0B",X"BF",X"0C",X"FF",X"0C",X"FF",
		X"CC",X"44",X"CF",X"44",X"BC",X"44",X"BC",X"4C",X"CC",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"BB",X"00",X"00",X"0B",X"00",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"00",X"B0",X"00",X"B0",X"00",X"BB",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"B0",X"00",X"BB",X"B0",X"00",X"B0",X"0B",X"BB",X"BB",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"8F",X"00",X"8F",X"00",X"8F",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"09",X"99",X"99",X"88",X"88",X"88",X"C8",X"8C",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"EE",
		X"E8",X"88",X"EE",X"88",X"EE",X"88",X"EE",X"89",X"E8",X"C9",X"CC",X"98",X"99",X"88",X"99",X"88",
		X"FF",X"EC",X"EE",X"C9",X"0C",X"09",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"88",X"98",X"88",X"88",X"8C",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"00",X"55",X"00",X"55",X"00",X"59",X"00",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"99",X"55",X"99",X"55",X"99",X"55",X"99",X"55",
		X"09",X"09",X"09",X"00",X"90",X"00",X"90",X"00",X"90",X"90",X"00",X"99",X"00",X"08",X"00",X"00",
		X"99",X"00",X"00",X"09",X"98",X"09",X"98",X"08",X"98",X"90",X"98",X"80",X"98",X"00",X"99",X"00",
		X"00",X"FE",X"00",X"CE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0F",X"FF",
		X"0F",X"00",X"0F",X"00",X"0F",X"E0",X"0F",X"E0",X"0F",X"E0",X"FF",X"E0",X"FF",X"E0",X"FF",X"FE",
		X"0F",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"E0",X"FE",X"00",X"00",X"00",X"FF",X"0F",X"FF",X"0F",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"B4",X"00",X"4F",X"00",X"FF",X"00",X"FF",X"00",X"11",
		X"00",X"00",X"44",X"00",X"44",X"C0",X"44",X"4C",X"4F",X"44",X"FF",X"44",X"FC",X"44",X"11",X"4C",
		X"00",X"41",X"0B",X"41",X"0B",X"CF",X"BB",X"C4",X"BC",X"4C",X"BC",X"41",X"11",X"11",X"1C",X"11",
		X"41",X"C4",X"11",X"C4",X"FD",X"44",X"44",X"4C",X"CC",X"C0",X"11",X"C0",X"11",X"4C",X"11",X"4C",
		X"00",X"0B",X"00",X"BB",X"00",X"B4",X"00",X"41",X"00",X"11",X"00",X"10",X"04",X"11",X"04",X"CF",
		X"44",X"00",X"44",X"00",X"44",X"40",X"41",X"40",X"11",X"40",X"11",X"44",X"11",X"14",X"11",X"F1",
		X"04",X"CF",X"00",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F1",X"FC",X"14",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"0B",X"00",X"0B",X"00",X"B0",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"04",X"BB",X"04",X"B0",X"44",X"B0",X"04",X"B0",X"04",
		X"0B",X"00",X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BF",X"00",X"FF",
		X"BB",X"04",X"BB",X"44",X"0B",X"40",X"B0",X"04",X"BB",X"44",X"FF",X"40",X"FF",X"44",X"FF",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"0B",X"00",X"0B",X"00",X"B0",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"04",X"BB",X"04",X"B0",X"44",X"B0",X"04",X"B0",X"04",
		X"0B",X"00",X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"0F",X"00",X"0F",
		X"BB",X"04",X"BB",X"44",X"0B",X"40",X"B0",X"00",X"BB",X"40",X"FF",X"44",X"FF",X"04",X"FF",X"F0",
		X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"AA",
		X"00",X"00",X"33",X"00",X"33",X"00",X"FF",X"00",X"CF",X"00",X"CF",X"00",X"AF",X"33",X"AA",X"33",
		X"00",X"3A",X"03",X"3F",X"03",X"3F",X"33",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"AA",X"00",X"AA",
		X"AA",X"33",X"FF",X"30",X"FF",X"30",X"FF",X"F0",X"FF",X"FA",X"FF",X"AA",X"FA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"88",X"08",X"89",X"90",X"DD",X"00",X"E5",X"08",X"5C",X"90",X"EE",
		X"00",X"00",X"80",X"09",X"98",X"80",X"88",X"88",X"8D",X"80",X"DE",X"D8",X"D5",X"D8",X"DE",X"D8",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DE",X"D0",X"FF",X"D0",X"CC",X"00",X"FF",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"28",X"22",X"88",X"22",X"88",X"22",X"68",X"22",X"58",X"22",X"88",X"22",X"88",X"22",X"88",
		X"88",X"22",X"88",X"C2",X"88",X"C2",X"88",X"C2",X"88",X"C2",X"88",X"C2",X"88",X"22",X"88",X"22",
		X"22",X"C8",X"22",X"8C",X"22",X"88",X"22",X"8A",X"28",X"8A",X"28",X"AA",X"2C",X"AA",X"28",X"AA",
		X"88",X"22",X"CC",X"22",X"A8",X"C2",X"AA",X"C2",X"AA",X"88",X"AA",X"88",X"AA",X"CC",X"AA",X"88",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FF",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"33",X"20",X"3F",X"20",X"3F",X"32",X"3F",X"32",
		X"00",X"FF",X"00",X"3F",X"03",X"FF",X"33",X"FF",X"30",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"BB",X"32",X"BF",X"32",X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"20",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"6F",X"00",X"FF",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"50",X"6F",X"50",X"6F",X"55",X"6F",X"55",
		X"00",X"FF",X"00",X"6F",X"06",X"FF",X"66",X"FF",X"60",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"AA",X"65",X"AC",X"65",X"CF",X"65",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"50",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"6F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"50",X"6F",X"50",X"6F",X"55",X"6C",X"55",
		X"00",X"FF",X"00",X"6F",X"06",X"FF",X"66",X"FF",X"60",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"AA",X"65",X"AC",X"65",X"CF",X"65",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"50",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"C0",X"00",X"C0",X"00",X"C5",X"00",X"C6",X"00",X"C6",X"50",X"66",X"50",X"6F",X"F5",X"6C",X"65",
		X"00",X"66",X"00",X"FF",X"06",X"FF",X"66",X"FF",X"66",X"FF",X"66",X"FF",X"60",X"FF",X"00",X"FF",
		X"AA",X"65",X"AC",X"65",X"CF",X"F5",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"00",X"00",X"00",X"AA",X"00",X"AA",X"00",X"5A",X"00",X"5A",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"00",X"00",X"AA",X"00",X"AA",X"60",X"AA",X"55",X"AA",X"55",X"AA",X"5A",X"AA",X"A0",X"AA",X"00",
		X"0A",X"BA",X"A0",X"BB",X"00",X"C4",X"0A",X"BC",X"A0",X"BB",X"00",X"C4",X"0A",X"BC",X"A0",X"BB",
		X"CC",X"AA",X"BA",X"A0",X"44",X"00",X"CC",X"AA",X"BB",X"A0",X"44",X"00",X"CC",X"AA",X"BB",X"A0",
		X"00",X"6F",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"8F",X"00",X"00",X"00",X"70",X"0E",X"5A",
		X"00",X"F0",X"F0",X"00",X"FF",X"0F",X"40",X"A0",X"00",X"00",X"5F",X"30",X"A0",X"0F",X"73",X"2A",
		X"F0",X"0F",X"78",X"A0",X"70",X"78",X"00",X"AF",X"53",X"80",X"00",X"70",X"00",X"2F",X"08",X"40",
		X"A0",X"00",X"83",X"87",X"71",X"05",X"58",X"05",X"14",X"A0",X"F0",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"FF",X"00",X"FF",X"60",X"FF",
		X"C0",X"00",X"C0",X"00",X"C5",X"00",X"C6",X"00",X"C6",X"50",X"66",X"50",X"6F",X"F5",X"6C",X"65",
		X"60",X"66",X"66",X"FA",X"66",X"FC",X"06",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"AA",X"65",X"CC",X"65",X"CA",X"F5",X"AC",X"F5",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C3",X"C0",X"2C",X"22",
		X"33",X"33",X"33",X"33",X"23",X"33",X"C2",X"33",X"0C",X"23",X"00",X"C2",X"00",X"0C",X"00",X"00",
		X"22",X"33",X"22",X"33",X"33",X"33",X"33",X"33",X"33",X"22",X"22",X"CC",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"2C",X"F3",X"F2",X"03",X"F2",X"F3",X"F2",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"20",X"2C",X"32",
		X"33",X"33",X"33",X"33",X"23",X"33",X"C2",X"33",X"0C",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"22",X"33",X"22",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"22",X"2C",X"CC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"FF",X"00",X"CF",X"00",X"FF",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"00",X"22",X"00",X"22",X"2C",X"22",X"32",
		X"33",X"33",X"33",X"33",X"23",X"33",X"C2",X"33",X"0C",X"33",X"00",X"22",X"00",X"CC",X"00",X"00",
		X"22",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"22",X"22",X"CC",X"CC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",X"BA",X"0A",X"CA",
		X"00",X"00",X"C0",X"00",X"BC",X"00",X"BA",X"C0",X"BC",X"C0",X"CA",X"BC",X"CA",X"BB",X"CA",X"BB",
		X"0A",X"CA",X"0A",X"CA",X"0A",X"CA",X"0A",X"CA",X"0C",X"CA",X"00",X"CA",X"00",X"0C",X"00",X"00",
		X"BC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"BB",X"C0",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"BB",X"0B",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"BB",X"4C",X"CC",X"44",
		X"BB",X"CC",X"BB",X"CF",X"CB",X"CC",X"0C",X"BB",X"00",X"CC",X"0B",X"BF",X"0B",X"CF",X"0C",X"CF",
		X"CC",X"44",X"CF",X"44",X"BC",X"44",X"BB",X"CC",X"CC",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"CC",X"0B",X"CC",X"BB",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"CC",X"4C",X"CC",X"44",X"CF",X"44",
		X"BC",X"CC",X"CB",X"BB",X"0B",X"BB",X"0B",X"CC",X"0B",X"BB",X"0C",X"BF",X"00",X"FF",X"00",X"FF",
		X"BC",X"44",X"BB",X"44",X"BB",X"CC",X"CC",X"44",X"BB",X"44",X"FF",X"CC",X"FF",X"4C",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"BC",X"0B",X"CC",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"4C",X"BB",X"4C",X"BC",X"4C",X"BC",X"C4",X"BC",X"C4",
		X"BB",X"CC",X"CB",X"BB",X"0C",X"BC",X"0B",X"CC",X"0B",X"BB",X"0C",X"BF",X"00",X"FF",X"00",X"FF",
		X"BB",X"C4",X"BB",X"44",X"CB",X"CC",X"BC",X"44",X"BB",X"44",X"FF",X"CC",X"FF",X"4C",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"00",X"4B",X"00",X"BB",X"0B",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"BB",X"4C",X"BB",X"4C",X"BC",X"44",
		X"BB",X"CC",X"BB",X"CC",X"CB",X"CC",X"0C",X"BB",X"00",X"CC",X"0B",X"CF",X"0C",X"BC",X"00",X"BB",
		X"BC",X"C4",X"BC",X"C4",X"BB",X"C4",X"CB",X"CC",X"FC",X"44",X"FF",X"44",X"FF",X"CC",X"FF",X"4C",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"CF",X"00",X"CC",X"0B",X"BB",X"BB",X"BC",X"BB",X"BB",X"CB",X"BF",
		X"00",X"00",X"00",X"00",X"CF",X"00",X"BC",X"4C",X"BB",X"44",X"CC",X"44",X"CB",X"44",X"FF",X"44",
		X"0B",X"FF",X"0C",X"FF",X"0B",X"FF",X"44",X"FF",X"44",X"FF",X"C4",X"FF",X"04",X"4F",X"0C",X"44",
		X"FF",X"44",X"FF",X"4C",X"FF",X"F4",X"FF",X"F4",X"FF",X"F4",X"FF",X"44",X"FF",X"44",X"44",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"6F",X"00",X"FF",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"50",X"6F",X"50",X"6F",X"55",X"6F",X"55",
		X"00",X"FF",X"00",X"6F",X"06",X"FF",X"66",X"FF",X"60",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"AA",X"65",X"AC",X"65",X"CF",X"65",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"50",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"6F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"50",X"6F",X"50",X"6F",X"55",X"6C",X"55",
		X"00",X"FF",X"00",X"6F",X"06",X"FF",X"66",X"FF",X"60",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"AA",X"65",X"AC",X"65",X"CF",X"65",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"50",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"C0",X"00",X"C0",X"00",X"C5",X"00",X"C6",X"00",X"C6",X"50",X"66",X"50",X"6F",X"F5",X"6C",X"65",
		X"00",X"66",X"00",X"FF",X"06",X"FF",X"66",X"FF",X"66",X"FF",X"66",X"FF",X"60",X"FF",X"00",X"FF",
		X"AA",X"65",X"AC",X"65",X"CF",X"F5",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"00",X"00",X"00",X"AA",X"00",X"AA",X"00",X"5A",X"00",X"5A",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"00",X"00",X"AA",X"00",X"AA",X"60",X"AA",X"55",X"AA",X"55",X"AA",X"5A",X"AA",X"A0",X"AA",X"00",
		X"0A",X"BA",X"A0",X"BB",X"00",X"C4",X"0A",X"BC",X"A0",X"BB",X"00",X"C4",X"0A",X"BC",X"A0",X"BB",
		X"CC",X"AA",X"BA",X"A0",X"44",X"00",X"CC",X"AA",X"BB",X"A0",X"44",X"00",X"CC",X"AA",X"BB",X"A0",
		X"00",X"6F",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"8F",X"00",X"00",X"00",X"70",X"0E",X"5A",
		X"00",X"F0",X"F0",X"00",X"FF",X"0F",X"40",X"A0",X"00",X"00",X"5F",X"30",X"A0",X"0F",X"73",X"2A",
		X"F0",X"0F",X"78",X"A0",X"70",X"78",X"00",X"AF",X"53",X"80",X"00",X"70",X"00",X"2F",X"08",X"40",
		X"A0",X"00",X"83",X"87",X"71",X"05",X"58",X"05",X"14",X"A0",X"F0",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"66",X"00",X"FF",X"00",X"FF",X"60",X"FF",
		X"C0",X"00",X"C0",X"00",X"C5",X"00",X"C6",X"00",X"C6",X"50",X"66",X"50",X"6F",X"F5",X"6C",X"65",
		X"60",X"66",X"66",X"FA",X"66",X"FC",X"06",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"AA",X"65",X"CC",X"65",X"CA",X"F5",X"AC",X"F5",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"00",X"0B",X"00",X"BB",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FF",X"00",X"BB",
		X"44",X"00",X"B4",X"C0",X"BB",X"FC",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BB",X"F4",X"CB",X"44",
		X"00",X"BC",X"0B",X"CB",X"BB",X"4C",X"BB",X"44",X"CB",X"4C",X"0C",X"C0",X"00",X"00",X"00",X"00",
		X"CB",X"CC",X"CC",X"B4",X"BB",X"BB",X"BC",X"BB",X"00",X"B4",X"00",X"4C",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"FB",X"00",X"FB",X"00",X"BB",X"00",X"CB",
		X"00",X"00",X"00",X"00",X"B4",X"00",X"BB",X"C0",X"BB",X"4C",X"BB",X"4C",X"BB",X"44",X"BB",X"44",
		X"00",X"CB",X"00",X"BB",X"0B",X"BB",X"0B",X"CB",X"0C",X"4C",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"BB",X"44",X"CB",X"44",X"CB",X"CB",X"BB",X"BB",X"CC",X"44",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"FB",X"00",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"00",X"BB",X"C0",X"BB",X"4C",X"BB",X"4C",
		X"00",X"BB",X"00",X"CB",X"00",X"CB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"44",X"BB",X"44",X"BB",X"44",X"CB",X"4C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"00",X"BB",X"C0",
		X"00",X"FB",X"00",X"FB",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"4C",X"BB",X"4C",X"BB",X"4C",X"BB",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BF",X"00",X"FB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B4",X"00",X"BB",X"C0",X"BB",X"4C",X"BB",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B4",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"C4",X"00",X"0C",X"00",X"0B",X"0B",X"BB",X"BB",X"BB",
		X"0F",X"00",X"FF",X"BC",X"FF",X"BB",X"BF",X"BF",X"BB",X"FC",X"CB",X"FF",X"BC",X"4F",X"BB",X"44",
		X"BB",X"BB",X"CB",X"BB",X"0B",X"BB",X"0C",X"BB",X"00",X"BB",X"00",X"44",X"0B",X"C4",X"BC",X"0C",
		X"BB",X"44",X"BB",X"44",X"BB",X"CC",X"44",X"C0",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"0F",X"FC",X"FF",X"CF",X"FF",X"CF",X"FF",X"CF",X"FF",X"CF",
		X"00",X"00",X"FF",X"00",X"FF",X"FF",X"CC",X"FF",X"FF",X"FC",X"CC",X"FC",X"FC",X"FC",X"FC",X"FF",
		X"0F",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"CC",X"FF",X"FF",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"BF",X"00",X"FB",X"00",X"FF",X"00",X"FF",X"00",X"CF",X"00",X"FF",
		X"00",X"00",X"B4",X"00",X"BB",X"C0",X"BB",X"C0",X"BB",X"4C",X"BF",X"FC",X"BF",X"FC",X"BB",X"4C",
		X"00",X"BB",X"00",X"CB",X"0B",X"4C",X"0B",X"44",X"0B",X"4C",X"0C",X"C0",X"00",X"00",X"00",X"00",
		X"CB",X"C0",X"CC",X"B4",X"CB",X"BB",X"BC",X"BB",X"C0",X"B4",X"00",X"4C",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"FB",X"00",X"BB",X"00",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"B4",X"C0",X"BB",X"C0",X"BB",X"4C",X"BB",X"4C",
		X"00",X"CB",X"00",X"BB",X"00",X"BB",X"00",X"CB",X"00",X"4C",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"BB",X"4C",X"CB",X"4C",X"CB",X"CB",X"BB",X"B4",X"CC",X"4C",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"BB",X"C0",X"BB",X"C0",
		X"00",X"BB",X"00",X"CB",X"00",X"CB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"4C",X"BB",X"4C",X"BB",X"4C",X"CB",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"00",
		X"00",X"BB",X"00",X"BF",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"C0",X"BB",X"C0",X"BB",X"C0",X"BB",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"FB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B4",X"00",X"BB",X"C0",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B4",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"0B",X"0B",X"BB",X"0B",X"BB",
		X"00",X"00",X"0F",X"BC",X"BF",X"B4",X"BF",X"44",X"BB",X"FF",X"CB",X"FC",X"CC",X"FF",X"CC",X"44",
		X"0B",X"BB",X"0C",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"44",X"00",X"C4",X"04",X"00",X"0C",X"00",
		X"BB",X"4C",X"BB",X"44",X"44",X"44",X"44",X"C4",X"4C",X"0C",X"4C",X"00",X"44",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"00",X"F0",X"00",X"00",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FB",
		X"32",X"00",X"33",X"00",X"33",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"2C",X"CF",X"22",X"BF",X"22",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"BB",X"FF",X"BC",X"CC",X"C0",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",
		X"33",X"00",X"33",X"C0",X"33",X"C0",X"3F",X"2C",X"3F",X"2C",X"3C",X"2C",X"BB",X"32",X"BF",X"32",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"33",X"00",X"3F",X"00",X"3F",X"00",X"3F",X"03",X"33",
		X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"F2",X"33",X"F2",X"33",X"F2",X"BB",X"32",
		X"33",X"3F",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"BB",X"00",X"CC",
		X"BB",X"F2",X"FF",X"FC",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"FF",X"00",X"CC",X"00",X"FC",X"30",X"BB",X"33",X"FF",
		X"32",X"00",X"33",X"00",X"33",X"00",X"33",X"C0",X"33",X"C0",X"33",X"2C",X"33",X"32",X"33",X"33",
		X"C3",X"FF",X"0C",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0B",X"FF",X"0C",X"BF",X"00",X"CC",
		X"33",X"32",X"F3",X"2C",X"F3",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"2C",X"BB",X"C0",X"BB",X"C0",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"3F",
		X"33",X"00",X"33",X"C0",X"33",X"C0",X"3F",X"2C",X"3C",X"2C",X"3F",X"2C",X"BB",X"32",X"BF",X"32",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"33",X"00",X"33",X"30",X"33",X"33",X"33",
		X"33",X"C0",X"33",X"2C",X"33",X"2C",X"3F",X"2F",X"FC",X"2C",X"FC",X"BB",X"FF",X"CC",X"33",X"BF",
		X"C3",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"3F",X"00",X"CF",X"00",X"0B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FB",X"BF",X"BB",X"BF",X"BB",X"CC",X"CC",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"3F",
		X"33",X"00",X"33",X"C0",X"33",X"C0",X"3F",X"2C",X"3C",X"2C",X"BF",X"2C",X"CB",X"32",X"BF",X"32",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"33",X"00",X"3F",X"00",X"F3",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"32",X"00",X"33",X"00",X"33",X"00",X"33",X"C0",X"33",X"C0",X"33",X"2C",X"33",X"22",X"33",X"22",
		X"03",X"33",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"0C",X"33",X"0C",X"BC",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"3C",X"CC",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",
		X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",
		X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"0B",X"33",X"0C",X"33",X"00",X"C3",
		X"33",X"22",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2C",X"22",X"BB",X"2C",X"BB",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",
		X"33",X"00",X"33",X"C0",X"33",X"C0",X"3F",X"2C",X"3F",X"2C",X"3C",X"2C",X"BB",X"32",X"BF",X"32",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FB",
		X"32",X"00",X"33",X"00",X"33",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"2C",X"CF",X"22",X"BF",X"22",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"22",X"FF",X"BB",X"FF",X"BC",X"CC",X"C0",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",
		X"33",X"00",X"33",X"C0",X"33",X"C0",X"3F",X"2C",X"3F",X"2C",X"3C",X"2C",X"BB",X"32",X"BF",X"32",
		X"03",X"FF",X"33",X"FF",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"33",X"00",X"3F",X"00",X"3F",X"00",X"3F",X"03",X"33",
		X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"F2",X"33",X"F2",X"33",X"F2",X"BB",X"32",
		X"33",X"3F",X"3C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"BB",X"00",X"CC",
		X"BB",X"F2",X"FF",X"FC",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"00",X"00",X"06",X"00",X"0F",X"00",X"66",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"06",X"66",
		X"66",X"C0",X"66",X"5C",X"66",X"5C",X"66",X"5C",X"66",X"F5",X"66",X"F5",X"66",X"F5",X"BB",X"65",
		X"66",X"6F",X"6C",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"BB",X"00",X"CC",
		X"BB",X"F5",X"FF",X"FC",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"5C",X"FF",X"BC",X"CC",X"BB",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"D1",X"11",X"ED",X"D1",X"EE",X"ED",X"FF",X"FE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"11",X"1F",X"DD",X"FF",X"EE",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"D1",X"11",X"ED",X"11",X"FE",X"11",X"FE",X"1E",X"FE",X"1E",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"D1",X"11",X"D1",X"11",
		X"FF",X"EF",X"EF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"DD",X"11",X"ED",X"11",X"ED",X"11",X"EE",X"11",X"FE",X"11",X"FF",X"D1",X"FF",X"DD",X"EF",X"ED",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"EE",X"FF",X"FE",X"FF",X"FF",X"FF",X"EF",X"FF",X"EF",X"FF",X"DD",X"FF",X"EF",X"FE",X"FE",X"EE",
		X"EE",X"DF",X"EE",X"ED",X"EF",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"DD",X"FE",X"EE",X"FF",X"EF",X"EE",X"EF",X"EF",X"FF",X"FF",X"EF",X"FF",X"EF",X"FF",X"FF",
		X"FF",X"EE",X"FF",X"FE",X"EE",X"FF",X"DD",X"FF",X"FD",X"EF",X"FE",X"DE",X"FF",X"DD",X"EF",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"EF",X"FF",X"DE",
		X"EE",X"FF",X"FE",X"FD",X"FF",X"DE",X"FD",X"FE",X"EE",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"EF",
		X"FF",X"EE",X"FE",X"FF",X"FF",X"FF",X"FD",X"FE",X"FF",X"FF",X"EE",X"FF",X"DD",X"EF",X"EE",X"DD",
		X"FF",X"FE",X"FE",X"FF",X"EF",X"FF",X"FF",X"FE",X"FF",X"EE",X"EF",X"FF",X"FF",X"EF",X"EE",X"FE",
		X"11",X"11",X"11",X"11",X"D1",X"11",X"DD",X"11",X"FE",X"11",X"FF",X"D1",X"FF",X"DD",X"FF",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",
		X"FF",X"EE",X"FF",X"EE",X"FF",X"FE",X"EE",X"FF",X"EF",X"FF",X"DD",X"FF",X"FF",X"FF",X"FF",X"DD",
		X"FF",X"DD",X"EF",X"FE",X"EE",X"FF",X"EE",X"EE",X"EE",X"EF",X"FE",X"EF",X"FF",X"EE",X"FF",X"FE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"D1",X"11",X"ED",X"FD",X"FE",X"EF",X"FD",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",
		X"11",X"11",X"FD",X"11",X"DE",X"FF",X"EE",X"DD",X"DE",X"EF",X"ED",X"EF",X"FF",X"EE",X"FE",X"DD",
		X"11",X"11",X"FD",X"11",X"FF",X"FE",X"FF",X"EF",X"FF",X"EF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FE",
		X"ED",X"11",X"FE",X"11",X"FE",X"D1",X"FF",X"ED",X"FF",X"EF",X"FF",X"EF",X"FF",X"EE",X"FF",X"DD",
		X"11",X"11",X"11",X"1F",X"11",X"FE",X"1F",X"EF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",
		X"ED",X"11",X"FE",X"11",X"FF",X"D1",X"FF",X"ED",X"FE",X"FE",X"FF",X"FF",X"FF",X"EF",X"EE",X"FE",
		X"11",X"11",X"11",X"11",X"11",X"FF",X"11",X"FF",X"DD",X"FF",X"FF",X"FF",X"FE",X"EE",X"EF",X"FF",
		X"11",X"11",X"D1",X"11",X"ED",X"11",X"FE",X"FF",X"FF",X"EE",X"FF",X"FE",X"FF",X"FF",X"EE",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"D1",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"FE",X"11",X"FE",X"11",X"FF",X"D1",X"EE",X"ED",X"FE",X"FE",X"FE",X"FF",X"FF",X"EF",
		X"11",X"11",X"11",X"D1",X"DF",X"FD",X"ED",X"FF",X"FE",X"FF",X"FF",X"DF",X"FF",X"ED",X"FF",X"FF",
		X"11",X"1D",X"11",X"FE",X"11",X"EF",X"1F",X"FE",X"DE",X"FF",X"FE",X"FF",X"FF",X"DD",X"FF",X"FE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"ED",X"EF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"D1",X"EE",X"ED",X"FD",X"FE",X"FE",X"FF",X"FF",X"DF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",X"FF",X"D1",X"FF",X"DD",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"1E",X"FE",X"FF",X"FF",X"FF",X"FE",X"EE",X"FF",X"FE",X"EF",
		X"11",X"11",X"11",X"11",X"11",X"1F",X"11",X"FF",X"11",X"FF",X"FF",X"EF",X"FF",X"EF",X"FF",X"FF",
		X"D1",X"11",X"ED",X"11",X"FD",X"11",X"EE",X"D1",X"FE",X"ED",X"FF",X"EE",X"FF",X"DD",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"FF",X"1F",X"FF",X"EF",X"DF",X"FF",X"ED",X"FE",X"FF",X"EE",X"FF",X"FF",X"FE",
		X"11",X"1F",X"11",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FE",X"FF",X"EF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",X"EE",X"D1",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"EE",
		X"FF",X"ED",X"FF",X"FE",X"FF",X"FD",X"FF",X"DE",X"FE",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1E",X"FF",X"DE",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"DD",X"FF",X"EE",X"FF",X"FE",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"11",X"FF",X"DE",X"EF",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"DD",X"FF",X"EF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"EE",X"EF",X"EF",X"FF",X"FF",X"DE",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",X"EE",X"1E",X"FE",X"EF",X"FF",X"EF",X"FE",X"FF",
		X"11",X"D1",X"11",X"DD",X"1F",X"ED",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"EF",X"FF",X"EF",X"FF",X"FF",X"FE",X"FF",
		X"FE",X"EF",X"FF",X"DD",X"FF",X"EE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"12",X"11",X"2F",X"11",X"FF",X"11",X"FF",X"12",X"FF",X"2F",X"FF",
		X"21",X"11",X"F2",X"11",X"FF",X"11",X"FF",X"11",X"FF",X"21",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",
		X"22",X"22",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",
		X"22",X"22",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"22",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"22",X"22",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"2E",X"EE",X"22",X"22",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"22",X"22",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"22",X"22",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"AB",X"00",X"AB",X"11",X"FE",X"11",X"FE",X"11",X"FE",X"11",X"FE",X"11",X"FE",X"11",X"FE",X"11",
		X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",
		X"FE",X"11",X"FE",X"11",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",
		X"11",X"10",X"11",X"10",X"11",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"5A",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"55",X"5A",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"AA",X"55",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"12",X"22",X"11",X"22",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"12",X"11",X"22",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"12",X"22",X"11",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"22",X"21",
		X"12",X"22",X"12",X"22",X"11",X"22",X"11",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0C",X"00",X"0C",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"3F",X"00",X"FF",X"00",X"FC",X"00",X"FF",X"00",X"3F",
		X"33",X"00",X"33",X"C0",X"33",X"C0",X"3F",X"2C",X"3F",X"2C",X"3F",X"2C",X"BB",X"32",X"BF",X"32",
		X"03",X"FF",X"33",X"FF",X"30",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BB",
		X"FF",X"32",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"2C",X"FF",X"BC",X"CC",X"BB",
		X"00",X"03",X"00",X"3F",X"00",X"F3",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"32",X"00",X"33",X"C0",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",
		X"03",X"33",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"0B",X"33",X"0C",X"33",X"00",X"C3",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"32",X"CC",
		X"00",X"33",X"00",X"3F",X"00",X"F3",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"32",X"00",X"33",X"00",X"33",X"00",X"33",X"C0",X"33",X"C0",X"33",X"2C",X"33",X"22",X"33",X"22",
		X"03",X"33",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"0C",X"33",X"0C",X"BC",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"3C",X"CC",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",
		X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",
		X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"0B",X"33",X"0C",X"33",X"00",X"C3",
		X"33",X"22",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2C",X"22",X"BB",X"2C",X"BB",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"4F",
		X"44",X"11",X"4F",X"11",X"EF",X"11",X"F1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"EF",X"44",X"F1",X"44",X"11",X"44",X"11",X"44",X"11",X"4F",X"11",X"EF",X"11",X"F1",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"4F",X"44",X"EF",X"44",X"F1",X"44",X"11",X"44",X"11",
		X"11",X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"44",X"FE",X"44",X"1F",X"44",X"11",X"44",
		X"F4",X"44",X"FE",X"44",X"1F",X"44",X"11",X"44",X"11",X"44",X"11",X"44",X"11",X"F4",X"11",X"FE",
		X"11",X"44",X"11",X"44",X"11",X"F4",X"11",X"FE",X"11",X"1F",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"4F",X"44",X"EF",X"44",X"FE",X"44",X"FE",X"44",X"EE",
		X"F4",X"44",X"FE",X"44",X"EF",X"44",X"EF",X"44",X"EE",X"44",X"EE",X"44",X"EE",X"F4",X"EE",X"FE",
		X"44",X"EE",X"4F",X"EE",X"EF",X"EE",X"FE",X"EE",X"FF",X"FF",X"FD",X"DD",X"FD",X"DD",X"FF",X"FF",
		X"EE",X"EF",X"EE",X"EF",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"4E",X"FF",X"4F",X"EE",X"FE",X"EE",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FD",X"DD",X"FD",X"DD",X"FD",X"DD",X"FD",X"DD",X"FF",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"EF",X"44",X"F1",X"44",X"11",X"44",X"11",X"44",X"11",X"4F",X"11",X"EF",X"FF",X"FF",X"FF",
		X"11",X"44",X"11",X"44",X"11",X"F4",X"11",X"FE",X"11",X"1F",X"11",X"11",X"FF",X"FF",X"FF",X"FF",
		X"44",X"22",X"44",X"22",X"44",X"22",X"42",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"22",X"24",X"22",X"22",X"22",X"22",X"22",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"44",X"44",X"44",X"44",X"44",X"42",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"24",X"44",X"22",X"44",X"22",X"44",
		X"44",X"42",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"22",X"44",X"22",X"44",X"22",X"24",X"22",X"24",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"44",X"F2",X"44",X"22",X"44",X"44",X"44",
		X"FE",X"11",X"FF",X"11",X"FF",X"EF",X"FF",X"FF",X"EF",X"EE",X"EF",X"FE",X"EE",X"FF",X"FE",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"FF",X"12",X"11",X"11",X"12",X"42",X"42",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"4F",X"12",X"4F",X"11",X"4F",X"42",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"4F",X"4F",X"2F",X"2F",X"4F",X"2F",X"24",X"24",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"4F",X"44",X"2F",X"2F",X"2F",X"2F",X"24",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"4F",X"4F",X"4F",X"4F",X"2F",X"24",X"24",X"24",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"24",X"44",X"24",X"F4",X"44",X"22",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"F4",X"FF",X"F2",X"F2",X"F2",X"42",X"42",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"F4",X"22",X"22",X"24",X"F4",X"24",X"22",X"44",X"44",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",
		X"FF",X"FF",X"FF",X"FF",X"22",X"22",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"22",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"88",X"AA",X"88",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"88",X"CC",X"88",X"F8",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"88",X"CC",
		X"88",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"88",X"8C",X"88",X"8F",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"8F",X"FF",X"CF",X"8C",X"CF",X"FF",
		X"88",X"F8",X"FF",X"FF",X"CC",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"8F",X"8C",X"8F",X"FF",X"C8",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"8F",X"8F",X"F8",X"8F",X"FF",X"CF",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"8F",X"FF",X"8F",X"8C",X"CF",X"FF",
		X"FC",X"CF",X"FC",X"C8",X"8C",X"C8",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"CF",X"CC",X"F8",X"C8",X"8C",X"C8",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",X"C8",X"88",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"CB",X"BC",X"CB",X"BC",X"CB",X"BC",X"BB",X"BB",X"BB",
		X"0B",X"00",X"BC",X"00",X"BC",X"00",X"C4",X"00",X"CC",X"C0",X"CC",X"4C",X"CC",X"4C",X"B4",X"C0",
		X"CB",X"BC",X"0C",X"CF",X"BB",X"FF",X"BC",X"FF",X"CB",X"FF",X"BF",X"FF",X"BB",X"FF",X"BB",X"FF",
		X"44",X"00",X"CC",X"00",X"B4",X"00",X"4C",X"00",X"F4",X"00",X"FF",X"00",X"FF",X"00",X"44",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"C0",X"0B",X"BB",X"0B",X"CC",X"BB",X"CC",X"BB",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"C0",X"BB",X"C0",X"CC",X"C0",X"CC",X"4C",X"FC",X"44",
		X"BB",X"CB",X"BB",X"BB",X"CC",X"BB",X"BB",X"CC",X"BB",X"BB",X"00",X"FF",X"0B",X"FF",X"0B",X"FF",
		X"CC",X"44",X"BB",X"4C",X"B4",X"C0",X"CC",X"4C",X"BB",X"44",X"F4",X"C0",X"FF",X"C0",X"FF",X"C0",
		X"00",X"00",X"0B",X"C0",X"0B",X"BB",X"0B",X"CC",X"BB",X"CC",X"BB",X"FC",X"BB",X"CB",X"BB",X"BB",
		X"00",X"00",X"0B",X"C0",X"BB",X"C0",X"CC",X"C0",X"CC",X"4C",X"FC",X"44",X"CC",X"44",X"BB",X"4C",
		X"CC",X"BB",X"00",X"CC",X"0B",X"FF",X"BB",X"FF",X"CC",X"FF",X"0B",X"FF",X"0B",X"FF",X"BB",X"FF",
		X"B4",X"C0",X"CC",X"00",X"FB",X"C0",X"F4",X"4C",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"F4",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"BB",X"BB",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"00",X"B4",X"00",X"CB",X"C0",
		X"BC",X"CB",X"BC",X"CB",X"BC",X"BB",X"CB",X"BC",X"BC",X"CF",X"BC",X"FF",X"BB",X"FF",X"BB",X"FF",
		X"CC",X"4C",X"CC",X"4C",X"CC",X"C0",X"44",X"00",X"CC",X"00",X"BC",X"C0",X"C4",X"C0",X"C4",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"CB",X"BC",X"CB",X"BC",X"CB",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"00",X"C4",X"00",X"CC",X"C0",X"CC",X"4C",
		X"BC",X"BB",X"CB",X"BB",X"BC",X"BC",X"BC",X"CB",X"BB",X"BB",X"BB",X"FF",X"BB",X"FF",X"BF",X"FF",
		X"CC",X"4C",X"B4",X"C0",X"44",X"00",X"CC",X"C0",X"B4",X"4C",X"44",X"00",X"F4",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"CC",X"BB",X"CC",X"BB",X"FC",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"B4",X"00",X"CC",X"00",X"CC",X"C0",X"FC",X"4C",
		X"BB",X"CB",X"CC",X"BB",X"BB",X"BB",X"BB",X"CC",X"BC",X"BB",X"BB",X"FF",X"BB",X"FF",X"BF",X"FF",
		X"CC",X"4C",X"B4",X"C0",X"44",X"00",X"CC",X"C0",X"B4",X"4C",X"44",X"C0",X"F4",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"BB",X"BB",X"BB",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BC",X"00",X"B4",X"00",X"CC",X"C0",
		X"BB",X"CC",X"BB",X"FC",X"BB",X"CB",X"CB",X"BB",X"BB",X"CC",X"BB",X"FF",X"BB",X"FF",X"CB",X"CF",
		X"CC",X"4C",X"FC",X"4C",X"CC",X"C0",X"44",X"00",X"CC",X"4C",X"F4",X"C0",X"FF",X"00",X"FF",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"CB",X"BC",X"BB",X"BB",X"BC",X"BB",X"CC",X"BB",X"CC",X"BB",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"CC",X"00",X"BB",X"C0",X"BB",X"4C",X"B4",X"4C",X"B4",X"C0",
		X"BB",X"FF",X"BF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"4F",X"FF",X"44",X"FF",X"CC",X"44",
		X"F4",X"C0",X"FF",X"00",X"FF",X"C0",X"FF",X"4C",X"FF",X"4C",X"FF",X"C0",X"44",X"C0",X"4C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BC",X"BC",X"BB",X"CC",X"BB",X"FF",X"BB",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"CC",X"00",X"B4",X"C0",X"B4",X"C0",X"F4",X"C0",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"FF",X"44",X"FF",X"CC",X"44",X"00",X"CC",
		X"FF",X"00",X"FF",X"C0",X"FF",X"4C",X"FF",X"4C",X"FF",X"C0",X"44",X"C0",X"4C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BC",X"BC",X"BB",X"FF",X"BB",X"FE",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"CC",X"00",X"B4",X"C0",X"F4",X"C0",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"44",X"FF",X"44",X"44",X"CC",X"CC",
		X"FF",X"00",X"FF",X"4C",X"FF",X"4C",X"FF",X"C0",X"FF",X"4C",X"44",X"4C",X"44",X"4C",X"CC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"BC",X"BB",X"BB",X"BB",X"BB",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"00",X"BC",X"00",X"B4",X"00",X"CB",X"C0",
		X"BC",X"CB",X"BC",X"CB",X"BB",X"BB",X"BB",X"BC",X"BC",X"CF",X"BC",X"FF",X"BB",X"FF",X"BF",X"FF",
		X"CC",X"4C",X"CC",X"4C",X"44",X"C0",X"44",X"00",X"C4",X"00",X"BC",X"C0",X"F4",X"C0",X"FF",X"00",
		X"00",X"BB",X"00",X"B0",X"00",X"B0",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"0B",X"B0",X"0B",
		X"00",X"00",X"B0",X"00",X"BB",X"00",X"0B",X"00",X"00",X"B0",X"00",X"BB",X"00",X"0B",X"00",X"0B",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"B0",X"0B",X"BB",X"BB",X"0B",X"B0",
		X"00",X"0B",X"BB",X"BB",X"BB",X"B0",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"FF",X"98",X"FF",X"98",X"FF",X"98",X"FF",X"88",X"FF",X"08",X"FF",X"08",X"8F",X"09",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"99",X"88",X"99",X"88",X"99",X"88",X"88",X"80",X"CC",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"EE",X"FF",X"EE",X"FF",X"CC",
		X"88",X"8C",X"88",X"8C",X"88",X"88",X"88",X"88",X"CC",X"88",X"99",X"88",X"98",X"88",X"88",X"88",
		X"FE",X"98",X"EE",X"89",X"00",X"89",X"00",X"89",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8C",X"89",X"8C",X"98",X"C0",X"98",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"0F",X"99",X"55",X"99",X"55",X"99",X"05",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"00",X"95",X"00",X"95",X"50",X"98",X"50",X"98",X"00",
		X"90",X"99",X"99",X"00",X"09",X"08",X"09",X"09",X"09",X"09",X"00",X"09",X"00",X"99",X"00",X"89",
		X"98",X"99",X"00",X"89",X"00",X"08",X"00",X"08",X"00",X"08",X"09",X"00",X"88",X"00",X"80",X"00",
		X"0F",X"00",X"0F",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FE",X"00",X"CE",X"00",X"CF",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"F6",X"00",
		X"F5",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"0F",X"00",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"F5",X"00",X"FF",X"00",X"FE",X"00",X"E0",X"00",X"00",X"00",X"F0",X"F0",X"EE",X"F0",X"EE",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"44",X"0B",X"44",X"BB",X"F4",X"B4",X"FF",X"44",X"CF",X"C4",X"11",
		X"00",X"00",X"C0",X"00",X"44",X"00",X"44",X"00",X"F4",X"C0",X"FF",X"C0",X"FF",X"C0",X"11",X"00",
		X"BC",X"14",X"BC",X"11",X"44",X"DF",X"C4",X"44",X"0C",X"CC",X"00",X"11",X"C4",X"11",X"04",X"11",
		X"14",X"C0",X"14",X"4C",X"FC",X"4C",X"4C",X"44",X"C4",X"B4",X"14",X"04",X"11",X"11",X"11",X"01",
		X"00",X"B4",X"00",X"44",X"0B",X"44",X"0B",X"14",X"0B",X"11",X"BB",X"11",X"41",X"11",X"1F",X"11",
		X"40",X"00",X"44",X"00",X"44",X"00",X"14",X"00",X"11",X"00",X"01",X"00",X"11",X"40",X"FC",X"40",
		X"1F",X"CF",X"41",X"CF",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"40",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",X"BB",X"0B",X"00",X"BB",X"00",X"BB",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"00",X"40",X"F0",X"44",
		X"BB",X"0B",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"FF",X"0B",X"FF",X"0B",X"FF",
		X"00",X"44",X"BB",X"40",X"B4",X"00",X"00",X"40",X"BB",X"40",X"F4",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",X"BB",X"0B",X"00",X"BB",X"00",X"BB",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"00",X"40",X"F0",X"44",
		X"BB",X"0B",X"BB",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"FF",X"BB",X"FF",X"00",X"FF",
		X"00",X"44",X"BB",X"40",X"B4",X"00",X"00",X"00",X"BB",X"00",X"F4",X"40",X"FF",X"40",X"FF",X"00",
		X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"F3",X"03",X"CF",X"03",X"CF",X"03",X"AA",X"33",X"AA",
		X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"F3",X"00",X"F3",X"00",X"F3",X"00",X"A3",X"30",
		X"33",X"AA",X"33",X"FF",X"33",X"FF",X"30",X"FF",X"00",X"FF",X"00",X"FF",X"0A",X"AF",X"AA",X"AA",
		X"33",X"33",X"F3",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"A0",X"FA",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"09",X"09",X"08",X"00",X"88",X"88",X"88",X"08",X"D8",X"8D",X"ED",X"88",X"5E",X"8E",X"EE",
		X"90",X"00",X"00",X"00",X"88",X"00",X"88",X"80",X"DD",X"09",X"5E",X"00",X"C5",X"80",X"EE",X"09",
		X"0E",X"EE",X"0E",X"FF",X"00",X"CC",X"00",X"FF",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"00",X"EE",X"00",X"ED",X"00",X"D0",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"88",X"28",X"88",X"26",X"88",X"26",X"88",X"25",X"88",X"28",X"88",X"2C",X"88",X"22",X"88",
		X"C2",X"22",X"88",X"22",X"86",X"22",X"66",X"22",X"55",X"22",X"88",X"22",X"8C",X"22",X"8C",X"22",
		X"22",X"88",X"22",X"CC",X"28",X"AA",X"28",X"AA",X"88",X"AA",X"8C",X"AA",X"C8",X"AA",X"88",X"AA",
		X"C2",X"22",X"8C",X"22",X"88",X"22",X"88",X"22",X"88",X"C2",X"AC",X"C8",X"A8",X"28",X"A8",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"03",X"33",X"03",X"F3",X"33",X"F3",X"33",X"F3",
		X"00",X"00",X"00",X"00",X"20",X"00",X"32",X"00",X"33",X"00",X"F3",X"00",X"FF",X"00",X"CF",X"00",
		X"33",X"BB",X"33",X"FB",X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"03",X"FF",
		X"FF",X"00",X"F3",X"00",X"FF",X"30",X"FF",X"23",X"FF",X"02",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"06",X"66",X"06",X"F6",X"66",X"F6",X"66",X"F6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"F6",X"00",X"FF",X"00",X"CF",X"00",
		X"66",X"AA",X"66",X"CA",X"66",X"FC",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"06",X"FF",
		X"FF",X"00",X"F6",X"00",X"FF",X"60",X"FF",X"56",X"FF",X"05",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"06",X"66",X"06",X"F6",X"66",X"F6",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"F6",X"00",X"FF",X"00",X"FF",X"00",
		X"66",X"AA",X"66",X"CA",X"66",X"FC",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"06",X"FF",
		X"FF",X"00",X"F6",X"00",X"FF",X"60",X"FF",X"56",X"FF",X"05",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"05",X"00",X"05",X"00",X"65",X"00",X"65",X"06",X"65",X"06",X"66",X"6F",X"F6",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"66",X"AA",X"66",X"CA",X"6F",X"FC",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",
		X"66",X"00",X"FF",X"00",X"FF",X"60",X"FF",X"66",X"FF",X"56",X"FF",X"55",X"FF",X"05",X"FF",X"00",
		X"00",X"00",X"00",X"AA",X"06",X"AA",X"F5",X"AA",X"55",X"AA",X"A5",X"AA",X"0A",X"AA",X"00",X"AA",
		X"00",X"00",X"AA",X"00",X"AA",X"00",X"AF",X"00",X"A5",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"CC",X"0A",X"AC",X"00",X"44",X"AA",X"CC",X"0A",X"BB",X"00",X"44",X"AA",X"CC",X"0A",X"BB",
		X"AC",X"A0",X"CB",X"0A",X"4C",X"00",X"CB",X"A0",X"BB",X"0A",X"4C",X"00",X"CB",X"A0",X"BB",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"F0",X"35",X"70",X"30",X"8A",X"30",X"F0",X"3D",X"7A",
		X"00",X"00",X"00",X"00",X"5F",X"00",X"A0",X"00",X"70",X"F0",X"76",X"00",X"50",X"00",X"80",X"F3",
		X"38",X"08",X"95",X"75",X"00",X"A0",X"A0",X"84",X"60",X"A1",X"05",X"FF",X"00",X"00",X"00",X"77",
		X"E5",X"F0",X"02",X"01",X"A2",X"30",X"70",X"76",X"3A",X"97",X"0A",X"00",X"DA",X"00",X"60",X"00",
		X"00",X"05",X"00",X"05",X"00",X"65",X"00",X"65",X"06",X"65",X"06",X"66",X"6F",X"F6",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"05",
		X"66",X"AA",X"66",X"CC",X"6F",X"AC",X"6F",X"CA",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",
		X"66",X"05",X"AF",X"55",X"CF",X"55",X"FF",X"50",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"C0",X"F3",X"FC",X"F3",X"F2",X"F3",X"F2",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"33",X"C0",
		X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"22",X"33",X"CC",X"22",X"00",X"CC",X"00",X"00",
		X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"2C",X"33",X"C0",X"22",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"FF",X"C0",X"CF",X"2C",X"FF",X"22",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"33",X"20",
		X"33",X"32",X"33",X"33",X"33",X"33",X"23",X"33",X"C2",X"23",X"0C",X"C2",X"00",X"0C",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"2C",X"F3",X"F2",X"C3",X"F2",X"F3",X"F2",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"32",X"00",X"23",X"2C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"23",X"33",X"22",X"33",X"CC",X"22",X"00",X"CC",X"00",X"00",
		X"23",X"32",X"33",X"32",X"33",X"32",X"33",X"2C",X"32",X"CC",X"2C",X"C0",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"AB",X"00",X"AB",X"0A",X"CB",X"0A",X"AB",X"0C",X"AB",X"CA",X"AB",
		X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"00",X"BB",X"00",X"AC",X"00",X"CA",X"C0",X"CA",X"C0",
		X"CA",X"AC",X"CA",X"CA",X"CA",X"CA",X"CA",X"CA",X"CA",X"CA",X"0C",X"CA",X"00",X"CC",X"00",X"00",
		X"CA",X"C0",X"CA",X"C0",X"CA",X"C0",X"CA",X"C0",X"CA",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"BB",X"BB",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"00",X"B4",X"00",X"CB",X"C0",
		X"BC",X"CB",X"BC",X"CB",X"BC",X"BB",X"CB",X"BC",X"BC",X"CF",X"BC",X"FF",X"BB",X"FF",X"BB",X"FF",
		X"CC",X"4C",X"CC",X"4C",X"CC",X"C0",X"44",X"00",X"CC",X"00",X"BC",X"C0",X"C4",X"C0",X"C4",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"CB",X"BC",X"CB",X"BC",X"CB",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"00",X"C4",X"00",X"CC",X"C0",X"CC",X"4C",
		X"BC",X"BB",X"CB",X"BB",X"BC",X"BC",X"BC",X"CB",X"BB",X"BB",X"BB",X"FF",X"BB",X"FF",X"BF",X"FF",
		X"CC",X"4C",X"B4",X"C0",X"44",X"00",X"CC",X"C0",X"B4",X"4C",X"44",X"00",X"F4",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"BC",X"BB",X"BB",X"CC",X"BB",X"CC",X"BB",X"FC",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"00",X"B4",X"00",X"CC",X"00",X"CC",X"C0",X"FC",X"4C",
		X"BB",X"CB",X"CC",X"BB",X"BB",X"BB",X"BB",X"CC",X"BC",X"BB",X"BB",X"FF",X"BB",X"FF",X"BF",X"FF",
		X"CC",X"4C",X"B4",X"C0",X"44",X"00",X"CC",X"C0",X"B4",X"4C",X"44",X"C0",X"F4",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BC",X"BB",X"BB",X"BB",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BC",X"00",X"B4",X"00",X"CC",X"C0",
		X"BB",X"CC",X"BB",X"FC",X"BB",X"CB",X"CB",X"BB",X"BB",X"CC",X"BB",X"FF",X"BB",X"FF",X"CB",X"CF",
		X"CC",X"4C",X"FC",X"4C",X"CC",X"C0",X"44",X"00",X"CC",X"4C",X"F4",X"C0",X"FF",X"00",X"FF",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"CB",X"BC",X"BB",X"BB",X"BC",X"BB",X"CC",X"BB",X"CC",X"BB",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"CC",X"00",X"BB",X"C0",X"BB",X"4C",X"B4",X"4C",X"B4",X"C0",
		X"BB",X"FF",X"BF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"4F",X"FF",X"44",X"FF",X"CC",X"44",
		X"F4",X"C0",X"FF",X"00",X"FF",X"C0",X"FF",X"4C",X"FF",X"4C",X"FF",X"C0",X"44",X"C0",X"4C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"06",X"66",X"06",X"F6",X"66",X"F6",X"66",X"F6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"F6",X"00",X"FF",X"00",X"CF",X"00",
		X"66",X"AA",X"66",X"CA",X"66",X"FC",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"06",X"FF",
		X"FF",X"00",X"F6",X"00",X"FF",X"60",X"FF",X"56",X"FF",X"05",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"06",X"66",X"06",X"F6",X"66",X"F6",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"F6",X"00",X"FF",X"00",X"FF",X"00",
		X"66",X"AA",X"66",X"CA",X"66",X"FC",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"06",X"FF",
		X"FF",X"00",X"F6",X"00",X"FF",X"60",X"FF",X"56",X"FF",X"05",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"05",X"00",X"05",X"00",X"65",X"00",X"65",X"06",X"65",X"06",X"66",X"6F",X"F6",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"66",X"AA",X"66",X"CA",X"6F",X"FC",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",
		X"66",X"00",X"FF",X"00",X"FF",X"60",X"FF",X"66",X"FF",X"56",X"FF",X"55",X"FF",X"05",X"FF",X"00",
		X"00",X"00",X"00",X"AA",X"06",X"AA",X"F5",X"AA",X"55",X"AA",X"A5",X"AA",X"0A",X"AA",X"00",X"AA",
		X"00",X"00",X"AA",X"00",X"AA",X"00",X"AF",X"00",X"A5",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"CC",X"0A",X"AC",X"00",X"44",X"AA",X"CC",X"0A",X"BB",X"00",X"44",X"AA",X"CC",X"0A",X"BB",
		X"AC",X"A0",X"CB",X"0A",X"4C",X"00",X"CB",X"A0",X"BB",X"0A",X"4C",X"00",X"CB",X"A0",X"BB",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"F0",X"35",X"70",X"30",X"8A",X"30",X"F0",X"3D",X"7A",
		X"00",X"00",X"00",X"00",X"5F",X"00",X"A0",X"00",X"70",X"F0",X"76",X"00",X"50",X"00",X"80",X"F3",
		X"38",X"08",X"95",X"75",X"00",X"A0",X"A0",X"84",X"60",X"A1",X"05",X"FF",X"00",X"00",X"00",X"77",
		X"E5",X"F0",X"02",X"01",X"A2",X"30",X"70",X"76",X"3A",X"97",X"0A",X"00",X"DA",X"00",X"60",X"00",
		X"00",X"05",X"00",X"05",X"00",X"65",X"00",X"65",X"06",X"65",X"06",X"66",X"6F",X"F6",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"65",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"05",
		X"66",X"AA",X"66",X"CC",X"6F",X"AC",X"6F",X"CA",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",
		X"66",X"05",X"AF",X"55",X"CF",X"55",X"FF",X"50",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"BB",X"00",X"BB",X"0F",X"BB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"BF",X"BB",X"BB",X"BC",
		X"4C",X"00",X"44",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"CF",X"C0",X"FF",X"C0",X"B4",X"C0",
		X"CC",X"BC",X"BB",X"CC",X"B4",X"BB",X"B4",X"CB",X"44",X"00",X"C4",X"00",X"0C",X"00",X"00",X"00",
		X"C4",X"00",X"BC",X"4C",X"CB",X"44",X"BB",X"B4",X"CB",X"4C",X"0C",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"0B",X"BB",X"0B",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"4C",X"00",X"44",X"00",X"B4",X"00",X"BB",X"00",X"BB",X"C0",X"BC",X"C0",
		X"BB",X"BB",X"BB",X"BC",X"BC",X"BC",X"B4",X"BB",X"44",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"BC",X"C0",X"BB",X"C0",X"BB",X"4C",X"BC",X"4C",X"CB",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"0B",X"BB",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"00",X"44",X"00",X"B4",X"00",X"BB",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"CB",X"BC",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"C0",X"BC",X"C0",X"BC",X"C0",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"00",X"44",X"00",
		X"0B",X"BB",X"0B",X"BB",X"0B",X"BB",X"0C",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B4",X"00",X"B4",X"00",X"B4",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"BB",X"0B",X"BB",X"0C",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4C",X"00",X"44",X"00",X"B4",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4C",X"00",X"4C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"4C",X"0B",X"4C",X"0C",X"4B",X"00",X"BB",X"00",X"BB",X"4C",X"BB",X"44",X"BB",
		X"F0",X"00",X"FF",X"00",X"CF",X"C0",X"FB",X"FC",X"BB",X"FF",X"CB",X"FF",X"BB",X"FC",X"C4",X"C0",
		X"B4",X"BB",X"B4",X"BB",X"B4",X"BB",X"BB",X"BB",X"CB",X"44",X"B4",X"44",X"4C",X"44",X"C0",X"C4",
		X"B4",X"44",X"44",X"44",X"44",X"44",X"44",X"CC",X"4C",X"00",X"C0",X"00",X"4C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"CF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"CF",X"F0",X"FF",X"CF",X"CC",X"CF",X"FF",X"CF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"0B",X"BB",X"0F",X"FB",X"0F",X"FB",X"0B",X"BB",
		X"00",X"00",X"4C",X"00",X"44",X"00",X"B4",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FF",X"00",
		X"0C",X"BC",X"BB",X"CC",X"B4",X"BC",X"B4",X"CB",X"44",X"0C",X"C4",X"00",X"0C",X"00",X"00",X"00",
		X"BB",X"00",X"BC",X"C0",X"CB",X"4C",X"BB",X"4C",X"CB",X"4C",X"0C",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"0B",X"BB",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"44",X"00",X"44",X"00",X"B4",X"00",X"BC",X"00",
		X"0B",X"BB",X"0B",X"BC",X"BC",X"BC",X"BB",X"BB",X"C4",X"CC",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"BC",X"00",X"B4",X"00",X"B4",X"C0",X"BC",X"C0",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"FB",X"00",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"44",X"00",X"44",X"00",
		X"0B",X"BB",X"0B",X"BB",X"0B",X"BB",X"0C",X"BC",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B4",X"00",X"BC",X"00",X"BC",X"00",X"B4",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"44",X"00",X"44",X"00",X"4C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"4C",X"00",X"44",X"00",X"4C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"4C",X"00",X"4C",X"00",X"4B",X"00",X"BB",X"00",X"BB",X"4C",X"BB",X"B4",X"BB",
		X"00",X"00",X"FF",X"00",X"CF",X"C0",X"FF",X"4C",X"BB",X"FC",X"C4",X"FC",X"B4",X"FC",X"C4",X"C0",
		X"B4",X"BB",X"B4",X"BB",X"BB",X"BB",X"CB",X"B4",X"04",X"44",X"4C",X"44",X"C0",X"C4",X"00",X"0C",
		X"44",X"00",X"44",X"4C",X"4C",X"4C",X"C0",X"4C",X"00",X"C0",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"33",X"03",X"33",X"0F",X"33",X"03",X"33",X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"BB",
		X"C0",X"00",X"2C",X"00",X"2C",X"00",X"32",X"00",X"F2",X"00",X"F2",X"00",X"F3",X"C0",X"33",X"2C",
		X"3F",X"BB",X"CF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"F3",X"22",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"C0",X"FB",X"C0",X"BB",X"00",X"CC",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"F3",X"03",X"F3",X"03",X"C3",X"33",X"BB",X"33",X"FB",
		X"2C",X"00",X"32",X"00",X"32",X"00",X"F3",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"F3",X"C0",
		X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"FF",X"00",X"FF",X"03",X"FF",X"33",X"FC",X"33",X"FB",
		X"22",X"00",X"32",X"00",X"33",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"CF",X"C0",X"BF",X"C0",
		X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"BB",X"FF",X"CB",X"FF",X"0C",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"33",X"03",X"33",X"03",X"33",X"F3",X"33",X"C3",X"F3",X"F3",X"F3",X"BB",X"F3",X"BB",X"33",
		X"C0",X"00",X"2C",X"00",X"2C",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"33",X"C2",X"33",X"32",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"0F",X"FF",X"BB",X"FF",X"BB",X"FF",X"CC",X"CC",
		X"33",X"2C",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"C0",X"F2",X"00",X"BC",X"00",X"BB",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"F3",X"03",X"C3",X"03",X"F3",X"33",X"BB",X"33",X"FB",
		X"2C",X"00",X"32",X"00",X"32",X"00",X"F3",X"00",X"CF",X"00",X"CF",X"00",X"FF",X"C0",X"F3",X"C0",
		X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",
		X"22",X"00",X"33",X"00",X"33",X"00",X"FF",X"C0",X"CF",X"C0",X"FB",X"C0",X"BC",X"C2",X"FB",X"22",
		X"33",X"33",X"C3",X"3F",X"33",X"3F",X"33",X"FF",X"33",X"FF",X"C3",X"FB",X"0C",X"BB",X"00",X"BB",
		X"FF",X"2C",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"BC",X"FF",X"BC",X"FB",X"C0",X"CC",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"F3",X"03",X"C3",X"03",X"FB",X"33",X"BC",X"33",X"FB",
		X"2C",X"00",X"32",X"00",X"32",X"00",X"F3",X"00",X"CF",X"00",X"CF",X"00",X"FF",X"C0",X"F3",X"C0",
		X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"2C",X"00",X"2C",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"33",X"C0",X"33",X"2C",
		X"33",X"33",X"C3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"C3",X"33",X"BB",X"33",X"BB",X"C3",
		X"33",X"22",X"33",X"C2",X"33",X"CC",X"33",X"C0",X"33",X"C0",X"32",X"BC",X"22",X"C0",X"2C",X"00",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",
		X"22",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"32",X"C0",X"33",X"C0",X"33",X"C0",X"33",X"C0",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"C2",
		X"33",X"2C",X"33",X"22",X"33",X"C2",X"32",X"0C",X"32",X"00",X"22",X"00",X"22",X"C0",X"CB",X"C0",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"F3",X"03",X"F3",X"03",X"C3",X"33",X"BB",X"33",X"FB",
		X"2C",X"00",X"32",X"00",X"32",X"00",X"F3",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"F3",X"C0",
		X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"33",X"03",X"33",X"0F",X"33",X"03",X"33",X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"BB",
		X"C0",X"00",X"2C",X"00",X"2C",X"00",X"32",X"00",X"F2",X"00",X"F2",X"00",X"F3",X"C0",X"33",X"2C",
		X"3F",X"BB",X"CF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"F3",X"22",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"C0",X"FB",X"C0",X"BB",X"00",X"CC",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"F3",X"03",X"F3",X"03",X"C3",X"33",X"BB",X"33",X"FB",
		X"2C",X"00",X"32",X"00",X"32",X"00",X"F3",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"F3",X"C0",
		X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"C3",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"FF",X"00",X"FF",X"03",X"FF",X"33",X"FC",X"33",X"FB",
		X"22",X"00",X"32",X"00",X"33",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"CF",X"C0",X"BF",X"C0",
		X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"BB",X"FF",X"CB",X"FF",X"0C",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"66",X"00",X"F6",X"00",X"66",X"00",X"FF",X"00",X"FF",X"06",X"FF",X"66",X"FC",X"66",X"FB",
		X"55",X"00",X"65",X"00",X"66",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"CF",X"C0",X"BF",X"C0",
		X"66",X"FF",X"66",X"FF",X"66",X"FF",X"66",X"FF",X"66",X"FF",X"BB",X"FF",X"CB",X"FF",X"0C",X"CC",
		X"FF",X"6C",X"FF",X"56",X"FF",X"C5",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",X"EE",X"DD",X"FF",X"EE",
		X"11",X"11",X"11",X"1F",X"11",X"1F",X"11",X"FF",X"11",X"FF",X"11",X"FF",X"11",X"FF",X"DD",X"FF",
		X"11",X"11",X"11",X"11",X"1F",X"11",X"1F",X"11",X"FF",X"D1",X"FF",X"DD",X"FE",X"ED",X"FF",X"ED",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FE",X"EE",X"FF",X"EE",X"EE",X"FE",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"D1",X"11",X"D1",X"11",X"DD",X"11",X"ED",X"11",X"FE",X"11",X"FF",X"D1",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"EE",X"EF",X"FE",X"EE",X"FE",X"FF",X"FF",X"FF",X"EE",X"EF",X"FF",X"DE",X"FF",X"FD",X"FF",
		X"ED",X"FF",X"EE",X"DF",X"FF",X"FD",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"EE",X"EF",X"FE",X"DE",X"EF",X"ED",X"EF",X"EE",X"EE",X"FF",X"FE",X"EF",X"FF",X"EE",X"FF",X"FE",
		X"EF",X"FF",X"FF",X"EF",X"FF",X"FF",X"EF",X"FF",X"DE",X"FF",X"DD",X"EE",X"EE",X"DD",X"FE",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"DE",X"FF",X"DE",X"FF",X"EF",
		X"FF",X"D1",X"FF",X"ED",X"FD",X"EE",X"DE",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"FE",X"EE",X"FF",
		X"FD",X"FF",X"DE",X"FF",X"DF",X"FE",X"FF",X"EF",X"FF",X"FF",X"FF",X"FE",X"EE",X"FF",X"DD",X"EE",
		X"FF",X"EE",X"EF",X"FF",X"FF",X"EE",X"FF",X"EE",X"FE",X"EE",X"FF",X"FF",X"FE",X"FF",X"FF",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"D1",X"11",X"DD",X"11",X"EE",X"DD",X"FE",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",
		X"FF",X"EF",X"FE",X"EE",X"EF",X"EE",X"EF",X"FE",X"FF",X"FF",X"EF",X"FF",X"DD",X"FF",X"FE",X"DF",
		X"FD",X"11",X"FF",X"DD",X"FF",X"EF",X"EF",X"FF",X"EE",X"FF",X"EE",X"FF",X"FE",X"EF",X"FF",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"DD",X"DD",X"EE",X"EE",X"FE",X"FF",X"EE",X"DF",X"FE",X"ED",X"FF",X"FE",X"EF",
		X"D1",X"11",X"DF",X"11",X"ED",X"DD",X"EF",X"FF",X"EE",X"FE",X"DE",X"EF",X"FD",X"EF",X"EF",X"EE",
		X"11",X"1F",X"11",X"EF",X"DF",X"FF",X"FF",X"FF",X"FD",X"FE",X"DE",X"FE",X"EF",X"EF",X"FF",X"FF",
		X"11",X"11",X"DD",X"11",X"EE",X"11",X"EF",X"D1",X"EE",X"ED",X"FE",X"EE",X"FD",X"EF",X"FF",X"EE",
		X"11",X"FF",X"11",X"FF",X"1F",X"EF",X"FF",X"FF",X"FF",X"EF",X"FE",X"EF",X"EF",X"EE",X"FF",X"FE",
		X"11",X"11",X"D1",X"11",X"ED",X"11",X"FF",X"D1",X"EF",X"ED",X"EE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"FE",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"EF",X"EF",X"FF",X"EE",
		X"11",X"11",X"11",X"11",X"D1",X"1F",X"ED",X"FF",X"FE",X"FF",X"FF",X"EF",X"FF",X"FE",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"1F",X"11",X"FF",X"11",X"FF",X"DF",X"FF",X"EE",X"FF",X"FF",X"FF",
		X"11",X"11",X"D1",X"11",X"ED",X"11",X"FE",X"11",X"FF",X"11",X"FF",X"DD",X"EE",X"EE",X"FE",X"FF",
		X"11",X"11",X"FE",X"11",X"FF",X"D1",X"FF",X"ED",X"DF",X"FE",X"ED",X"FF",X"FF",X"DF",X"FF",X"ED",
		X"11",X"11",X"11",X"D1",X"FF",X"ED",X"FF",X"FE",X"FF",X"FF",X"DD",X"FF",X"FE",X"FF",X"FF",X"DD",
		X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"11",X"FF",X"DD",X"EF",X"FE",X"EE",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"FE",X"11",X"FF",X"D1",X"FF",X"ED",X"DD",X"EE",X"FE",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"EE",X"FF",X"EF",X"FF",X"EE",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"EE",X"D1",X"FF",X"FD",X"FF",X"FF",X"FF",X"EF",X"EE",X"EF",
		X"11",X"1F",X"11",X"FE",X"11",X"FF",X"11",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FE",X"FF",
		X"11",X"11",X"11",X"11",X"D1",X"11",X"DD",X"1E",X"EE",X"ED",X"DE",X"DF",X"FD",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"11",X"FF",
		X"11",X"11",X"11",X"11",X"EF",X"FF",X"FE",X"EE",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"11",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FF",X"FF",X"EE",X"FE",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"1E",X"FF",
		X"EE",X"DD",X"FF",X"ED",X"FF",X"DE",X"FD",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FE",X"FF",X"EF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"ED",X"11",X"FE",X"11",X"FE",X"DD",X"FF",X"EE",X"FF",X"ED",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"11",X"FF",X"EF",X"FF",X"FE",X"FF",X"EF",X"EE",
		X"FF",X"DE",X"FF",X"EF",X"FE",X"FF",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FD",X"FF",X"DE",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"D1",X"EF",X"EF",X"FF",X"FE",X"FF",X"EF",X"FF",
		X"1E",X"11",X"FF",X"11",X"FF",X"D1",X"FF",X"DD",X"FF",X"ED",X"FF",X"EE",X"FF",X"FE",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",
		X"DD",X"FF",X"FE",X"FF",X"FF",X"DF",X"FF",X"DF",X"FF",X"ED",X"FF",X"EE",X"FF",X"FE",X"FF",X"FF",
		X"11",X"12",X"11",X"2F",X"11",X"FF",X"11",X"FF",X"12",X"FF",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"21",X"11",X"F2",X"11",X"FF",X"11",X"FF",X"11",X"FF",X"21",X"FF",X"F2",
		X"22",X"22",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",
		X"22",X"22",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",
		X"22",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"22",X"22",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",
		X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",
		X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",
		X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",
		X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"22",X"22",
		X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"EE",X"E2",X"22",X"22",
		X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EF",X"22",X"22",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"11",X"11",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"A5",X"55",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"AA",X"AA",
		X"A5",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"55",X"AA",X"55",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"22",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"12",X"22",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"22",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"21",X"11",X"22",X"11",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"12",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"21",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"12",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"11",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"21",X"22",X"21",X"22",X"11",X"22",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",
		X"00",X"BA",X"00",X"BA",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"F3",X"03",X"F3",X"03",X"F3",X"33",X"BB",X"33",X"FB",
		X"2C",X"00",X"32",X"00",X"32",X"00",X"F3",X"00",X"FF",X"00",X"CF",X"00",X"FF",X"C0",X"F3",X"C0",
		X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"03",X"FF",X"0B",X"FF",X"BB",X"CC",
		X"FF",X"3C",X"FF",X"23",X"FF",X"C2",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"BB",X"00",X"BB",X"C0",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",
		X"2C",X"00",X"22",X"00",X"22",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"33",X"C0",X"33",X"C0",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"3C",
		X"33",X"3C",X"33",X"23",X"33",X"C2",X"33",X"CC",X"32",X"C0",X"32",X"BC",X"22",X"C0",X"2C",X"00",
		X"00",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"2C",X"00",X"2C",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"33",X"C0",X"33",X"2C",
		X"33",X"33",X"C3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"C3",X"33",X"BB",X"33",X"BB",X"C3",
		X"33",X"22",X"33",X"C2",X"33",X"CC",X"33",X"C0",X"33",X"C0",X"32",X"BC",X"22",X"C0",X"2C",X"00",
		X"00",X"33",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",
		X"22",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"32",X"C0",X"33",X"C0",X"33",X"C0",X"33",X"C0",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"C2",
		X"33",X"2C",X"33",X"22",X"33",X"C2",X"32",X"0C",X"32",X"00",X"22",X"00",X"22",X"C0",X"CB",X"C0",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"4F",X"44",X"EF",X"44",X"F1",X"44",X"11",
		X"F1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"11",X"44",X"11",X"4F",X"11",X"EF",X"11",X"F1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"4F",X"44",X"EF",X"44",X"F1",X"44",X"11",X"44",X"11",X"44",X"11",X"4F",X"11",X"EF",X"11",
		X"11",X"44",X"11",X"F4",X"11",X"FE",X"11",X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"44",X"FE",X"44",X"1F",X"44",X"11",X"44",X"11",X"44",
		X"FE",X"44",X"1F",X"44",X"11",X"44",X"11",X"44",X"11",X"44",X"11",X"F4",X"11",X"FE",X"11",X"1F",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"44",X"4F",X"44",X"EF",X"44",X"FE",X"44",X"FE",X"44",X"EE",X"44",X"EE",X"4F",X"EE",X"EF",X"EE",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"44",X"FE",X"44",X"EF",X"44",X"EF",X"44",X"EE",X"44",
		X"FE",X"EE",X"FE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"EE",X"44",X"EE",X"F4",X"EE",X"FE",X"EE",X"EF",X"FF",X"FF",X"DD",X"DF",X"DD",X"DF",X"FF",X"FF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"E4",X"EE",X"F4",X"EE",X"EF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"DF",X"DD",X"DF",X"DD",X"DF",X"DD",X"DF",X"FF",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"11",X"44",X"11",X"4F",X"11",X"EF",X"11",X"F1",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"44",X"1F",X"44",X"11",X"44",X"11",X"44",X"11",X"44",X"11",X"F4",X"FF",X"FE",X"FF",X"FF",
		X"42",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"22",X"44",X"22",X"44",X"22",X"44",X"22",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"44",X"42",X"44",X"22",X"44",X"22",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"44",X"44",X"44",X"44",X"24",X"44",
		X"44",X"22",X"44",X"22",X"42",X"22",X"42",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"24",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"E1",X"11",X"EE",X"11",X"FE",X"11",X"FF",X"F1",X"FE",X"FF",X"FF",X"EF",X"FF",X"EF",X"EE",X"EF",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"F4",X"12",X"12",X"12",X"22",X"22",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"44",X"22",X"14",X"FF",X"22",X"22",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"2F",X"FF",X"FF",X"2F",X"22",X"24",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"F4",X"FF",X"FF",X"22",X"2F",X"24",X"24",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"4F",X"2F",X"FF",X"2F",X"F2",X"24",X"42",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"F4",X"F2",X"F2",X"FF",X"F2",X"42",X"42",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"FF",X"F2",X"4F",X"F2",X"4F",X"42",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",X"42",X"42",X"44",X"44",
		X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",
		X"FF",X"FF",X"FF",X"FF",X"22",X"22",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"22",X"22",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AC",X"CC",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"8F",X"FC",X"CF",X"FF",X"8F",
		X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"AA",X"AA",X"8C",X"CC",
		X"FC",X"8F",X"FC",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"F8",X"FF",X"FC",X"CF",X"FC",X"F8",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"F8",X"CF",X"CC",X"C8",X"88",
		X"FC",X"CC",X"8C",X"FF",X"C8",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"C8",X"F8",X"CF",X"8C",X"C8",X"C8",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"F8",X"88",X"CF",X"CF",X"FF",X"CF",
		X"AA",X"AA",X"CC",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"CF",X"F8",X"CF",X"FC",
		X"CF",X"CF",X"8F",X"F8",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"CF",X"FC",X"CF",X"FC",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"AA",X"CC",X"CA",X"88",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"8A",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"8A",X"AA",X"AA",X"CC",X"CC",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
