library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd_prg is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd_prg is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"01",X"80",X"40",X"02",X"B0",X"82",X"F0",X"01",X"B0",X"84",X"A0",X"01",X"50",
		X"85",X"F0",X"10",X"00",X"95",X"F0",X"18",X"80",X"AE",X"70",X"03",X"A0",X"B2",X"10",X"08",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"AA",X"98",X"26",X"10",X"80",X"28",X"8B",X"BA",X"10",X"0A",X"8B",X"AA",X"22",X"71",X"19",X"10",
		X"10",X"AC",X"B1",X"00",X"CB",X"E9",X"25",X"31",X"80",X"01",X"0A",X"C8",X"00",X"AD",X"DA",X"04",
		X"42",X"18",X"00",X"08",X"D9",X"88",X"9E",X"A8",X"17",X"21",X"98",X"11",X"0B",X"C8",X"AB",X"E9",
		X"14",X"71",X"89",X"81",X"19",X"B9",X"9B",X"E9",X"25",X"51",X"99",X"82",X"0B",X"BC",X"AB",X"25",
		X"53",X"09",X"98",X"0A",X"CB",X"AD",X"05",X"53",X"8A",X"A0",X"19",X"CA",X"BB",X"37",X"61",X"99",
		X"A1",X"09",X"AB",X"C2",X"73",X"08",X"AA",X"88",X"89",X"CA",X"47",X"20",X"AA",X"89",X"98",X"AA",
		X"37",X"78",X"99",X"89",X"80",X"A8",X"46",X"19",X"A9",X"89",X"88",X"A2",X"73",X"9A",X"99",X"A1",
		X"2E",X"06",X"29",X"99",X"99",X"11",X"D0",X"71",X"99",X"89",X"81",X"0C",X"17",X"0A",X"88",X"98",
		X"49",X"B3",X"69",X"A0",X"0B",X"14",X"C8",X"50",X"A8",X"0A",X"84",X"8B",X"62",X"C9",X"18",X"A3",
		X"1E",X"25",X"AA",X"10",X"B2",X"3E",X"05",X"8C",X"10",X"A1",X"2B",X"87",X"8B",X"11",X"B0",X"3C",
		X"06",X"8B",X"10",X"A1",X"1C",X"35",X"C9",X"39",X"A3",X"AB",X"72",X"D0",X"2A",X"03",X"F0",X"58",
		X"C2",X"8A",X"48",X"D4",X"2D",X"03",X"C0",X"3E",X"05",X"9B",X"49",X"96",X"CB",X"51",X"C3",X"A9",
		X"7B",X"C4",X"1B",X"3C",X"96",X"8D",X"11",X"12",X"DB",X"51",X"B8",X"02",X"00",X"F0",X"48",X"B0",
		X"18",X"5B",X"B6",X"8B",X"03",X"A3",X"9F",X"31",X"B8",X"4A",X"11",X"E1",X"2A",X"81",X"09",X"4D",
		X"03",X"A9",X"84",X"80",X"9B",X"58",X"A8",X"59",X"81",X"D2",X"1A",X"A7",X"A0",X"0A",X"20",X"9C",
		X"7A",X"82",X"B2",X"92",X"D5",X"A8",X"3C",X"19",X"2B",X"31",X"C5",X"C2",X"A2",X"90",X"2C",X"5C",
		X"3C",X"3A",X"3A",X"83",X"D4",X"C2",X"93",X"B1",X"1B",X"3B",X"3C",X"2A",X"31",X"C1",X"A6",X"C2",
		X"A3",X"89",X"89",X"4A",X"81",X"4C",X"1B",X"86",X"98",X"3C",X"2C",X"01",X"39",X"9C",X"3B",X"26",
		X"A1",X"D1",X"95",X"88",X"A8",X"11",X"82",X"A0",X"E1",X"A7",X"91",X"B2",X"A8",X"97",X"91",X"D3",
		X"90",X"87",X"C0",X"A1",X"88",X"41",X"BA",X"18",X"2C",X"7B",X"3D",X"39",X"09",X"7D",X"18",X"82",
		X"B5",X"88",X"D4",X"A2",X"C5",X"B1",X"99",X"2C",X"7A",X"1E",X"4A",X"3C",X"5B",X"91",X"A4",X"C2",
		X"2A",X"A2",X"01",X"C2",X"3B",X"B1",X"22",X"F4",X"B3",X"D3",X"A2",X"D5",X"B1",X"A2",X"08",X"A7",
		X"9B",X"3A",X"4E",X"49",X"2D",X"4B",X"3E",X"5A",X"2C",X"20",X"99",X"6B",X"80",X"04",X"C9",X"59",
		X"99",X"13",X"C8",X"30",X"C2",X"A4",X"D1",X"28",X"B3",X"92",X"F0",X"30",X"C1",X"01",X"D2",X"01",
		X"C2",X"81",X"BA",X"78",X"A0",X"12",X"C8",X"15",X"BA",X"6B",X"1D",X"33",X"9C",X"28",X"1E",X"15",
		X"AA",X"01",X"2D",X"85",X"89",X"C4",X"88",X"B0",X"7A",X"9A",X"51",X"D0",X"06",X"D8",X"06",X"BB",
		X"21",X"6D",X"94",X"0D",X"84",X"3C",X"C3",X"5B",X"D2",X"25",X"DA",X"34",X"CB",X"48",X"5D",X"82",
		X"3F",X"85",X"B5",X"D1",X"28",X"F2",X"5D",X"4D",X"5A",X"0C",X"40",X"C1",X"10",X"A0",X"A7",X"B8",
		X"97",X"AA",X"05",X"AA",X"04",X"B5",X"D2",X"81",X"98",X"1C",X"7A",X"98",X"39",X"B2",X"0A",X"7D",
		X"4A",X"2B",X"3A",X"12",X"9D",X"22",X"9C",X"13",X"D5",X"B0",X"02",X"B8",X"12",X"AE",X"7C",X"01",
		X"19",X"A2",X"09",X"95",X"B3",X"A8",X"81",X"3F",X"A7",X"99",X"11",X"A8",X"3B",X"A0",X"7E",X"32",
		X"8D",X"15",X"D0",X"2A",X"5D",X"48",X"A8",X"21",X"D1",X"19",X"00",X"B3",X"80",X"A2",X"2C",X"A5",
		X"9D",X"7B",X"02",X"90",X"B7",X"A8",X"01",X"B2",X"2F",X"39",X"09",X"12",X"F2",X"09",X"84",X"D3",
		X"88",X"91",X"3E",X"10",X"89",X"10",X"2E",X"12",X"C1",X"01",X"A9",X"5A",X"08",X"08",X"4C",X"95",
		X"A0",X"82",X"8C",X"38",X"90",X"83",X"9F",X"5A",X"93",X"90",X"A2",X"0A",X"03",X"AA",X"23",X"F2",
		X"0B",X"20",X"8A",X"25",X"E0",X"29",X"80",X"97",X"D2",X"1B",X"10",X"88",X"83",X"C8",X"5A",X"92",
		X"83",X"F1",X"3E",X"12",X"A0",X"82",X"B0",X"3B",X"02",X"C1",X"2A",X"93",X"9A",X"4A",X"18",X"81",
		X"99",X"49",X"A3",X"A1",X"99",X"2B",X"7F",X"32",X"E0",X"28",X"A2",X"90",X"09",X"18",X"1A",X"89",
		X"7B",X"B7",X"A1",X"1B",X"49",X"81",X"A2",X"90",X"00",X"A1",X"80",X"0A",X"42",X"F6",X"AA",X"4A",
		X"00",X"91",X"08",X"92",X"A1",X"80",X"91",X"93",X"D3",X"B9",X"7F",X"41",X"F2",X"0A",X"10",X"88",
		X"00",X"91",X"09",X"81",X"88",X"82",X"A8",X"6B",X"97",X"B8",X"39",X"90",X"2A",X"00",X"09",X"18",
		X"00",X"B3",X"91",X"99",X"7B",X"81",X"87",X"F4",X"0E",X"38",X"A1",X"08",X"88",X"29",X"92",X"89",
		X"10",X"99",X"38",X"C4",X"90",X"89",X"16",X"F1",X"3E",X"11",X"A1",X"09",X"18",X"80",X"80",X"80",
		X"E7",X"F0",X"79",X"F3",X"1B",X"18",X"83",X"AA",X"39",X"82",X"93",X"F0",X"5B",X"93",X"91",X"9A",
		X"48",X"98",X"7A",X"D5",X"8A",X"18",X"10",X"B1",X"2A",X"97",X"AB",X"68",X"A1",X"81",X"8A",X"49",
		X"A3",X"4F",X"03",X"B0",X"80",X"2C",X"11",X"B5",X"8E",X"38",X"80",X"A3",X"99",X"2A",X"59",X"F4",
		X"89",X"1A",X"28",X"A3",X"82",X"F0",X"28",X"8A",X"22",X"D1",X"4E",X"11",X"91",X"C3",X"0B",X"22",
		X"E1",X"00",X"0C",X"38",X"92",X"9B",X"40",X"8A",X"97",X"A8",X"4D",X"28",X"00",X"B4",X"91",X"9C",
		X"59",X"1A",X"01",X"82",X"E2",X"92",X"99",X"3A",X"88",X"12",X"D1",X"01",X"0E",X"29",X"3B",X"82",
		X"2C",X"81",X"82",X"E2",X"02",X"E1",X"93",X"99",X"11",X"98",X"93",X"A0",X"1B",X"3A",X"4B",X"95",
		X"0D",X"95",X"88",X"A2",X"2A",X"8A",X"22",X"AA",X"24",X"B9",X"03",X"B0",X"91",X"7A",X"92",X"89",
		X"D4",X"19",X"A0",X"49",X"8C",X"22",X"8C",X"22",X"8B",X"81",X"08",X"A1",X"27",X"BC",X"34",X"CA",
		X"15",X"98",X"90",X"20",X"BD",X"41",X"8B",X"13",X"AB",X"28",X"29",X"18",X"2B",X"A1",X"5E",X"08",
		X"78",X"A9",X"14",X"BA",X"38",X"5D",X"01",X"80",X"A1",X"03",X"BE",X"58",X"8D",X"59",X"1B",X"10",
		X"2B",X"01",X"0B",X"A1",X"79",X"00",X"A9",X"A5",X"7C",X"2B",X"2B",X"17",X"8A",X"90",X"1A",X"70",
		X"B9",X"03",X"B3",X"6E",X"09",X"4A",X"21",X"E0",X"02",X"B2",X"2C",X"88",X"3A",X"05",X"B9",X"85",
		X"A8",X"5C",X"1A",X"39",X"83",X"9C",X"85",X"99",X"39",X"B1",X"38",X"AC",X"7B",X"19",X"6B",X"02",
		X"C2",X"80",X"A0",X"7C",X"A4",X"1B",X"97",X"C0",X"84",X"A9",X"23",X"F0",X"38",X"E5",X"A1",X"A0",
		X"2A",X"5B",X"B7",X"8B",X"06",X"AB",X"05",X"AA",X"6D",X"20",X"8A",X"25",X"D9",X"58",X"A8",X"30",
		X"E3",X"89",X"96",X"8D",X"31",X"AB",X"44",X"D9",X"5A",X"94",X"8D",X"30",X"0D",X"5B",X"A6",X"9A",
		X"32",X"F3",X"8A",X"01",X"7D",X"95",X"AB",X"69",X"D5",X"98",X"97",X"AD",X"42",X"CA",X"50",X"D1",
		X"39",X"E5",X"1D",X"38",X"9B",X"7A",X"B4",X"3D",X"A5",X"2D",X"95",X"A9",X"5D",X"5D",X"29",X"69",
		X"D2",X"5D",X"B5",X"0C",X"85",X"8D",X"59",X"89",X"39",X"A7",X"D3",X"81",X"F5",X"3D",X"A5",X"8D",
		X"41",X"D1",X"18",X"B4",X"2F",X"12",X"0E",X"5A",X"80",X"08",X"97",X"BA",X"33",X"DA",X"5A",X"0A",
		X"7B",X"B6",X"8A",X"94",X"0B",X"4D",X"4A",X"3E",X"42",X"D8",X"23",X"F3",X"1C",X"81",X"3E",X"13",
		X"C0",X"02",X"D4",X"9A",X"03",X"8E",X"59",X"A8",X"20",X"C7",X"B9",X"84",X"A9",X"59",X"A1",X"19",
		X"A7",X"A9",X"83",X"9A",X"7B",X"08",X"2A",X"87",X"B0",X"92",X"98",X"5C",X"00",X"1A",X"03",X"B1",
		X"A2",X"A1",X"4E",X"28",X"0A",X"11",X"A2",X"89",X"95",X"9B",X"30",X"8C",X"59",X"93",X"99",X"96",
		X"A9",X"38",X"99",X"4B",X"84",X"8B",X"05",X"A9",X"11",X"A0",X"3D",X"02",X"0A",X"A4",X"88",X"08",
		X"01",X"9D",X"31",X"8D",X"12",X"A1",X"80",X"A4",X"0C",X"18",X"3B",X"8B",X"63",X"CC",X"41",X"C1",
		X"81",X"91",X"80",X"91",X"91",X"80",X"00",X"81",X"80",X"81",X"90",X"80",X"80",X"81",X"80",X"08",
		X"A9",X"2A",X"57",X"CD",X"5A",X"94",X"92",X"2F",X"00",X"B2",X"28",X"4C",X"93",X"D0",X"39",X"21",
		X"F2",X"AA",X"50",X"83",X"F0",X"1B",X"13",X"A4",X"8E",X"29",X"A3",X"00",X"6A",X"B3",X"BB",X"58",
		X"16",X"AA",X"2B",X"A2",X"83",X"78",X"A0",X"A9",X"98",X"25",X"40",X"B8",X"AC",X"98",X"15",X"51",
		X"99",X"9D",X"89",X"93",X"43",X"5A",X"88",X"DA",X"89",X"03",X"44",X"3B",X"88",X"EA",X"90",X"91",
		X"62",X"20",X"A0",X"BD",X"A8",X"88",X"36",X"22",X"89",X"8C",X"BA",X"A0",X"12",X"74",X"00",X"0A",
		X"AB",X"C9",X"91",X"03",X"72",X"00",X"8B",X"AB",X"BA",X"82",X"25",X"72",X"01",X"0B",X"BB",X"CA",
		X"91",X"22",X"65",X"18",X"09",X"CA",X"B9",X"98",X"24",X"35",X"30",X"A9",X"AD",X"BA",X"99",X"14",
		X"34",X"35",X"89",X"9A",X"CB",X"A8",X"90",X"33",X"36",X"48",X"90",X"9A",X"C9",X"89",X"14",X"32",
		X"46",X"89",X"89",X"BC",X"B9",X"98",X"13",X"33",X"73",X"88",X"89",X"CB",X"A9",X"B1",X"33",X"46",
		X"40",X"08",X"AB",X"BC",X"C9",X"81",X"22",X"44",X"31",X"88",X"BC",X"BC",X"A9",X"91",X"42",X"34",
		X"41",X"88",X"9C",X"C8",X"BB",X"08",X"13",X"43",X"43",X"30",X"9A",X"CC",X"CA",X"A8",X"09",X"25",
		X"21",X"44",X"18",X"08",X"BD",X"99",X"BA",X"00",X"04",X"42",X"24",X"28",X"99",X"BD",X"B9",X"9A",
		X"02",X"0A",X"43",X"19",X"43",X"9B",X"89",X"FB",X"18",X"D2",X"2A",X"14",X"01",X"42",X"12",X"18",
		X"9C",X"BC",X"B9",X"BA",X"89",X"B9",X"9A",X"A2",X"51",X"55",X"34",X"22",X"41",X"11",X"19",X"9C",
		X"CB",X"CB",X"AA",X"99",X"01",X"11",X"12",X"1B",X"98",X"9A",X"82",X"26",X"23",X"42",X"20",X"1A",
		X"CA",X"CB",X"B1",X"13",X"53",X"43",X"10",X"9A",X"BB",X"BA",X"92",X"23",X"34",X"11",X"9A",X"CC",
		X"BB",X"AA",X"03",X"31",X"43",X"18",X"18",X"9A",X"9A",X"8A",X"98",X"08",X"08",X"08",X"19",X"00",
		X"10",X"08",X"18",X"8A",X"08",X"89",X"08",X"08",X"10",X"80",X"08",X"8A",X"88",X"00",X"11",X"11",
		X"08",X"09",X"9A",X"89",X"00",X"00",X"30",X"20",X"18",X"0A",X"8A",X"8A",X"08",X"02",X"10",X"30",
		X"19",X"89",X"9A",X"89",X"80",X"00",X"11",X"18",X"08",X"09",X"88",X"09",X"08",X"89",X"18",X"08",
		X"98",X"91",X"91",X"88",X"10",X"08",X"80",X"90",X"00",X"01",X"01",X"00",X"B8",X"A9",X"90",X"A0",
		X"89",X"80",X"81",X"72",X"48",X"8D",X"0C",X"88",X"29",X"50",X"08",X"0C",X"89",X"88",X"40",X"22",
		X"3D",X"1B",X"B9",X"1B",X"10",X"E9",X"99",X"76",X"12",X"0B",X"AB",X"C9",X"20",X"34",X"29",X"1C",
		X"BB",X"8B",X"44",X"41",X"29",X"CC",X"BC",X"8A",X"16",X"70",X"38",X"AB",X"9C",X"80",X"11",X"51",
		X"88",X"8D",X"98",X"81",X"52",X"81",X"AD",X"AA",X"B1",X"27",X"34",X"09",X"B9",X"E8",X"81",X"14",
		X"10",X"98",X"C9",X"98",X"32",X"31",X"0F",X"BB",X"99",X"73",X"31",X"1D",X"8B",X"AA",X"20",X"43",
		X"28",X"8B",X"E9",X"00",X"14",X"89",X"BC",X"B4",X"23",X"72",X"A9",X"9C",X"A1",X"81",X"25",X"81",
		X"9A",X"B3",X"C0",X"21",X"E0",X"BB",X"71",X"22",X"1D",X"0A",X"A9",X"29",X"34",X"19",X"19",X"D0",
		X"88",X"92",X"D9",X"C4",X"22",X"62",X"C8",X"9A",X"B2",X"82",X"26",X"90",X"89",X"A0",X"99",X"09",
		X"EA",X"70",X"23",X"2E",X"0A",X"9A",X"39",X"23",X"2A",X"28",X"E8",X"89",X"B3",X"DA",X"71",X"03",
		X"2E",X"09",X"A9",X"39",X"14",X"09",X"29",X"D0",X"8A",X"91",X"C5",X"21",X"15",X"C9",X"89",X"B3",
		X"01",X"23",X"98",X"0D",X"98",X"9D",X"0A",X"71",X"21",X"2D",X"8A",X"A8",X"11",X"16",X"88",X"80",
		X"C8",X"8A",X"8A",X"61",X"23",X"4F",X"09",X"8A",X"20",X"02",X"00",X"90",X"E0",X"89",X"A9",X"70",
		X"21",X"3F",X"0A",X"09",X"28",X"13",X"90",X"A0",X"E1",X"99",X"98",X"70",X"20",X"0C",X"0B",X"93",
		X"82",X"06",X"A0",X"9A",X"89",X"9C",X"17",X"01",X"30",X"F0",X"A8",X"11",X"82",X"3C",X"08",X"AA",
		X"1A",X"B0",X"71",X"23",X"8F",X"89",X"93",X"10",X"23",X"E8",X"0B",X"81",X"AB",X"47",X"82",X"1E",
		X"80",X"A8",X"40",X"83",X"A9",X"88",X"C1",X"1C",X"87",X"80",X"29",X"B0",X"9C",X"51",X"92",X"0A",
		X"A1",X"B8",X"1A",X"B7",X"48",X"2B",X"B8",X"0C",X"53",X"A1",X"0A",X"B2",X"BB",X"3D",X"70",X"10",
		X"1D",X"A1",X"92",X"21",X"88",X"0F",X"00",X"98",X"96",X"93",X"01",X"E9",X"09",X"31",X"00",X"0A",
		X"D2",X"99",X"8A",X"71",X"10",X"C8",X"90",X"95",X"2A",X"3C",X"A1",X"89",X"B1",X"70",X"10",X"BA",
		X"09",X"87",X"19",X"1B",X"B3",X"8C",X"96",X"10",X"28",X"F8",X"19",X"22",X"A1",X"8B",X"B3",X"AD",
		X"54",X"91",X"1F",X"93",X"A1",X"39",X"A1",X"AB",X"38",X"E7",X"09",X"18",X"D0",X"29",X"24",X"C9",
		X"19",X"80",X"93",X"48",X"A2",X"EA",X"40",X"02",X"AB",X"00",X"A8",X"87",X"29",X"0D",X"81",X"01",
		X"28",X"C8",X"8A",X"09",X"73",X"C1",X"9A",X"11",X"12",X"2F",X"90",X"90",X"87",X"0A",X"1C",X"82",
		X"01",X"29",X"E0",X"0A",X"03",X"49",X"80",X"F8",X"48",X"11",X"D9",X"29",X"A0",X"71",X"C3",X"D9",
		X"58",X"02",X"BC",X"10",X"B8",X"73",X"D4",X"DA",X"41",X"82",X"AE",X"11",X"B8",X"72",X"D4",X"D9",
		X"42",X"A3",X"BE",X"11",X"B2",X"79",X"B4",X"D8",X"52",X"C4",X"DA",X"29",X"97",X"3D",X"2A",X"C0",
		X"58",X"01",X"F9",X"4B",X"16",X"9C",X"3D",X"85",X"4C",X"3D",X"B1",X"09",X"73",X"D0",X"9B",X"54",
		X"B0",X"AC",X"02",X"B7",X"3D",X"09",X"B1",X"79",X"08",X"E0",X"1A",X"73",X"C8",X"AA",X"27",X"08",
		X"AE",X"10",X"91",X"78",X"C4",X"CA",X"54",X"D2",X"CA",X"10",X"97",X"3D",X"19",X"C4",X"4D",X"19",
		X"C1",X"08",X"44",X"B9",X"0B",X"15",X"99",X"0C",X"83",X"18",X"18",X"D2",X"5A",X"92",X"A9",X"30",
		X"C1",X"9C",X"21",X"07",X"2E",X"80",X"A2",X"3C",X"30",X"D1",X"29",X"99",X"C8",X"37",X"2A",X"B9",
		X"92",X"48",X"8C",X"93",X"39",X"3C",X"C8",X"81",X"58",X"B0",X"58",X"18",X"A8",X"0A",X"83",X"C9",
		X"3C",X"14",X"90",X"11",X"C2",X"88",X"A9",X"5A",X"82",X"01",X"B0",X"F4",X"8B",X"10",X"8A",X"72",
		X"08",X"B0",X"8D",X"10",X"90",X"05",X"8C",X"10",X"C1",X"59",X"3A",X"C2",X"89",X"12",X"D0",X"08",
		X"38",X"B4",X"AD",X"32",X"D2",X"18",X"91",X"81",X"B9",X"48",X"B9",X"83",X"A9",X"79",X"03",X"82",
		X"A0",X"AA",X"AA",X"86",X"8B",X"25",X"08",X"A0",X"B8",X"93",X"4D",X"4A",X"23",X"C2",X"0A",X"0A",
		X"0B",X"88",X"B4",X"B1",X"49",X"55",X"1D",X"20",X"B0",X"90",X"AD",X"94",X"88",X"68",X"09",X"03",
		X"B9",X"19",X"98",X"3A",X"1E",X"B7",X"8A",X"78",X"90",X"08",X"80",X"80",X"9E",X"28",X"B6",X"08",
		X"20",X"90",X"89",X"19",X"D2",X"9A",X"09",X"8A",X"44",X"23",X"99",X"6E",X"02",X"A1",X"A9",X"08",
		X"B1",X"5B",X"84",X"10",X"81",X"09",X"B1",X"3D",X"81",X"C8",X"90",X"6A",X"95",X"92",X"92",X"09",
		X"99",X"19",X"89",X"9A",X"D1",X"28",X"87",X"2A",X"30",X"91",X"92",X"9F",X"90",X"1C",X"02",X"C1",
		X"93",X"40",X"F3",X"1D",X"21",X"98",X"91",X"88",X"91",X"1C",X"12",X"B9",X"4B",X"40",X"B3",X"1E",
		X"28",X"92",X"98",X"20",X"D5",X"9B",X"49",X"92",X"99",X"29",X"94",X"99",X"4B",X"01",X"82",X"A8",
		X"1B",X"10",X"2A",X"2A",X"F2",X"80",X"5A",X"91",X"B4",X"29",X"A8",X"D2",X"1A",X"48",X"A8",X"81",
		X"30",X"91",X"F3",X"2B",X"2D",X"88",X"5A",X"01",X"C2",X"09",X"12",X"F8",X"3B",X"59",X"A3",X"9A",
		X"48",X"B0",X"19",X"5A",X"11",X"B1",X"82",X"A0",X"0A",X"89",X"78",X"98",X"80",X"82",X"04",X"D8",
		X"89",X"5A",X"00",X"D0",X"22",X"91",X"AA",X"A3",X"28",X"2C",X"2A",X"B3",X"01",X"0C",X"2A",X"30",
		X"98",X"4B",X"91",X"09",X"18",X"92",X"88",X"2A",X"93",X"89",X"5C",X"92",X"A3",X"89",X"A3",X"89",
		X"30",X"A3",X"B9",X"4B",X"20",X"D1",X"1A",X"93",X"88",X"4B",X"21",X"D1",X"3B",X"4A",X"E2",X"98",
		X"38",X"88",X"AA",X"48",X"11",X"8A",X"0B",X"35",X"BB",X"48",X"B0",X"22",X"99",X"00",X"10",X"18",
		X"BB",X"69",X"81",X"80",X"9D",X"79",X"92",X"9A",X"6B",X"11",X"9A",X"30",X"95",X"F1",X"09",X"20",
		X"8B",X"39",X"90",X"32",X"E1",X"D2",X"1A",X"10",X"1C",X"83",X"00",X"A6",X"AB",X"14",X"92",X"99",
		X"B9",X"27",X"0B",X"0A",X"81",X"5C",X"4B",X"84",X"C0",X"3B",X"02",X"91",X"99",X"97",X"C1",X"3F",
		X"21",X"A8",X"3B",X"00",X"08",X"89",X"02",X"3E",X"88",X"39",X"11",X"D1",X"81",X"84",X"E1",X"91",
		X"2D",X"22",X"E3",X"0B",X"94",X"C4",X"0C",X"29",X"95",X"89",X"90",X"83",X"0E",X"3A",X"02",X"89",
		X"8A",X"17",X"B0",X"81",X"08",X"B8",X"51",X"B0",X"8D",X"68",X"B6",X"A8",X"29",X"90",X"02",X"08",
		X"E1",X"19",X"10",X"08",X"AB",X"7A",X"11",X"A0",X"83",X"BB",X"7A",X"11",X"B3",X"9A",X"A7",X"91",
		X"08",X"A8",X"28",X"F7",X"A8",X"3D",X"29",X"18",X"82",X"C3",X"98",X"0A",X"5C",X"38",X"91",X"D4",
		X"A2",X"8B",X"49",X"88",X"2A",X"39",X"D4",X"91",X"8D",X"48",X"90",X"10",X"9A",X"83",X"2A",X"A0",
		X"49",X"B8",X"43",X"A9",X"F4",X"2E",X"1A",X"48",X"B1",X"21",X"D0",X"93",X"1B",X"19",X"4A",X"C2",
		X"31",X"F0",X"10",X"09",X"A1",X"3D",X"04",X"B3",X"AA",X"28",X"3B",X"2B",X"94",X"92",X"E4",X"8A",
		X"81",X"85",X"9B",X"A7",X"89",X"80",X"5D",X"02",X"A3",X"AA",X"15",X"A9",X"82",X"08",X"A8",X"20",
		X"9A",X"58",X"93",X"B4",X"99",X"18",X"0A",X"00",X"3F",X"E9",X"30",X"9A",X"37",X"21",X"41",X"C0",
		X"CA",X"0A",X"9D",X"DB",X"27",X"63",X"9C",X"98",X"02",X"09",X"AB",X"A0",X"83",X"77",X"A8",X"98",
		X"22",X"99",X"9D",X"9A",X"87",X"7A",X"9A",X"B4",X"69",X"99",X"C8",X"80",X"73",X"C0",X"C9",X"45",
		X"B0",X"AD",X"08",X"07",X"3D",X"0C",X"84",X"4A",X"1D",X"A8",X"19",X"73",X"D0",X"B9",X"55",X"B3",
		X"DC",X"03",X"C1",X"50",X"D5",X"D9",X"58",X"13",X"FA",X"3A",X"A1",X"70",X"A3",X"F9",X"58",X"23",
		X"FA",X"2B",X"85",X"5C",X"00",X"E0",X"59",X"30",X"F9",X"3C",X"85",X"4D",X"1A",X"B5",X"3B",X"4A",
		X"D0",X"2C",X"05",X"2D",X"3D",X"95",X"19",X"5C",X"C3",X"9A",X"17",X"0B",X"4D",X"95",X"88",X"5D",
		X"B4",X"A9",X"37",X"C0",X"1E",X"05",X"A1",X"4D",X"B5",X"B9",X"63",X"D0",X"0D",X"34",X"C3",X"1E",
		X"A4",X"B9",X"64",X"D2",X"BB",X"52",X"A4",X"9D",X"01",X"C0",X"53",X"D2",X"D9",X"51",X"95",X"AD",
		X"00",X"A0",X"71",X"D2",X"BA",X"61",X"94",X"AD",X"10",X"A0",X"70",X"B1",X"9B",X"25",X"A3",X"8F",
		X"01",X"A0",X"17",X"9A",X"1C",X"95",X"82",X"2F",X"91",X"90",X"01",X"69",X"A3",X"C8",X"40",X"98",
		X"B9",X"28",X"80",X"71",X"B0",X"B8",X"61",X"89",X"AA",X"00",X"88",X"72",X"C1",X"9A",X"34",X"99",
		X"8C",X"10",X"98",X"97",X"2C",X"28",X"B2",X"2B",X"28",X"E1",X"08",X"19",X"93",X"2A",X"38",X"C1",
		X"8A",X"48",X"A1",X"B1",X"4C",X"82",X"F0",X"11",X"84",X"01",X"9C",X"08",X"90",X"0A",X"8A",X"17",
		X"3C",X"10",X"B8",X"1A",X"01",X"92",X"2A",X"72",X"B0",X"88",X"A8",X"8B",X"99",X"25",X"AB",X"11",
		X"22",X"75",X"99",X"99",X"81",X"1A",X"9D",X"92",X"81",X"02",X"90",X"13",X"1E",X"40",X"A2",X"9B",
		X"19",X"A6",X"8A",X"1A",X"90",X"93",X"71",X"A8",X"9A",X"24",X"C0",X"09",X"0A",X"A6",X"2A",X"10",
		X"B0",X"10",X"29",X"C1",X"82",X"E8",X"2B",X"72",X"D0",X"80",X"38",X"B1",X"BE",X"51",X"90",X"8C",
		X"40",X"A0",X"89",X"78",X"98",X"98",X"40",X"B2",X"AC",X"60",X"91",X"9A",X"31",X"A0",X"9D",X"60",
		X"A0",X"89",X"21",X"90",X"9B",X"40",X"82",X"C8",X"3A",X"10",X"D8",X"58",X"80",X"C0",X"59",X"81",
		X"B0",X"3B",X"10",X"98",X"4C",X"14",X"D1",X"2B",X"01",X"B1",X"5C",X"83",X"C2",X"4C",X"81",X"91",
		X"3D",X"82",X"A1",X"3B",X"C2",X"00",X"5A",X"B2",X"B2",X"59",X"A9",X"81",X"78",X"B1",X"A3",X"4A",
		X"B9",X"95",X"5A",X"B1",X"91",X"59",X"98",X"B3",X"69",X"99",X"B2",X"78",X"A0",X"B2",X"79",X"90",
		X"A1",X"49",X"90",X"B0",X"79",X"81",X"C0",X"49",X"80",X"A0",X"30",X"A9",X"90",X"50",X"A8",X"B3",
		X"38",X"8A",X"B0",X"69",X"10",X"F2",X"09",X"3B",X"B5",X"81",X"0B",X"A5",X"0A",X"3C",X"96",X"A0",
		X"2C",X"12",X"C0",X"29",X"83",X"D0",X"3C",X"12",X"C2",X"0C",X"30",X"C2",X"1C",X"40",X"D2",X"98",
		X"5A",X"91",X"91",X"2B",X"94",X"A1",X"3E",X"82",X"92",X"0B",X"88",X"14",X"8C",X"80",X"17",X"AA",
		X"1A",X"51",X"D1",X"90",X"49",X"A1",X"99",X"78",X"B2",X"98",X"49",X"90",X"A2",X"39",X"B8",X"82",
		X"5A",X"A0",X"C5",X"2B",X"8A",X"06",X"0A",X"0A",X"04",X"89",X"0B",X"B6",X"1B",X"3A",X"B7",X"39",
		X"0A",X"B9",X"2A",X"CD",X"B1",X"67",X"18",X"8B",X"02",X"19",X"89",X"E8",X"8B",X"A9",X"87",X"72",
		X"9A",X"C2",X"11",X"1A",X"D8",X"8A",X"08",X"76",X"A8",X"8A",X"13",X"00",X"AD",X"81",X"B9",X"75",
		X"B0",X"8B",X"26",X"98",X"0C",X"82",X"9A",X"37",X"A9",X"2D",X"85",X"89",X"2C",X"A4",X"89",X"86",
		X"9A",X"2A",X"A3",X"3A",X"28",X"F0",X"19",X"0A",X"17",X"98",X"2C",X"94",X"89",X"3B",X"A3",X"89",
		X"90",X"78",X"92",X"C9",X"48",X"82",X"AB",X"49",X"89",X"B7",X"2A",X"2B",X"C3",X"19",X"49",X"C1",
		X"09",X"98",X"70",X"92",X"CA",X"48",X"83",X"AC",X"20",X"A8",X"33",X"B0",X"2F",X"84",X"90",X"2D",
		X"82",X"99",X"84",X"1A",X"08",X"C1",X"59",X"02",X"E8",X"29",X"98",X"78",X"A1",X"AA",X"34",X"91",
		X"0F",X"82",X"98",X"97",X"0A",X"0A",X"A3",X"30",X"2A",X"F8",X"19",X"0A",X"71",X"A8",X"9A",X"25",
		X"00",X"9D",X"81",X"80",X"93",X"4A",X"90",X"B0",X"70",X"90",X"D8",X"18",X"08",X"70",X"C0",X"09",
		X"23",X"AA",X"0C",X"01",X"A9",X"63",X"B1",X"1C",X"83",X"99",X"3E",X"91",X"01",X"48",X"B9",X"00",
		X"28",X"99",X"A0",X"63",X"09",X"BB",X"05",X"09",X"99",X"A0",X"D3",X"6C",X"24",X"B1",X"1B",X"82",
		X"D8",X"3C",X"04",X"A0",X"39",X"B2",X"8A",X"39",X"B2",X"20",X"83",X"AA",X"4C",X"08",X"97",X"89",
		X"89",X"01",X"B1",X"0A",X"40",X"B8",X"50",X"24",X"9C",X"09",X"A0",X"29",X"99",X"A9",X"61",X"11",
		X"BA",X"10",X"25",X"99",X"1A",X"91",X"B9",X"69",X"1A",X"D8",X"25",X"2B",X"B8",X"25",X"A9",X"09",
		X"15",X"AA",X"91",X"71",X"D9",X"01",X"3A",X"90",X"03",X"9D",X"01",X"84",X"8B",X"8B",X"63",X"AA",
		X"0B",X"51",X"D0",X"81",X"4A",X"99",X"85",X"0A",X"01",X"D3",X"1D",X"10",X"B6",X"8A",X"2A",X"84",
		X"0A",X"90",X"96",X"0D",X"18",X"03",X"A8",X"98",X"13",X"9C",X"2A",X"97",X"99",X"2B",X"04",X"99",
		X"1C",X"05",X"09",X"9A",X"97",X"1A",X"89",X"95",X"1A",X"89",X"82",X"28",X"C0",X"90",X"78",X"B2",
		X"9A",X"68",X"90",X"A0",X"21",X"89",X"90",X"82",X"59",X"C8",X"88",X"60",X"B8",X"8A",X"62",X"A9",
		X"8A",X"33",X"8A",X"BB",X"16",X"18",X"9C",X"84",X"28",X"8A",X"C2",X"49",X"09",X"B0",X"22",X"19",
		X"AC",X"42",X"98",X"AA",X"33",X"C1",X"88",X"94",X"1C",X"09",X"11",X"90",X"29",X"90",X"1B",X"20",
		X"A1",X"1C",X"33",X"F8",X"29",X"01",X"8A",X"09",X"41",X"8A",X"98",X"40",X"C4",X"99",X"89",X"02",
		X"29",X"81",X"A8",X"3B",X"01",X"0A",X"10",X"81",X"99",X"4A",X"90",X"A2",X"2B",X"83",X"9A",X"49",
		X"80",X"A0",X"3A",X"88",X"80",X"82",X"99",X"01",X"0B",X"04",X"9B",X"11",X"98",X"29",X"80",X"19",
		X"3B",X"A4",X"98",X"11",X"99",X"09",X"39",X"19",X"08",X"92",X"92",X"8A",X"19",X"82",X"0A",X"29",
		X"92",X"1B",X"91",X"90",X"5A",X"81",X"80",X"88",X"1A",X"00",X"8A",X"5A",X"A3",X"89",X"29",X"00",
		X"09",X"2A",X"92",X"80",X"2D",X"20",X"90",X"2D",X"03",X"A9",X"38",X"B4",X"8A",X"11",X"82",X"C0",
		X"09",X"11",X"A4",X"AC",X"15",X"A8",X"1B",X"12",X"90",X"A6",X"8A",X"89",X"03",X"30",X"B0",X"AF",
		X"00",X"A9",X"E2",X"74",X"18",X"99",X"80",X"BA",X"9F",X"C9",X"A3",X"77",X"88",X"A9",X"22",X"29",
		X"BC",X"00",X"19",X"DD",X"97",X"58",X"A8",X"A0",X"42",X"9A",X"A9",X"22",X"0A",X"FB",X"47",X"88",
		X"8B",X"84",X"18",X"0C",X"91",X"20",X"1D",X"C1",X"78",X"80",X"C8",X"30",X"83",X"DA",X"21",X"82",
		X"AF",X"85",X"08",X"0B",X"B3",X"31",X"1B",X"F8",X"30",X"18",X"DA",X"16",X"00",X"9D",X"83",X"10",
		X"1C",X"B3",X"10",X"2D",X"C0",X"50",X"01",X"E9",X"30",X"03",X"CB",X"21",X"83",X"BF",X"13",X"92",
		X"0F",X"83",X"81",X"2D",X"A3",X"88",X"3D",X"A7",X"8A",X"4B",X"B3",X"2A",X"48",X"D1",X"1A",X"18",
		X"D4",X"3C",X"18",X"D1",X"48",X"82",X"D8",X"28",X"80",X"E2",X"4A",X"01",X"D8",X"40",X"92",X"C9",
		X"20",X"80",X"E2",X"3A",X"01",X"D8",X"48",X"82",X"C9",X"28",X"80",X"C6",X"1B",X"3B",X"C3",X"19",
		X"39",X"D1",X"08",X"0C",X"15",X"98",X"3C",X"A5",X"09",X"1B",X"A3",X"08",X"8D",X"70",X"B3",X"AB",
		X"32",X"B3",X"9E",X"21",X"A0",X"C4",X"4A",X"92",X"BA",X"70",X"B2",X"AA",X"28",X"B7",X"3C",X"82",
		X"B0",X"39",X"92",X"C8",X"2A",X"04",X"A9",X"68",X"B2",X"1B",X"01",X"92",X"8B",X"11",X"B1",X"1B",
		X"01",X"09",X"42",X"00",X"82",X"3D",X"E1",X"0A",X"90",X"9B",X"4A",X"A4",X"15",X"41",X"91",X"BD",
		X"00",X"A9",X"89",X"04",X"80",X"39",X"A4",X"28",X"0A",X"F8",X"20",X"80",X"82",X"8B",X"03",X"C2",
		X"3C",X"81",X"AA",X"34",X"B9",X"2C",X"90",X"24",X"10",X"98",X"0B",X"E2",X"31",X"9F",X"91",X"12",
		X"09",X"99",X"14",X"3F",X"92",X"82",X"0D",X"A1",X"86",X"1D",X"01",X"A2",X"3C",X"92",X"08",X"2B",
		X"B3",X"88",X"5C",X"83",X"90",X"88",X"91",X"38",X"A2",X"9C",X"19",X"B6",X"1B",X"5A",X"A4",X"B3",
		X"1A",X"10",X"F0",X"2A",X"12",X"A9",X"1C",X"40",X"A5",X"98",X"1A",X"89",X"1A",X"25",X"B9",X"2E",
		X"13",X"89",X"10",X"C8",X"95",X"0B",X"31",X"BD",X"50",X"C1",X"3B",X"84",X"AA",X"3A",X"22",X"BB",
		X"01",X"B7",X"0A",X"19",X"81",X"9A",X"69",X"94",X"9A",X"81",X"A0",X"31",X"9B",X"03",X"81",X"0A",
		X"90",X"81",X"3C",X"A4",X"98",X"1E",X"13",X"08",X"1C",X"82",X"09",X"8B",X"03",X"08",X"0C",X"12",
		X"38",X"9B",X"11",X"08",X"0C",X"02",X"80",X"1C",X"21",X"81",X"80",X"91",X"A9",X"19",X"3A",X"88",
		X"2B",X"58",X"A3",X"AD",X"40",X"A3",X"9C",X"30",X"B4",X"8C",X"58",X"A2",X"0C",X"03",X"A8",X"88",
		X"21",X"98",X"89",X"83",X"1A",X"08",X"19",X"08",X"91",X"18",X"88",X"A1",X"29",X"00",X"99",X"29",
		X"20",X"8A",X"29",X"80",X"8A",X"39",X"81",X"0B",X"31",X"A2",X"0D",X"20",X"B1",X"2A",X"83",X"B8",
		X"4A",X"82",X"98",X"19",X"01",X"89",X"28",X"91",X"19",X"1B",X"00",X"80",X"1C",X"13",X"90",X"09",
		X"09",X"00",X"09",X"08",X"19",X"82",X"88",X"88",X"81",X"08",X"09",X"92",X"09",X"18",X"09",X"20",
		X"C2",X"0A",X"00",X"08",X"11",X"A0",X"80",X"1A",X"91",X"88",X"18",X"92",X"99",X"11",X"A1",X"01",
		X"90",X"91",X"88",X"1A",X"03",X"98",X"88",X"18",X"A3",X"90",X"00",X"A0",X"81",X"09",X"92",X"91",
		X"08",X"80",X"80",X"90",X"98",X"28",X"93",X"AA",X"3A",X"84",X"99",X"3A",X"B6",X"99",X"18",X"82",
		X"80",X"1A",X"18",X"08",X"19",X"A1",X"8A",X"68",X"90",X"1B",X"81",X"02",X"8A",X"31",X"C1",X"68",
		X"C9",X"BF",X"C9",X"96",X"73",X"C0",X"BA",X"63",X"8A",X"BA",X"12",X"9A",X"FA",X"74",X"B2",X"BB",
		X"52",X"91",X"9D",X"12",X"80",X"9C",X"B0",X"74",X"A0",X"C9",X"33",X"80",X"BC",X"13",X"81",X"AF",
		X"A7",X"19",X"1B",X"B2",X"40",X"19",X"F0",X"28",X"01",X"DA",X"51",X"92",X"BC",X"22",X"82",X"0F",
		X"82",X"80",X"1D",X"96",X"89",X"3C",X"B4",X"08",X"39",X"D1",X"19",X"00",X"D1",X"49",X"83",X"D9",
		X"38",X"84",X"BB",X"40",X"91",X"9E",X"33",X"B1",X"0E",X"04",X"90",X"2D",X"94",X"89",X"2C",X"A6",
		X"1B",X"3B",X"D2",X"28",X"20",X"F0",X"3A",X"82",X"F0",X"58",X"93",X"DA",X"58",X"94",X"AB",X"30",
		X"A3",X"CB",X"72",X"C2",X"9D",X"23",X"91",X"1F",X"12",X"A0",X"1F",X"05",X"89",X"4D",X"94",X"09",
		X"3B",X"B4",X"0A",X"3C",X"B6",X"2B",X"28",X"F1",X"49",X"02",X"D8",X"29",X"01",X"CA",X"71",X"B4",
		X"BB",X"32",X"94",X"9E",X"11",X"90",X"8C",X"61",X"B1",X"8C",X"23",X"A1",X"0D",X"82",X"98",X"8B",
		X"73",X"B0",X"8C",X"14",X"89",X"0B",X"83",X"89",X"0C",X"17",X"08",X"8A",X"92",X"10",X"0A",X"C1",
		X"08",X"20",X"C0",X"20",X"31",X"BA",X"0A",X"22",X"B9",X"09",X"B3",X"1B",X"63",X"A3",X"0E",X"01",
		X"B1",X"9A",X"21",X"95",X"1B",X"A5",X"29",X"8A",X"A8",X"11",X"88",X"C9",X"40",X"28",X"F9",X"41",
		X"02",X"8D",X"82",X"90",X"3C",X"92",X"A9",X"9C",X"27",X"09",X"29",X"A2",X"8B",X"13",X"B3",X"8C",
		X"BB",X"07",X"38",X"08",X"A8",X"18",X"B1",X"20",X"3A",X"FC",X"03",X"78",X"91",X"AA",X"31",X"99",
		X"2B",X"31",X"F8",X"0A",X"45",X"B1",X"1D",X"02",X"99",X"1A",X"23",X"B8",X"9D",X"16",X"89",X"3B",
		X"B6",X"8A",X"18",X"93",X"8A",X"1B",X"B7",X"2B",X"00",X"A4",X"3D",X"A3",X"A2",X"3C",X"90",X"A3",
		X"7A",X"B2",X"91",X"69",X"B1",X"80",X"39",X"91",X"D8",X"59",X"A1",X"88",X"58",X"A1",X"89",X"29",
		X"B4",X"0D",X"31",X"C0",X"3B",X"22",X"BA",X"49",X"94",X"BA",X"5A",X"94",X"9D",X"30",X"A3",X"0B",
		X"10",X"C2",X"2C",X"21",X"C1",X"3A",X"A3",X"C8",X"50",X"80",X"0B",X"18",X"92",X"8D",X"23",X"A2",
		X"0E",X"11",X"93",X"0A",X"A0",X"92",X"1C",X"94",X"A1",X"28",X"00",X"AA",X"58",X"A1",X"99",X"20",
		X"A1",X"89",X"21",X"A2",X"0A",X"02",X"B8",X"08",X"01",X"99",X"10",X"01",X"98",X"00",X"93",X"9A",
		X"01",X"92",X"0A",X"92",X"A2",X"08",X"91",X"91",X"19",X"98",X"01",X"08",X"80",X"00",X"91",X"80",
		X"89",X"01",X"A0",X"08",X"83",X"B0",X"81",X"90",X"82",X"98",X"91",X"08",X"00",X"A3",X"9A",X"20",
		X"90",X"92",X"08",X"80",X"81",X"89",X"91",X"80",X"01",X"98",X"01",X"09",X"91",X"92",X"88",X"80",
		X"08",X"80",X"91",X"91",X"08",X"88",X"81",X"91",X"A0",X"01",X"80",X"98",X"00",X"00",X"90",X"90",
		X"18",X"88",X"02",X"90",X"90",X"80",X"18",X"88",X"81",X"00",X"80",X"80",X"09",X"90",X"80",X"11",
		X"90",X"90",X"88",X"08",X"98",X"10",X"00",X"90",X"92",X"00",X"99",X"08",X"02",X"9A",X"10",X"91",
		X"81",X"80",X"88",X"81",X"90",X"08",X"81",X"90",X"08",X"00",X"90",X"18",X"08",X"91",X"92",X"A1",
		X"99",X"38",X"92",X"A8",X"3A",X"93",X"88",X"80",X"82",X"89",X"08",X"A1",X"0A",X"11",X"91",X"90",
		X"08",X"91",X"80",X"81",X"88",X"82",X"80",X"08",X"80",X"AA",X"AE",X"91",X"E7",X"78",X"A8",X"A1",
		X"50",X"99",X"BB",X"0A",X"D4",X"72",X"C2",X"D8",X"40",X"91",X"BA",X"42",X"88",X"BD",X"98",X"75",
		X"A9",X"8A",X"06",X"09",X"8A",X"94",X"11",X"9D",X"98",X"07",X"2B",X"8A",X"93",X"48",X"8A",X"C1",
		X"32",X"0B",X"F8",X"05",X"2A",X"9B",X"92",X"60",X"8A",X"B0",X"32",X"3C",X"D9",X"05",X"28",X"AB",
		X"A2",X"51",X"0B",X"B8",X"24",X"2B",X"D9",X"05",X"39",X"9D",X"92",X"22",X"0C",X"B0",X"25",X"0B",
		X"BA",X"36",X"18",X"AC",X"83",X"21",X"8E",X"91",X"13",X"8C",X"A9",X"61",X"08",X"C9",X"12",X"12",
		X"AD",X"81",X"21",X"AC",X"A2",X"61",X"89",X"C8",X"22",X"10",X"E9",X"11",X"28",X"BC",X"97",X"18",
		X"0B",X"B2",X"31",X"3B",X"F8",X"20",X"18",X"BC",X"07",X"18",X"8C",X"92",X"21",X"1C",X"B1",X"28",
		X"28",X"F8",X"84",X"39",X"AA",X"B2",X"61",X"89",X"C8",X"20",X"10",X"CA",X"02",X"70",X"A9",X"89",
		X"42",X"99",X"9A",X"11",X"00",X"BB",X"97",X"48",X"89",X"A8",X"22",X"09",X"C9",X"10",X"00",X"AA",
		X"07",X"31",X"AA",X"89",X"02",X"8C",X"99",X"01",X"11",X"1A",X"26",X"89",X"19",X"90",X"A9",X"0A",
		X"85",X"80",X"08",X"21",X"09",X"8B",X"A7",X"1A",X"8C",X"91",X"10",X"08",X"92",X"03",X"38",X"8B",
		X"A2",X"22",X"DF",X"81",X"11",X"98",X"99",X"14",X"40",X"99",X"CA",X"12",X"9B",X"98",X"41",X"82",
		X"8A",X"23",X"18",X"2D",X"9B",X"A0",X"28",X"11",X"1A",X"11",X"02",X"91",X"8A",X"10",X"0D",X"9A",
		X"23",X"05",X"9A",X"2A",X"11",X"8A",X"3E",X"04",X"9B",X"99",X"35",X"82",X"9B",X"A2",X"93",X"8A",
		X"89",X"84",X"0C",X"99",X"26",X"01",X"9D",X"01",X"82",X"0C",X"19",X"14",X"9B",X"88",X"24",X"8A",
		X"8C",X"96",X"19",X"09",X"88",X"80",X"09",X"29",X"21",X"9B",X"1B",X"04",X"08",X"98",X"09",X"19",
		X"88",X"21",X"28",X"B9",X"89",X"41",X"9A",X"00",X"03",X"9E",X"00",X"04",X"2C",X"09",X"91",X"30",
		X"AB",X"80",X"40",X"8A",X"98",X"51",X"88",X"BB",X"03",X"00",X"0C",X"82",X"01",X"99",X"A2",X"04",
		X"0A",X"99",X"A2",X"38",X"99",X"B4",X"11",X"98",X"B8",X"33",X"88",X"BA",X"04",X"80",X"8C",X"83",
		X"02",X"89",X"B0",X"22",X"08",X"AA",X"95",X"19",X"99",X"A3",X"20",X"09",X"A9",X"04",X"89",X"99",
		X"82",X"39",X"0A",X"A3",X"00",X"08",X"B0",X"02",X"89",X"A0",X"82",X"01",X"88",X"90",X"01",X"A0",
		X"80",X"94",X"89",X"08",X"90",X"29",X"92",X"A1",X"18",X"90",X"98",X"01",X"81",X"98",X"80",X"01",
		X"89",X"80",X"82",X"98",X"08",X"80",X"00",X"88",X"80",X"00",X"90",X"80",X"80",X"01",X"98",X"81",
		X"A2",X"88",X"80",X"00",X"00",X"90",X"80",X"81",X"90",X"88",X"81",X"90",X"09",X"10",X"00",X"80",
		X"A0",X"81",X"90",X"80",X"00",X"81",X"90",X"88",X"81",X"89",X"18",X"08",X"81",X"90",X"80",X"80",
		X"08",X"00",X"90",X"08",X"00",X"A2",X"80",X"08",X"88",X"81",X"92",X"89",X"00",X"91",X"08",X"80",
		X"92",X"80",X"90",X"88",X"01",X"88",X"90",X"81",X"91",X"91",X"A1",X"00",X"88",X"90",X"81",X"80",
		X"90",X"81",X"18",X"91",X"88",X"00",X"88",X"80",X"00",X"00",X"98",X"00",X"01",X"99",X"00",X"01",
		X"A8",X"80",X"00",X"08",X"89",X"02",X"A1",X"98",X"10",X"92",X"A8",X"00",X"81",X"90",X"80",X"81",
		X"80",X"90",X"80",X"80",X"00",X"80",X"08",X"88",X"80",X"82",X"80",X"90",X"00",X"90",X"91",X"80",
		X"08",X"A2",X"89",X"18",X"81",X"98",X"10",X"91",X"88",X"81",X"88",X"09",X"81",X"80",X"90",X"82",
		X"01",X"89",X"88",X"82",X"98",X"08",X"10",X"A2",X"89",X"88",X"A0",X"BC",X"F2",X"77",X"A9",X"99",
		X"35",X"89",X"BA",X"88",X"B0",X"77",X"B1",X"AA",X"43",X"90",X"AE",X"13",X"00",X"8D",X"02",X"A8",
		X"AA",X"74",X"A0",X"AC",X"42",X"80",X"AC",X"03",X"11",X"9B",X"A9",X"BA",X"77",X"A1",X"BA",X"52",
		X"90",X"9C",X"03",X"00",X"1C",X"90",X"AA",X"74",X"C1",X"A9",X"41",X"91",X"9C",X"03",X"80",X"1C",
		X"80",X"A9",X"72",X"C2",X"BA",X"51",X"91",X"9C",X"13",X"90",X"1C",X"80",X"99",X"71",X"B2",X"BB",
		X"61",X"90",X"8C",X"13",X"88",X"1C",X"92",X"AA",X"72",X"C1",X"9A",X"42",X"A0",X"8C",X"04",X"88",
		X"1B",X"A2",X"9B",X"73",X"D1",X"8A",X"24",X"A8",X"0C",X"04",X"88",X"1B",X"A3",X"9B",X"64",X"B8",
		X"1C",X"05",X"99",X"2B",X"95",X"89",X"2A",X"A2",X"8A",X"15",X"19",X"99",X"A2",X"41",X"9B",X"C1",
		X"21",X"29",X"E9",X"18",X"02",X"1A",X"48",X"B3",X"1C",X"21",X"C0",X"2D",X"82",X"A0",X"2C",X"82",
		X"99",X"53",X"82",X"AC",X"28",X"83",X"9E",X"98",X"02",X"09",X"B9",X"11",X"25",X"31",X"AB",X"18",
		X"37",X"9C",X"A9",X"83",X"08",X"9C",X"83",X"02",X"21",X"A8",X"98",X"43",X"19",X"E9",X"2B",X"13",
		X"8E",X"80",X"91",X"40",X"80",X"D8",X"20",X"20",X"B9",X"39",X"B4",X"1D",X"81",X"A0",X"39",X"01",
		X"89",X"30",X"88",X"D8",X"60",X"88",X"B9",X"04",X"08",X"1C",X"A1",X"21",X"28",X"09",X"C9",X"33",
		X"19",X"8A",X"A3",X"18",X"2A",X"A9",X"18",X"21",X"18",X"AC",X"12",X"80",X"2B",X"B3",X"18",X"29",
		X"90",X"19",X"89",X"12",X"0D",X"01",X"92",X"29",X"C1",X"20",X"19",X"D0",X"12",X"0A",X"80",X"19",
		X"11",X"0B",X"00",X"90",X"18",X"89",X"19",X"21",X"09",X"A8",X"29",X"08",X"09",X"11",X"80",X"89",
		X"09",X"00",X"18",X"09",X"81",X"18",X"A1",X"8A",X"20",X"91",X"00",X"09",X"88",X"18",X"08",X"89",
		X"10",X"08",X"08",X"08",X"08",X"08",X"19",X"09",X"00",X"09",X"18",X"00",X"0A",X"08",X"19",X"19",
		X"08",X"00",X"89",X"10",X"09",X"08",X"10",X"08",X"B8",X"10",X"20",X"99",X"88",X"20",X"89",X"89",
		X"10",X"28",X"19",X"90",X"80",X"18",X"98",X"29",X"18",X"08",X"90",X"88",X"00",X"00",X"89",X"09",
		X"10",X"09",X"19",X"08",X"00",X"88",X"08",X"18",X"10",X"90",X"98",X"19",X"09",X"28",X"18",X"89",
		X"00",X"08",X"88",X"29",X"08",X"00",X"09",X"08",X"80",X"19",X"88",X"00",X"08",X"80",X"08",X"09",
		X"08",X"19",X"08",X"08",X"18",X"80",X"88",X"00",X"08",X"88",X"18",X"00",X"09",X"88",X"10",X"08",
		X"88",X"09",X"19",X"80",X"08",X"10",X"09",X"09",X"80",X"08",X"18",X"09",X"19",X"18",X"89",X"18",
		X"00",X"80",X"09",X"00",X"09",X"28",X"0A",X"00",X"19",X"1A",X"08",X"10",X"88",X"09",X"00",X"08",
		X"08",X"08",X"19",X"08",X"88",X"08",X"09",X"18",X"18",X"88",X"00",X"08",X"08",X"88",X"00",X"08",
		X"19",X"08",X"08",X"09",X"00",X"88",X"08",X"08",X"19",X"18",X"08",X"09",X"19",X"00",X"08",X"18",
		X"88",X"88",X"08",X"00",X"08",X"09",X"19",X"18",X"88",X"00",X"08",X"18",X"88",X"88",X"10",X"08",
		X"89",X"00",X"08",X"88",X"08",X"10",X"09",X"88",X"09",X"39",X"08",X"08",X"19",X"80",X"88",X"10",
		X"09",X"08",X"09",X"19",X"08",X"08",X"00",X"80",X"88",X"08",X"00",X"08",X"08",X"88",X"08",X"00",
		X"80",X"91",X"08",X"08",X"08",X"08",X"80",X"08",X"09",X"18",X"08",X"88",X"18",X"08",X"80",X"88",
		X"08",X"00",X"00",X"08",X"88",X"08",X"08",X"89",X"18",X"18",X"88",X"08",X"18",X"08",X"08",X"08",
		X"09",X"00",X"80",X"08",X"08",X"88",X"19",X"00",X"08",X"19",X"08",X"88",X"18",X"08",X"88",X"18",
		X"80",X"88",X"19",X"00",X"09",X"29",X"08",X"08",X"80",X"08",X"09",X"18",X"08",X"09",X"18",X"08",
		X"88",X"99",X"B9",X"B7",X"71",X"B0",X"BB",X"72",X"90",X"8D",X"82",X"89",X"E9",X"72",X"90",X"AC",
		X"14",X"00",X"8C",X"92",X"10",X"3B",X"D1",X"00",X"39",X"CA",X"D9",X"75",X"A1",X"BB",X"34",X"92",
		X"9E",X"82",X"01",X"2C",X"A2",X"88",X"4A",X"F4",X"0A",X"20",X"C0",X"29",X"03",X"CA",X"38",X"95",
		X"8B",X"11",X"B2",X"1E",X"93",X"38",X"19",X"F0",X"10",X"11",X"C9",X"18",X"14",X"9B",X"08",X"02",
		X"9E",X"A3",X"70",X"88",X"C9",X"31",X"02",X"CB",X"11",X"04",X"0C",X"80",X"91",X"0D",X"97",X"1A",
		X"18",X"C1",X"39",X"01",X"D9",X"38",X"04",X"BA",X"2A",X"83",X"AF",X"27",X"98",X"1C",X"83",X"80",
		X"1A",X"B2",X"19",X"21",X"D8",X"19",X"02",X"D9",X"37",X"88",X"8B",X"82",X"11",X"0B",X"B0",X"10",
		X"31",X"CB",X"88",X"22",X"A9",X"85",X"70",X"80",X"AA",X"10",X"01",X"BC",X"08",X"83",X"0C",X"90",
		X"83",X"3A",X"06",X"19",X"51",X"A8",X"8B",X"92",X"89",X"9F",X"92",X"98",X"38",X"93",X"09",X"51",
		X"91",X"00",X"38",X"CB",X"A0",X"40",X"A9",X"98",X"89",X"28",X"20",X"9A",X"21",X"19",X"08",X"0A",
		X"08",X"A1",X"49",X"9A",X"19",X"2A",X"30",X"90",X"09",X"10",X"89",X"00",X"09",X"88",X"80",X"38",
		X"8A",X"2C",X"4A",X"3A",X"88",X"85",X"B2",X"2E",X"80",X"11",X"B6",X"C1",X"90",X"88",X"48",X"9A",
		X"11",X"8D",X"32",X"2F",X"10",X"82",X"0C",X"10",X"8A",X"01",X"88",X"0C",X"94",X"2D",X"19",X"92",
		X"12",X"B4",X"A9",X"3B",X"31",X"C1",X"A3",X"A5",X"E1",X"19",X"10",X"91",X"93",X"BC",X"A2",X"79",
		X"91",X"D4",X"A2",X"08",X"91",X"B4",X"03",X"9E",X"1A",X"11",X"83",X"9B",X"3E",X"3B",X"20",X"59",
		X"B0",X"97",X"B3",X"C0",X"21",X"B1",X"C5",X"D1",X"1A",X"3A",X"11",X"8B",X"20",X"2C",X"58",X"D1",
		X"A4",X"90",X"A4",X"D1",X"92",X"28",X"88",X"A9",X"30",X"3C",X"9A",X"59",X"08",X"95",X"B0",X"91",
		X"2D",X"5F",X"11",X"08",X"A8",X"2A",X"20",X"38",X"CA",X"10",X"A7",X"82",X"9D",X"28",X"12",X"0A",
		X"CC",X"03",X"28",X"08",X"F9",X"22",X"3B",X"2F",X"2A",X"2E",X"48",X"92",X"92",X"19",X"1D",X"20",
		X"00",X"8E",X"A9",X"06",X"12",X"AA",X"A3",X"56",X"89",X"EB",X"90",X"13",X"90",X"D0",X"84",X"12",
		X"88",X"80",X"12",X"3A",X"1B",X"05",X"73",X"93",X"80",X"80",X"88",X"FF",X"F8",X"08",X"08",X"08",
		X"00",X"73",X"AA",X"99",X"17",X"90",X"B9",X"03",X"78",X"80",X"88",X"E2",X"92",X"AA",X"08",X"01",
		X"07",X"B1",X"A3",X"11",X"99",X"E1",X"32",X"90",X"80",X"80",X"F3",X"88",X"F8",X"08",X"08",X"60",
		X"8C",X"80",X"06",X"90",X"C1",X"80",X"38",X"08",X"A9",X"A2",X"80",X"B1",X"88",X"07",X"30",X"A0",
		X"F5",X"88",X"08",X"08",X"BB",X"70",X"80",X"D0",X"08",X"31",X"88",X"F1",X"80",X"49",X"0C",X"08",
		X"04",X"80",X"C8",X"08",X"03",X"B8",X"00",X"70",X"88",X"08",X"08",X"08",X"BF",X"13",X"19",X"AB",
		X"80",X"62",X"91",X"F8",X"08",X"24",X"D8",X"08",X"04",X"80",X"C8",X"08",X"12",X"A1",X"D2",X"48",
		X"08",X"08",X"E8",X"14",X"90",X"E1",X"82",X"18",X"80",X"F1",X"80",X"49",X"8B",X"18",X"15",X"99",
		X"B1",X"80",X"7B",X"80",X"83",X"29",X"08",X"0D",X"A1",X"33",X"AE",X"91",X"24",X"90",X"8F",X"00",
		X"84",X"80",X"C8",X"08",X"31",X"F1",X"80",X"12",X"D1",X"02",X"90",X"80",X"8F",X"10",X"39",X"0A",
		X"C5",X"08",X"08",X"D0",X"08",X"48",X"0C",X"08",X"08",X"19",X"08",X"03",X"59",X"00",X"80",X"88",
		X"8F",X"89",X"78",X"08",X"C4",X"80",X"89",X"B1",X"80",X"41",X"8F",X"00",X"80",X"80",X"80",X"41",
		X"D2",X"18",X"08",X"8A",X"E1",X"14",X"90",X"8E",X"13",X"90",X"AB",X"18",X"07",X"08",X"C8",X"00",
		X"80",X"1A",X"01",X"97",X"00",X"80",X"80",X"9F",X"01",X"49",X"08",X"80",X"80",X"8F",X"08",X"80",
		X"07",X"B8",X"08",X"08",X"08",X"83",X"59",X"18",X"80",X"80",X"8D",X"D1",X"50",X"88",X"08",X"81",
		X"AF",X"08",X"00",X"80",X"80",X"84",X"59",X"E0",X"08",X"23",X"90",X"80",X"88",X"08",X"0D",X"48",
		X"80",X"80",X"80",X"FB",X"19",X"00",X"80",X"80",X"80",X"47",X"E0",X"08",X"06",X"88",X"08",X"08",
		X"08",X"08",X"0F",X"48",X"80",X"80",X"8F",X"00",X"80",X"80",X"80",X"80",X"80",X"7B",X"80",X"84",
		X"83",X"90",X"80",X"80",X"80",X"80",X"88",X"08",X"08",X"08",X"FF",X"A0",X"80",X"80",X"80",X"80",
		X"80",X"08",X"7B",X"70",X"18",X"4A",X"18",X"08",X"80",X"80",X"80",X"88",X"08",X"0A",X"FF",X"A4",
		X"C0",X"08",X"08",X"08",X"08",X"08",X"08",X"27",X"78",X"0F",X"03",X"80",X"88",X"08",X"08",X"08",
		X"08",X"08",X"08",X"F2",X"F5",X"98",X"B2",X"90",X"08",X"08",X"08",X"08",X"02",X"97",X"B6",X"98",
		X"02",X"90",X"08",X"80",X"F4",X"88",X"A9",X"15",X"90",X"80",X"F3",X"A3",X"C1",X"B2",X"90",X"08",
		X"08",X"08",X"08",X"08",X"65",X"B9",X"20",X"3A",X"18",X"A1",X"F1",X"49",X"08",X"BA",X"7D",X"49",
		X"00",X"88",X"A8",X"84",X"82",X"E0",X"88",X"08",X"19",X"08",X"08",X"03",X"3E",X"12",X"82",X"E2",
		X"28",X"08",X"90",X"19",X"D1",X"B7",X"8B",X"3C",X"14",X"99",X"0F",X"11",X"29",X"0E",X"18",X"2B",
		X"19",X"01",X"0A",X"3C",X"6A",X"18",X"3B",X"2C",X"39",X"1B",X"79",X"00",X"9C",X"20",X"2A",X"1A",
		X"3E",X"1A",X"59",X"1C",X"09",X"49",X"10",X"AA",X"58",X"10",X"CA",X"18",X"39",X"09",X"79",X"99",
		X"80",X"32",X"0D",X"A8",X"25",X"18",X"AA",X"00",X"28",X"09",X"80",X"89",X"41",X"3A",X"1F",X"9D",
		X"11",X"3A",X"08",X"04",X"B9",X"BC",X"32",X"8B",X"0B",X"61",X"14",X"9C",X"8A",X"48",X"08",X"40",
		X"49",X"99",X"98",X"83",X"90",X"C8",X"32",X"0E",X"AA",X"19",X"41",X"A0",X"A8",X"14",X"21",X"BB",
		X"9B",X"87",X"00",X"A5",X"87",X"8A",X"B0",X"17",X"91",X"A0",X"B3",X"C2",X"8A",X"0B",X"21",X"8E",
		X"02",X"61",X"0B",X"A9",X"11",X"13",X"B0",X"92",X"68",X"8E",X"00",X"02",X"B2",X"91",X"80",X"B2",
		X"DB",X"96",X"B8",X"D1",X"17",X"00",X"A0",X"A4",X"A2",X"B2",X"93",X"04",X"AA",X"0B",X"28",X"2F",
		X"28",X"08",X"A4",X"B2",X"A1",X"98",X"8F",X"1B",X"4A",X"68",X"2B",X"0B",X"01",X"58",X"09",X"82",
		X"12",X"4D",X"AC",X"28",X"69",X"1B",X"1C",X"2A",X"82",X"93",X"C1",X"B1",X"10",X"0A",X"4A",X"29",
		X"E2",X"16",X"00",X"8A",X"8C",X"48",X"49",X"A9",X"08",X"69",X"0A",X"88",X"A9",X"83",X"80",X"08",
		X"32",X"C2",X"6C",X"1F",X"91",X"22",X"28",X"0A",X"0B",X"80",X"97",X"A1",X"2B",X"2C",X"49",X"3D",
		X"0B",X"89",X"21",X"83",X"D4",X"92",X"A2",X"B2",X"E5",X"88",X"1C",X"29",X"11",X"19",X"C1",X"A2",
		X"84",X"82",X"DA",X"81",X"F7",X"B4",X"B1",X"99",X"4B",X"5A",X"88",X"01",X"28",X"0A",X"AA",X"50",
		X"28",X"9B",X"88",X"71",X"0B",X"A9",X"20",X"20",X"B8",X"A0",X"11",X"0C",X"8C",X"50",X"1B",X"93",
		X"04",X"A0",X"4A",X"29",X"BF",X"3C",X"7A",X"5B",X"0A",X"21",X"10",X"D9",X"00",X"68",X"99",X"80",
		X"18",X"69",X"BC",X"10",X"59",X"00",X"80",X"BB",X"25",X"11",X"BB",X"08",X"84",X"11",X"D8",X"B3",
		X"04",X"83",X"AA",X"97",X"79",X"20",X"88",X"8F",X"C9",X"13",X"19",X"9C",X"90",X"80",X"08",X"00",
		X"62",X"18",X"4E",X"0C",X"71",X"90",X"0C",X"A7",X"88",X"08",X"00",X"9B",X"91",X"08",X"18",X"B2",
		X"23",X"02",X"FA",X"84",X"18",X"E0",X"07",X"80",X"88",X"D1",X"21",X"90",X"80",X"80",X"8F",X"80",
		X"81",X"3E",X"5A",X"1A",X"09",X"2A",X"2B",X"18",X"52",X"90",X"8F",X"00",X"49",X"00",X"80",X"80",
		X"F0",X"80",X"48",X"A1",X"C1",X"91",X"85",X"B1",X"B1",X"87",X"80",X"8A",X"A1",X"32",X"90",X"80",
		X"08",X"AF",X"88",X"78",X"0D",X"18",X"80",X"10",X"2F",X"18",X"84",X"80",X"8A",X"A1",X"06",X"90",
		X"08",X"08",X"D8",X"01",X"49",X"0E",X"18",X"80",X"5B",X"3D",X"18",X"85",X"90",X"8C",X"18",X"13",
		X"90",X"80",X"BD",X"18",X"50",X"90",X"C0",X"80",X"86",X"80",X"D1",X"88",X"59",X"00",X"B8",X"03",
		X"18",X"08",X"8E",X"90",X"16",X"D0",X"00",X"91",X"93",X"29",X"B9",X"80",X"27",X"80",X"8E",X"08",
		X"69",X"08",X"08",X"9B",X"18",X"4A",X"3C",X"91",X"81",X"79",X"8B",X"19",X"17",X"90",X"09",X"C1",
		X"04",X"90",X"80",X"9D",X"18",X"14",X"9B",X"91",X"80",X"78",X"0A",X"B1",X"87",X"80",X"89",X"B1",
		X"58",X"80",X"08",X"9E",X"18",X"40",X"9C",X"18",X"80",X"58",X"0C",X"80",X"05",X"90",X"08",X"E1",
		X"11",X"80",X"88",X"BA",X"18",X"78",X"0D",X"18",X"80",X"58",X"8B",X"80",X"87",X"88",X"08",X"B8",
		X"04",X"08",X"08",X"9F",X"18",X"31",X"99",X"C1",X"88",X"35",X"90",X"F0",X"02",X"19",X"08",X"08",
		X"F3",X"08",X"08",X"08",X"F0",X"08",X"48",X"C1",X"80",X"80",X"30",X"8C",X"88",X"17",X"90",X"80",
		X"80",X"91",X"08",X"08",X"80",X"FA",X"08",X"18",X"80",X"80",X"80",X"07",X"28",X"D8",X"16",X"88",
		X"08",X"08",X"08",X"08",X"08",X"08",X"0F",X"D0",X"87",X"99",X"91",X"88",X"01",X"7A",X"98",X"00",
		X"22",X"88",X"92",X"88",X"08",X"08",X"92",X"90",X"9F",X"F8",X"81",X"90",X"08",X"08",X"00",X"70",
		X"A8",X"B7",X"20",X"80",X"C4",X"90",X"08",X"08",X"80",X"80",X"91",X"F6",X"F1",X"80",X"80",X"90",
		X"08",X"08",X"06",X"C1",X"93",X"84",X"90",X"A1",X"A4",X"A2",X"80",X"88",X"08",X"08",X"A8",X"4F",
		X"2F",X"09",X"15",X"8C",X"08",X"08",X"2A",X"08",X"03",X"4F",X"2A",X"20",X"19",X"99",X"05",X"80",
		X"89",X"C6",X"90",X"08",X"9A",X"A7",X"0B",X"80",X"02",X"B9",X"18",X"02",X"C3",X"99",X"40",X"33",
		X"E2",X"09",X"2B",X"86",X"90",X"8E",X"12",X"80",X"8A",X"A3",X"09",X"F0",X"85",X"1B",X"B0",X"80",
		X"01",X"31",X"E2",X"91",X"3D",X"20",X"B2",X"94",X"20",X"8A",X"AE",X"98",X"70",X"0A",X"0A",X"3C",
		X"02",X"92",X"80",X"08",X"D0",X"AB",X"73",X"90",X"D2",X"29",X"BA",X"80",X"78",X"28",X"B0",X"99",
		X"95",X"83",X"92",X"B9",X"03",X"80",X"FA",X"22",X"41",X"9A",X"C9",X"C2",X"02",X"52",X"9C",X"AC",
		X"13",X"11",X"B0",X"97",X"80",X"B1",X"A9",X"83",X"37",X"08",X"BB",X"E1",X"05",X"01",X"99",X"B9",
		X"82",X"41",X"8A",X"B1",X"23",X"00",X"CF",X"98",X"51",X"38",X"BA",X"C8",X"20",X"51",X"99",X"98",
		X"A0",X"94",X"21",X"C0",X"A1",X"83",X"08",X"9D",X"94",X"51",X"9B",X"A2",X"90",X"A8",X"71",X"2C",
		X"BA",X"02",X"50",X"0C",X"90",X"31",X"8A",X"A9",X"20",X"12",X"4A",X"3F",X"A0",X"82",X"06",X"A0",
		X"D0",X"01",X"01",X"90",X"99",X"10",X"51",X"BA",X"9C",X"04",X"40",X"08",X"D9",X"81",X"52",X"8A",
		X"F8",X"01",X"28",X"0A",X"89",X"A1",X"53",X"89",X"C8",X"A4",X"05",X"18",X"CB",X"A8",X"53",X"38",
		X"8E",X"AA",X"12",X"40",X"89",X"AB",X"81",X"50",X"0C",X"98",X"43",X"29",X"9C",X"B9",X"34",X"70",
		X"89",X"99",X"C8",X"86",X"10",X"B9",X"A2",X"08",X"92",X"8A",X"39",X"35",X"1C",X"0D",X"00",X"27",
		X"01",X"C8",X"A0",X"91",X"41",X"0E",X"80",X"0A",X"88",X"13",X"A0",X"A2",X"25",X"A9",X"C9",X"46",
		X"10",X"A9",X"A2",X"98",X"20",X"80",X"B2",X"1D",X"F0",X"13",X"9A",X"A3",X"59",X"A9",X"92",X"13",
		X"41",X"0F",X"99",X"30",X"6B",X"01",X"C8",X"10",X"19",X"98",X"1C",X"1A",X"70",X"2E",X"09",X"02",
		X"28",X"3E",X"2C",X"88",X"32",X"0A",X"AC",X"11",X"81",X"38",X"8D",X"2F",X"3C",X"59",X"1A",X"18",
		X"88",X"31",X"1D",X"BA",X"52",X"18",X"AB",X"98",X"33",X"9C",X"09",X"32",X"BC",X"F4",X"20",X"BC",
		X"95",X"31",X"9A",X"9D",X"40",X"00",X"9A",X"40",X"4B",X"99",X"13",X"13",X"C9",X"C9",X"88",X"EB",
		X"19",X"21",X"C8",X"A8",X"09",X"F7",X"30",X"9D",X"82",X"63",X"90",X"8E",X"D2",X"59",X"00",X"80",
		X"9E",X"18",X"1A",X"08",X"02",X"59",X"A8",X"A0",X"80",X"4A",X"92",X"70",X"08",X"F0",X"85",X"88",
		X"08",X"08",X"0A",X"D1",X"05",X"B9",X"02",X"28",X"0D",X"90",X"08",X"08",X"04",X"59",X"0A",X"E1",
		X"05",X"90",X"80",X"80",X"89",X"E1",X"84",X"0A",X"80",X"20",X"D9",X"08",X"08",X"00",X"83",X"78",
		X"09",X"F1",X"03",X"90",X"81",X"90",X"0B",X"F1",X"84",X"08",X"98",X"82",X"F0",X"00",X"09",X"80",
		X"85",X"29",X"0B",X"D1",X"24",X"98",X"82",X"90",X"0F",X"A1",X"87",X"89",X"92",X"18",X"D0",X"80",
		X"80",X"80",X"07",X"80",X"8D",X"00",X"48",X"89",X"28",X"80",X"8F",X"08",X"31",X"BA",X"78",X"8A",
		X"91",X"88",X"08",X"00",X"78",X"00",X"F1",X"83",X"08",X"08",X"80",X"80",X"F0",X"88",X"19",X"17",
		X"90",X"C0",X"08",X"81",X"90",X"07",X"91",X"8D",X"18",X"38",X"08",X"08",X"08",X"CB",X"18",X"07",
		X"B4",X"08",X"9B",X"08",X"87",X"B0",X"83",X"29",X"0B",X"D1",X"07",X"90",X"80",X"0D",X"08",X"59",
		X"0A",X"88",X"1A",X"78",X"8C",X"2A",X"2A",X"18",X"58",X"08",X"8D",X"10",X"49",X"08",X"09",X"E1",
		X"85",X"90",X"9A",X"08",X"06",X"89",X"92",X"C1",X"90",X"15",X"90",X"0D",X"80",X"59",X"00",X"80",
		X"D0",X"80",X"48",X"09",X"C1",X"88",X"41",X"A2",X"F0",X"08",X"14",X"90",X"89",X"D1",X"22",X"90",
		X"80",X"BE",X"18",X"33",X"9A",X"E1",X"80",X"86",X"80",X"9B",X"08",X"26",X"90",X"80",X"8E",X"04",
		X"88",X"08",X"0B",X"B2",X"96",X"19",X"C0",X"80",X"80",X"78",X"0A",X"A1",X"10",X"39",X"00",X"80",
		X"88",X"E3",X"00",X"88",X"0F",X"B1",X"80",X"78",X"C0",X"08",X"08",X"34",X"99",X"E1",X"83",X"18",
		X"81",X"88",X"08",X"08",X"9F",X"82",X"12",X"99",X"EA",X"00",X"80",X"80",X"80",X"08",X"43",X"4F",
		X"08",X"41",X"09",X"8A",X"40",X"80",X"80",X"8A",X"AF",X"78",X"80",X"8E",X"00",X"80",X"59",X"B0",
		X"08",X"08",X"10",X"29",X"D2",X"84",X"28",X"89",X"9A",X"78",X"08",X"08",X"08",X"0D",X"C1",X"79",
		X"1D",X"00",X"88",X"08",X"00",X"91",X"01",X"0B",X"84",X"12",X"09",X"48",X"A2",X"1B",X"2E",X"B2",
		X"25",X"90",X"AF",X"00",X"20",X"9E",X"1A",X"59",X"1A",X"0A",X"08",X"22",X"2A",X"2E",X"01",X"12",
		X"3D",X"09",X"04",X"8E",X"00",X"12",X"9A",X"A9",X"24",X"01",X"D9",X"1A",X"3B",X"48",X"3F",X"08",
		X"00",X"18",X"3D",X"88",X"82",X"1A",X"38",X"A1",X"A0",X"2A",X"72",X"E0",X"89",X"21",X"23",X"E9",
		X"91",X"20",X"A4",X"A0",X"AE",X"14",X"A2",X"8B",X"A8",X"87",X"80",X"08",X"91",X"B1",X"C3",X"32",
		X"02",X"DA",X"9A",X"36",X"13",X"BF",X"A1",X"04",X"08",X"A9",X"A2",X"01",X"01",X"21",X"CC",X"A8",
		X"50",X"40",X"8B",X"A9",X"84",X"14",X"8A",X"CC",X"11",X"59",X"2C",X"0A",X"08",X"30",X"4B",X"1B",
		X"4B",X"8B",X"14",X"52",X"BB",X"A0",X"51",X"00",X"FA",X"81",X"34",X"80",X"D9",X"A2",X"83",X"20",
		X"89",X"A3",X"C8",X"90",X"52",X"B9",X"10",X"51",X"99",X"DA",X"C8",X"37",X"20",X"D9",X"90",X"21",
		X"00",X"98",X"20",X"0D",X"A8",X"43",X"0B",X"B2",X"07",X"1A",X"AB",X"B9",X"14",X"72",X"0C",X"C9",
		X"01",X"31",X"91",X"92",X"08",X"BC",X"03",X"69",X"B9",X"32",X"7A",X"9A",X"89",X"8A",X"33",X"71",
		X"9E",X"98",X"02",X"10",X"00",X"10",X"BB",X"A4",X"44",X"AE",X"00",X"40",X"89",X"AB",X"81",X"02",
		X"23",X"9C",X"D9",X"03",X"83",X"A3",X"13",X"CA",X"D1",X"42",X"0C",X"C3",X"14",X"91",X"F0",X"91",
		X"81",X"93",X"01",X"DC",X"98",X"41",X"00",X"81",X"8C",X"A8",X"45",X"19",X"C9",X"13",X"38",X"CC",
		X"98",X"43",X"09",X"90",X"9A",X"E0",X"14",X"1B",X"18",X"38",X"E8",X"91",X"59",X"0A",X"02",X"38",
		X"1E",X"9B",X"96",X"11",X"89",X"0B",X"A9",X"07",X"81",X"90",X"11",X"AB",X"A0",X"71",X"A8",X"A2",
		X"20",X"2A",X"FA",X"93",X"50",X"1B",X"1B",X"0A",X"93",X"79",X"1D",X"81",X"48",X"1D",X"88",X"92",
		X"10",X"20",X"B0",X"1F",X"0B",X"30",X"78",X"0B",X"88",X"29",X"31",X"BA",X"F2",X"22",X"90",X"E3",
		X"C0",X"A1",X"16",X"B8",X"A1",X"11",X"A0",X"10",X"9E",X"DA",X"52",X"73",X"90",X"09",X"FC",X"03",
		X"48",X"08",X"0A",X"F8",X"80",X"83",X"18",X"8A",X"B0",X"08",X"04",X"72",X"80",X"8F",X"90",X"50",
		X"80",X"88",X"08",X"DA",X"18",X"85",X"02",X"88",X"08",X"F8",X"80",X"79",X"09",X"81",X"9A",X"08",
		X"42",X"90",X"19",X"18",X"9D",X"C0",X"33",X"A3",X"D2",X"02",X"9F",X"90",X"80",X"60",X"B8",X"90",
		X"80",X"08",X"08",X"72",X"80",X"BF",X"18",X"40",X"A3",X"88",X"08",X"F0",X"88",X"08",X"34",X"90",
		X"8F",X"08",X"04",X"88",X"08",X"A8",X"A1",X"87",X"08",X"0C",X"80",X"6A",X"2E",X"48",X"00",X"8D",
		X"00",X"21",X"9C",X"30",X"08",X"F1",X"00",X"2A",X"B2",X"90",X"27",X"90",X"8E",X"10",X"11",X"99",
		X"59",X"08",X"AB",X"18",X"51",X"91",X"89",X"2F",X"90",X"02",X"3F",X"08",X"03",X"08",X"0C",X"A1",
		X"05",X"8D",X"31",X"90",X"0F",X"18",X"85",X"98",X"18",X"08",X"E1",X"82",X"0D",X"18",X"01",X"39",
		X"08",X"F1",X"91",X"4B",X"84",X"90",X"8A",X"A1",X"86",X"0A",X"02",X"88",X"D8",X"00",X"1B",X"18",
		X"81",X"70",X"08",X"F0",X"00",X"39",X"A5",X"90",X"89",X"C1",X"86",X"9A",X"05",X"90",X"9C",X"18",
		X"00",X"88",X"00",X"78",X"08",X"D0",X"02",X"19",X"B7",X"90",X"89",X"C1",X"85",X"8C",X"14",X"90",
		X"AA",X"18",X"31",X"F1",X"91",X"49",X"08",X"D1",X"84",X"98",X"A5",X"90",X"0B",X"90",X"86",X"C3",
		X"19",X"08",X"D1",X"82",X"B1",X"90",X"07",X"80",X"8D",X"18",X"38",X"0D",X"5A",X"18",X"8D",X"18",
		X"80",X"13",X"80",X"8F",X"08",X"3C",X"4C",X"18",X"59",X"08",X"C1",X"85",X"90",X"80",X"80",X"88",
		X"F1",X"88",X"31",X"90",X"0F",X"08",X"04",X"9B",X"00",X"15",X"90",X"8C",X"80",X"32",X"90",X"80",
		X"9F",X"48",X"0D",X"00",X"80",X"38",X"19",X"8D",X"08",X"08",X"08",X"05",X"39",X"08",X"CD",X"14",
		X"19",X"18",X"8D",X"A1",X"07",X"8C",X"00",X"80",X"30",X"08",X"AE",X"18",X"19",X"50",X"80",X"80",
		X"9F",X"31",X"90",X"08",X"0F",X"08",X"48",X"8C",X"18",X"08",X"23",X"90",X"D9",X"02",X"2A",X"59",
		X"08",X"08",X"0F",X"49",X"00",X"80",X"8E",X"08",X"11",X"9A",X"18",X"08",X"37",X"9A",X"A0",X"06",
		X"08",X"88",X"18",X"08",X"08",X"08",X"EC",X"51",X"88",X"09",X"E1",X"88",X"08",X"08",X"08",X"00",
		X"58",X"0C",X"15",X"81",X"9A",X"81",X"04",X"90",X"80",X"80",X"80",X"BB",X"78",X"BF",X"08",X"08",
		X"01",X"A8",X"08",X"08",X"75",X"AA",X"A1",X"83",X"51",X"88",X"8A",X"04",X"90",X"08",X"88",X"D4",
		X"91",X"88",X"FA",X"91",X"85",X"98",X"B1",X"80",X"08",X"12",X"92",X"18",X"73",X"98",X"29",X"18",
		X"4A",X"9E",X"80",X"79",X"8B",X"10",X"39",X"8B",X"9F",X"08",X"35",X"9A",X"AA",X"20",X"3B",X"83",
		X"58",X"2E",X"11",X"92",X"91",X"0C",X"81",X"42",X"19",X"BE",X"AA",X"16",X"48",X"8B",X"89",X"2A",
		X"8B",X"52",X"3B",X"8F",X"0A",X"22",X"10",X"9F",X"00",X"13",X"29",X"C9",X"B0",X"14",X"60",X"8A",
		X"C0",X"02",X"81",X"19",X"98",X"99",X"91",X"44",X"A9",X"BB",X"88",X"53",X"2A",X"8D",X"AB",X"14",
		X"70",X"8B",X"80",X"21",X"89",X"90",X"80",X"8A",X"B7",X"23",X"B9",X"B9",X"E0",X"05",X"15",X"99",
		X"CA",X"83",X"60",X"0B",X"09",X"28",X"8E",X"00",X"32",X"AB",X"B1",X"13",X"0A",X"8A",X"78",X"1B",
		X"0B",X"49",X"29",X"38",X"19",X"B2",X"52",X"0C",X"FC",X"30",X"69",X"8B",X"90",X"43",X"0C",X"AA",
		X"52",X"A8",X"A1",X"28",X"39",X"9C",X"A1",X"30",X"23",X"29",X"FF",X"01",X"20",X"98",X"A8",X"29",
		X"28",X"84",X"79",X"AB",X"B3",X"26",X"1A",X"A8",X"80",X"80",X"12",X"2D",X"CA",X"31",X"39",X"C9",
		X"B0",X"22",X"70",X"20",X"0F",X"8B",X"32",X"59",X"88",X"00",X"8C",X"A9",X"21",X"22",X"08",X"AC",
		X"C9",X"91",X"94",X"87",X"04",X"98",X"D9",X"92",X"38",X"03",X"30",X"2D",X"AF",X"88",X"83",X"42",
		X"09",X"E9",X"A8",X"20",X"82",X"33",X"4E",X"9B",X"01",X"39",X"88",X"44",X"1A",X"BB",X"A0",X"92",
		X"15",X"42",X"9B",X"E8",X"A2",X"91",X"B6",X"13",X"8C",X"A8",X"09",X"00",X"22",X"11",X"33",X"D3",
		X"F8",X"CA",X"15",X"11",X"2D",X"0B",X"89",X"49",X"39",X"39",X"8C",X"12",X"90",X"F9",X"32",X"29",
		X"90",X"28",X"0F",X"99",X"86",X"11",X"8A",X"B9",X"A2",X"07",X"00",X"A1",X"90",X"29",X"BC",X"B7",
		X"03",X"B2",X"E2",X"80",X"1A",X"9B",X"35",X"18",X"0B",X"B0",X"93",X"27",X"B9",X"A2",X"35",X"99",
		X"D8",X"02",X"89",X"1A",X"12",X"07",X"AC",X"9A",X"42",X"90",X"89",X"29",X"87",X"8A",X"0B",X"24",
		X"00",X"11",X"C3",X"D9",X"83",X"04",X"88",X"1B",X"0F",X"80",X"1D",X"89",X"B3",X"C5",X"08",X"99",
		X"A2",X"83",X"29",X"FF",X"51",X"17",X"08",X"08",X"EE",X"10",X"59",X"19",X"18",X"8E",X"08",X"08",
		X"30",X"09",X"3A",X"BC",X"18",X"52",X"89",X"90",X"2A",X"8A",X"83",X"40",X"8C",X"83",X"22",X"CE",
		X"98",X"10",X"08",X"18",X"98",X"C8",X"42",X"08",X"A2",X"21",X"10",X"81",X"5A",X"1E",X"88",X"88",
		X"2B",X"99",X"29",X"4C",X"19",X"9C",X"B0",X"07",X"32",X"9A",X"90",X"85",X"C1",X"02",X"58",X"88",
		X"94",X"7E",X"9D",X"11",X"3B",X"24",X"29",X"18",X"FD",X"00",X"48",X"1A",X"49",X"0A",X"F1",X"80",
		X"22",X"B9",X"28",X"B8",X"81",X"54",X"F8",X"31",X"90",X"AC",X"18",X"68",X"B5",X"90",X"08",X"D0",
		X"00",X"20",X"08",X"0B",X"C0",X"08",X"52",X"B9",X"A1",X"60",X"88",X"C2",X"B8",X"27",X"90",X"0E",
		X"00",X"20",X"0B",X"59",X"00",X"9E",X"18",X"08",X"21",X"08",X"1E",X"80",X"01",X"2E",X"08",X"01",
		X"59",X"08",X"C8",X"02",X"39",X"80",X"08",X"0D",X"D1",X"82",X"5A",X"80",X"28",X"BD",X"18",X"42",
		X"AD",X"00",X"80",X"07",X"80",X"8A",X"B1",X"84",X"28",X"80",X"80",X"8F",X"90",X"81",X"68",X"08",
		X"09",X"F1",X"81",X"28",X"D0",X"08",X"08",X"07",X"90",X"0A",X"B1",X"87",X"88",X"08",X"08",X"0F",
		X"18",X"82",X"3A",X"18",X"8B",X"C0",X"80",X"68",X"C1",X"88",X"08",X"70",X"80",X"8E",X"18",X"13",
		X"90",X"80",X"80",X"F8",X"08",X"06",X"88",X"08",X"0D",X"80",X"01",X"3E",X"08",X"08",X"00",X"69",
		X"08",X"B8",X"08",X"60",X"80",X"88",X"08",X"F0",X"80",X"31",X"91",X"88",X"F0",X"80",X"48",X"C0",
		X"08",X"08",X"16",X"90",X"8D",X"00",X"02",X"18",X"08",X"08",X"8F",X"09",X"07",X"90",X"80",X"8A",
		X"B2",X"92",X"7D",X"00",X"80",X"13",X"80",X"88",X"F0",X"80",X"58",X"80",X"80",X"8C",X"90",X"80",
		X"60",X"80",X"8A",X"C1",X"84",X"9A",X"80",X"08",X"17",X"00",X"80",X"F0",X"84",X"80",X"80",X"80",
		X"89",X"F1",X"88",X"01",X"30",X"B4",X"98",X"A9",X"B1",X"80",X"80",X"74",X"90",X"08",X"0F",X"88",
		X"41",X"90",X"80",X"8F",X"09",X"18",X"19",X"00",X"68",X"19",X"0A",X"B9",X"18",X"82",X"71",X"80",
		X"80",X"80",X"CF",X"10",X"59",X"08",X"08",X"E0",X"08",X"00",X"88",X"80",X"36",X"90",X"9C",X"80",
		X"82",X"68",X"80",X"80",X"80",X"80",X"F9",X"24",X"90",X"80",X"0F",X"80",X"82",X"A8",X"08",X"01",
		X"70",X"8A",X"B0",X"00",X"70",X"88",X"00",X"88",X"08",X"08",X"8F",X"95",X"08",X"08",X"8F",X"00",
		X"80",X"18",X"A0",X"08",X"04",X"28",X"E8",X"00",X"60",X"88",X"08",X"91",X"80",X"08",X"00",X"80",
		X"8D",X"1F",X"3B",X"4D",X"09",X"00",X"80",X"09",X"00",X"80",X"82",X"71",X"8D",X"21",X"28",X"0C",
		X"93",X"02",X"90",X"B4",X"F2",X"82",X"99",X"C1",X"28",X"1F",X"98",X"00",X"7C",X"19",X"08",X"00",
		X"00",X"03",X"A8",X"90",X"61",X"89",X"89",X"28",X"81",X"B0",X"18",X"2B",X"F1",X"93",X"04",X"92",
		X"FB",X"91",X"28",X"88",X"7B",X"A8",X"84",X"19",X"88",X"82",X"58",X"1A",X"18",X"88",X"A3",X"23",
		X"3F",X"A8",X"35",X"B1",X"D9",X"82",X"01",X"96",X"98",X"B8",X"B2",X"A4",X"80",X"30",X"F9",X"B5",
		X"81",X"94",X"B1",X"A1",X"11",X"20",X"06",X"C8",X"9B",X"68",X"01",X"89",X"2C",X"94",X"B3",X"9C",
		X"21",X"95",X"B1",X"9C",X"12",X"81",X"C9",X"10",X"20",X"D2",X"7A",X"0A",X"A0",X"18",X"51",X"01",
		X"C8",X"9A",X"50",X"80",X"A8",X"20",X"3A",X"D2",X"80",X"B1",X"B4",X"B4",X"14",X"01",X"DA",X"C0",
		X"04",X"93",X"C3",X"9A",X"02",X"89",X"E0",X"01",X"29",X"11",X"A8",X"05",X"9A",X"90",X"68",X"AB",
		X"45",X"39",X"BE",X"80",X"20",X"09",X"28",X"00",X"F8",X"83",X"18",X"E8",X"82",X"19",X"A2",X"13",
		X"E8",X"91",X"82",X"31",X"03",X"AD",X"BA",X"60",X"59",X"8A",X"88",X"49",X"1C",X"09",X"1A",X"29",
		X"2E",X"01",X"42",X"9D",X"98",X"21",X"1C",X"10",X"50",X"A9",X"A9",X"13",X"1A",X"6A",X"2B",X"2A",
		X"3C",X"0F",X"2A",X"12",X"0A",X"29",X"5C",X"0B",X"58",X"2B",X"90",X"29",X"52",X"C8",X"B1",X"11",
		X"E3",X"83",X"09",X"A0",X"B0",X"A9",X"09",X"28",X"34",X"8C",X"B8",X"23",X"B2",X"23",X"B3",X"95",
		X"2C",X"7A",X"2E",X"09",X"00",X"70",X"1A",X"9A",X"B9",X"34",X"00",X"A9",X"09",X"8C",X"86",X"03",
		X"0F",X"0A",X"22",X"01",X"89",X"80",X"0C",X"A2",X"36",X"A5",X"98",X"AD",X"18",X"10",X"2B",X"1C",
		X"49",X"2D",X"29",X"2A",X"A8",X"96",X"22",X"C9",X"90",X"58",X"8A",X"A2",X"18",X"51",X"A2",X"A9",
		X"BC",X"B8",X"73",X"19",X"AD",X"22",X"11",X"DB",X"01",X"32",X"22",X"9F",X"C8",X"03",X"B3",X"B2",
		X"A3",X"91",X"B1",X"C3",X"B1",X"E3",X"17",X"89",X"B3",X"30",X"0B",X"04",X"74",X"18",X"8D",X"BA",
		X"98",X"1A",X"4A",X"C8",X"99",X"AB",X"22",X"43",X"9D",X"E8",X"73",X"2C",X"87",X"11",X"8B",X"F9",
		X"87",X"00",X"91",X"90",X"E8",X"08",X"03",X"18",X"81",X"89",X"F8",X"00",X"50",X"09",X"88",X"0A",
		X"A9",X"14",X"21",X"9A",X"00",X"8A",X"BA",X"36",X"30",X"AB",X"08",X"1A",X"B9",X"23",X"58",X"AB",
		X"01",X"3E",X"09",X"43",X"09",X"AD",X"08",X"40",X"88",X"08",X"0A",X"AC",X"30",X"69",X"0C",X"28",
		X"2B",X"18",X"39",X"91",X"40",X"0A",X"AD",X"03",X"09",X"D1",X"13",X"5A",X"A9",X"E0",X"03",X"80",
		X"86",X"90",X"A0",X"8A",X"8D",X"24",X"A2",X"03",X"20",X"FA",X"B5",X"11",X"8B",X"A7",X"0F",X"9C",
		X"71",X"89",X"98",X"10",X"02",X"C6",X"9A",X"BA",X"14",X"70",X"08",X"8B",X"E1",X"81",X"58",X"08",
		X"0A",X"BA",X"03",X"7C",X"1B",X"12",X"4A",X"0E",X"10",X"09",X"88",X"06",X"08",X"0D",X"80",X"30",
		X"1D",X"49",X"08",X"0E",X"18",X"01",X"1B",X"59",X"08",X"C0",X"08",X"58",X"8A",X"0A",X"2A",X"00",
		X"07",X"80",X"8E",X"18",X"21",X"A8",X"49",X"08",X"AC",X"18",X"13",X"01",X"08",X"0F",X"98",X"87",
		X"08",X"8D",X"18",X"80",X"40",X"80",X"9E",X"18",X"31",X"90",X"08",X"80",X"F8",X"08",X"03",X"29",
		X"18",X"CD",X"18",X"07",X"80",X"C8",X"00",X"83",X"29",X"08",X"F0",X"80",X"48",X"08",X"08",X"0C",
		X"B2",X"90",X"17",X"80",X"89",X"D1",X"80",X"69",X"0C",X"18",X"80",X"05",X"90",X"0B",X"A1",X"82",
		X"69",X"08",X"08",X"0F",X"08",X"00",X"59",X"08",X"C0",X"80",X"06",X"90",X"C0",X"08",X"08",X"68",
		X"80",X"9B",X"18",X"24",X"90",X"80",X"80",X"F8",X"80",X"50",X"88",X"8B",X"90",X"80",X"70",X"8E",
		X"18",X"08",X"11",X"29",X"08",X"F0",X"80",X"58",X"80",X"80",X"8C",X"80",X"87",X"88",X"0A",X"A2",
		X"A1",X"07",X"99",X"A1",X"80",X"12",X"D6",X"90",X"0C",X"00",X"84",X"88",X"08",X"08",X"C8",X"08",
		X"50",X"80",X"C9",X"19",X"51",X"9B",X"91",X"88",X"17",X"09",X"18",X"08",X"9F",X"08",X"58",X"08",
		X"08",X"E1",X"80",X"20",X"B9",X"19",X"07",X"80",X"8D",X"18",X"00",X"49",X"0A",X"84",X"88",X"08",
		X"D8",X"04",X"08",X"08",X"0E",X"80",X"87",X"9A",X"08",X"08",X"32",X"99",X"D1",X"88",X"50",X"89",
		X"91",X"39",X"08",X"00",X"FA",X"06",X"08",X"80",X"AC",X"18",X"33",X"CC",X"18",X"08",X"78",X"0C",
		X"00",X"82",X"29",X"1A",X"B8",X"51",X"80",X"80",X"80",X"DD",X"23",X"08",X"08",X"F8",X"80",X"03",
		X"C0",X"80",X"80",X"07",X"98",X"A8",X"25",X"08",X"08",X"B0",X"13",X"90",X"88",X"08",X"08",X"0E",
		X"BF",X"16",X"80",X"8F",X"00",X"80",X"81",X"89",X"00",X"80",X"68",X"0C",X"81",X"13",X"19",X"08",
		X"E3",X"89",X"38",X"89",X"F1",X"03",X"91",X"E1",X"A4",X"A3",X"D1",X"A0",X"80",X"05",X"98",X"A9",
		X"18",X"13",X"1C",X"19",X"38",X"89",X"23",X"2C",X"A8",X"61",X"9A",X"A7",X"A2",X"A2",X"C9",X"B3",
		X"32",X"11",X"A0",X"FD",X"81",X"50",X"88",X"C8",X"00",X"20",X"98",X"B1",X"69",X"09",X"12",X"10",
		X"8D",X"19",X"3A",X"80",X"24",X"01",X"F9",X"91",X"83",X"93",X"D2",X"B3",X"A1",X"82",X"C0",X"F1",
		X"00",X"00",X"B5",X"02",X"0F",X"99",X"03",X"09",X"12",X"31",X"CC",X"AA",X"25",X"30",X"AB",X"11",
		X"28",X"A9",X"8B",X"32",X"8E",X"95",X"35",X"AA",X"B9",X"A2",X"94",X"04",X"A1",X"A1",X"BB",X"88",
		X"33",X"B8",X"DC",X"38",X"76",X"0B",X"9B",X"10",X"B4",X"34",X"5A",X"9B",X"C0",X"22",X"08",X"A3",
		X"82",X"8A",X"F2",X"B2",X"A0",X"14",X"BA",X"E1",X"44",X"0A",X"D8",X"91",X"12",X"13",X"29",X"DE",
		X"80",X"30",X"3B",X"89",X"11",X"2F",X"09",X"00",X"11",X"1C",X"AB",X"36",X"20",X"9E",X"98",X"20",
		X"29",X"20",X"2C",X"99",X"09",X"58",X"00",X"39",X"0E",X"89",X"20",X"0D",X"90",X"20",X"00",X"6A",
		X"1C",X"09",X"10",X"21",X"B2",X"05",X"1B",X"E9",X"B3",X"13",X"36",X"88",X"F8",X"93",X"02",X"B0",
		X"C1",X"C1",X"86",X"02",X"B9",X"C1",X"11",X"09",X"A4",X"31",X"9E",X"0A",X"19",X"20",X"30",X"28",
		X"8E",X"89",X"8A",X"13",X"49",X"DC",X"83",X"40",X"A0",X"93",X"BA",X"C3",X"17",X"48",X"C9",X"92",
		X"81",X"90",X"12",X"02",X"C9",X"BA",X"39",X"06",X"09",X"8D",X"28",X"5C",X"29",X"82",X"D9",X"01",
		X"60",X"89",X"98",X"19",X"09",X"82",X"58",X"81",X"0C",X"8E",X"91",X"42",X"8A",X"C8",X"24",X"18",
		X"C1",X"A1",X"B5",X"91",X"11",X"BB",X"93",X"80",X"4D",X"5B",X"19",X"19",X"38",X"4B",X"B4",X"B8",
		X"D3",X"03",X"B6",X"99",X"89",X"0A",X"04",X"93",X"08",X"83",X"9F",X"09",X"31",X"69",X"1F",X"0A",
		X"49",X"1A",X"82",X"90",X"9A",X"01",X"39",X"7A",X"08",X"2B",X"28",X"6A",X"8D",X"39",X"5B",X"8A",
		X"31",X"39",X"AF",X"98",X"70",X"1B",X"92",X"98",X"A8",X"12",X"59",X"9B",X"84",X"01",X"91",X"B4",
		X"B1",X"41",X"11",X"B1",X"71",X"8D",X"D9",X"82",X"2A",X"9A",X"08",X"9C",X"B2",X"17",X"09",X"99",
		X"CD",X"47",X"10",X"78",X"08",X"0F",X"B0",X"36",X"90",X"80",X"AB",X"A1",X"90",X"47",X"91",X"A1",
		X"C8",X"91",X"87",X"08",X"08",X"A0",X"9A",X"80",X"53",X"80",X"AC",X"09",X"08",X"02",X"51",X"0B",
		X"C9",X"00",X"10",X"20",X"2A",X"AD",X"90",X"21",X"10",X"20",X"1B",X"EA",X"84",X"02",X"01",X"89",
		X"9F",X"90",X"14",X"0A",X"88",X"10",X"0B",X"8B",X"71",X"2D",X"09",X"31",X"0B",X"0A",X"08",X"1A",
		X"31",X"50",X"CA",X"9A",X"4D",X"48",X"11",X"A9",X"81",X"83",X"90",X"E0",X"21",X"AA",X"27",X"80",
		X"8C",X"A2",X"01",X"B6",X"B3",X"B3",X"B7",X"A9",X"FA",X"44",X"81",X"B0",X"71",X"FA",X"08",X"53",
		X"A1",X"88",X"0C",X"E1",X"82",X"59",X"09",X"A9",X"90",X"08",X"17",X"00",X"0D",X"90",X"80",X"16",
		X"80",X"9C",X"08",X"12",X"B9",X"71",X"90",X"C9",X"18",X"41",X"91",X"80",X"8A",X"F0",X"85",X"08",
		X"92",X"91",X"BD",X"18",X"07",X"90",X"C1",X"81",X"A1",X"88",X"07",X"88",X"0D",X"18",X"03",X"88",
		X"08",X"08",X"E8",X"08",X"68",X"80",X"08",X"0E",X"00",X"84",X"88",X"0D",X"18",X"80",X"80",X"40",
		X"80",X"AD",X"18",X"16",X"90",X"80",X"88",X"E1",X"80",X"59",X"08",X"08",X"8E",X"18",X"04",X"90",
		X"9B",X"18",X"08",X"00",X"61",X"90",X"8F",X"19",X"05",X"88",X"08",X"09",X"D1",X"80",X"48",X"08",
		X"08",X"C9",X"08",X"43",X"90",X"F8",X"08",X"01",X"98",X"27",X"90",X"9C",X"18",X"40",X"80",X"80",
		X"8A",X"E1",X"80",X"69",X"00",X"89",X"C1",X"80",X"79",X"0A",X"91",X"88",X"21",X"C0",X"87",X"88",
		X"0D",X"18",X"38",X"80",X"08",X"08",X"F0",X"80",X"59",X"00",X"8D",X"18",X"03",X"09",X"0F",X"18",
		X"01",X"29",X"D1",X"84",X"88",X"0D",X"18",X"38",X"80",X"80",X"0D",X"90",X"80",X"78",X"08",X"D1",
		X"80",X"12",X"91",X"E0",X"80",X"30",X"88",X"E1",X"83",X"08",X"08",X"F2",X"82",X"88",X"08",X"08",
		X"F0",X"80",X"22",X"D2",X"B0",X"80",X"25",X"99",X"C1",X"81",X"11",X"08",X"BA",X"04",X"A0",X"4F",
		X"69",X"08",X"B1",X"03",X"88",X"08",X"F0",X"80",X"58",X"9B",X"18",X"00",X"69",X"0C",X"00",X"82",
		X"39",X"0A",X"B9",X"70",X"80",X"80",X"08",X"88",X"F0",X"49",X"18",X"80",X"F0",X"08",X"10",X"B1",
		X"80",X"82",X"40",X"E8",X"08",X"34",X"90",X"89",X"9A",X"24",X"08",X"0D",X"85",X"90",X"09",X"F1",
		X"20",X"80",X"BB",X"08",X"00",X"17",X"B9",X"08",X"00",X"30",X"8D",X"83",X"61",X"88",X"D0",X"02",
		X"08",X"10",X"89",X"F9",X"13",X"10",X"8A",X"8F",X"19",X"21",X"11",X"A9",X"F8",X"80",X"31",X"AC",
		X"00",X"41",X"2E",X"88",X"01",X"21",X"39",X"8A",X"F8",X"12",X"49",X"0B",X"D1",X"39",X"8A",X"97",
		X"00",X"98",X"99",X"A0",X"50",X"3A",X"A8",X"98",X"C3",X"18",X"9C",X"A7",X"28",X"9E",X"11",X"11",
		X"98",X"2A",X"18",X"C0",X"01",X"53",X"C2",X"E0",X"A0",X"05",X"81",X"A9",X"00",X"98",X"19",X"1A",
		X"25",X"98",X"AE",X"19",X"13",X"94",X"9B",X"1A",X"8B",X"97",X"48",X"1C",X"09",X"90",X"20",X"68",
		X"00",X"BA",X"09",X"38",X"09",X"79",X"2C",X"AA",X"81",X"62",X"80",X"9B",X"0D",X"81",X"04",X"12",
		X"8D",X"AB",X"83",X"25",X"01",X"98",X"D8",X"A2",X"13",X"02",X"F3",X"A2",X"BA",X"E1",X"05",X"20",
		X"0B",X"CA",X"A2",X"42",X"39",X"0A",X"BD",X"99",X"34",X"41",X"8A",X"BA",X"80",X"3A",X"38",X"72",
		X"8C",X"BD",X"82",X"23",X"10",X"8A",X"CB",X"82",X"31",X"10",X"43",X"AE",X"EA",X"83",X"63",X"0B",
		X"D9",X"82",X"38",X"09",X"02",X"10",X"FA",X"A2",X"34",X"0A",X"B9",X"12",X"A3",X"A3",X"09",X"B5",
		X"A2",X"BC",X"A4",X"37",X"0A",X"CB",X"02",X"40",X"09",X"32",X"9D",X"D9",X"14",X"22",X"CB",X"B0",
		X"43",X"93",X"F0",X"80",X"01",X"91",X"8A",X"03",X"05",X"A9",X"D8",X"01",X"11",X"88",X"10",X"88",
		X"FA",X"83",X"72",X"AB",X"B9",X"32",X"12",X"A2",X"8C",X"98",X"A1",X"07",X"31",X"C9",X"9A",X"08",
		X"48",X"49",X"B2",X"41",X"AF",X"A8",X"36",X"00",X"B9",X"C2",X"02",X"A0",X"15",X"88",X"C9",X"91",
		X"15",X"10",X"8A",X"CA",X"93",X"23",X"0A",X"2F",X"29",X"81",X"8B",X"03",X"73",X"B0",X"F0",X"88",
		X"A3",X"97",X"18",X"9C",X"98",X"13",X"30",X"AA",X"91",X"8B",X"00",X"01",X"59",X"3C",X"1B",X"1E",
		X"88",X"61",X"2A",X"A8",X"90",X"E2",X"05",X"01",X"AA",X"BB",X"13",X"53",X"9A",X"8B",X"49",X"AC",
		X"02",X"40",X"0D",X"90",X"19",X"3B",X"43",X"21",X"D8",X"D1",X"90",X"05",X"40",X"AB",X"CA",X"02",
		X"44",X"8A",X"1B",X"1A",X"2C",X"98",X"71",X"0A",X"9B",X"8A",X"30",X"54",X"90",X"C1",X"D2",X"A5",
		X"95",X"88",X"A8",X"90",X"82",X"A3",X"82",X"88",X"E8",X"B2",X"04",X"40",X"0D",X"89",X"B2",X"20",
		X"51",X"91",X"BC",X"AC",X"61",X"81",X"A1",X"99",X"A8",X"86",X"82",X"9A",X"91",X"84",X"C0",X"02",
		X"39",X"2A",X"EA",X"39",X"68",X"29",X"2C",X"8E",X"03",X"11",X"99",X"0B",X"C8",X"01",X"49",X"01",
		X"90",X"FB",X"04",X"01",X"00",X"88",X"99",X"0B",X"24",X"77",X"23",X"FA",X"B0",X"86",X"82",X"90",
		X"BA",X"C0",X"04",X"11",X"08",X"90",X"AA",X"11",X"44",X"09",X"9A",X"02",X"9A",X"0B",X"23",X"25",
		X"BB",X"F9",X"03",X"11",X"A6",X"A0",X"DA",X"12",X"48",X"3C",X"0A",X"99",X"20",X"4A",X"19",X"A2",
		X"B0",X"71",X"99",X"F8",X"12",X"39",X"89",X"B2",X"92",X"02",X"19",X"CA",X"A4",X"44",X"99",X"B9",
		X"C2",X"32",X"0A",X"F2",X"E1",X"11",X"30",X"CA",X"80",X"11",X"91",X"E2",X"38",X"BA",X"88",X"79",
		X"1B",X"16",X"99",X"90",X"23",X"89",X"9C",X"01",X"07",X"B9",X"08",X"79",X"80",X"A0",X"0A",X"40",
		X"79",X"AB",X"C3",X"23",X"0C",X"9C",X"81",X"42",X"F5",X"E3",X"88",X"D4",X"03",X"90",X"DD",X"10",
		X"32",X"88",X"99",X"9D",X"08",X"06",X"29",X"0E",X"80",X"80",X"41",X"9A",X"9A",X"18",X"08",X"64",
		X"90",X"9F",X"19",X"58",X"08",X"08",X"88",X"E1",X"80",X"59",X"08",X"9B",X"4B",X"11",X"49",X"0D",
		X"80",X"04",X"89",X"0C",X"18",X"08",X"87",X"80",X"8C",X"00",X"05",X"90",X"80",X"80",X"D8",X"08",
		X"24",X"90",X"89",X"A9",X"90",X"87",X"29",X"0E",X"80",X"80",X"08",X"08",X"70",X"80",X"AC",X"18",
		X"68",X"08",X"08",X"0C",X"A1",X"81",X"79",X"00",X"B1",X"8C",X"29",X"25",X"90",X"AB",X"19",X"06",
		X"9A",X"08",X"78",X"08",X"AA",X"18",X"78",X"80",X"80",X"8C",X"80",X"83",X"4A",X"18",X"BB",X"08",
		X"03",X"78",X"0B",X"C1",X"82",X"79",X"A9",X"08",X"78",X"80",X"C0",X"01",X"28",X"08",X"80",X"8F",
		X"08",X"85",X"80",X"88",X"D1",X"80",X"30",X"80",X"F0",X"08",X"30",X"80",X"F1",X"88",X"48",X"80",
		X"D1",X"82",X"18",X"88",X"E1",X"10",X"B1",X"86",X"88",X"0B",X"91",X"86",X"88",X"0D",X"00",X"03",
		X"88",X"0E",X"00",X"49",X"00",X"88",X"BA",X"15",X"19",X"00",X"E8",X"02",X"10",X"80",X"AF",X"18",
		X"05",X"88",X"AA",X"18",X"25",X"9B",X"82",X"03",X"D8",X"01",X"12",X"AC",X"06",X"90",X"09",X"F1",
		X"03",X"90",X"8C",X"91",X"84",X"A9",X"80",X"80",X"60",X"89",X"B0",X"80",X"71",X"80",X"C9",X"23",
		X"08",X"88",X"CA",X"07",X"08",X"08",X"9F",X"01",X"20",X"80",X"8F",X"00",X"82",X"2D",X"80",X"80",
		X"18",X"1A",X"38",X"00",X"08",X"3B",X"28",X"83",X"9F",X"21",X"10",X"F9",X"08",X"10",X"86",X"08",
		X"8F",X"91",X"11",X"2B",X"2C",X"A8",X"00",X"09",X"11",X"A0",X"03",X"7B",X"3C",X"00",X"18",X"43",
		X"08",X"EA",X"01",X"32",X"B3",X"F1",X"B0",X"04",X"09",X"9D",X"85",X"84",X"AA",X"98",X"30",X"98",
		X"B2",X"4A",X"2C",X"1C",X"0B",X"40",X"49",X"00",X"B3",X"E1",X"11",X"20",X"A0",X"A2",X"2A",X"1F",
		X"82",X"50",X"BC",X"00",X"12",X"BA",X"A0",X"52",X"68",X"8E",X"99",X"20",X"22",X"89",X"89",X"BB",
		X"B1",X"55",X"01",X"A1",X"A9",X"C8",X"27",X"02",X"B9",X"A1",X"84",X"99",X"C1",X"17",X"18",X"AC",
		X"89",X"13",X"02",X"29",X"8C",X"E9",X"92",X"44",X"09",X"99",X"99",X"89",X"33",X"71",X"BA",X"C8",
		X"21",X"00",X"90",X"05",X"10",X"DA",X"98",X"31",X"22",X"48",X"DB",X"D8",X"12",X"52",X"9A",X"9A",
		X"09",X"10",X"41",X"4C",X"8B",X"00",X"3D",X"88",X"25",X"01",X"BA",X"AA",X"84",X"23",X"41",X"1F",
		X"D9",X"83",X"25",X"09",X"BC",X"00",X"31",X"80",X"89",X"1A",X"08",X"A8",X"8B",X"02",X"57",X"10",
		X"EA",X"90",X"33",X"81",X"20",X"AD",X"E9",X"23",X"23",X"99",X"F9",X"01",X"18",X"90",X"22",X"2D",
		X"B0",X"92",X"01",X"89",X"26",X"9A",X"9A",X"20",X"90",X"13",X"74",X"8F",X"B8",X"13",X"31",X"9D",
		X"98",X"22",X"9B",X"A2",X"63",X"1D",X"BA",X"15",X"1A",X"99",X"24",X"2B",X"D9",X"82",X"20",X"18",
		X"39",X"1F",X"AA",X"26",X"28",X"9D",X"90",X"22",X"1A",X"B9",X"33",X"2D",X"90",X"01",X"CA",X"86",
		X"42",X"9D",X"B9",X"13",X"38",X"08",X"88",X"8B",X"D9",X"37",X"19",X"B8",X"95",X"10",X"9D",X"90",
		X"23",X"29",X"CA",X"11",X"8A",X"1A",X"73",X"0B",X"E9",X"11",X"31",X"08",X"B1",X"AB",X"D0",X"46",
		X"0A",X"B9",X"14",X"1A",X"9B",X"13",X"32",X"FA",X"20",X"19",X"B2",X"15",X"1B",X"AE",X"92",X"13",
		X"59",X"A9",X"93",X"8C",X"01",X"17",X"B0",X"A9",X"12",X"4A",X"0D",X"3B",X"38",X"A9",X"23",X"93",
		X"96",X"C9",X"93",X"BA",X"A6",X"23",X"1E",X"C9",X"03",X"10",X"08",X"33",X"DC",X"90",X"42",X"88",
		X"C1",X"21",X"AC",X"A9",X"24",X"43",X"AB",X"D0",X"11",X"9A",X"B5",X"32",X"CD",X"80",X"28",X"89",
		X"08",X"40",X"3D",X"89",X"21",X"08",X"1A",X"70",X"51",X"0C",X"B8",X"31",X"DB",X"A4",X"50",X"9F",
		X"98",X"12",X"08",X"00",X"18",X"B9",X"34",X"05",X"98",X"A8",X"12",X"80",X"92",X"2B",X"8F",X"B0",
		X"22",X"AB",X"F0",X"94",X"99",X"9B",X"84",X"35",X"A8",X"13",X"03",X"E0",X"A2",X"31",X"28",X"89",
		X"AB",X"AE",X"41",X"29",X"EB",X"BA",X"35",X"29",X"B8",X"10",X"90",X"09",X"74",X"30",X"CB",X"02",
		X"50",X"99",X"D8",X"20",X"32",X"8B",X"F9",X"B0",X"84",X"13",X"BB",X"E8",X"12",X"20",X"91",X"52",
		X"28",X"B9",X"B9",X"83",X"73",X"B0",X"46",X"AE",X"F8",X"84",X"12",X"9A",X"A3",X"89",X"AF",X"01",
		X"51",X"0C",X"0B",X"28",X"21",X"28",X"1D",X"A7",X"00",X"9F",X"08",X"23",X"98",X"9B",X"08",X"99",
		X"30",X"71",X"8A",X"A9",X"28",X"82",X"87",X"18",X"AB",X"C2",X"27",X"AB",X"90",X"27",X"88",X"D0",
		X"01",X"00",X"93",X"00",X"9F",X"03",X"08",X"8D",X"82",X"21",X"AC",X"90",X"31",X"A9",X"83",X"78",
		X"AE",X"18",X"22",X"0B",X"99",X"00",X"5D",X"19",X"02",X"31",X"80",X"DE",X"18",X"79",X"00",X"80",
		X"8C",X"80",X"08",X"79",X"00",X"A9",X"08",X"08",X"17",X"90",X"80",X"D0",X"00",X"21",X"88",X"8B",
		X"B1",X"84",X"48",X"99",X"84",X"09",X"C1",X"03",X"80",X"F9",X"32",X"89",X"F8",X"00",X"5A",X"88",
		X"83",X"88",X"9A",X"84",X"82",X"8A",X"18",X"09",X"AA",X"78",X"19",X"D8",X"80",X"17",X"10",X"0E",
		X"A1",X"07",X"90",X"08",X"08",X"E0",X"08",X"14",X"90",X"9B",X"08",X"08",X"07",X"80",X"8E",X"18",
		X"59",X"08",X"99",X"00",X"88",X"09",X"07",X"08",X"09",X"D1",X"85",X"88",X"08",X"08",X"AC",X"18",
		X"07",X"88",X"0B",X"88",X"08",X"22",X"39",X"08",X"F9",X"05",X"08",X"0A",X"9A",X"09",X"00",X"82",
		X"71",X"08",X"0F",X"90",X"15",X"90",X"08",X"09",X"F1",X"88",X"31",X"80",X"BC",X"19",X"00",X"37",
		X"90",X"8F",X"18",X"21",X"90",X"9B",X"08",X"04",X"0B",X"95",X"3A",X"1B",X"F1",X"86",X"90",X"08",
		X"08",X"C8",X"08",X"07",X"90",X"8B",X"18",X"84",X"19",X"09",X"E1",X"83",X"18",X"0B",X"D1",X"05",
		X"80",X"C8",X"05",X"90",X"8D",X"18",X"22",X"90",X"AC",X"10",X"04",X"D0",X"38",X"00",X"E1",X"81",
		X"29",X"A2",X"C1",X"09",X"23",X"91",X"EB",X"22",X"21",X"E9",X"80",X"41",X"08",X"08",X"F8",X"84",
		X"19",X"00",X"CA",X"18",X"14",X"0A",X"AA",X"18",X"63",X"98",X"D9",X"00",X"40",X"09",X"90",X"80",
		X"30",X"0E",X"AA",X"22",X"43",X"90",X"C1",X"39",X"0F",X"D0",X"23",X"19",X"0E",X"A1",X"80",X"58",
		X"AA",X"00",X"06",X"18",X"B9",X"A1",X"06",X"18",X"A8",X"88",X"21",X"29",X"E9",X"03",X"31",X"AA",
		X"C9",X"20",X"49",X"81",X"A0",X"C1",X"13",X"CB",X"BA",X"07",X"83",X"CA",X"08",X"41",X"99",X"A1",
		X"43",X"08",X"B8",X"58",X"9A",X"B4",X"71",X"1C",X"B9",X"12",X"48",X"98",X"A8",X"A5",X"82",X"0D",
		X"89",X"18",X"21",X"89",X"A9",X"19",X"94",X"DA",X"03",X"15",X"8D",X"9A",X"62",X"8A",X"B8",X"53",
		X"18",X"D9",X"11",X"20",X"B2",X"92",X"0D",X"90",X"12",X"20",X"BF",X"B8",X"41",X"19",X"A8",X"31",
		X"CA",X"D0",X"43",X"38",X"FA",X"82",X"20",X"A9",X"83",X"4B",X"A8",X"06",X"0A",X"89",X"59",X"19",
		X"00",X"99",X"38",X"3B",X"1B",X"0D",X"1A",X"13",X"53",X"2F",X"D9",X"82",X"40",X"08",X"B0",X"91",
		X"A8",X"A7",X"15",X"AA",X"B8",X"14",X"01",X"09",X"E8",X"11",X"00",X"B1",X"10",X"69",X"1B",X"9E",
		X"81",X"33",X"4A",X"9F",X"91",X"21",X"00",X"B0",X"11",X"0A",X"CD",X"03",X"33",X"2A",X"BF",X"99",
		X"13",X"24",X"18",X"DA",X"B1",X"23",X"39",X"B9",X"C0",X"90",X"84",X"83",X"81",X"BA",X"09",X"00",
		X"41",X"6A",X"8D",X"A1",X"96",X"91",X"83",X"80",X"E9",X"00",X"23",X"00",X"4C",X"BC",X"03",X"38",
		X"2E",X"9A",X"84",X"30",X"BB",X"B0",X"45",X"2A",X"AE",X"11",X"21",X"9B",X"A0",X"52",X"99",X"B0",
		X"30",X"90",X"B2",X"24",X"D8",X"91",X"21",X"AA",X"96",X"08",X"AE",X"81",X"58",X"9A",X"08",X"22",
		X"8C",X"08",X"38",X"20",X"D9",X"05",X"28",X"BF",X"00",X"31",X"8C",X"80",X"21",X"9A",X"80",X"41",
		X"1D",X"09",X"10",X"2D",X"11",X"30",X"EA",X"93",X"34",X"AB",X"AB",X"15",X"28",X"BB",X"22",X"81",
		X"B8",X"C5",X"18",X"0A",X"02",X"19",X"AA",X"14",X"21",X"AC",X"0D",X"4A",X"3A",X"09",X"20",X"2B",
		X"D0",X"14",X"92",X"C1",X"A0",X"38",X"8B",X"12",X"08",X"0C",X"80",X"33",X"A9",X"91",X"28",X"A0",
		X"C3",X"23",X"98",X"C9",X"31",X"80",X"98",X"21",X"AE",X"10",X"10",X"11",X"AC",X"1A",X"38",X"40",
		X"8A",X"80",X"8B",X"19",X"43",X"92",X"BA",X"A8",X"81",X"12",X"29",X"0A",X"C1",X"83",X"2B",X"02",
		X"A4",X"A9",X"8B",X"02",X"28",X"91",X"91",X"A9",X"91",X"51",X"8A",X"D9",X"00",X"60",X"80",X"88",
		X"B9",X"82",X"30",X"2B",X"2A",X"18",X"C8",X"12",X"01",X"B2",X"00",X"B8",X"91",X"01",X"82",X"81",
		X"C8",X"B3",X"14",X"90",X"F1",X"A3",X"80",X"A1",X"30",X"0C",X"B9",X"33",X"32",X"AB",X"88",X"91",
		X"2A",X"A8",X"41",X"39",X"CB",X"A1",X"25",X"80",X"A8",X"88",X"B3",X"12",X"0A",X"AA",X"21",X"08",
		X"1D",X"20",X"19",X"A9",X"03",X"00",X"A2",X"89",X"09",X"2A",X"29",X"80",X"30",X"8C",X"80",X"02",
		X"0A",X"18",X"82",X"D8",X"12",X"11",X"B8",X"A0",X"13",X"98",X"91",X"29",X"9A",X"A3",X"13",X"A8",
		X"B1",X"00",X"19",X"09",X"A3",X"02",X"98",X"99",X"20",X"00",X"A1",X"81",X"8A",X"91",X"32",X"A0",
		X"B2",X"A1",X"92",X"D3",X"02",X"A9",X"99",X"12",X"09",X"01",X"98",X"A3",X"88",X"80",X"10",X"88",
		X"B0",X"95",X"81",X"A1",X"A0",X"B2",X"81",X"38",X"88",X"D3",X"A3",X"88",X"91",X"80",X"90",X"19",
		X"80",X"80",X"91",X"80",X"80",X"80",X"80",X"01",X"D8",X"12",X"34",X"52",X"13",X"77",X"20",X"11",
		X"47",X"50",X"CE",X"DB",X"01",X"13",X"43",X"8B",X"99",X"89",X"00",X"44",X"8D",X"B9",X"01",X"12",
		X"22",X"10",X"99",X"84",X"49",X"DC",X"BA",X"A8",X"13",X"33",X"42",X"0A",X"9A",X"37",X"61",X"8A",
		X"AB",X"BA",X"98",X"11",X"21",X"B1",X"76",X"08",X"89",X"AA",X"C9",X"14",X"29",X"C8",X"23",X"33",
		X"21",X"8A",X"83",X"8F",X"FE",X"80",X"13",X"21",X"99",X"AB",X"AB",X"C9",X"27",X"62",X"09",X"A8",
		X"90",X"80",X"10",X"00",X"89",X"99",X"9A",X"89",X"80",X"01",X"57",X"19",X"EB",X"81",X"18",X"00",
		X"08",X"01",X"0B",X"D8",X"47",X"33",X"32",X"9E",X"C9",X"08",X"AB",X"03",X"30",X"90",X"23",X"58",
		X"DA",X"99",X"80",X"02",X"12",X"00",X"08",X"99",X"98",X"90",X"02",X"77",X"50",X"BE",X"B0",X"11",
		X"01",X"08",X"CB",X"16",X"42",X"10",X"9A",X"AB",X"BB",X"99",X"B8",X"73",X"03",X"61",X"88",X"9E",
		X"A9",X"81",X"33",X"9B",X"A9",X"00",X"24",X"32",X"20",X"0A",X"AB",X"05",X"AF",X"D8",X"80",X"02",
		X"22",X"21",X"10",X"89",X"80",X"82",X"BF",X"AE",X"B0",X"54",X"09",X"CB",X"90",X"13",X"43",X"54",
		X"28",X"9C",X"DC",X"A8",X"21",X"18",X"01",X"25",X"31",X"8A",X"DD",X"A8",X"00",X"35",X"21",X"09",
		X"BB",X"AA",X"99",X"81",X"12",X"32",X"32",X"12",X"00",X"88",X"99",X"99",X"99",X"A8",X"98",X"90",
		X"98",X"88",X"89",X"9F",X"F1",X"32",X"DC",X"80",X"23",X"53",X"22",X"09",X"9B",X"DA",X"BB",X"AA",
		X"88",X"00",X"22",X"22",X"23",X"13",X"11",X"11",X"01",X"07",X"75",X"19",X"AC",X"BC",X"AA",X"88",
		X"22",X"43",X"33",X"2A",X"B3",X"2B",X"B1",X"53",X"44",X"21",X"8A",X"BD",X"DA",X"BB",X"BA",X"A8",
		X"88",X"11",X"13",X"23",X"32",X"46",X"76",X"08",X"9A",X"BC",X"9A",X"AB",X"A2",X"64",X"44",X"23",
		X"18",X"80",X"BD",X"BA",X"B9",X"98",X"80",X"01",X"12",X"42",X"20",X"BE",X"CC",X"AA",X"98",X"03",
		X"20",X"92",X"75",X"43",X"51",X"01",X"8A",X"DB",X"89",X"99",X"89",X"88",X"80",X"80",X"00",X"11",
		X"20",X"20",X"11",X"00",X"0C",X"FC",X"16",X"22",X"11",X"89",X"AD",X"CC",X"A0",X"26",X"42",X"11",
		X"99",X"BB",X"CA",X"AA",X"88",X"08",X"AA",X"25",X"53",X"53",X"21",X"18",X"8A",X"BB",X"CB",X"BA",
		X"B9",X"A8",X"80",X"10",X"21",X"21",X"20",X"21",X"11",X"28",X"20",X"10",X"00",X"11",X"32",X"76",
		X"19",X"BD",X"BA",X"EA",X"98",X"13",X"73",X"21",X"18",X"9A",X"AB",X"BA",X"A9",X"00",X"8A",X"36",
		X"41",X"19",X"AB",X"B9",X"37",X"22",X"12",X"20",X"82",X"9F",X"BB",X"AB",X"AA",X"91",X"29",X"17",
		X"61",X"09",X"AB",X"CA",X"BD",X"BA",X"45",X"20",X"45",X"21",X"8A",X"99",X"98",X"80",X"10",X"10",
		X"08",X"A0",X"42",X"AF",X"BD",X"CA",X"BA",X"99",X"B8",X"55",X"33",X"23",X"11",X"00",X"89",X"98",
		X"98",X"80",X"8B",X"FD",X"91",X"13",X"64",X"30",X"9A",X"BB",X"CA",X"9A",X"88",X"02",X"34",X"0D",
		X"DB",X"99",X"90",X"23",X"43",X"43",X"22",X"23",X"15",X"30",X"9A",X"FE",X"BA",X"98",X"11",X"44",
		X"21",X"33",X"1B",X"BA",X"BF",X"A9",X"89",X"98",X"8B",X"E9",X"02",X"64",X"22",X"20",X"89",X"AB",
		X"BB",X"A9",X"98",X"01",X"21",X"30",X"88",X"A8",X"02",X"71",X"35",X"21",X"89",X"BC",X"CA",X"BD",
		X"CA",X"98",X"23",X"43",X"43",X"31",X"10",X"89",X"9B",X"CB",X"AB",X"AA",X"A8",X"98",X"80",X"81",
		X"01",X"81",X"01",X"01",X"10",X"01",X"81",X"81",X"83",X"73",X"08",X"9B",X"FA",X"BA",X"BA",X"91",
		X"14",X"43",X"41",X"21",X"8A",X"83",X"01",X"81",X"98",X"99",X"A9",X"99",X"99",X"90",X"90",X"80",
		X"90",X"A9",X"00",X"13",X"23",X"01",X"80",X"AA",X"FB",X"03",X"33",X"33",X"AE",X"BA",X"80",X"13",
		X"53",X"43",X"41",X"AB",X"CA",X"BB",X"B9",X"98",X"80",X"81",X"80",X"81",X"80",X"81",X"81",X"81",
		X"82",X"46",X"0A",X"BA",X"88",X"AB",X"80",X"21",X"32",X"32",X"21",X"10",X"88",X"89",X"8A",X"99",
		X"8A",X"8A",X"89",X"88",X"09",X"08",X"08",X"00",X"13",X"62",X"08",X"9B",X"FC",X"B9",X"81",X"31",
		X"24",X"33",X"23",X"31",X"38",X"12",X"38",X"AC",X"CC",X"CB",X"AB",X"B9",X"99",X"10",X"31",X"32",
		X"39",X"9A",X"12",X"34",X"62",X"33",X"53",X"19",X"9B",X"CD",X"BA",X"CB",X"A8",X"00",X"11",X"9B",
		X"01",X"23",X"53",X"44",X"12",X"11",X"00",X"03",X"00",X"BB",X"DC",X"BC",X"AA",X"99",X"98",X"11",
		X"22",X"32",X"22",X"22",X"11",X"20",X"10",X"00",X"08",X"88",X"89",X"09",X"89",X"89",X"89",X"89",
		X"89",X"BD",X"99",X"23",X"23",X"13",X"12",X"35",X"12",X"9D",X"BC",X"BB",X"A8",X"02",X"35",X"10",
		X"13",X"29",X"BB",X"9A",X"00",X"41",X"09",X"11",X"32",X"28",X"8A",X"9A",X"BB",X"AA",X"8A",X"08",
		X"09",X"A9",X"02",X"54",X"42",X"10",X"9A",X"A9",X"A9",X"18",X"20",X"18",X"18",X"01",X"29",X"AE",
		X"A8",X"89",X"99",X"BB",X"91",X"09",X"91",X"12",X"24",X"33",X"44",X"32",X"18",X"9A",X"9A",X"AA",
		X"9A",X"00",X"29",X"0A",X"99",X"BA",X"9A",X"89",X"08",X"10",X"18",X"00",X"01",X"10",X"22",X"51",
		X"00",X"10",X"81",X"80",X"88",X"90",X"A8",X"99",X"A8",X"A8",X"A8",X"98",X"90",X"80",X"80",X"81",
		X"81",X"01",X"81",X"01",X"01",X"00",X"01",X"80",X"00",X"81",X"13",X"8A",X"A8",X"81",X"98",X"99",
		X"98",X"AA",X"BA",X"82",X"11",X"21",X"01",X"01",X"88",X"B9",X"91",X"02",X"25",X"33",X"11",X"0A",
		X"AA",X"BB",X"9B",X"9A",X"98",X"88",X"88",X"18",X"10",X"10",X"18",X"10",X"10",X"18",X"18",X"18",
		X"00",X"08",X"08",X"88",X"09",X"08",X"88",X"09",X"08",X"88",X"09",X"08",X"88",X"09",X"80",X"18",
		X"8A",X"09",X"10",X"21",X"21",X"20",X"10",X"08",X"89",X"89",X"88",X"99",X"09",X"89",X"88",X"88",
		X"08",X"08",X"08",X"00",X"00",X"08",X"10",X"00",X"08",X"18",X"18",X"08",X"08",X"08",X"10",X"10",
		X"08",X"09",X"9C",X"BB",X"9A",X"02",X"32",X"31",X"18",X"0B",X"A8",X"00",X"10",X"18",X"0A",X"9A",
		X"09",X"10",X"21",X"21",X"10",X"18",X"08",X"89",X"89",X"88",X"89",X"98",X"89",X"09",X"08",X"09",
		X"00",X"08",X"18",X"02",X"21",X"18",X"9A",X"AA",X"89",X"01",X"11",X"20",X"20",X"10",X"08",X"08",
		X"09",X"09",X"88",X"10",X"09",X"89",X"9B",X"99",X"99",X"89",X"89",X"01",X"21",X"31",X"10",X"10",
		X"08",X"10",X"08",X"08",X"08",X"88",X"08",X"09",X"08",X"09",X"08",X"09",X"08",X"88",X"08",X"08",
		X"81",X"A8",X"00",X"81",X"A2",X"B0",X"09",X"28",X"00",X"81",X"80",X"3A",X"A2",X"B3",X"B0",X"18",
		X"98",X"01",X"A2",X"89",X"92",X"92",X"A2",X"89",X"28",X"94",X"A8",X"89",X"91",X"09",X"11",X"90",
		X"84",X"89",X"80",X"0A",X"10",X"B1",X"88",X"80",X"02",X"88",X"1A",X"19",X"03",X"A9",X"18",X"09",
		X"29",X"A1",X"A1",X"93",X"88",X"A1",X"18",X"80",X"19",X"92",X"89",X"30",X"A8",X"A1",X"89",X"81",
		X"3A",X"82",X"4C",X"92",X"0C",X"27",X"DA",X"68",X"C1",X"49",X"80",X"88",X"98",X"15",X"1F",X"03",
		X"BC",X"52",X"BC",X"41",X"C8",X"58",X"C1",X"29",X"B4",X"2D",X"83",X"8C",X"24",X"BB",X"41",X"D0",
		X"49",X"B2",X"2B",X"96",X"8C",X"13",X"B9",X"40",X"D1",X"2A",X"94",X"8C",X"22",X"B9",X"69",X"B3",
		X"2D",X"04",X"AB",X"58",X"B2",X"3D",X"84",X"9A",X"30",X"E1",X"3B",X"84",X"9D",X"32",X"D1",X"3C",
		X"95",X"9B",X"40",X"D2",X"3C",X"84",X"AC",X"41",X"C2",X"2C",X"94",X"99",X"30",X"C0",X"08",X"11",
		X"98",X"A0",X"49",X"02",X"F8",X"5A",X"02",X"BC",X"41",X"B3",X"1D",X"93",X"1A",X"39",X"D8",X"22",
		X"08",X"8D",X"B6",X"2A",X"00",X"D0",X"59",X"92",X"BC",X"51",X"A1",X"8E",X"05",X"88",X"0B",X"A1",
		X"61",X"AA",X"09",X"87",X"1D",X"00",X"B4",X"5C",X"A1",X"A8",X"72",X"D9",X"09",X"37",X"BC",X"19",
		X"87",X"2D",X"B3",X"98",X"71",X"DB",X"48",X"03",X"BE",X"21",X"01",X"0E",X"82",X"94",X"2E",X"A5",
		X"A8",X"68",X"D0",X"11",X"8A",X"28",X"D3",X"3C",X"B1",X"79",X"B2",X"80",X"0F",X"35",X"DA",X"59",
		X"81",X"E3",X"5D",X"94",X"A0",X"2F",X"35",X"D8",X"5D",X"13",X"E8",X"50",X"A3",X"E0",X"5D",X"95",
		X"9C",X"5A",X"84",X"BB",X"63",X"D8",X"19",X"28",X"98",X"7D",X"85",X"C1",X"4D",X"95",X"0B",X"18",
		X"81",X"88",X"E6",X"2D",X"A5",X"99",X"2E",X"15",X"AC",X"5A",X"85",X"CA",X"42",X"B9",X"10",X"08",
		X"0F",X"15",X"BA",X"38",X"83",X"B8",X"07",X"D9",X"59",X"83",X"CA",X"32",X"1D",X"A3",X"3B",X"8A",
		X"C7",X"4D",X"B5",X"81",X"8F",X"05",X"3D",X"B3",X"20",X"9C",X"A6",X"00",X"BB",X"62",X"AA",X"89",
		X"34",X"2F",X"84",X"0C",X"08",X"91",X"26",X"D1",X"12",X"F0",X"09",X"49",X"A3",X"B1",X"5B",X"A4",
		X"0C",X"84",X"0C",X"12",X"A0",X"3A",X"E8",X"53",X"D5",X"D3",X"A8",X"B9",X"78",X"92",X"C9",X"60",
		X"C8",X"28",X"98",X"69",X"D3",X"4B",X"A2",X"19",X"B9",X"71",X"2E",X"4C",X"82",X"B0",X"5B",X"95",
		X"A9",X"49",X"A2",X"1A",X"98",X"35",X"CA",X"31",X"A1",X"8B",X"88",X"73",X"F9",X"58",X"B2",X"98",
		X"39",X"C4",X"1C",X"11",X"B1",X"3B",X"A0",X"87",X"3F",X"A5",X"1B",X"80",X"00",X"A2",X"3F",X"85",
		X"9B",X"20",X"A4",X"8D",X"14",X"AB",X"30",X"91",X"1C",X"01",X"C4",X"4D",X"A5",X"0C",X"11",X"91",
		X"A8",X"30",X"A0",X"88",X"49",X"C2",X"3D",X"92",X"4B",X"A4",X"0A",X"08",X"06",X"AD",X"13",X"0C",
		X"81",X"20",X"BA",X"33",X"B8",X"D0",X"70",X"C0",X"29",X"82",X"8A",X"1B",X"87",X"8B",X"31",X"B0",
		X"89",X"60",X"C8",X"13",X"8E",X"03",X"A9",X"30",X"B2",X"9F",X"35",X"BA",X"20",X"80",X"80",X"2C",
		X"90",X"97",X"2F",X"02",X"90",X"3B",X"B4",X"0E",X"25",X"CB",X"40",X"93",X"9E",X"21",X"90",X"81",
		X"0D",X"03",X"08",X"0E",X"84",X"09",X"90",X"08",X"84",X"0B",X"A8",X"33",X"19",X"FB",X"45",X"A8",
		X"0A",X"A7",X"0B",X"11",X"D0",X"4A",X"01",X"B9",X"51",X"A8",X"98",X"23",X"AC",X"20",X"B3",X"2B",
		X"12",X"F9",X"78",X"98",X"88",X"14",X"AD",X"22",X"88",X"C0",X"48",X"98",X"82",X"0C",X"11",X"A1",
		X"18",X"1E",X"85",X"8B",X"18",X"34",X"F9",X"5A",X"93",X"B9",X"79",X"B4",X"8C",X"59",X"D4",X"2D",
		X"12",X"D2",X"2B",X"12",X"D9",X"69",X"B2",X"19",X"3C",X"D5",X"1D",X"11",X"A1",X"4B",X"C3",X"2A",
		X"81",X"A0",X"7B",X"A5",X"8B",X"30",X"D3",X"1E",X"22",X"C1",X"2B",X"03",X"AC",X"34",X"C9",X"38",
		X"A3",X"0F",X"22",X"C1",X"0A",X"06",X"AD",X"42",X"C1",X"0A",X"14",X"AB",X"12",X"0B",X"10",X"A5",
		X"3F",X"A5",X"8A",X"19",X"04",X"9C",X"84",X"1B",X"80",X"01",X"1C",X"80",X"23",X"DA",X"03",X"4A",
		X"C0",X"84",X"3F",X"92",X"18",X"80",X"AD",X"62",X"DA",X"58",X"80",X"A8",X"49",X"88",X"92",X"2B",
		X"10",X"99",X"04",X"AB",X"33",X"F0",X"51",X"EB",X"53",X"CA",X"20",X"10",X"B9",X"38",X"10",X"C9",
		X"31",X"09",X"A2",X"C1",X"7A",X"D3",X"2A",X"92",X"19",X"F1",X"6B",X"B4",X"09",X"18",X"A3",X"0D",
		X"20",X"B1",X"28",X"A0",X"31",X"DB",X"51",X"A8",X"08",X"11",X"89",X"D2",X"7A",X"A2",X"09",X"19",
		X"83",X"0D",X"02",X"A9",X"69",X"C2",X"49",X"9A",X"97",X"1C",X"93",X"09",X"88",X"39",X"D4",X"0C",
		X"12",X"A8",X"2B",X"15",X"AC",X"31",X"98",X"90",X"10",X"88",X"1B",X"C7",X"1D",X"02",X"99",X"39",
		X"92",X"0B",X"11",X"90",X"09",X"28",X"E4",X"0C",X"12",X"B9",X"58",X"92",X"BB",X"71",X"AA",X"84",
		X"1C",X"82",X"80",X"1B",X"83",X"2B",X"E0",X"50",X"C1",X"1C",X"05",X"A8",X"3B",X"94",X"9A",X"38",
		X"92",X"BA",X"70",X"B1",X"88",X"3A",X"82",X"AC",X"68",X"95",X"AE",X"23",X"B8",X"3C",X"83",X"A0",
		X"39",X"8D",X"86",X"0A",X"81",X"A0",X"59",X"B5",X"8E",X"23",X"B9",X"2A",X"04",X"9A",X"18",X"91",
		X"01",X"0B",X"A1",X"07",X"1D",X"92",X"18",X"80",X"8D",X"04",X"08",X"8A",X"A2",X"52",X"BF",X"11",
		X"81",X"2E",X"93",X"0B",X"40",X"C1",X"09",X"22",X"CA",X"21",X"01",X"BD",X"25",X"A9",X"39",X"B2",
		X"88",X"68",X"D0",X"28",X"00",X"9C",X"34",X"B9",X"09",X"51",X"D0",X"18",X"09",X"94",X"8A",X"10",
		X"8A",X"06",X"0D",X"02",X"80",X"AC",X"61",X"D1",X"1A",X"12",X"F1",X"3B",X"83",X"C0",X"4A",X"A4",
		X"9A",X"49",X"91",X"09",X"11",X"C0",X"39",X"A1",X"A3",X"7D",X"82",X"88",X"19",X"A3",X"3C",X"91",
		X"08",X"18",X"E3",X"3E",X"83",X"9A",X"4A",X"A7",X"9A",X"38",X"A2",X"89",X"12",X"AC",X"32",X"B8",
		X"2C",X"07",X"AA",X"30",X"A2",X"0F",X"15",X"B9",X"38",X"92",X"9B",X"23",X"9A",X"93",X"09",X"1C",
		X"C7",X"2E",X"02",X"90",X"89",X"03",X"1D",X"93",X"09",X"09",X"A4",X"19",X"9B",X"43",X"9B",X"C2",
		X"59",X"1C",X"B7",X"1A",X"91",X"88",X"14",X"DB",X"61",X"B8",X"18",X"10",X"A0",X"00",X"1A",X"A4",
		X"99",X"21",X"8C",X"13",X"AA",X"40",X"F8",X"44",X"CB",X"33",X"B8",X"89",X"32",X"C0",X"89",X"41",
		X"B9",X"00",X"2A",X"21",X"F0",X"6A",X"A1",X"2A",X"90",X"78",X"E1",X"3A",X"92",X"98",X"3B",X"95",
		X"A9",X"48",X"A0",X"10",X"AA",X"35",X"BB",X"40",X"91",X"9A",X"11",X"49",X"F1",X"3A",X"91",X"91",
		X"2C",X"94",X"0A",X"11",X"C8",X"79",X"B0",X"30",X"2F",X"A5",X"1A",X"90",X"10",X"A8",X"5A",X"A5",
		X"8B",X"21",X"B2",X"1E",X"05",X"9A",X"10",X"08",X"88",X"81",X"80",X"4D",X"95",X"8A",X"02",X"B0",
		X"3B",X"83",X"8A",X"10",X"81",X"9A",X"7A",X"B5",X"0B",X"13",X"AB",X"38",X"87",X"BC",X"32",X"0B",
		X"B4",X"3B",X"90",X"93",X"2D",X"A1",X"70",X"C9",X"30",X"B3",X"3F",X"01",X"A1",X"3D",X"03",X"AA",
		X"3A",X"13",X"E8",X"38",X"80",X"B1",X"2A",X"06",X"BA",X"4D",X"07",X"8C",X"11",X"90",X"1A",X"10",
		X"B1",X"04",X"1E",X"93",X"0A",X"30",X"E8",X"4A",X"97",X"8C",X"11",X"91",X"0B",X"03",X"A0",X"19",
		X"89",X"02",X"29",X"8D",X"B7",X"19",X"90",X"08",X"84",X"0D",X"80",X"11",X"2B",X"BC",X"37",X"8A",
		X"08",X"B6",X"2C",X"82",X"AA",X"68",X"91",X"9A",X"33",X"B9",X"98",X"35",X"AD",X"22",X"C1",X"29",
		X"91",X"B9",X"70",X"A8",X"08",X"13",X"AF",X"12",X"81",X"C9",X"40",X"A0",X"81",X"2C",X"83",X"99",
		X"02",X"0E",X"96",X"8A",X"00",X"14",X"DA",X"68",X"A2",X"9A",X"68",X"D2",X"1A",X"20",X"D2",X"1B",
		X"12",X"B0",X"3B",X"82",X"AA",X"60",X"C1",X"18",X"08",X"E3",X"2C",X"01",X"90",X"3B",X"C3",X"2A",
		X"81",X"A8",X"6A",X"C4",X"1C",X"12",X"B1",X"3F",X"03",X"B8",X"3A",X"83",X"AB",X"35",X"BB",X"40",
		X"A3",X"0F",X"13",X"B9",X"3A",X"85",X"9E",X"22",X"B0",X"19",X"04",X"AB",X"12",X"1B",X"82",X"A3",
		X"4F",X"A7",X"8A",X"18",X"01",X"8B",X"95",X"1B",X"80",X"10",X"1B",X"A2",X"14",X"CB",X"23",X"3B",
		X"E1",X"83",X"4E",X"A3",X"2A",X"08",X"9D",X"53",X"E9",X"30",X"90",X"98",X"38",X"98",X"92",X"2B",
		X"02",X"B9",X"05",X"9B",X"23",X"C9",X"71",X"DB",X"45",X"BA",X"21",X"81",X"B9",X"38",X"01",X"CA",
		X"41",X"89",X"91",X"98",X"79",X"C1",X"49",X"A2",X"08",X"D0",X"79",X"B3",X"1A",X"00",X"A2",X"2E",
		X"11",X"B1",X"28",X"A8",X"31",X"CB",X"52",X"B9",X"18",X"21",X"A9",X"C1",X"79",X"B2",X"2A",X"18",
		X"B4",X"1D",X"83",X"8A",X"40",X"E1",X"39",X"AA",X"97",X"2D",X"93",X"19",X"98",X"20",X"D2",X"3E",
		X"02",X"99",X"29",X"95",X"9C",X"13",X"99",X"80",X"02",X"8A",X"19",X"C7",X"1D",X"02",X"8A",X"20",
		X"B2",X"1C",X"02",X"98",X"19",X"11",X"D2",X"3D",X"83",X"9B",X"23",X"C0",X"0C",X"53",X"CA",X"83",
		X"3C",X"A3",X"08",X"1B",X"93",X"3A",X"F9",X"60",X"A8",X"2A",X"A7",X"8A",X"3A",X"B6",X"8A",X"20",
		X"A1",X"99",X"41",X"C0",X"80",X"29",X"A3",X"8D",X"32",X"B6",X"AF",X"14",X"9A",X"29",X"93",X"98",
		X"39",X"8C",X"A7",X"2C",X"81",X"98",X"40",X"C2",X"1F",X"04",X"9A",X"18",X"84",X"9A",X"10",X"91",
		X"00",X"0A",X"A1",X"14",X"2F",X"91",X"29",X"80",X"0B",X"86",X"08",X"9A",X"93",X"41",X"BF",X"03",
		X"90",X"4D",X"A4",X"1A",X"11",X"D0",X"19",X"22",X"CA",X"21",X"01",X"BC",X"25",X"9B",X"30",X"C1",
		X"19",X"31",X"F8",X"20",X"88",X"8B",X"17",X"9A",X"19",X"33",X"F8",X"28",X"09",X"93",X"0B",X"02",
		X"8B",X"05",X"2F",X"83",X"98",X"0C",X"36",X"D8",X"3A",X"03",X"E8",X"59",X"A3",X"A9",X"59",X"A3",
		X"8B",X"48",X"A1",X"09",X"12",X"C9",X"58",X"A0",X"80",X"5B",X"B5",X"0A",X"18",X"A2",X"4B",X"A2",
		X"08",X"18",X"C2",X"6C",X"83",X"9A",X"4A",X"A7",X"9A",X"38",X"A2",X"8A",X"22",X"BC",X"34",X"B9",
		X"3B",X"87",X"9B",X"31",X"B2",X"0E",X"16",X"AA",X"38",X"91",X"8C",X"23",X"9A",X"82",X"0A",X"1A",
		X"B7",X"3F",X"83",X"98",X"0A",X"13",X"1E",X"93",X"19",X"98",X"94",X"19",X"AA",X"43",X"AC",X"A3",
		X"59",X"0C",X"A7",X"1B",X"92",X"80",X"13",X"FA",X"50",X"B0",X"18",X"10",X"B0",X"11",X"0B",X"94",
		X"99",X"21",X"9C",X"13",X"BA",X"58",X"C8",X"73",X"EA",X"32",X"A9",X"08",X"30",X"B0",X"89",X"41",
		X"C9",X"02",X"09",X"28",X"F1",X"5A",X"B3",X"1A",X"80",X"69",X"F2",X"2A",X"92",X"90",X"2B",X"95",
		X"A9",X"49",X"A1",X"18",X"A8",X"34",X"D9",X"30",X"90",X"99",X"21",X"3A",X"F1",X"4A",X"A2",X"90",
		X"2B",X"96",X"0B",X"02",X"C8",X"59",X"C2",X"20",X"1F",X"95",X"0A",X"91",X"01",X"A8",X"5A",X"B6",
		X"8A",X"10",X"91",X"0C",X"15",X"AA",X"11",X"08",X"98",X"01",X"81",X"3F",X"95",X"8B",X"12",X"B0",
		X"3A",X"A4",X"8A",X"18",X"81",X"A9",X"69",X"B5",X"0B",X"13",X"BA",X"38",X"85",X"DB",X"51",X"89",
		X"B4",X"2B",X"80",X"82",X"0A",X"B2",X"70",X"D9",X"30",X"B4",X"0D",X"12",X"B2",X"2D",X"03",X"B9",
		X"3A",X"13",X"F8",X"38",X"08",X"A0",X"2B",X"14",X"C9",X"3D",X"27",X"9D",X"12",X"A1",X"1B",X"01",
		X"A0",X"23",X"2F",X"B5",X"09",X"18",X"C0",X"4A",X"97",X"9C",X"21",X"91",X"8B",X"13",X"A0",X"19",
		X"98",X"03",X"2B",X"9E",X"97",X"1A",X"A1",X"19",X"03",X"8F",X"00",X"11",X"0A",X"B8",X"54",X"9C",
		X"08",X"A6",X"1B",X"93",X"B8",X"78",X"90",X"9A",X"42",X"AA",X"09",X"33",X"BE",X"21",X"A0",X"4A",
		X"81",X"B8",X"70",X"B8",X"00",X"03",X"AF",X"21",X"80",X"BA",X"70",X"A0",X"81",X"1B",X"84",X"99",
		X"01",X"0C",X"97",X"8A",X"10",X"02",X"BF",X"58",X"A2",X"8B",X"58",X"D2",X"2B",X"20",X"D2",X"2C",
		X"02",X"B1",X"3A",X"91",X"9A",X"50",X"B0",X"39",X"09",X"F4",X"1B",X"82",X"A1",X"3B",X"D3",X"2A",
		X"81",X"89",X"4A",X"F4",X"0B",X"12",X"B1",X"2F",X"13",X"B8",X"3A",X"93",X"AA",X"25",X"BB",X"41",
		X"B2",X"0F",X"23",X"B9",X"3A",X"84",X"9F",X"23",X"C0",X"1A",X"03",X"AB",X"13",X"1B",X"93",X"91",
		X"4F",X"A7",X"0B",X"01",X"92",X"8B",X"95",X"1B",X"91",X"28",X"1B",X"A3",X"13",X"DC",X"23",X"1A",
		X"E1",X"83",X"4E",X"A3",X"29",X"88",X"9B",X"64",X"D9",X"30",X"90",X"99",X"38",X"98",X"82",X"3C",
		X"83",X"B8",X"13",X"8D",X"12",X"BB",X"71",X"EA",X"44",X"BB",X"22",X"08",X"A9",X"30",X"81",X"BA",
		X"35",X"9B",X"82",X"99",X"78",X"E2",X"3A",X"A1",X"18",X"E1",X"59",X"D2",X"19",X"00",X"A1",X"2C",
		X"12",X"B0",X"38",X"A8",X"21",X"BF",X"23",X"C9",X"28",X"01",X"9A",X"90",X"78",X"C3",X"1A",X"18",
		X"B4",X"0C",X"94",X"89",X"22",X"F1",X"28",X"B0",X"95",X"2E",X"93",X"19",X"A0",X"11",X"C1",X"4D",
		X"83",X"9A",X"39",X"95",X"8D",X"13",X"99",X"80",X"00",X"0A",X"08",X"C6",X"2D",X"84",X"8A",X"28",
		X"A0",X"2B",X"83",X"98",X"10",X"01",X"B2",X"4D",X"94",X"0D",X"12",X"A8",X"8B",X"62",X"D8",X"82",
		X"19",X"B2",X"10",X"0C",X"03",X"2A",X"E8",X"52",X"C8",X"19",X"A6",X"8B",X"28",X"B5",X"89",X"21",
		X"B1",X"8B",X"42",X"E8",X"08",X"38",X"A3",X"8A",X"41",X"B3",X"9F",X"06",X"9B",X"28",X"B5",X"99",
		X"3A",X"9A",X"87",X"2C",X"81",X"98",X"40",X"D1",X"2E",X"14",X"AA",X"29",X"03",X"9B",X"10",X"91",
		X"38",X"99",X"B3",X"23",X"4F",X"C2",X"29",X"91",X"8B",X"07",X"09",X"98",X"82",X"31",X"EC",X"05",
		X"89",X"3C",X"A4",X"1A",X"11",X"E0",X"29",X"11",X"BB",X"41",X"01",X"BD",X"24",X"AA",X"38",X"C2",
		X"08",X"13",X"F9",X"31",X"89",X"8A",X"17",X"AA",X"18",X"23",X"F8",X"20",X"88",X"94",X"8B",X"02",
		X"9A",X"05",X"8D",X"02",X"88",X"8A",X"37",X"C8",X"3A",X"03",X"E9",X"79",X"91",X"89",X"39",X"C3",
		X"1C",X"30",X"C1",X"19",X"01",X"A9",X"48",X"A8",X"18",X"6B",X"C4",X"09",X"18",X"A2",X"4B",X"A2",
		X"09",X"10",X"B0",X"7A",X"B5",X"8B",X"30",X"C5",X"8C",X"21",X"B1",X"1A",X"12",X"9C",X"24",X"B9",
		X"29",X"A7",X"9C",X"30",X"91",X"0B",X"17",X"AB",X"40",X"A1",X"8B",X"24",X"9B",X"83",X"1A",X"00",
		X"A7",X"2F",X"83",X"99",X"19",X"83",X"2F",X"82",X"1A",X"90",X"82",X"19",X"9A",X"36",X"BA",X"01",
		X"4A",X"99",X"C6",X"2B",X"B3",X"01",X"12",X"ED",X"51",X"B8",X"18",X"10",X"B8",X"10",X"2B",X"94",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"87",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E0",X"04",
		X"ED",X"00",X"7C",X"BA",X"C0",X"7D",X"BB",X"C9",X"A7",X"ED",X"52",X"23",X"C9",X"23",X"7C",X"B5",
		X"2B",X"C9",X"7D",X"02",X"03",X"7C",X"02",X"03",X"C9",X"1A",X"6F",X"13",X"1A",X"67",X"C9",X"DB",
		X"04",X"E6",X"80",X"32",X"FD",X"FE",X"C9",X"31",X"00",X"F6",X"CD",X"60",X"F0",X"CD",X"23",X"EB",
		X"31",X"00",X"F6",X"21",X"03",X"E0",X"06",X"5F",X"AF",X"77",X"23",X"10",X"FC",X"CD",X"CA",X"E0",
		X"AF",X"32",X"FD",X"FE",X"32",X"FE",X"FE",X"3A",X"04",X"E0",X"A7",X"CC",X"84",X"F2",X"06",X"01",
		X"CD",X"43",X"F3",X"CD",X"B8",X"F2",X"06",X"01",X"CD",X"43",X"F3",X"CD",X"B8",X"F2",X"0E",X"00",
		X"CD",X"86",X"F3",X"0E",X"00",X"CD",X"86",X"F3",X"18",X"C6",X"AF",X"32",X"03",X"E0",X"32",X"FD",
		X"FE",X"32",X"01",X"F6",X"21",X"05",X"E0",X"22",X"5D",X"E0",X"21",X"04",X"ED",X"22",X"5F",X"E0",
		X"06",X"4D",X"36",X"20",X"23",X"10",X"FB",X"21",X"3D",X"EB",X"CD",X"50",X"F2",X"CD",X"1E",X"F1",
		X"FE",X"01",X"CA",X"36",X"E1",X"FE",X"02",X"CA",X"96",X"E1",X"FE",X"03",X"CA",X"36",X"E2",X"FE",
		X"04",X"CA",X"47",X"E2",X"FE",X"06",X"CA",X"D0",X"F0",X"FE",X"07",X"20",X"BD",X"21",X"85",X"EB",
		X"CD",X"50",X"F2",X"CD",X"1E",X"F1",X"FE",X"01",X"CA",X"C3",X"EE",X"FE",X"02",X"CA",X"00",X"F7",
		X"FE",X"03",X"CA",X"00",X"F4",X"FE",X"04",X"CA",X"94",X"ED",X"FE",X"05",X"CA",X"00",X"FB",X"FE",
		X"07",X"C2",X"0D",X"E1",X"18",X"94",X"21",X"3F",X"EB",X"0E",X"05",X"CD",X"FE",X"EA",X"CD",X"75",
		X"E2",X"CD",X"84",X"F2",X"21",X"20",X"EC",X"CD",X"50",X"F2",X"CD",X"45",X"F1",X"CD",X"D3",X"EA",
		X"20",X"F8",X"21",X"22",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"2D",X"EC",
		X"CD",X"50",X"F2",X"CD",X"45",X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"38",X"26",X"21",X"2F",X"EC",
		X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"47",X"EC",X"CD",X"50",X"F2",X"CD",X"45",
		X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"38",X"0B",X"21",X"4F",X"EC",X"0E",X"02",X"CD",X"FE",X"EA",
		X"CD",X"12",X"EB",X"C3",X"19",X"E9",X"21",X"49",X"EB",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"75",
		X"E2",X"CD",X"84",X"F2",X"21",X"5C",X"EC",X"CD",X"50",X"F2",X"CD",X"45",X"F1",X"CD",X"D3",X"EA",
		X"20",X"EF",X"21",X"5E",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"69",X"EC",
		X"CD",X"50",X"F2",X"CD",X"1E",X"F1",X"FE",X"01",X"28",X"5F",X"FE",X"03",X"20",X"F5",X"21",X"7D",
		X"EC",X"0E",X"0C",X"CD",X"FE",X"EA",X"CD",X"84",X"F2",X"21",X"8A",X"EC",X"CD",X"50",X"F2",X"CD",
		X"45",X"F1",X"CD",X"D3",X"EA",X"20",X"F8",X"CD",X"12",X"EB",X"CD",X"84",X"F2",X"21",X"93",X"EC",
		X"CD",X"50",X"F2",X"CD",X"45",X"F1",X"3A",X"04",X"F8",X"CD",X"DD",X"EA",X"20",X"F5",X"38",X"26",
		X"21",X"22",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"A9",X"EC",X"CD",X"50",
		X"F2",X"CD",X"45",X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"38",X"0B",X"21",X"2F",X"EC",X"0E",X"04",
		X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"C3",X"99",X"E8",X"21",X"6B",X"EC",X"0E",X"0A",X"CD",X"FE",
		X"EA",X"CD",X"04",X"E3",X"18",X"B4",X"21",X"52",X"EB",X"0E",X"0A",X"CD",X"FE",X"EA",X"CD",X"75",
		X"E2",X"CD",X"04",X"E3",X"C3",X"19",X"E9",X"21",X"5D",X"EB",X"0E",X"07",X"CD",X"FE",X"EA",X"CD",
		X"75",X"E2",X"CD",X"04",X"E3",X"CD",X"84",X"F2",X"21",X"8A",X"EC",X"CD",X"50",X"F2",X"CD",X"45",
		X"F1",X"CD",X"D3",X"EA",X"20",X"F8",X"21",X"7D",X"EC",X"01",X"0C",X"00",X"CD",X"FE",X"EA",X"CD",
		X"12",X"EB",X"C3",X"EA",X"E1",X"21",X"CD",X"EB",X"CD",X"50",X"F2",X"CD",X"1E",X"F1",X"FE",X"07",
		X"28",X"1A",X"FE",X"06",X"28",X"23",X"FE",X"05",X"28",X"2C",X"FE",X"04",X"28",X"35",X"FE",X"03",
		X"28",X"3E",X"FE",X"02",X"28",X"47",X"FE",X"01",X"28",X"50",X"18",X"D9",X"3E",X"00",X"01",X"09",
		X"00",X"11",X"0B",X"EC",X"21",X"00",X"08",X"18",X"4C",X"3E",X"32",X"01",X"06",X"00",X"11",X"02",
		X"EC",X"21",X"20",X"00",X"18",X"3F",X"3E",X"34",X"01",X"06",X"00",X"11",X"F8",X"EB",X"21",X"00",
		X"02",X"18",X"32",X"3E",X"54",X"01",X"04",X"00",X"11",X"EE",X"EB",X"21",X"00",X"10",X"18",X"25",
		X"3E",X"54",X"01",X"04",X"10",X"11",X"E4",X"EB",X"21",X"00",X"20",X"18",X"18",X"3E",X"49",X"01",
		X"04",X"00",X"11",X"DA",X"EB",X"21",X"00",X"10",X"18",X"0B",X"3E",X"49",X"01",X"04",X"10",X"11",
		X"D0",X"EB",X"21",X"00",X"20",X"32",X"41",X"E0",X"22",X"45",X"E0",X"21",X"40",X"E0",X"70",X"EB",
		X"CD",X"FE",X"EA",X"C9",X"11",X"FF",X"FF",X"2A",X"5D",X"E0",X"73",X"23",X"72",X"23",X"22",X"5D",
		X"E0",X"21",X"03",X"E0",X"34",X"C9",X"21",X"00",X"00",X"22",X"4D",X"E0",X"7D",X"32",X"3F",X"E0",
		X"2A",X"05",X"E0",X"22",X"49",X"E0",X"22",X"4F",X"E0",X"3A",X"03",X"E0",X"C9",X"CD",X"33",X"E3",
		X"C3",X"B8",X"E3",X"CD",X"16",X"E3",X"FE",X"01",X"20",X"23",X"2A",X"49",X"E0",X"11",X"00",X"E0",
		X"CD",X"62",X"E0",X"38",X"07",X"21",X"FF",X"FF",X"22",X"49",X"E0",X"23",X"EB",X"2A",X"45",X"E0",
		X"22",X"47",X"E0",X"2B",X"19",X"22",X"4B",X"E0",X"3E",X"01",X"D8",X"AF",X"C9",X"FE",X"02",X"20",
		X"21",X"EB",X"2A",X"07",X"E0",X"22",X"4B",X"E0",X"CD",X"68",X"E0",X"38",X"EB",X"22",X"47",X"E0",
		X"EB",X"2A",X"45",X"E0",X"1B",X"CD",X"62",X"E0",X"3E",X"00",X"30",X"01",X"3C",X"32",X"3F",X"E0",
		X"AF",X"C9",X"EB",X"2A",X"07",X"E0",X"22",X"4B",X"E0",X"CD",X"68",X"E0",X"38",X"CA",X"22",X"47",
		X"E0",X"2A",X"09",X"E0",X"22",X"4D",X"E0",X"EB",X"2A",X"45",X"E0",X"2B",X"CD",X"62",X"E0",X"3E",
		X"01",X"38",X"DA",X"2A",X"47",X"E0",X"19",X"EB",X"2A",X"45",X"E0",X"CD",X"62",X"E0",X"3E",X"00",
		X"30",X"CB",X"3C",X"18",X"C8",X"CD",X"92",X"E4",X"A7",X"C0",X"21",X"05",X"E0",X"06",X"3A",X"36",
		X"00",X"23",X"10",X"FB",X"3A",X"3F",X"E0",X"A7",X"28",X"2E",X"2A",X"45",X"E0",X"11",X"00",X"10",
		X"CD",X"62",X"E0",X"3E",X"00",X"30",X"61",X"ED",X"5B",X"45",X"E0",X"2A",X"47",X"E0",X"2B",X"CD",
		X"62",X"E0",X"D2",X"F9",X"E4",X"44",X"4D",X"2A",X"4D",X"E0",X"09",X"DA",X"58",X"E3",X"CD",X"62",
		X"E0",X"3E",X"01",X"D0",X"AF",X"32",X"3F",X"E0",X"D5",X"2A",X"45",X"E0",X"11",X"00",X"10",X"CD",
		X"62",X"E0",X"D1",X"21",X"56",X"E0",X"3E",X"01",X"38",X"02",X"3E",X"07",X"77",X"01",X"05",X"E0",
		X"2A",X"47",X"E0",X"CD",X"72",X"E0",X"2A",X"4D",X"E0",X"CD",X"72",X"E0",X"EB",X"2A",X"45",X"E0",
		X"19",X"22",X"4D",X"E0",X"2A",X"49",X"E0",X"CD",X"72",X"E0",X"2A",X"4F",X"E0",X"CD",X"72",X"E0",
		X"21",X"56",X"E0",X"35",X"20",X"DA",X"AF",X"C9",X"01",X"05",X"E0",X"ED",X"5B",X"45",X"E0",X"2A",
		X"4D",X"E0",X"A7",X"ED",X"52",X"30",X"FC",X"7D",X"2F",X"5F",X"7C",X"2F",X"57",X"13",X"2A",X"47",
		X"E0",X"CD",X"62",X"E0",X"F5",X"28",X"08",X"38",X"06",X"ED",X"52",X"22",X"47",X"E0",X"EB",X"CD",
		X"72",X"E0",X"EB",X"2A",X"4D",X"E0",X"CD",X"72",X"E0",X"19",X"22",X"4D",X"E0",X"2A",X"49",X"E0",
		X"CD",X"72",X"E0",X"CD",X"6D",X"E0",X"28",X"01",X"19",X"22",X"49",X"E0",X"2A",X"4F",X"E0",X"CD",
		X"72",X"E0",X"CD",X"6D",X"E0",X"28",X"01",X"19",X"22",X"4F",X"E0",X"F1",X"3E",X"00",X"C8",X"30",
		X"AA",X"C9",X"CD",X"16",X"E3",X"11",X"FF",X"FF",X"ED",X"53",X"4F",X"E0",X"FE",X"01",X"20",X"0C",
		X"11",X"00",X"E0",X"CD",X"62",X"E0",X"DA",X"4C",X"E3",X"3E",X"01",X"C9",X"47",X"11",X"00",X"E0",
		X"CD",X"62",X"E0",X"38",X"07",X"21",X"FF",X"FF",X"22",X"49",X"E0",X"23",X"78",X"FE",X"02",X"EB",
		X"2A",X"07",X"E0",X"22",X"4F",X"E0",X"CA",X"4D",X"E3",X"2A",X"09",X"E0",X"22",X"4D",X"E0",X"3E",
		X"01",X"32",X"3F",X"E0",X"78",X"FE",X"03",X"CA",X"4D",X"E3",X"EB",X"2A",X"0B",X"E0",X"CD",X"68",
		X"E0",X"DA",X"58",X"E3",X"22",X"47",X"E0",X"EB",X"2A",X"49",X"E0",X"CD",X"6D",X"E0",X"C8",X"19",
		X"22",X"4B",X"E0",X"11",X"00",X"E0",X"CD",X"62",X"E0",X"3E",X"01",X"D0",X"AF",X"C9",X"3A",X"41",
		X"E0",X"FE",X"32",X"28",X"04",X"FE",X"34",X"20",X"03",X"AF",X"18",X"10",X"A7",X"20",X"04",X"3E",
		X"10",X"18",X"09",X"06",X"30",X"FE",X"49",X"28",X"02",X"06",X"20",X"78",X"32",X"43",X"E0",X"C9",
		X"3A",X"3F",X"E0",X"A7",X"28",X"14",X"21",X"07",X"E0",X"7E",X"23",X"66",X"6F",X"ED",X"5B",X"45",
		X"E0",X"06",X"FF",X"A7",X"ED",X"52",X"04",X"30",X"FA",X"78",X"32",X"51",X"E0",X"C9",X"CD",X"5E",
		X"E5",X"D5",X"11",X"10",X"27",X"1B",X"7A",X"B3",X"20",X"FB",X"D1",X"C9",X"11",X"C0",X"C0",X"3A",
		X"43",X"E0",X"E6",X"30",X"FE",X"20",X"30",X"03",X"50",X"18",X"01",X"58",X"B2",X"C9",X"F5",X"32",
		X"44",X"E0",X"06",X"82",X"FE",X"00",X"20",X"02",X"06",X"80",X"78",X"D3",X"03",X"F1",X"E6",X"C0",
		X"47",X"D5",X"CD",X"4C",X"E5",X"D3",X"02",X"3A",X"3F",X"E0",X"A7",X"3E",X"0E",X"28",X"01",X"AF",
		X"47",X"3A",X"40",X"E0",X"E6",X"10",X"B0",X"32",X"40",X"E0",X"B3",X"D3",X"05",X"D1",X"C9",X"3A",
		X"44",X"E0",X"E6",X"C0",X"47",X"D5",X"CD",X"4C",X"E5",X"47",X"7C",X"E6",X"0F",X"B0",X"D3",X"02",
		X"7D",X"D3",X"00",X"3A",X"40",X"E0",X"E6",X"0E",X"FE",X"0E",X"7C",X"28",X"17",X"E6",X"F0",X"47",
		X"3A",X"43",X"E0",X"E6",X"20",X"28",X"0A",X"3A",X"40",X"E0",X"E6",X"10",X"20",X"03",X"78",X"17",
		X"47",X"78",X"18",X"04",X"E6",X"10",X"F6",X"E0",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"40",X"E0",
		X"E6",X"10",X"B0",X"E6",X"1F",X"32",X"40",X"E0",X"B3",X"D1",X"D3",X"05",X"C9",X"D5",X"C5",X"06",
		X"80",X"CD",X"4C",X"E5",X"47",X"7C",X"E6",X"0F",X"B0",X"D3",X"02",X"47",X"3A",X"40",X"E0",X"B3",
		X"D3",X"05",X"4F",X"ED",X"5B",X"58",X"E0",X"1B",X"7A",X"B3",X"20",X"FB",X"78",X"CD",X"0B",X"E6",
		X"D3",X"02",X"79",X"CD",X"0B",X"E6",X"D3",X"05",X"C1",X"D1",X"C9",X"CB",X"77",X"C0",X"E6",X"7F",
		X"C9",X"21",X"05",X"E0",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",
		X"EB",X"C9",X"3A",X"03",X"E0",X"FE",X"03",X"3E",X"00",X"C8",X"D5",X"E5",X"2A",X"45",X"E0",X"11",
		X"00",X"10",X"CD",X"62",X"E0",X"E1",X"D1",X"01",X"01",X"01",X"38",X"02",X"0E",X"07",X"C5",X"3E",
		X"40",X"CD",X"3E",X"E5",X"3A",X"40",X"E0",X"E6",X"10",X"32",X"40",X"E0",X"11",X"00",X"00",X"C1",
		X"3E",X"00",X"F5",X"C5",X"D5",X"CD",X"8B",X"E6",X"D1",X"C1",X"28",X"01",X"C5",X"04",X"0D",X"28",
		X"07",X"2A",X"45",X"E0",X"19",X"EB",X"18",X"EB",X"3E",X"C0",X"CD",X"3E",X"E5",X"F1",X"A7",X"C8",
		X"CD",X"DB",X"E7",X"21",X"C5",X"EC",X"CD",X"54",X"F2",X"F1",X"A7",X"28",X"0B",X"CD",X"DB",X"E7",
		X"21",X"C5",X"EC",X"CD",X"54",X"F2",X"18",X"F1",X"3E",X"80",X"C9",X"ED",X"4B",X"45",X"E0",X"EB",
		X"50",X"59",X"CD",X"8F",X"E5",X"23",X"3A",X"43",X"E0",X"E6",X"30",X"06",X"FF",X"20",X"01",X"04",
		X"DB",X"01",X"B8",X"C0",X"1B",X"7A",X"B3",X"20",X"E9",X"C9",X"3E",X"C0",X"CD",X"3E",X"E5",X"3E",
		X"40",X"CD",X"3E",X"E5",X"3A",X"40",X"E0",X"E6",X"10",X"32",X"40",X"E0",X"AF",X"32",X"5B",X"E0",
		X"21",X"00",X"00",X"22",X"56",X"E0",X"22",X"52",X"E0",X"21",X"51",X"E0",X"34",X"2A",X"4B",X"E0",
		X"7E",X"4F",X"23",X"B6",X"F5",X"3E",X"C0",X"CC",X"3E",X"E5",X"F1",X"C8",X"46",X"23",X"EB",X"CD",
		X"79",X"E0",X"22",X"4D",X"E0",X"13",X"CD",X"79",X"E0",X"22",X"49",X"E0",X"13",X"CD",X"79",X"E0",
		X"22",X"4F",X"E0",X"13",X"EB",X"22",X"4B",X"E0",X"C5",X"2A",X"4D",X"E0",X"CD",X"8F",X"E5",X"EB",
		X"2A",X"49",X"E0",X"CD",X"6D",X"E0",X"DB",X"01",X"28",X"0D",X"47",X"3A",X"54",X"E0",X"A7",X"78",
		X"28",X"05",X"77",X"23",X"22",X"49",X"E0",X"21",X"5B",X"E0",X"FE",X"FF",X"28",X"05",X"35",X"28",
		X"01",X"34",X"34",X"F5",X"2A",X"52",X"E0",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"22",X"52",X"E0",
		X"F1",X"2A",X"4F",X"E0",X"BE",X"C4",X"19",X"E8",X"C1",X"28",X"04",X"AF",X"32",X"55",X"E0",X"2A",
		X"4D",X"E0",X"23",X"22",X"4D",X"E0",X"2A",X"4F",X"E0",X"CD",X"6D",X"E0",X"28",X"04",X"23",X"22",
		X"4F",X"E0",X"0B",X"78",X"B1",X"20",X"A1",X"3E",X"C0",X"CD",X"3E",X"E5",X"3A",X"5C",X"E0",X"A7",
		X"20",X"05",X"3A",X"5B",X"E0",X"A7",X"C0",X"F5",X"F5",X"CD",X"D8",X"E7",X"F1",X"21",X"BF",X"EC",
		X"CC",X"54",X"F2",X"F1",X"C8",X"3A",X"61",X"E0",X"A7",X"28",X"2B",X"06",X"02",X"CD",X"43",X"F3",
		X"CD",X"B8",X"F2",X"06",X"02",X"CD",X"43",X"F3",X"CD",X"B8",X"F2",X"06",X"02",X"CD",X"43",X"F3",
		X"CD",X"B8",X"F2",X"AF",X"32",X"61",X"E0",X"0E",X"80",X"CD",X"86",X"F3",X"0E",X"80",X"CD",X"86",
		X"F3",X"0E",X"80",X"CD",X"86",X"F3",X"CD",X"D8",X"E7",X"CD",X"0E",X"F2",X"2A",X"4F",X"E0",X"CD",
		X"6D",X"E0",X"28",X"12",X"2A",X"56",X"E0",X"7C",X"B5",X"28",X"0B",X"21",X"CE",X"EC",X"CD",X"57",
		X"F2",X"2A",X"56",X"E0",X"18",X"09",X"21",X"D3",X"EC",X"CD",X"57",X"F2",X"2A",X"52",X"E0",X"CD",
		X"E6",X"E7",X"2A",X"56",X"E0",X"7C",X"B5",X"C9",X"3A",X"51",X"E0",X"47",X"3E",X"F8",X"C6",X"0A",
		X"10",X"FC",X"57",X"1E",X"11",X"C9",X"7C",X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",X"0D",X"E8",X"CD",
		X"2C",X"F2",X"F1",X"CD",X"0D",X"E8",X"CD",X"2C",X"F2",X"7D",X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",
		X"0D",X"E8",X"CD",X"2C",X"F2",X"F1",X"CD",X"0D",X"E8",X"CD",X"2C",X"F2",X"C9",X"E6",X"0F",X"FE",
		X"0A",X"30",X"03",X"F6",X"30",X"C9",X"C6",X"37",X"C9",X"4F",X"2A",X"4F",X"E0",X"CD",X"6D",X"E0",
		X"C8",X"2A",X"56",X"E0",X"23",X"22",X"56",X"E0",X"3A",X"55",X"E0",X"A7",X"C8",X"C5",X"3E",X"01",
		X"32",X"61",X"E0",X"3A",X"FE",X"FE",X"FE",X"12",X"38",X"23",X"CD",X"45",X"F1",X"C1",X"3A",X"04",
		X"F8",X"FE",X"0D",X"28",X"52",X"C5",X"AF",X"32",X"FE",X"FE",X"21",X"D8",X"EC",X"CD",X"74",X"F1",
		X"3A",X"51",X"E0",X"F6",X"30",X"CD",X"BA",X"F2",X"CD",X"B8",X"F2",X"18",X"0A",X"2B",X"7C",X"B5",
		X"20",X"05",X"CD",X"B8",X"F2",X"18",X"E3",X"06",X"02",X"CD",X"43",X"F3",X"2A",X"4D",X"E0",X"CD",
		X"26",X"F3",X"06",X"02",X"CD",X"43",X"F3",X"C1",X"79",X"CD",X"2B",X"F3",X"06",X"03",X"CD",X"43",
		X"F3",X"2A",X"4F",X"E0",X"7E",X"F5",X"CD",X"26",X"F3",X"06",X"02",X"CD",X"43",X"F3",X"F1",X"CD",
		X"2B",X"F3",X"CD",X"B8",X"F2",X"AF",X"C9",X"A7",X"C9",X"CD",X"B5",X"E3",X"A7",X"C0",X"CD",X"FE",
		X"E4",X"11",X"11",X"01",X"CD",X"87",X"F2",X"11",X"12",X"01",X"CD",X"87",X"F2",X"3E",X"01",X"32",
		X"5C",X"E0",X"32",X"54",X"E0",X"32",X"55",X"E0",X"21",X"05",X"E0",X"22",X"4B",X"E0",X"CD",X"20",
		X"E5",X"3A",X"3F",X"E0",X"A7",X"28",X"0C",X"2A",X"4B",X"E0",X"7E",X"23",X"B6",X"C8",X"CD",X"AA",
		X"E6",X"18",X"F4",X"06",X"07",X"D5",X"E5",X"2A",X"45",X"E0",X"11",X"00",X"10",X"CD",X"62",X"E0",
		X"E1",X"D1",X"30",X"02",X"06",X"01",X"C5",X"AF",X"32",X"5C",X"E0",X"32",X"54",X"E0",X"32",X"55",
		X"E0",X"CD",X"AA",X"E6",X"3A",X"5B",X"E0",X"A7",X"28",X"1A",X"32",X"5C",X"E0",X"32",X"54",X"E0",
		X"00",X"00",X"00",X"01",X"A0",X"40",X"02",X"B0",X"A2",X"F0",X"01",X"B0",X"A4",X"A0",X"01",X"50",
		X"A5",X"F0",X"10",X"00",X"B5",X"F0",X"18",X"80",X"CE",X"70",X"03",X"A0",X"D2",X"10",X"08",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"F0",X"E5",X"F1",X"0A",X"F1",X"AF",X"F1",X"DD",X"F2",X"6D",X"F2",X"C8",
		X"F3",X"FE",X"F4",X"1C",X"F4",X"36",X"F3",X"63",X"F1",X"81",X"E9",X"D9",X"E9",X"D9",X"E9",X"D9",
		X"E9",X"D9",X"E9",X"D9",X"E9",X"7E",X"EA",X"2F",X"EA",X"F2",X"EB",X"CB",X"ED",X"26",X"40",X"00",
		X"41",X"00",X"42",X"00",X"43",X"00",X"44",X"00",X"48",X"00",X"49",X"00",X"4A",X"00",X"45",X"00",
		X"4B",X"00",X"4C",X"00",X"4D",X"00",X"6C",X"00",X"6D",X"00",X"6E",X"00",X"66",X"BC",X"6C",X"14",
		X"6D",X"14",X"FE",X"E9",X"DA",X"FE",X"EA",X"1B",X"FE",X"E9",X"DA",X"FE",X"EA",X"1B",X"FE",X"E9",
		X"DA",X"40",X"8E",X"48",X"0D",X"69",X"0D",X"02",X"7A",X"40",X"69",X"0D",X"02",X"7A",X"20",X"48",
		X"00",X"40",X"9F",X"68",X"0D",X"69",X"0D",X"02",X"1C",X"40",X"40",X"8E",X"68",X"0D",X"69",X"0D",
		X"02",X"1C",X"20",X"6C",X"00",X"6D",X"00",X"67",X"03",X"FF",X"42",X"38",X"43",X"02",X"49",X"0D",
		X"68",X"0D",X"00",X"47",X"20",X"68",X"0D",X"00",X"4F",X"20",X"49",X"00",X"68",X"0D",X"69",X"0D",
		X"00",X"5E",X"20",X"42",X"DD",X"43",X"01",X"49",X"0D",X"68",X"0D",X"00",X"6A",X"20",X"68",X"0D",
		X"00",X"77",X"20",X"49",X"00",X"68",X"0D",X"69",X"0D",X"00",X"8E",X"20",X"40",X"77",X"48",X"0D",
		X"69",X"0D",X"02",X"A9",X"40",X"69",X"0D",X"02",X"A9",X"20",X"FD",X"40",X"8E",X"48",X"0D",X"69",
		X"0D",X"02",X"7A",X"20",X"69",X"0D",X"02",X"3E",X"20",X"69",X"0D",X"02",X"1C",X"20",X"FD",X"66",
		X"BC",X"6C",X"10",X"6D",X"10",X"41",X"00",X"43",X"01",X"40",X"6A",X"68",X"0D",X"69",X"0D",X"02",
		X"7A",X"20",X"40",X"5E",X"68",X"0D",X"69",X"0D",X"02",X"7A",X"20",X"40",X"4F",X"48",X"0D",X"69",
		X"0D",X"02",X"C1",X"20",X"69",X"0D",X"02",X"C1",X"20",X"48",X"00",X"40",X"5E",X"68",X"0D",X"69",
		X"0D",X"02",X"A9",X"20",X"40",X"6A",X"68",X"0D",X"69",X"0D",X"02",X"A9",X"20",X"40",X"7E",X"48",
		X"0D",X"69",X"0D",X"02",X"90",X"20",X"69",X"0D",X"02",X"90",X"20",X"40",X"6A",X"48",X"0D",X"69",
		X"0D",X"02",X"7A",X"20",X"69",X"0D",X"02",X"7A",X"20",X"40",X"7E",X"48",X"0D",X"69",X"0D",X"02",
		X"C1",X"20",X"69",X"0D",X"02",X"C1",X"20",X"40",X"8E",X"48",X"0D",X"69",X"0D",X"02",X"A9",X"20",
		X"69",X"0D",X"02",X"A9",X"20",X"40",X"9F",X"48",X"0D",X"69",X"0D",X"02",X"90",X"20",X"69",X"0D",
		X"02",X"90",X"20",X"42",X"7A",X"49",X"0D",X"68",X"0D",X"00",X"8E",X"20",X"68",X"0D",X"00",X"9F",
		X"20",X"49",X"00",X"40",X"BD",X"68",X"0D",X"69",X"0D",X"02",X"C1",X"40",X"40",X"D4",X"43",X"01",
		X"68",X"0D",X"69",X"0D",X"02",X"1C",X"20",X"40",X"C8",X"68",X"0D",X"69",X"0D",X"02",X"0C",X"20",
		X"40",X"BD",X"43",X"00",X"68",X"0D",X"69",X"0D",X"02",X"FD",X"80",X"67",X"03",X"6C",X"00",X"6D",
		X"00",X"FF",X"66",X"BC",X"6C",X"10",X"6D",X"10",X"40",X"38",X"41",X"02",X"48",X"0D",X"43",X"00",
		X"69",X"0D",X"02",X"EE",X"20",X"69",X"0D",X"02",X"E1",X"20",X"48",X"00",X"40",X"C1",X"41",X"01",
		X"68",X"0D",X"69",X"0D",X"02",X"8E",X"40",X"40",X"7A",X"68",X"0D",X"69",X"0D",X"02",X"9F",X"40",
		X"40",X"51",X"68",X"0D",X"69",X"0D",X"02",X"A8",X"40",X"40",X"3E",X"48",X"0D",X"69",X"0D",X"02",
		X"BD",X"20",X"69",X"0D",X"02",X"D4",X"20",X"48",X"00",X"40",X"51",X"68",X"0D",X"69",X"0D",X"02",
		X"EE",X"40",X"40",X"7A",X"48",X"0D",X"69",X"0D",X"02",X"EE",X"20",X"69",X"0D",X"02",X"E1",X"20",
		X"48",X"00",X"40",X"C1",X"68",X"0D",X"69",X"0D",X"02",X"D4",X"40",X"40",X"A7",X"41",X"02",X"68",
		X"0D",X"69",X"0D",X"02",X"E1",X"20",X"40",X"51",X"41",X"01",X"68",X"0D",X"69",X"0D",X"02",X"8E",
		X"20",X"40",X"7D",X"41",X"02",X"68",X"0D",X"69",X"0D",X"02",X"D4",X"20",X"40",X"3E",X"41",X"01",
		X"68",X"0D",X"69",X"0D",X"02",X"7E",X"20",X"40",X"58",X"41",X"02",X"68",X"0D",X"69",X"0D",X"02",
		X"C8",X"20",X"40",X"2C",X"41",X"01",X"68",X"0D",X"69",X"0D",X"02",X"77",X"20",X"40",X"38",X"41",
		X"02",X"68",X"0D",X"69",X"0D",X"02",X"BD",X"20",X"40",X"1C",X"41",X"01",X"68",X"0D",X"69",X"0D",
		X"02",X"70",X"20",X"40",X"38",X"41",X"02",X"68",X"0D",X"69",X"0D",X"02",X"70",X"40",X"67",X"03",
		X"6C",X"00",X"6D",X"00",X"48",X"00",X"49",X"00",X"4A",X"00",X"FF",X"66",X"B8",X"6C",X"14",X"6D",
		X"14",X"6E",X"14",X"FE",X"EC",X"62",X"FE",X"EC",X"62",X"FE",X"EC",X"62",X"40",X"3F",X"42",X"54",
		X"45",X"01",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"68",X"0D",X"69",X"0D",X"6A",
		X"0D",X"04",X"7A",X"2D",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"68",X"0D",X"69",
		X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"68",
		X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",
		X"2D",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"40",X"3C",X"42",X"4F",X"68",X"0D",
		X"69",X"0D",X"6A",X"0D",X"04",X"A9",X"5A",X"40",X"3F",X"42",X"54",X"68",X"0D",X"69",X"0D",X"6A",
		X"0D",X"04",X"C1",X"2D",X"40",X"47",X"42",X"5E",X"45",X"02",X"68",X"0D",X"69",X"0D",X"6A",X"0D",
		X"04",X"38",X"5A",X"67",X"07",X"6C",X"00",X"6D",X"00",X"6E",X"00",X"48",X"00",X"49",X"00",X"4A",
		X"00",X"FF",X"4A",X"00",X"41",X"00",X"43",X"00",X"45",X"02",X"40",X"8E",X"42",X"BD",X"48",X"0D",
		X"49",X"0D",X"6A",X"0D",X"04",X"38",X"2D",X"45",X"01",X"6A",X"0D",X"04",X"C1",X"2D",X"48",X"00",
		X"49",X"00",X"40",X"70",X"42",X"8E",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"7A",X"2D",X"40",
		X"5E",X"44",X"38",X"45",X"02",X"4A",X"0D",X"68",X"0D",X"69",X"0D",X"02",X"70",X"2D",X"40",X"6A",
		X"68",X"0D",X"69",X"0D",X"02",X"8E",X"2D",X"4A",X"00",X"40",X"54",X"42",X"6A",X"45",X"01",X"68",
		X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"C1",X"2D",X"6A",X"0D",X"04",X"7A",X"2D",X"40",X"4F",X"42",
		X"6A",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"A9",X"5A",X"40",X"54",X"42",X"6A",X"68",X"0D",
		X"69",X"0D",X"6A",X"0D",X"04",X"51",X"2D",X"40",X"5E",X"42",X"70",X"68",X"0D",X"69",X"0D",X"6A",
		X"0D",X"04",X"1C",X"2D",X"40",X"77",X"44",X"EE",X"45",X"00",X"4A",X"0D",X"68",X"0D",X"69",X"0D",
		X"02",X"9F",X"2D",X"40",X"70",X"68",X"0D",X"69",X"0D",X"02",X"8E",X"2D",X"4A",X"00",X"40",X"9F",
		X"42",X"D4",X"68",X"0D",X"69",X"0D",X"6A",X"0D",X"04",X"FD",X"2D",X"40",X"9F",X"44",X"1C",X"45",
		X"01",X"4A",X"0D",X"68",X"0D",X"69",X"0D",X"02",X"D4",X"2D",X"40",X"8E",X"68",X"0D",X"69",X"0D",
		X"02",X"BD",X"2D",X"4A",X"00",X"FD",X"66",X"B5",X"6D",X"14",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"46",X"01",X"43",X"02",X"FE",X"EF",X"27",X"FE",X"EF",X"27",X"FE",X"EF",X"27",X"FE",X"EF",X"27",
		X"43",X"00",X"FE",X"F0",X"09",X"FE",X"F0",X"09",X"43",X"01",X"FE",X"EF",X"27",X"FE",X"EF",X"27",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"7A",X"30",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"69",X"0E",X"02",X"7A",X"16",X"43",X"00",X"02",X"00",
		X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",X"69",X"0E",X"02",X"A9",X"16",
		X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",
		X"0E",X"02",X"7A",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"69",X"0E",X"02",X"7A",
		X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",
		X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"7A",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",
		X"10",X"69",X"0E",X"02",X"7A",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"48",X"10",X"43",X"01",X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"69",X"0E",X"43",X"01",X"02",X"7A",X"16",X"43",X"00",
		X"02",X"00",X"02",X"43",X"01",X"69",X"0E",X"02",X"3E",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",
		X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"7A",X"16",X"43",X"00",
		X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",
		X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",
		X"01",X"69",X"0E",X"02",X"A9",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",
		X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"DD",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",
		X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",X"69",X"0E",X"02",X"A9",X"30",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"48",X"10",X"43",X"01",X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",
		X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"DD",X"16",
		X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",X"69",
		X"0E",X"02",X"A9",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",X"69",X"0E",
		X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",
		X"48",X"10",X"69",X"0E",X"02",X"DD",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",
		X"43",X"01",X"69",X"0E",X"02",X"65",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"48",X"10",X"43",X"01",X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"43",X"01",X"69",X"0E",X"02",X"DD",X"16",X"43",
		X"00",X"02",X"00",X"02",X"FE",X"ED",X"26",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"02",X"48",
		X"10",X"69",X"0E",X"02",X"38",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"69",X"0E",
		X"02",X"38",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"02",
		X"48",X"10",X"69",X"0E",X"02",X"7D",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"43",X"02",X"48",X"10",X"69",X"0E",X"02",X"38",X"30",X"48",X"10",X"69",X"0E",X"02",
		X"38",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"02",X"48",
		X"10",X"69",X"0E",X"02",X"7D",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",
		X"09",X"43",X"02",X"48",X"10",X"69",X"0E",X"02",X"38",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",
		X"48",X"10",X"69",X"0E",X"02",X"38",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"43",X"02",X"48",X"10",X"69",X"0E",X"02",X"7D",X"16",X"43",X"00",X"02",X"00",X"02",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"02",X"48",X"10",X"69",X"0E",X"02",X"38",X"16",X"43",
		X"00",X"02",X"00",X"02",X"43",X"01",X"69",X"0E",X"02",X"DD",X"16",X"43",X"00",X"02",X"00",X"02",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"02",X"48",X"10",X"69",X"0E",X"02",X"38",X"16",X"43",
		X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"02",X"48",X"10",X"69",X"0E",
		X"02",X"7D",X"16",X"43",X"00",X"02",X"00",X"02",X"FD",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",
		X"01",X"48",X"10",X"69",X"0E",X"02",X"A9",X"30",X"48",X"10",X"69",X"0E",X"02",X"A9",X"16",X"43",
		X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",
		X"02",X"DD",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",
		X"48",X"10",X"69",X"0E",X"02",X"A9",X"30",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"69",
		X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",
		X"01",X"48",X"10",X"69",X"0E",X"02",X"DD",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",
		X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"A9",X"30",X"48",X"10",X"69",X"0E",
		X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",
		X"48",X"10",X"69",X"0E",X"02",X"DD",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",
		X"43",X"01",X"69",X"0E",X"02",X"65",X"16",X"43",X"00",X"02",X"00",X"02",X"4B",X"03",X"4C",X"02",
		X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"A9",X"16",X"43",X"00",X"02",X"00",X"02",
		X"4B",X"03",X"4C",X"02",X"4D",X"09",X"43",X"01",X"48",X"10",X"69",X"0E",X"02",X"DD",X"16",X"43",
		X"00",X"02",X"00",X"02",X"FD",X"76",X"AE",X"50",X"00",X"51",X"00",X"52",X"00",X"53",X"00",X"58",
		X"10",X"59",X"10",X"5B",X"00",X"5C",X"02",X"5D",X"00",X"70",X"00",X"08",X"16",X"0C",X"10",X"58",
		X"00",X"59",X"00",X"5B",X"00",X"5C",X"00",X"77",X"11",X"FF",X"76",X"A7",X"58",X"0F",X"59",X"0F",
		X"51",X"01",X"53",X"01",X"16",X"16",X"05",X"58",X"05",X"59",X"00",X"30",X"00",X"00",X"04",X"58",
		X"0F",X"59",X"0F",X"16",X"08",X"05",X"58",X"0E",X"59",X"0E",X"16",X"07",X"05",X"58",X"0D",X"59",
		X"0D",X"16",X"09",X"05",X"58",X"0C",X"59",X"0C",X"16",X"0A",X"05",X"58",X"0B",X"59",X"0B",X"16",
		X"08",X"05",X"58",X"0A",X"59",X"0A",X"16",X"09",X"05",X"58",X"09",X"59",X"09",X"16",X"06",X"05",
		X"58",X"08",X"59",X"09",X"16",X"07",X"05",X"58",X"07",X"59",X"07",X"16",X"0A",X"05",X"58",X"06",
		X"59",X"06",X"16",X"08",X"05",X"58",X"05",X"59",X"05",X"16",X"06",X"05",X"58",X"04",X"59",X"04",
		X"16",X"08",X"05",X"58",X"02",X"59",X"02",X"16",X"0A",X"05",X"58",X"00",X"59",X"00",X"77",X"18",
		X"FF",X"66",X"AF",X"46",X"09",X"89",X"20",X"01",X"09",X"0A",X"0B",X"0D",X"0D",X"0E",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",
		X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"49",X"00",X"67",X"10",X"46",X"00",X"FF",X"66",
		X"97",X"46",X"09",X"8A",X"20",X"01",X"09",X"0A",X"0B",X"0D",X"0D",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",
		X"05",X"04",X"03",X"02",X"01",X"00",X"4A",X"00",X"67",X"20",X"46",X"01",X"FF",X"76",X"A4",X"58",
		X"0F",X"59",X"0F",X"56",X"18",X"70",X"12",X"00",X"31",X"25",X"01",X"02",X"70",X"18",X"00",X"31",
		X"28",X"00",X"02",X"70",X"1A",X"00",X"31",X"22",X"02",X"03",X"70",X"2C",X"00",X"31",X"2A",X"01",
		X"03",X"70",X"2D",X"00",X"31",X"22",X"00",X"02",X"70",X"2F",X"00",X"31",X"25",X"00",X"01",X"59",
		X"03",X"18",X"03",X"02",X"76",X"AC",X"58",X"0F",X"59",X"0F",X"56",X"02",X"5B",X"F0",X"5C",X"0A",
		X"FE",X"F2",X"34",X"58",X"10",X"59",X"10",X"FE",X"F2",X"34",X"FE",X"F2",X"34",X"58",X"00",X"59",
		X"00",X"77",X"1B",X"FF",X"70",X"18",X"00",X"31",X"10",X"00",X"05",X"70",X"1D",X"00",X"31",X"13",
		X"00",X"04",X"70",X"1C",X"00",X"31",X"0E",X"00",X"05",X"70",X"0A",X"00",X"31",X"10",X"00",X"04",
		X"70",X"08",X"00",X"31",X"10",X"00",X"04",X"70",X"0E",X"00",X"31",X"13",X"00",X"05",X"70",X"15",
		X"00",X"31",X"0E",X"00",X"04",X"70",X"1A",X"00",X"31",X"0A",X"00",X"04",X"FD",X"76",X"BB",X"66",
		X"B3",X"4A",X"0F",X"5A",X"0F",X"FE",X"F2",X"8F",X"0A",X"00",X"08",X"FE",X"F2",X"8F",X"44",X"00",
		X"45",X"00",X"55",X"00",X"54",X"00",X"48",X"A0",X"5A",X"00",X"77",X"04",X"67",X"04",X"FF",X"62",
		X"20",X"00",X"32",X"18",X"00",X"02",X"62",X"25",X"00",X"32",X"1A",X"00",X"01",X"62",X"23",X"00",
		X"32",X"15",X"00",X"02",X"62",X"0B",X"00",X"32",X"12",X"00",X"01",X"62",X"09",X"00",X"32",X"16",
		X"00",X"01",X"62",X"0E",X"00",X"32",X"1A",X"00",X"02",X"62",X"20",X"00",X"32",X"0E",X"00",X"01",
		X"62",X"29",X"00",X"32",X"0D",X"00",X"01",X"FD",X"66",X"97",X"46",X"00",X"4A",X"05",X"5A",X"05",
		X"76",X"BB",X"14",X"60",X"01",X"4A",X"07",X"5A",X"06",X"14",X"5C",X"01",X"4A",X"08",X"5A",X"07",
		X"14",X"58",X"01",X"4A",X"09",X"5A",X"08",X"14",X"54",X"01",X"4A",X"0A",X"5A",X"09",X"14",X"50",
		X"01",X"4A",X"0B",X"5A",X"0A",X"14",X"4C",X"01",X"4A",X"0C",X"5A",X"0B",X"14",X"48",X"01",X"4A",
		X"0D",X"5A",X"0C",X"14",X"44",X"01",X"4A",X"0E",X"5A",X"0D",X"14",X"40",X"01",X"4A",X"0F",X"5A",
		X"0E",X"14",X"3C",X"01",X"4A",X"0F",X"5A",X"0E",X"14",X"38",X"01",X"4A",X"0E",X"5A",X"0E",X"14",
		X"34",X"01",X"4A",X"0D",X"5A",X"0E",X"14",X"30",X"01",X"4A",X"0B",X"5A",X"0D",X"14",X"40",X"01",
		X"5A",X"0B",X"14",X"45",X"01",X"5A",X"09",X"14",X"4A",X"01",X"5A",X"08",X"14",X"4F",X"01",X"5A",
		X"06",X"14",X"53",X"01",X"5A",X"05",X"14",X"57",X"01",X"5A",X"04",X"14",X"5B",X"01",X"5A",X"03",
		X"14",X"60",X"01",X"5A",X"02",X"14",X"64",X"01",X"4A",X"00",X"5A",X"00",X"77",X"20",X"67",X"20",
		X"46",X"01",X"FF",X"66",X"9F",X"46",X"00",X"4A",X"05",X"5A",X"05",X"76",X"BB",X"14",X"60",X"01",
		X"4A",X"07",X"5A",X"06",X"14",X"5C",X"01",X"4A",X"08",X"5A",X"07",X"14",X"58",X"01",X"4A",X"09",
		X"5A",X"08",X"14",X"54",X"01",X"4A",X"0A",X"5A",X"09",X"14",X"50",X"01",X"4A",X"0B",X"5A",X"0A",
		X"14",X"4C",X"01",X"4A",X"0C",X"5A",X"0B",X"14",X"48",X"01",X"4A",X"0D",X"5A",X"0C",X"14",X"44",
		X"01",X"4A",X"0E",X"5A",X"0D",X"14",X"40",X"01",X"4A",X"0F",X"5A",X"0E",X"14",X"3C",X"01",X"4A",
		X"0F",X"5A",X"0E",X"14",X"38",X"01",X"4A",X"0E",X"5A",X"0E",X"14",X"34",X"01",X"4A",X"0D",X"5A",
		X"0E",X"14",X"30",X"01",X"4A",X"0B",X"5A",X"0D",X"14",X"40",X"01",X"5A",X"0B",X"14",X"45",X"01",
		X"5A",X"09",X"14",X"4A",X"01",X"5A",X"08",X"14",X"4F",X"01",X"5A",X"06",X"14",X"53",X"01",X"5A",
		X"05",X"14",X"57",X"01",X"5A",X"04",X"14",X"5B",X"01",X"5A",X"03",X"14",X"60",X"01",X"5A",X"02",
		X"14",X"64",X"01",X"4A",X"00",X"5A",X"00",X"77",X"04",X"67",X"20",X"46",X"00",X"FF",X"76",X"BC",
		X"58",X"10",X"59",X"10",X"5B",X"80",X"5C",X"02",X"5D",X"00",X"70",X"30",X"00",X"31",X"60",X"00",
		X"0C",X"30",X"30",X"00",X"04",X"58",X"00",X"59",X"00",X"77",X"03",X"FF",X"66",X"BE",X"41",X"00",
		X"6C",X"09",X"68",X"0F",X"00",X"77",X"22",X"68",X"0F",X"00",X"77",X"22",X"68",X"0F",X"00",X"77",
		X"22",X"6C",X"00",X"67",X"01",X"FF",X"66",X"B3",X"45",X"00",X"6E",X"14",X"6A",X"0F",X"04",X"43",
		X"30",X"6A",X"0F",X"04",X"53",X"E0",X"67",X"04",X"6E",X"00",X"FF",X"47",X"BF",X"57",X"BF",X"40",
		X"00",X"41",X"00",X"42",X"00",X"43",X"00",X"44",X"00",X"45",X"00",X"46",X"00",X"48",X"00",X"49",
		X"00",X"4A",X"00",X"4B",X"00",X"4C",X"00",X"4D",X"00",X"51",X"00",X"50",X"00",X"52",X"00",X"53",
		X"00",X"54",X"00",X"55",X"00",X"56",X"00",X"58",X"00",X"59",X"00",X"5A",X"00",X"5B",X"00",X"5C",
		X"00",X"5D",X"00",X"FF",X"73",X"F4",X"2A",X"07",X"E0",X"ED",X"5B",X"05",X"E0",X"09",X"2B",X"EB",
		X"09",X"2B",X"EB",X"ED",X"B8",X"C9",X"21",X"46",X"FF",X"CD",X"74",X"F1",X"C9",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"F7",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FD",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"99",X"E5",X"01",X"00",X"75",X"E5",X"75",X"E5",X"05",X"E8",
		X"0C",X"E8",X"D2",X"E7",X"80",X"EA",X"00",X"01",X"00",X"20",X"00",X"00",X"F0",X"E0",X"A0",X"E0",
		X"00",X"45",X"77",X"72",X"69",X"74",X"65",X"20",X"20",X"20",X"20",X"20",X"72",X"65",X"61",X"64",
		X"20",X"20",X"20",X"20",X"20",X"65",X"72",X"61",X"73",X"65",X"63",X"68",X"65",X"63",X"6B",X"20",
		X"63",X"6F",X"6D",X"70",X"61",X"72",X"65",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"65",X"6E",X"64",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"2D",X"2D",
		X"2D",X"45",X"54",X"43",X"2D",X"2D",X"2D",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"0D",X"0A",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"40",X"01",X"00",
		X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"02",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"F7",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"3E",X"01",X"32",X"FD",X"FE",X"21",X"91",X"EB",X"0E",X"05",X"CD",X"FE",X"EA",X"CD",X"5F",X"F7",
		X"CD",X"CE",X"EE",X"C3",X"4B",X"F3",X"D9",X"01",X"4B",X"00",X"11",X"89",X"FF",X"21",X"88",X"FF",
		X"3E",X"20",X"77",X"ED",X"B0",X"3E",X"0D",X"77",X"23",X"3E",X"00",X"77",X"D9",X"C9",X"13",X"79",
		X"1F",X"1F",X"1F",X"1F",X"CD",X"38",X"F7",X"79",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"07",
		X"C6",X"30",X"12",X"13",X"C9",X"13",X"CD",X"4E",X"F7",X"3E",X"2D",X"12",X"13",X"C9",X"4C",X"CD",
		X"2F",X"F7",X"4D",X"C3",X"2F",X"F7",X"7E",X"E6",X"7F",X"FE",X"20",X"D0",X"3E",X"20",X"C9",X"CD",
		X"84",X"F2",X"21",X"20",X"EC",X"CD",X"50",X"F2",X"CD",X"45",X"F1",X"CD",X"D3",X"EA",X"20",X"F8",
		X"21",X"22",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"2D",X"EC",X"CD",X"50",
		X"F2",X"CD",X"45",X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"D8",X"21",X"2F",X"EC",X"0E",X"04",X"CD",
		X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"3A",X"EC",X"CD",X"50",X"F2",X"CD",X"45",X"F1",X"CD",X"DD",
		X"EA",X"20",X"F8",X"D8",X"21",X"3C",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"C9",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"06",X"20",X"00",X"0D",X"46",X"46",X"46",X"0D",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",X"BF",X"00",X"FD",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FE",X"00",X"FF",X"00",X"EE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FD",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",
		X"EF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"7F",X"00",
		X"0F",X"8E",X"00",X"FF",X"BD",X"FA",X"93",X"86",X"BF",X"C6",X"07",X"BD",X"FA",X"D5",X"86",X"13",
		X"C6",X"0F",X"BD",X"FA",X"D5",X"86",X"3F",X"C6",X"17",X"BD",X"FA",X"D5",X"BD",X"FA",X"A8",X"7F",
		X"08",X"00",X"0F",X"BD",X"FA",X"43",X"96",X"BC",X"2B",X"07",X"BD",X"FC",X"C7",X"86",X"FF",X"97",
		X"BC",X"0E",X"CE",X"00",X"00",X"DF",X"D1",X"96",X"80",X"26",X"0B",X"DE",X"84",X"D6",X"8C",X"BD",
		X"FB",X"DB",X"DF",X"84",X"97",X"80",X"7C",X"00",X"D2",X"96",X"81",X"26",X"0B",X"DE",X"86",X"D6",
		X"8D",X"BD",X"FB",X"DB",X"DF",X"86",X"97",X"81",X"7C",X"00",X"D2",X"96",X"82",X"26",X"0B",X"DE",
		X"88",X"D6",X"8E",X"BD",X"FB",X"DB",X"DF",X"88",X"97",X"82",X"7C",X"00",X"D2",X"96",X"83",X"26",
		X"0B",X"DE",X"8A",X"D6",X"8F",X"BD",X"FB",X"DB",X"DF",X"8A",X"97",X"83",X"96",X"A8",X"27",X"08",
		X"7F",X"00",X"A8",X"C6",X"08",X"BD",X"FB",X"37",X"96",X"A9",X"27",X"08",X"7F",X"00",X"A9",X"C6",
		X"09",X"BD",X"FB",X"37",X"96",X"AA",X"27",X"08",X"7F",X"00",X"AA",X"C6",X"0A",X"BD",X"FB",X"37",
		X"96",X"AB",X"27",X"08",X"7F",X"00",X"AB",X"C6",X"18",X"BD",X"FB",X"50",X"96",X"AC",X"27",X"08",
		X"7F",X"00",X"AC",X"C6",X"19",X"BD",X"FB",X"50",X"96",X"AD",X"27",X"08",X"7F",X"00",X"AD",X"C6",
		X"1A",X"BD",X"FB",X"50",X"96",X"BE",X"16",X"9A",X"D8",X"0F",X"97",X"D8",X"C6",X"0F",X"BD",X"FA",
		X"DB",X"7E",X"F9",X"22",X"96",X"C1",X"B7",X"08",X"01",X"96",X"C2",X"B7",X"08",X"02",X"7C",X"00",
		X"BD",X"96",X"BF",X"4C",X"97",X"BF",X"44",X"24",X"32",X"DE",X"C3",X"09",X"27",X"1E",X"DF",X"C3",
		X"DE",X"C7",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C1",X"DE",X"C5",X"09",X"27",X"15",X"DF",
		X"C5",X"DE",X"C9",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C2",X"3B",X"86",X"01",X"9A",X"BE",
		X"97",X"BE",X"20",X"E6",X"86",X"02",X"9A",X"BE",X"97",X"BE",X"3B",X"96",X"C7",X"81",X"20",X"25",
		X"09",X"DE",X"C7",X"A6",X"00",X"97",X"C1",X"08",X"DF",X"C7",X"96",X"C9",X"81",X"20",X"25",X"09",
		X"DE",X"C9",X"A6",X"00",X"97",X"C2",X"08",X"DF",X"C9",X"96",X"BF",X"84",X"0E",X"26",X"CC",X"7C",
		X"00",X"C0",X"3B",X"96",X"C0",X"27",X"3E",X"7A",X"00",X"C0",X"96",X"80",X"27",X"06",X"4C",X"27",
		X"03",X"7A",X"00",X"80",X"96",X"81",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"81",X"96",X"82",
		X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"82",X"96",X"83",X"27",X"06",X"4C",X"27",X"03",X"7A",
		X"00",X"83",X"CE",X"00",X"06",X"A6",X"AD",X"27",X"09",X"4A",X"26",X"04",X"6C",X"A7",X"A6",X"B3",
		X"A7",X"AD",X"09",X"26",X"F0",X"39",X"B7",X"08",X"00",X"C6",X"0E",X"BD",X"FB",X"1D",X"84",X"3F",
		X"97",X"BC",X"3B",X"CE",X"FF",X"FF",X"DF",X"00",X"C6",X"4F",X"08",X"86",X"00",X"A7",X"80",X"08",
		X"5A",X"26",X"FA",X"86",X"13",X"97",X"D8",X"39",X"BD",X"FA",X"C0",X"86",X"BF",X"97",X"BB",X"C6",
		X"FF",X"D7",X"82",X"D7",X"83",X"D7",X"B1",X"D7",X"B2",X"D7",X"B3",X"C6",X"17",X"7E",X"FA",X"DB",
		X"86",X"BF",X"97",X"BA",X"C6",X"FF",X"D7",X"80",X"D7",X"81",X"D7",X"AE",X"D7",X"AF",X"D7",X"B0",
		X"C6",X"07",X"7E",X"FA",X"DB",X"7C",X"00",X"BD",X"20",X"04",X"0F",X"7F",X"00",X"BD",X"37",X"36",
		X"C1",X"10",X"2A",X"19",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"08",X"D7",X"03",X"5C",X"32",
		X"97",X"02",X"96",X"BD",X"27",X"FC",X"D7",X"03",X"5A",X"D7",X"03",X"33",X"39",X"86",X"15",X"97",
		X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"10",X"20",X"E3",X"37",X"20",X"E4",X"37",X"86",X"15",X"97",
		X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"14",X"20",X"0D",X"C1",X"10",X"2A",X"EF",X"37",X"86",X"0D",
		X"97",X"03",X"D7",X"02",X"C6",X"0C",X"4F",X"97",X"03",X"97",X"00",X"D7",X"03",X"96",X"02",X"5F",
		X"D7",X"03",X"5A",X"D7",X"00",X"33",X"39",X"0F",X"BD",X"FB",X"1D",X"C6",X"09",X"7F",X"00",X"BD",
		X"84",X"1F",X"81",X"10",X"2A",X"08",X"4A",X"81",X"07",X"2B",X"03",X"BD",X"FB",X"09",X"0E",X"39",
		X"0F",X"BD",X"FB",X"0C",X"C6",X"11",X"20",X"E5",X"17",X"84",X"0F",X"81",X"0D",X"2A",X"08",X"A6",
		X"94",X"AB",X"98",X"A7",X"94",X"20",X"69",X"5A",X"58",X"C4",X"17",X"DE",X"CD",X"A6",X"05",X"36",
		X"DE",X"D1",X"AB",X"94",X"A7",X"94",X"32",X"2B",X"0C",X"24",X"02",X"6C",X"98",X"BD",X"FA",X"DA",
		X"5C",X"A6",X"94",X"20",X"4B",X"25",X"F6",X"6A",X"98",X"20",X"F2",X"6F",X"8C",X"DE",X"CD",X"C1",
		X"A0",X"2B",X"02",X"08",X"08",X"08",X"08",X"08",X"C1",X"C0",X"2B",X"08",X"17",X"84",X"0F",X"81",
		X"08",X"2B",X"01",X"08",X"86",X"00",X"39",X"DF",X"CD",X"DE",X"D1",X"6A",X"90",X"27",X"DC",X"C1",
		X"A0",X"2A",X"10",X"C4",X"1F",X"A6",X"94",X"36",X"DE",X"CD",X"A6",X"03",X"BD",X"FA",X"DA",X"0E",
		X"32",X"08",X"39",X"C1",X"C0",X"2A",X"91",X"A6",X"90",X"44",X"A6",X"94",X"25",X"02",X"A6",X"98",
		X"C4",X"1F",X"BD",X"FA",X"DA",X"0E",X"DE",X"CD",X"A6",X"04",X"39",X"26",X"CA",X"DF",X"CD",X"E6",
		X"00",X"2A",X"03",X"7E",X"FC",X"79",X"C4",X"3F",X"C1",X"20",X"2A",X"11",X"A6",X"01",X"BD",X"FA",
		X"DA",X"0E",X"E6",X"00",X"08",X"08",X"58",X"2B",X"E4",X"A6",X"00",X"08",X"39",X"C4",X"1F",X"17",
		X"84",X"0F",X"81",X"06",X"2A",X"16",X"48",X"C4",X"10",X"1B",X"16",X"A6",X"01",X"97",X"CE",X"A6",
		X"02",X"97",X"CD",X"BD",X"FC",X"BA",X"0E",X"E6",X"00",X"08",X"20",X"D8",X"80",X"08",X"2B",X"29",
		X"DD",X"CF",X"84",X"03",X"C1",X"10",X"2B",X"02",X"8B",X"03",X"16",X"A6",X"01",X"CE",X"00",X"00",
		X"3A",X"D6",X"CF",X"C1",X"04",X"2A",X"0B",X"A6",X"B4",X"A7",X"AE",X"DE",X"CD",X"D6",X"D0",X"7E",
		X"FB",X"EC",X"A7",X"B4",X"DE",X"CD",X"7E",X"FB",X"F2",X"4C",X"27",X"17",X"5C",X"C1",X"10",X"2A",
		X"09",X"96",X"BA",X"A4",X"01",X"97",X"BA",X"7E",X"FB",X"EE",X"96",X"BB",X"A4",X"01",X"97",X"BB",
		X"7E",X"FB",X"EE",X"C1",X"10",X"2A",X"09",X"96",X"BA",X"AA",X"01",X"97",X"BA",X"7E",X"FB",X"EE",
		X"96",X"BB",X"AA",X"01",X"97",X"BB",X"7E",X"FB",X"EE",X"C1",X"F0",X"2A",X"17",X"A6",X"01",X"EE",
		X"02",X"3C",X"DE",X"D1",X"E7",X"8C",X"4C",X"A7",X"90",X"32",X"A7",X"94",X"32",X"A7",X"98",X"DE",
		X"CD",X"86",X"00",X"39",X"5C",X"27",X"12",X"DE",X"D1",X"5C",X"26",X"10",X"DC",X"CD",X"A7",X"9C",
		X"E7",X"A0",X"DE",X"CD",X"EE",X"01",X"86",X"00",X"39",X"86",X"FF",X"39",X"A6",X"9C",X"E6",X"A0",
		X"DD",X"CD",X"DE",X"CD",X"08",X"08",X"08",X"86",X"00",X"39",X"96",X"CE",X"BD",X"FA",X"DA",X"5C",
		X"96",X"CD",X"BD",X"FA",X"DB",X"5C",X"39",X"26",X"03",X"7E",X"FD",X"BD",X"81",X"10",X"2B",X"03",
		X"7E",X"FD",X"41",X"81",X"03",X"2A",X"35",X"97",X"CB",X"96",X"D8",X"8A",X"01",X"16",X"C4",X"FE",
		X"D7",X"D8",X"C6",X"0F",X"BD",X"FA",X"DB",X"86",X"05",X"7F",X"00",X"BD",X"D6",X"BD",X"27",X"FC",
		X"4A",X"26",X"F6",X"D6",X"CB",X"58",X"58",X"CE",X"E9",X"00",X"3A",X"3C",X"EE",X"00",X"DF",X"C7",
		X"38",X"EE",X"02",X"DF",X"C3",X"96",X"BE",X"84",X"02",X"97",X"BE",X"39",X"97",X"CC",X"96",X"D8",
		X"8A",X"02",X"16",X"C4",X"FD",X"D7",X"D8",X"C6",X"0F",X"BD",X"FA",X"DB",X"86",X"05",X"7F",X"00",
		X"BD",X"D6",X"BD",X"27",X"FC",X"4A",X"26",X"F6",X"D6",X"CC",X"58",X"58",X"CE",X"E9",X"00",X"3A",
		X"3C",X"EE",X"00",X"DF",X"C9",X"38",X"EE",X"02",X"DF",X"C5",X"96",X"BE",X"84",X"01",X"97",X"BE",
		X"39",X"16",X"58",X"CE",X"E9",X"34",X"3A",X"EE",X"00",X"81",X"20",X"2B",X"1F",X"81",X"24",X"27",
		X"0A",X"3C",X"36",X"BD",X"FA",X"93",X"BD",X"FA",X"A8",X"32",X"38",X"97",X"A4",X"DF",X"84",X"7F",
		X"00",X"80",X"7F",X"00",X"8C",X"C6",X"B8",X"DA",X"BA",X"D7",X"BA",X"39",X"81",X"12",X"2A",X"11",
		X"DF",X"88",X"97",X"A6",X"7F",X"00",X"82",X"7F",X"00",X"8E",X"86",X"78",X"9A",X"BB",X"97",X"BB",
		X"39",X"81",X"13",X"27",X"EB",X"81",X"16",X"27",X"E7",X"81",X"17",X"2A",X"17",X"DF",X"8A",X"97",
		X"A7",X"7F",X"00",X"83",X"7F",X"00",X"8F",X"86",X"B8",X"9A",X"BB",X"97",X"BB",X"86",X"B8",X"9A",
		X"BA",X"97",X"BA",X"39",X"81",X"17",X"27",X"B3",X"81",X"19",X"27",X"E1",X"DF",X"86",X"97",X"A5",
		X"7F",X"00",X"81",X"7F",X"00",X"8D",X"86",X"78",X"9A",X"BA",X"97",X"BA",X"39",X"CE",X"F4",X"4B",
		X"4F",X"3C",X"36",X"BD",X"FA",X"93",X"BD",X"FA",X"A8",X"32",X"38",X"97",X"A4",X"DF",X"84",X"7F",
		X"00",X"80",X"7F",X"00",X"8C",X"C6",X"B8",X"DA",X"BA",X"D7",X"BA",X"C6",X"B8",X"DA",X"BB",X"D7",
		X"BB",X"39",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"1D",X"4E",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"40",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"40",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"02",X"00",
		X"09",X"0A",X"0C",X"0D",X"0F",X"10",X"12",X"13",X"15",X"16",X"18",X"19",X"1B",X"1C",X"1E",X"1F",
		X"23",X"24",X"26",X"27",X"29",X"2A",X"2C",X"2D",X"2F",X"30",X"32",X"33",X"35",X"36",X"38",X"39",
		X"22",X"5A",X"38",X"30",X"22",X"3B",X"3B",X"20",X"20",X"64",X"65",X"74",X"61",X"20",X"69",X"73",
		X"20",X"20",X"2D",X"2D",X"2D",X"2D",X"48",X"20",X"74",X"6F",X"20",X"2D",X"2D",X"2D",X"2D",X"48",
		X"45",X"4E",X"44",X"48",X"45",X"58",X"3E",X"3E",X"20",X"50",X"61",X"72",X"61",X"6D",X"74",X"65",
		X"72",X"20",X"65",X"72",X"72",X"6F",X"72",X"20",X"3C",X"3C",X"0D",X"00",X"44",X"55",X"4D",X"50",
		X"20",X"4C",X"49",X"53",X"54",X"20",X"50",X"41",X"47",X"45",X"20",X"3D",X"20",X"FF",X"00",X"0D",
		X"0D",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"D1",X"AE",X"02",X"00",X"4D",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"35",X"00",X"FE",X"FF",X"08",X"2E",X"E4",X"41",X"0C",X"00",
		X"F9",X"00",X"F9",X"00",X"F9",X"00",X"F9",X"00",X"FA",X"86",X"F9",X"00",X"F9",X"D4",X"F9",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
