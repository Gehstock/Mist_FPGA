library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tapper_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tapper_bg_bits_2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"BB",X"0A",X"EE",X"26",X"AA",X"26",X"AA",X"0A",X"66",X"02",X"66",X"00",X"A8",
		X"00",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"3F",X"00",X"3F",X"00",X"0F",X"00",X"0F",X"00",X"03",
		X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"05",X"55",X"05",X"55",X"05",X"FF",X"05",X"7F",X"05",X"7F",X"05",X"7F",
		X"05",X"7F",X"05",X"7F",X"05",X"7F",X"05",X"7F",X"15",X"7F",X"FF",X"FF",X"05",X"55",X"05",X"7F",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"FF",X"FF",X"55",X"55",X"55",X"7F",
		X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"D5",X"FF",X"55",X"7F",X"55",X"7F",X"55",X"7F",
		X"9A",X"00",X"96",X"80",X"95",X"A8",X"9A",X"5A",X"99",X"96",X"99",X"65",X"99",X"55",X"95",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F6",X"BF",
		X"FE",X"AB",X"FA",X"AA",X"EA",X"AA",X"FF",X"EA",X"FF",X"FA",X"55",X"7E",X"FF",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AB",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F5",X"6F",X"F5",X"5F",X"F5",X"5B",X"D5",X"5B",X"D5",X"5B",X"D5",X"5B",X"D5",X"5B",X"D5",X"5B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FE",X"EB",X"FA",X"EA",X"EA",X"EA",X"AA",
		X"AB",X"FF",X"EB",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",
		X"FA",X"BF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"F6",X"FF",X"F6",
		X"FF",X"F6",X"FF",X"D6",X"FF",X"D6",X"FF",X"D6",X"FF",X"56",X"FF",X"56",X"FF",X"56",X"FD",X"56",
		X"FD",X"56",X"FD",X"56",X"F5",X"56",X"F5",X"56",X"F5",X"56",X"D5",X"56",X"D5",X"56",X"D5",X"56",
		X"A9",X"55",X"9A",X"55",X"96",X"95",X"95",X"A5",X"9A",X"6A",X"99",X"96",X"99",X"65",X"99",X"55",
		X"95",X"55",X"9A",X"A9",X"9A",X"55",X"99",X"55",X"99",X"55",X"99",X"55",X"99",X"55",X"99",X"55",
		X"95",X"55",X"95",X"55",X"AA",X"AA",X"54",X"05",X"54",X"15",X"50",X"FF",X"50",X"00",X"50",X"05",
		X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",X"00",X"00",
		X"0A",X"A0",X"28",X"A8",X"00",X"28",X"00",X"A0",X"02",X"80",X"0A",X"00",X"2A",X"A8",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"00",X"28",X"02",X"A0",X"00",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"02",X"28",X"0A",X"28",X"08",X"28",X"28",X"28",X"2A",X"A8",X"00",X"28",X"00",X"28",X"00",X"00",
		X"2A",X"A8",X"28",X"00",X"2A",X"A0",X"00",X"28",X"00",X"28",X"2A",X"A8",X"2A",X"A0",X"00",X"00",
		X"02",X"A0",X"0A",X"08",X"28",X"00",X"2A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"2A",X"A8",X"20",X"28",X"00",X"A0",X"02",X"80",X"0A",X"80",X"0A",X"00",X"0A",X"00",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"0A",X"A8",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"00",
		X"2A",X"A0",X"80",X"08",X"8A",X"88",X"88",X"08",X"8A",X"88",X"80",X"08",X"2A",X"A0",X"00",X"00",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A0",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"08",X"0A",X"A0",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"08",X"28",X"08",X"28",X"08",X"28",X"28",X"2A",X"A0",X"00",X"00",
		X"2A",X"A8",X"28",X"00",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",X"2A",X"A8",X"00",X"00",
		X"2A",X"A8",X"28",X"00",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",X"28",X"00",X"00",X"00",
		X"0A",X"A8",X"28",X"00",X"28",X"00",X"28",X"A8",X"28",X"08",X"2A",X"A8",X"0A",X"88",X"00",X"00",
		X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",
		X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",X"00",X"00",
		X"0A",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A0",X"2A",X"A0",X"0A",X"80",X"00",X"00",
		X"28",X"08",X"28",X"28",X"28",X"A0",X"2A",X"A0",X"28",X"28",X"28",X"08",X"28",X"08",X"00",X"00",
		X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"08",X"2A",X"A8",X"00",X"00",
		X"28",X"28",X"28",X"28",X"22",X"88",X"22",X"88",X"20",X"08",X"20",X"08",X"20",X"08",X"00",X"00",
		X"28",X"08",X"2A",X"08",X"2A",X"08",X"22",X"88",X"20",X"88",X"20",X"A8",X"20",X"28",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"08",X"2A",X"A8",X"28",X"00",X"28",X"00",X"28",X"00",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"20",X"08",X"20",X"08",X"20",X"88",X"28",X"A0",X"0A",X"A8",X"00",X"00",
		X"2A",X"A0",X"28",X"28",X"28",X"08",X"2A",X"A8",X"28",X"20",X"28",X"28",X"28",X"08",X"00",X"00",
		X"0A",X"A8",X"28",X"08",X"28",X"00",X"2A",X"A8",X"00",X"28",X"20",X"28",X"2A",X"A0",X"00",X"00",
		X"2A",X"A8",X"2A",X"A8",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"00",X"00",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",X"00",X"00",
		X"20",X"08",X"20",X"08",X"28",X"28",X"08",X"20",X"0A",X"A0",X"02",X"80",X"02",X"80",X"00",X"00",
		X"20",X"08",X"20",X"08",X"20",X"08",X"22",X"88",X"22",X"88",X"2A",X"A8",X"08",X"20",X"00",X"00",
		X"20",X"08",X"28",X"28",X"0A",X"A0",X"02",X"80",X"0A",X"A0",X"28",X"28",X"20",X"08",X"00",X"00",
		X"20",X"08",X"20",X"08",X"28",X"28",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",X"00",X"00",
		X"2A",X"A8",X"20",X"28",X"00",X"A0",X"02",X"80",X"0A",X"00",X"28",X"08",X"2A",X"A8",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"AB",X"F0",
		X"9A",X"F0",X"96",X"80",X"95",X"A8",X"9A",X"5A",X"99",X"96",X"99",X"65",X"99",X"55",X"95",X"55",
		X"95",X"55",X"95",X"55",X"9A",X"A9",X"9A",X"55",X"99",X"55",X"99",X"55",X"99",X"55",X"99",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"A5",X"55",X"65",X"55",
		X"6A",X"AA",X"6A",X"AA",X"65",X"55",X"60",X"00",X"6F",X"57",X"6D",X"55",X"6D",X"55",X"6D",X"55",
		X"6D",X"55",X"6D",X"55",X"AD",X"55",X"FD",X"55",X"FD",X"55",X"FF",X"FF",X"00",X"00",X"FD",X"55",
		X"9A",X"00",X"96",X"80",X"95",X"A8",X"9A",X"5A",X"99",X"96",X"99",X"65",X"99",X"55",X"95",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",
		X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"FE",X"FF",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"3F",X"EA",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"3F",X"0F",X"FA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"03",X"FB",X"FF",X"AB",
		X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FB",X"AF",X"FB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AB",X"FE",X"AB",X"FF",X"AB",X"FF",
		X"00",X"3F",X"0F",X"FA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BE",X"AA",X"FF",X"AA",X"FF",X"AA",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FB",X"AF",X"FB",X"AF",X"FF",X"BF",X"FF",
		X"FE",X"AA",X"FB",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"FB",X"FB",X"FF",X"FF",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"FB",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",
		X"BE",X"AA",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"EB",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BE",X"EB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"EB",X"FF",X"AB",X"FF",X"AB",X"FF",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",
		X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EF",X"FF",X"AB",X"FB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AF",X"AA",X"FF",X"AF",X"FF",X"FF",X"F0",X"FF",X"00",
		X"FF",X"FF",X"BE",X"BF",X"AA",X"AA",X"FA",X"AA",X"FF",X"AA",X"FF",X"FE",X"0F",X"FF",X"00",X"3F",
		X"BF",X"FF",X"AF",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FF",X"EA",
		X"FF",X"FF",X"FF",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"EF",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"BB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0E",
		X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FF",X"AF",X"FF",X"FF",X"F0",X"FC",X"00",
		X"AA",X"FF",X"AF",X"FF",X"FF",X"F0",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"03",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"FE",X"AA",X"FF",X"FA",X"3F",X"FF",X"00",X"FF",X"00",X"03",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FF",X"AA",X"FF",X"FE",X"0F",X"FF",X"00",X"3F",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"FA",X"AB",X"FF",X"EB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"56",X"BF",X"56",X"F5",X"56",X"D5",X"56",X"D5",
		X"56",X"D5",X"56",X"D5",X"56",X"D5",X"56",X"D5",X"56",X"D5",X"56",X"D5",X"56",X"D5",X"56",X"D5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"FB",X"FF",X"EB",X"FF",X"AF",X"FF",X"BD",
		X"AF",X"55",X"BD",X"55",X"B5",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"1B",X"55",X"1B",X"55",X"1B",X"55",X"1B",X"55",X"1B",X"55",X"1B",X"55",X"5B",X"55",X"5B",
		X"D0",X"1B",X"40",X"1B",X"40",X"1B",X"00",X"1B",X"14",X"1B",X"54",X"1B",X"55",X"1B",X"55",X"1B",
		X"FF",X"FB",X"FF",X"EB",X"FF",X"AF",X"FF",X"BD",X"FE",X"B4",X"FA",X"F4",X"FB",X"D0",X"EB",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",
		X"FE",X"BB",X"FA",X"FB",X"FB",X"DB",X"EB",X"5B",X"AF",X"5B",X"BD",X"1B",X"B4",X"1B",X"F4",X"1B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FB",X"FF",X"EB",X"FF",X"AB",X"FF",X"BB",
		X"FE",X"B5",X"FA",X"F5",X"FB",X"D5",X"EB",X"55",X"AF",X"55",X"BD",X"55",X"B5",X"55",X"F5",X"55",
		X"55",X"55",X"55",X"54",X"55",X"04",X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"55",X"5B",X"05",X"5B",X"05",X"5B",X"05",X"5B",X"15",X"5B",X"15",X"5B",X"55",X"5B",X"55",X"5B",
		X"55",X"5B",X"55",X"5B",X"55",X"5B",X"55",X"5B",X"55",X"5B",X"55",X"5B",X"55",X"5B",X"55",X"5B",
		X"54",X"05",X"50",X"05",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",X"05",X"55",
		X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"50",X"55",X"50",
		X"FF",X"FB",X"FF",X"EB",X"FF",X"AF",X"FF",X"BD",X"FE",X"B5",X"FA",X"F5",X"FB",X"D5",X"EB",X"55",
		X"AF",X"55",X"BD",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",
		X"55",X"50",X"55",X"00",X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"05",
		X"05",X"55",X"05",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"6B",X"55",X"6F",X"55",X"AF",X"55",X"BF",X"56",X"BF",X"56",X"FF",X"5A",X"FF",X"5B",X"FF",
		X"6B",X"FF",X"6F",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"5A",X"55",X"5B",
		X"54",X"05",X"50",X"05",X"00",X"05",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"15",X"55",
		X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"54",X"B5",X"54",X"B5",X"50",X"B5",X"50",
		X"B5",X"50",X"B5",X"50",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"6B",X"55",X"6F",X"55",X"AF",X"55",X"BF",X"56",X"BF",X"56",X"FF",X"5A",X"FF",X"5B",X"FF",
		X"6B",X"FF",X"6F",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"46",X"55",X"1A",X"55",X"1B",
		X"B5",X"55",X"B4",X"55",X"B4",X"55",X"B4",X"55",X"B4",X"55",X"B4",X"55",X"B4",X"55",X"B4",X"15",
		X"B4",X"15",X"B4",X"15",X"B4",X"15",X"B4",X"05",X"B4",X"05",X"B4",X"00",X"B4",X"00",X"B4",X"00",
		X"B4",X"00",X"B4",X"00",X"B4",X"01",X"B4",X"01",X"B4",X"06",X"B4",X"06",X"B4",X"1A",X"B4",X"1B",
		X"B4",X"6B",X"B4",X"6F",X"B5",X"AF",X"B5",X"BF",X"B6",X"BF",X"B6",X"FF",X"BA",X"FF",X"BB",X"FF",
		X"BB",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"6B",X"FF",X"6F",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"54",X"6B",X"50",X"6F",X"41",X"AF",X"41",X"BF",X"06",X"BF",X"06",X"FF",X"1A",X"FF",X"1B",X"FF",
		X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",
		X"AB",X"A5",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"95",
		X"56",X"AE",X"5A",X"BE",X"5A",X"BA",X"5A",X"B9",X"6A",X"F9",X"6A",X"E9",X"6A",X"E5",X"AB",X"E5",
		X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"AB",X"55",X"AB",X"55",X"AB",X"56",X"AF",X"56",X"AE",
		X"F9",X"5E",X"E9",X"5E",X"E5",X"5E",X"E5",X"5E",X"A5",X"5E",X"95",X"5E",X"95",X"5E",X"95",X"5E",
		X"AB",X"AE",X"AB",X"9E",X"AF",X"9E",X"AE",X"9E",X"AE",X"5E",X"BE",X"5E",X"BA",X"5E",X"B9",X"5E",
		X"56",X"AE",X"5A",X"BE",X"5A",X"BA",X"5A",X"BA",X"6A",X"FA",X"6A",X"EE",X"6A",X"EE",X"AB",X"EE",
		X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"6A",
		X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",
		X"55",X"AA",X"56",X"A9",X"56",X"A9",X"56",X"A9",X"5A",X"A5",X"5A",X"A5",X"5A",X"A5",X"6A",X"95",
		X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"56",X"A9",X"56",X"A9",X"56",X"A9",
		X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"56",
		X"6A",X"95",X"6A",X"95",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",
		X"5A",X"A5",X"5A",X"A5",X"5A",X"A5",X"6A",X"95",X"6A",X"95",X"6A",X"95",X"AA",X"55",X"AA",X"55",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"AA",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"AB",X"95",X"AB",X"95",X"AB",X"95",X"AB",X"97",X"AB",X"97",X"AB",X"97",X"AB",X"9F",X"AB",X"9E",
		X"AB",X"9E",X"AB",X"BE",X"AB",X"BA",X"AB",X"B8",X"AB",X"F8",X"AB",X"E8",X"AB",X"E0",X"57",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"E8",X"00",X"E0",X"00",X"E0",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"57",X"A0",X"57",X"80",X"5F",X"80",X"5E",X"80",X"5E",X"00",X"7E",X"00",X"7A",X"00",X"78",X"00",
		X"55",X"5E",X"55",X"7E",X"55",X"7A",X"55",X"78",X"55",X"F8",X"55",X"E8",X"55",X"E0",X"57",X"E0",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"5C",X"05",X"F0",X"07",X"F0",X"17",X"C0",X"14",X"80",X"50",X"A0",X"50",X"A8",X"50",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"28",X"00",X"A8",X"00",X"A8",X"00",
		X"A8",X"00",X"A8",X"00",X"28",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"AA",X"50",X"A8",X"50",X"A0",X"10",X"80",X"14",X"00",X"04",X"00",X"05",X"00",X"01",X"40",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5C",X"55",X"F0",X"57",X"F0",X"57",X"C0",X"54",X"80",X"50",X"A0",X"50",X"A8",X"50",X"AA",
		X"A9",X"5C",X"A5",X"F0",X"A7",X"F0",X"97",X"C0",X"94",X"80",X"50",X"A0",X"50",X"A8",X"50",X"AA",
		X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"01",X"08",X"01",X"28",X"00",X"A8",X"00",X"A8",X"00",
		X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"01",X"08",X"01",X"28",X"00",X"A8",X"00",X"A8",X"00",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"0A",X"55",X"02",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"01",X"55",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"80",X"55",X"00",
		X"00",X"01",X"00",X"05",X"00",X"14",X"01",X"50",X"55",X"40",X"54",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"11",
		X"40",X"00",X"50",X"00",X"14",X"00",X"05",X"40",X"01",X"55",X"00",X"15",X"00",X"05",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"3C",X"00",X"7C",X"00",X"40",X"00",X"50",X"00",
		X"40",X"44",X"11",X"10",X"04",X"40",X"04",X"10",X"04",X"40",X"04",X"10",X"04",X"40",X"04",X"10",
		X"03",X"80",X"03",X"00",X"00",X"00",X"0F",X"00",X"3C",X"00",X"7C",X"00",X"40",X"00",X"50",X"00",
		X"40",X"00",X"50",X"00",X"14",X"00",X"05",X"40",X"01",X"55",X"03",X"95",X"03",X"95",X"03",X"81",
		X"03",X"80",X"03",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"05",X"00",X"14",X"01",X"50",X"55",X"40",X"57",X"80",X"43",X"80",X"13",X"80",
		X"40",X"44",X"10",X"10",X"04",X"40",X"04",X"10",X"04",X"40",X"55",X"55",X"00",X"00",X"00",X"00",
		X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"02",X"80",X"55",X"55",X"00",X"00",X"00",X"00",
		X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"02",X"80",X"25",X"55",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",
		X"1F",X"FD",X"1F",X"FD",X"1F",X"FD",X"DF",X"FD",X"D7",X"FD",X"F7",X"F4",X"F5",X"D4",X"FD",X"50",
		X"A9",X"50",X"A5",X"D4",X"A7",X"F4",X"97",X"FD",X"9F",X"FD",X"1F",X"FD",X"1F",X"FD",X"1F",X"FD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"00",X"40",X"00",X"40",X"00",X"7F",X"FF",X"7F",X"FF",X"1F",X"FF",X"1F",X"FF",X"07",X"FF",
		X"05",X"AA",X"16",X"AA",X"1A",X"AA",X"5A",X"AA",X"6A",X"AA",X"40",X"00",X"40",X"00",X"40",X"00",
		X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"28",X"02",X"08",X"08",X"0A",X"28",X"02",X"A0",
		X"56",X"A0",X"5A",X"28",X"58",X"08",X"68",X"02",X"60",X"02",X"20",X"02",X"20",X"02",X"20",X"02",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"20",X"00",X"20",X"00",X"08",X"00",
		X"09",X"55",X"25",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"AF",
		X"02",X"80",X"02",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
		X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
		X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"02",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5E",X"AA",X"5E",X"AA",X"5E",X"AA",X"5E",X"AA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AF",X"AA",X"BD",X"AA",X"B5",X"AA",X"B5",X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"95",X"5E",X"55",X"5E",X"55",X"5E",X"55",X"5E",X"FF",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AF",X"D5",X"BD",X"55",X"B5",X"55",X"B5",X"55",X"BF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FA",X"AA",X"BE",X"9A",X"AE",
		X"FF",X"FF",X"FF",X"FE",X"BF",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",
		X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",X"FA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"3F",X"EA",X"FA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"03",X"FE",X"FF",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",X"AB",X"F0",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"3F",X"EA",X"FA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",X"FA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"03",X"FE",X"FF",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"AB",X"FF",X"AA",X"FF",X"AB",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",
		X"AB",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FB",X"FF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"BF",X"FE",X"BF",X"FE",X"AF",X"FE",X"AF",X"FE",X"AF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"FF",X"EB",X"FF",X"EF",X"FF",X"EF",X"FB",X"EF",X"EA",
		X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"BF",X"FE",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"BF",X"FF",X"AF",X"EB",X"BF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FE",X"FF",X"FE",X"FF",X"FB",X"FE",X"FB",X"FF",X"FB",X"FF",
		X"AA",X"BF",X"AA",X"AF",X"FE",X"AF",X"FF",X"BF",X"FF",X"FF",X"BF",X"EF",X"FF",X"EF",X"FE",X"AF",
		X"EA",X"AA",X"EA",X"AA",X"AB",X"FF",X"EF",X"FF",X"EF",X"FF",X"EF",X"EF",X"EF",X"FF",X"EB",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"EA",X"FF",X"EB",X"FF",X"EB",X"FF",X"EF",X"FA",X"EF",X"FF",X"EF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"FA",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FA",X"BF",
		X"AA",X"AB",X"AA",X"AB",X"FE",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"BF",X"AB",X"AA",X"AB",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"EB",X"EB",X"EB",X"EB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EF",X"EA",X"EF",X"FA",X"EF",X"FF",X"EB",X"FF",X"AA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EB",X"FF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"EF",X"AF",X"EF",X"FF",X"EF",X"FF",X"BF",X"FE",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EB",X"FA",X"EB",X"FE",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FE",X"AF",X"FE",X"AF",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EF",X"EB",X"EF",X"FB",X"FF",X"FF",X"FB",X"FF",X"FA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FE",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",X"AB",X"F0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"EA",X"F0",X"FF",X"00",X"03",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"0F",X"FA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3B",X"00",X"3F",X"00",X"00",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",X"AB",X"F0",X"BF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",X"AB",X"F0",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",X"AB",X"F0",X"BF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"AA",X"FF",X"AA",X"03",X"FE",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"3F",X"EA",X"00",X"FF",X"00",X"03",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"0F",X"FA",
		X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"AA",X"FF",X"AA",X"03",X"FE",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"3F",X"EA",X"00",X"FF",X"00",X"03",X"00",X"00",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"FE",X"AB",X"0F",X"FB",
		X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"EB",X"FA",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"3B",X"00",X"3A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",
		X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FD",X"55",X"FD",X"55",X"FD",X"55",
		X"FD",X"95",X"FD",X"97",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",
		X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",
		X"FD",X"9F",X"F5",X"9F",X"D5",X"9F",X"55",X"9F",X"FF",X"FF",X"D5",X"55",X"FD",X"55",X"FD",X"55",
		X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"7D",X"9F",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",
		X"56",X"A5",X"F5",X"97",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",X"FD",X"9F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FC",X"7F",X"FC",X"5F",X"F0",X"5F",X"F0",X"57",X"C0",X"57",X"C0",X"55",X"00",X"55",X"00",
		X"55",X"40",X"55",X"40",X"55",X"50",X"95",X"50",X"95",X"54",X"A5",X"54",X"E5",X"55",X"E9",X"55",
		X"F9",X"55",X"7A",X"55",X"7E",X"55",X"5E",X"95",X"5F",X"95",X"57",X"A5",X"57",X"E5",X"55",X"E9",
		X"40",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"00",
		X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",
		X"55",X"F9",X"55",X"FA",X"55",X"FE",X"55",X"FE",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"EA",
		X"AD",X"55",X"BD",X"55",X"B5",X"45",X"B5",X"01",X"B0",X"00",X"F0",X"00",X"C0",X"C0",X"CC",X"F3",
		X"55",X"55",X"45",X"55",X"55",X"55",X"50",X"54",X"00",X"00",X"3F",X"F0",X"FA",X"B0",X"EA",X"BF",
		X"55",X"55",X"51",X"55",X"15",X"55",X"05",X"01",X"00",X"00",X"0C",X"00",X"00",X"0C",X"C0",X"FC",
		X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"54",X"00",X"00",X"3F",X"F0",X"3A",X"BF",X"FA",X"AB",
		X"55",X"EA",X"55",X"FA",X"15",X"7A",X"01",X"7A",X"00",X"3A",X"0C",X"3E",X"00",X"0E",X"FC",X"CE",
		X"EA",X"AA",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AA",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FB",X"FA",X"AA",X"EA",X"AB",X"AA",X"FF",X"AA",X"AA",X"AA",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",
		X"FF",X"EF",X"FF",X"BF",X"EF",X"FF",X"EB",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"96",X"96",
		X"EA",X"AB",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"AA",X"AD",X"AA",X"AD",X"AA",X"AD",X"AA",X"AD",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",
		X"55",X"55",X"51",X"55",X"55",X"45",X"44",X"15",X"00",X"00",X"00",X"C0",X"C0",X"03",X"F3",X"CF",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"AB",X"FA",X"AA",X"EA",X"AA",X"AA",X"6A",X"AA",X"9A",X"5A",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"AA",X"BD",X"AA",X"B5",X"AA",X"F5",X"AF",X"D4",X"FC",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"55",X"55",X"55",X"55",X"14",X"55",X"05",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"AA",X"7A",X"AA",X"7E",X"AA",X"5F",X"EA",X"00",X"FE",X"00",X"0E",X"00",X"0E",X"00",X"0E",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"AE",X"AB",X"AF",X"AB",X"AB",X"FF",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"FF",X"FF",X"96",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FA",X"AA",X"BF",
		X"AA",X"AF",X"AA",X"BD",X"AA",X"B5",X"AA",X"B4",X"AA",X"B0",X"AA",X"B0",X"AA",X"B0",X"AA",X"BC",
		X"D5",X"55",X"55",X"55",X"55",X"55",X"41",X"FF",X"00",X"EA",X"03",X"EA",X"03",X"AF",X"0E",X"F0",
		X"69",X"57",X"55",X"55",X"54",X"55",X"D5",X"05",X"F0",X"00",X"BC",X"00",X"EC",X"00",X"3C",X"CF",
		X"EA",X"AA",X"FA",X"AA",X"7E",X"AA",X"5E",X"AA",X"0E",X"AA",X"0E",X"AA",X"CE",X"AA",X"0F",X"AA",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"E9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"FE",X"AA",X"FA",X"AA",X"EA",X"9B",X"EA",X"6B",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"BF",X"AF",X"AE",X"AA",X"AE",X"AA",X"AE",X"99",X"AE",X"96",
		X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"5B",X"AA",
		X"AA",X"D5",X"AA",X"D5",X"AA",X"D4",X"AA",X"C1",X"AA",X"C1",X"AA",X"F0",X"AA",X"B0",X"AA",X"BC",
		X"57",X"EA",X"55",X"EA",X"55",X"FA",X"41",X"7E",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AD",X"55",X"AD",X"55",X"BD",X"51",X"F5",X"14",X"C0",X"10",X"00",X"00",X"3C",X"00",X"FC",X"00",
		X"57",X"AA",X"57",X"AA",X"57",X"AA",X"07",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F0",X"0F",X"BF",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"FA",X"AF",X"BA",X"BE",X"BB",X"FA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"FA",X"AA",X"AA",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"AF",X"FA",X"6A",X"BE",
		X"56",X"5F",X"55",X"57",X"51",X"57",X"40",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"3C",
		X"55",X"55",X"55",X"55",X"5F",X"54",X"FF",X"F5",X"EA",X"BC",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",
		X"56",X"75",X"55",X"55",X"15",X"55",X"50",X"15",X"00",X"07",X"00",X"0F",X"00",X"0E",X"3C",X"0E",
		X"BF",X"FF",X"B5",X"55",X"B5",X"55",X"B5",X"41",X"BF",X"00",X"AB",X"C0",X"AA",X"F3",X"AA",X"B0",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BE",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",
		X"FF",X"CE",X"FF",X"FE",X"FB",X"FE",X"FE",X"BE",X"AA",X"AE",X"AA",X"AE",X"9A",X"AE",X"56",X"AF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"AE",X"EA",X"AA",X"EA",X"AA",X"AA",X"9A",X"A6",X"6A",
		X"55",X"55",X"55",X"55",X"54",X"55",X"15",X"07",X"00",X"0F",X"00",X"3E",X"03",X"FA",X"FF",X"AA",
		X"AA",X"AF",X"EA",X"BD",X"FE",X"F5",X"5F",X"D4",X"00",X"00",X"00",X"00",X"00",X"30",X"FC",X"FC",
		X"55",X"97",X"55",X"57",X"55",X"55",X"05",X"15",X"00",X"00",X"00",X"00",X"30",X"0F",X"0F",X"0F",
		X"AA",X"B5",X"AA",X"B5",X"AA",X"B5",X"AA",X"B5",X"AA",X"B0",X"AA",X"B0",X"AA",X"B0",X"AA",X"B0",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BA",X"AA",X"FA",X"AA",X"EA",X"AA",X"E5",
		X"FF",X"FE",X"FB",X"FE",X"FF",X"FE",X"AF",X"FE",X"AB",X"AE",X"6A",X"AE",X"AA",X"AE",X"A9",X"AE",
		X"AF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"BF",X"AA",X"B5",X"EA",X"B5",X"EA",X"B5",X"EA",X"BF",X"FA",X"AB",X"3A",X"AA",X"3A",X"AA",
		X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"FA",X"AA",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"55",X"55",X"55",X"55",X"41",X"01",X"40",X"00",X"00",X"C3",X"00",X"F0",X"30",X"B0",X"3F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"BE",X"AB",X"FA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"BA",X"BF",X"BB",X"FA",X"BF",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FE",X"6A",X"AF",X"A5",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"BE",X"AA",
		X"5F",X"AA",X"57",X"AA",X"57",X"EA",X"55",X"EA",X"00",X"EA",X"00",X"FA",X"30",X"3A",X"C0",X"3A",
		X"55",X"55",X"55",X"55",X"55",X"15",X"F5",X"40",X"BC",X"00",X"AF",X"00",X"AB",X"00",X"AB",X"C3",
		X"B5",X"55",X"55",X"55",X"51",X"5F",X"55",X"FF",X"03",X"EA",X"0F",X"AA",X"0E",X"AA",X"0E",X"AA",
		X"BC",X"FF",X"BF",X"FE",X"BF",X"FF",X"BF",X"BE",X"BA",X"AA",X"BA",X"9A",X"BA",X"AA",X"BA",X"56",
		X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"BE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"EA",X"AB",X"EA",X"AB",X"AA",X"AB",X"A5",
		X"FF",X"FA",X"FE",X"FA",X"BF",X"FA",X"AF",X"FA",X"AB",X"BA",X"6A",X"BA",X"AA",X"BA",X"A6",X"FA",
		X"55",X"EA",X"55",X"EA",X"45",X"EA",X"17",X"EA",X"0F",X"AA",X"3E",X"AA",X"FA",X"AA",X"AA",X"AA",
		X"AF",X"55",X"BD",X"55",X"F5",X"55",X"D5",X"14",X"00",X"00",X"0C",X"00",X"00",X"03",X"3C",X"FF",
		X"5F",X"AA",X"57",X"EA",X"15",X"FE",X"05",X"5F",X"00",X"00",X"00",X"00",X"0F",X"00",X"CF",X"FC",
		X"B5",X"55",X"B5",X"51",X"B5",X"55",X"B5",X"04",X"B0",X"00",X"B3",X"00",X"B0",X"00",X"B0",X"30",
		X"BC",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"EB",X"BA",X"AA",X"FA",X"AA",X"EA",X"9A",X"E9",X"6A",
		X"FE",X"AF",X"FE",X"AA",X"BE",X"AA",X"FE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"6E",X"AA",
		X"AA",X"F5",X"AB",X"D5",X"AF",X"51",X"AD",X"54",X"BC",X"00",X"B0",X"00",X"B0",X"03",X"B0",X"F0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"FF",X"FE",X"AA",X"AA",X"AA",
		X"65",X"55",X"55",X"55",X"55",X"FF",X"17",X"EB",X"0F",X"AA",X"0E",X"AA",X"0E",X"AA",X"CF",X"FF",
		X"55",X"5F",X"55",X"57",X"51",X"57",X"D4",X"15",X"F0",X"00",X"B3",X"00",X"B0",X"F0",X"F0",X"FC",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"A7",X"FE",X"5A",X"AE",
		X"FF",X"FF",X"FF",X"EF",X"EA",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",
		X"BF",X"FF",X"BF",X"BF",X"BF",X"FF",X"BF",X"AA",X"BA",X"AA",X"BA",X"6A",X"BA",X"A9",X"BA",X"56",
		X"B5",X"55",X"B5",X"55",X"BD",X"45",X"AD",X"50",X"AC",X"00",X"AF",X"00",X"AB",X"C0",X"AA",X"F0",
		X"5F",X"AA",X"57",X"AA",X"57",X"EA",X"05",X"FE",X"00",X"0F",X"00",X"00",X"0C",X"00",X"00",X"30",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"FD",X"AF",X"D5",X"FC",X"04",X"00",X"00",X"00",X"03",X"00",X"CF",
		X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"C3",X"FC",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"0F",X"FE",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AF",X"EA",X"AD",X"EA",X"AD",X"FA",X"AC",X"3A",X"AF",X"3A",X"AA",X"3E",X"AA",
		X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",
		X"7E",X"AA",X"5E",X"AA",X"5E",X"AA",X"5E",X"AA",X"3E",X"BF",X"FA",X"B0",X"EA",X"B0",X"AA",X"B0",
		X"AD",X"55",X"AD",X"55",X"BD",X"54",X"F5",X"41",X"C0",X"00",X"00",X"00",X"0C",X"00",X"F0",X"00",
		X"AF",X"FF",X"AF",X"FF",X"AF",X"EF",X"AF",X"FA",X"AE",X"AA",X"AE",X"AA",X"AE",X"A9",X"AE",X"5A",
		X"AB",X"F5",X"FF",X"55",X"55",X"55",X"55",X"04",X"00",X"00",X"F0",X"00",X"BC",X"00",X"AC",X"F3",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AB",X"EB",X"BF",X"AB",X"FA",
		X"67",X"55",X"55",X"55",X"15",X"7F",X"05",X"FF",X"03",X"EC",X"03",X"AC",X"33",X"AF",X"C3",X"AB",
		X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"6B",X"AA",
		X"57",X"AA",X"57",X"AA",X"57",X"AA",X"17",X"EA",X"00",X"FF",X"00",X"03",X"3C",X"03",X"FC",X"03",
		X"55",X"9F",X"54",X"57",X"55",X"55",X"41",X"05",X"00",X"00",X"00",X"00",X"00",X"C3",X"0F",X"03",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"78",X"01",X"78",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"78",X"01",X"78",X"01",X"7B",X"01",X"7B",X"01",X"7B",X"01",X"FB",X"01",X"E6",X"01",X"E6",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"C1",X"40",X"C1",X"40",X"C1",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"02",X"80",X"09",X"A0",X"05",X"60",X"05",X"60",
		X"03",X"E6",X"03",X"96",X"03",X"96",X"0F",X"96",X"0E",X"56",X"0E",X"56",X"3E",X"56",X"39",X"56",
		X"C1",X"0C",X"C1",X"3F",X"C0",X"F5",X"CA",X"D5",X"CB",X"D5",X"CB",X"57",X"CF",X"5F",X"CD",X"5D",
		X"00",X"00",X"F0",X"00",X"FF",X"00",X"5F",X"F0",X"55",X"FF",X"D5",X"5F",X"FD",X"57",X"FF",X"57",
		X"C0",X"0B",X"C0",X"2F",X"C0",X"2F",X"C0",X"BF",X"C5",X"BE",X"C6",X"FE",X"C2",X"F5",X"CB",X"F9",
		X"E0",X"00",X"F8",X"00",X"FE",X"00",X"AF",X"80",X"57",X"E0",X"55",X"F9",X"55",X"7E",X"55",X"7E",
		X"55",X"5B",X"F5",X"67",X"FF",X"6F",X"5F",X"FF",X"55",X"FF",X"D5",X"5F",X"FD",X"57",X"FF",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"68",X"05",X"7A",X"09",X"BE",X"02",X"8E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"43",X"01",X"43",X"01",X"43",X"01",X"4F",
		X"39",X"56",X"F9",X"56",X"E5",X"56",X"E5",X"5A",X"E5",X"5B",X"95",X"5B",X"95",X"5F",X"FD",X"5D",
		X"FD",X"7F",X"F5",X"7D",X"F5",X"7F",X"D5",X"5F",X"D7",X"D5",X"57",X"FD",X"5F",X"FF",X"5F",X"FF",
		X"5F",X"5C",X"5F",X"5C",X"7D",X"70",X"FD",X"70",X"F5",X"C0",X"55",X"C0",X"D7",X"00",X"D7",X"00",
		X"EF",X"F5",X"EF",X"FE",X"FF",X"BF",X"FE",X"AF",X"FE",X"5B",X"F9",X"55",X"E5",X"55",X"E5",X"55",
		X"55",X"7E",X"55",X"78",X"95",X"F8",X"EB",X"E0",X"0F",X"80",X"0E",X"00",X"5E",X"00",X"B8",X"00",
		X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",
		X"01",X"4F",X"01",X"4D",X"01",X"75",X"01",X"D4",X"03",X"53",X"0D",X"4F",X"35",X"3F",X"35",X"F7",
		X"5F",X"AA",X"57",X"EA",X"15",X"FA",X"C5",X"7E",X"F1",X"5F",X"5C",X"57",X"D7",X"15",X"5F",X"35",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"7E",X"AA",
		X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",
		X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"0E",X"00",X"0E",X"00",X"5E",X"05",X"5F",X"15",X"55",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"51",X"40",X"55",X"40",X"55",X"40",
		X"35",X"7F",X"0D",X"5F",X"03",X"57",X"01",X"D5",X"01",X"B5",X"01",X"AD",X"01",X"4F",X"01",X"4E",
		X"DC",X"DA",X"F3",X"5A",X"FD",X"55",X"F5",X"4F",X"55",X"3D",X"57",X"F5",X"57",X"FD",X"D5",X"FF",
		X"5F",X"FF",X"D7",X"EA",X"15",X"FA",X"C5",X"7E",X"71",X"5F",X"FC",X"57",X"5F",X"D5",X"7F",X"D5",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"D5",X"55",X"F5",X"55",X"7F",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"54",X"55",X"50",X"FF",X"F0",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"15",X"55",X"15",X"55",X"41",X"55",X"50",X"55",X"54",X"00",X"56",X"55",X"16",X"95",X"06",X"A6",
		X"55",X"40",X"55",X"40",X"54",X"10",X"50",X"50",X"01",X"50",X"65",X"50",X"A5",X"40",X"A5",X"00",
		X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",X"01",X"4E",
		X"35",X"7F",X"0D",X"5F",X"0F",X"57",X"0E",X"D5",X"0E",X"B5",X"0E",X"AD",X"0F",X"AB",X"0F",X"FF",
		X"FF",X"55",X"FD",X"55",X"F5",X"57",X"D5",X"5F",X"55",X"7B",X"55",X"EB",X"57",X"AF",X"DF",X"FF",
		X"5A",X"AF",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"FA",X"AF",X"FF",X"FF",
		X"EA",X"F0",X"AA",X"B0",X"AA",X"B0",X"AA",X"B0",X"AA",X"B0",X"AA",X"B0",X"EA",X"F0",X"FF",X"F0",
		X"FA",X"AF",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"FA",X"AF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"03",X"FD",
		X"42",X"AA",X"56",X"A6",X"56",X"95",X"56",X"55",X"55",X"55",X"05",X"55",X"40",X"55",X"14",X"00",
		X"A0",X"10",X"A5",X"50",X"A5",X"50",X"65",X"50",X"55",X"50",X"55",X"00",X"50",X"00",X"01",X"40",
		X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"00",X"FF",X"00",X"03",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"D5",X"55",X"F5",X"55",X"FF",X"FF",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"55",X"40",X"57",X"40",X"FF",X"C0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"45",X"01",X"45",X"01",X"45",X"01",X"55",X"01",X"59",X"01",X"59",X"01",X"59",X"01",X"69",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"69",X"01",X"69",X"01",X"A9",X"01",X"89",X"05",X"89",X"06",X"89",X"06",X"49",X"16",X"49",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"41",X"01",X"41",X"01",X"41",
		X"1A",X"49",X"1B",X"49",X"5B",X"49",X"69",X"49",X"6F",X"49",X"6F",X"49",X"AF",X"49",X"BF",X"49",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"02",X"A0",X"0A",X"54",X"09",X"45",X"09",X"15",X"09",X"45",X"0A",X"54",X"02",X"A0",X"00",X"00",
		X"01",X"40",X"51",X"40",X"75",X"40",X"55",X"40",X"55",X"40",X"51",X"40",X"01",X"40",X"01",X"40",
		X"01",X"45",X"01",X"46",X"01",X"46",X"01",X"56",X"01",X"5A",X"01",X"5B",X"01",X"5B",X"01",X"6B",
		X"BF",X"59",X"BF",X"49",X"F7",X"49",X"F5",X"49",X"D7",X"59",X"DF",X"59",X"7F",X"59",X"7D",X"49",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"6F",X"01",X"6F",X"01",X"AF",X"01",X"B7",X"05",X"B5",X"06",X"BD",X"06",X"FD",X"16",X"DE",
		X"57",X"49",X"DD",X"49",X"5D",X"49",X"DD",X"59",X"D5",X"49",X"DF",X"59",X"5D",X"49",X"95",X"49",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"41",X"01",X"41",X"01",X"41",
		X"1A",X"D5",X"1B",X"55",X"5B",X"55",X"6B",X"D5",X"6F",X"F5",X"6F",X"75",X"AD",X"55",X"AF",X"55",
		X"55",X"49",X"57",X"49",X"55",X"49",X"55",X"49",X"57",X"49",X"55",X"59",X"55",X"49",X"55",X"49",
		X"01",X"45",X"01",X"46",X"01",X"46",X"01",X"56",X"01",X"5A",X"01",X"58",X"01",X"58",X"01",X"68",
		X"AF",X"55",X"AD",X"55",X"65",X"75",X"6D",X"D5",X"6F",X"D5",X"6F",X"55",X"6D",X"75",X"6D",X"D5",
		X"55",X"49",X"5D",X"49",X"57",X"59",X"55",X"49",X"55",X"49",X"5F",X"49",X"55",X"49",X"77",X"49",
		X"01",X"6C",X"01",X"6C",X"01",X"AC",X"01",X"BC",X"05",X"BC",X"06",X"BC",X"06",X"F4",X"16",X"D4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"54",X"FD",X"40",X"F5",X"00",X"C4",X"00",X"C4",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"FF",X"3F",X"F5",
		X"FF",X"F5",X"F7",X"F5",X"F5",X"F5",X"F5",X"D5",X"F5",X"55",X"F5",X"55",X"D5",X"5F",X"55",X"FF",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"7F",X"F5",X"5F",X"F5",X"5F",X"F5",X"57",X"F5",X"57",X"F5",X"55",
		X"D0",X"3F",X"D0",X"FF",X"D0",X"FF",X"D7",X"FD",X"D7",X"D5",X"D5",X"55",X"55",X"5E",X"55",X"FE",
		X"FA",X"BD",X"EA",X"AD",X"AA",X"AB",X"AA",X"AF",X"6A",X"FB",X"AB",X"DF",X"AB",X"FF",X"BA",X"FA",
		X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"FF",
		X"FD",X"55",X"FF",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"FA",X"D4",X"3A",X"04",X"3E",X"C5",X"0F",X"F1",X"03",X"F1",X"40",X"FC",X"50",X"FF",X"D5",
		X"FA",X"AA",X"BA",X"AA",X"BE",X"AA",X"BE",X"AA",X"FB",X"AA",X"FB",X"EA",X"3B",X"BA",X"7B",X"AF",
		X"BF",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",X"A6",X"6B",X"A6",X"6B",X"A6",X"6B",X"AA",X"AB",
		X"FB",X"BF",X"FA",X"BF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"AF",X"FA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"FC",X"1B",X"FC",X"5B",X"F4",X"6B",X"D4",X"6D",X"DC",X"6D",X"5C",X"6F",X"5C",X"6F",X"DC",
		X"6F",X"F7",X"6F",X"57",X"6D",X"5F",X"6F",X"D5",X"6F",X"57",X"6D",X"5F",X"6F",X"57",X"67",X"D5",
		X"55",X"09",X"57",X"09",X"DF",X"29",X"D7",X"25",X"DC",X"24",X"5C",X"A4",X"5C",X"94",X"54",X"90",
		X"6F",X"D5",X"6D",X"55",X"6F",X"54",X"6D",X"5C",X"6D",X"54",X"65",X"54",X"6D",X"54",X"65",X"54",
		X"65",X"55",X"65",X"57",X"65",X"D7",X"6F",X"D5",X"6F",X"D5",X"6F",X"5D",X"67",X"5F",X"65",X"57",
		X"72",X"90",X"72",X"50",X"C2",X"40",X"CA",X"40",X"49",X"40",X"09",X"40",X"29",X"40",X"25",X"40",
		X"65",X"54",X"6D",X"54",X"6F",X"54",X"6D",X"5C",X"65",X"7C",X"65",X"5C",X"65",X"7C",X"65",X"5C",
		X"6D",X"7C",X"6F",X"7C",X"6F",X"5C",X"6F",X"70",X"6D",X"72",X"6D",X"F2",X"6F",X"C2",X"6F",X"CA",
		X"25",X"40",X"A5",X"40",X"95",X"40",X"91",X"40",X"91",X"40",X"51",X"40",X"41",X"40",X"41",X"40",
		X"6D",X"5C",X"6D",X"54",X"6F",X"54",X"6F",X"5C",X"6F",X"5C",X"6D",X"54",X"65",X"D4",X"65",X"D4",
		X"6F",X"C9",X"6F",X"09",X"6F",X"29",X"6F",X"25",X"6C",X"24",X"6C",X"A4",X"6C",X"94",X"60",X"90",
		X"41",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"65",X"40",X"65",X"40",X"55",X"40",X"51",X"40",X"51",X"40",X"51",X"40",X"41",X"40",X"41",X"40",
		X"62",X"90",X"62",X"50",X"62",X"40",X"6A",X"40",X"69",X"40",X"69",X"40",X"69",X"40",X"65",X"40",
		X"67",X"DC",X"6F",X"5C",X"6F",X"7C",X"6D",X"7C",X"6F",X"7C",X"6F",X"DC",X"6F",X"5C",X"6F",X"74",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"10",X"00",X"50",X"04",X"54",X"05",X"54",X"05",X"54",
		X"15",X"50",X"04",X"50",X"00",X"10",X"00",X"10",X"00",X"50",X"04",X"50",X"00",X"10",X"00",X"00",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"02",X"AA",
		X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"A1",X"40",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AB",X"00",X"03",
		X"BD",X"40",X"BD",X"40",X"BD",X"40",X"FD",X"40",X"FD",X"40",X"FD",X"40",X"DD",X"40",X"FD",X"40",
		X"00",X"03",X"04",X"03",X"05",X"03",X"01",X"43",X"05",X"03",X"15",X"03",X"01",X"03",X"00",X"03",
		X"DD",X"40",X"7D",X"40",X"DD",X"40",X"7D",X"40",X"DD",X"40",X"7D",X"40",X"DD",X"40",X"7D",X"40",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"FD",X"40",X"7D",X"40",X"F1",X"40",X"F1",X"40",X"F1",X"40",X"C1",X"40",X"C1",X"40",X"C1",X"40",
		X"AA",X"AA",X"80",X"00",X"8F",X"33",X"8C",X"33",X"8C",X"33",X"8C",X"33",X"8F",X"3F",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"3C",X"FC",X"30",X"30",X"3C",X"30",X"0C",X"30",X"3C",X"30",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"FC",X"C3",X"CC",X"FF",X"CC",X"FF",X"CC",X"C3",X"FC",X"C3",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"3C",X"FC",X"30",X"CC",X"3C",X"FC",X"30",X"CC",X"3C",X"CC",X"AA",X"AA",
		X"AA",X"AA",X"02",X"00",X"F2",X"00",X"C2",X"00",X"F2",X"00",X"32",X"00",X"F2",X"00",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"AA",X"AA",
		X"AA",X"AA",X"02",X"00",X"F2",X"3C",X"C2",X"0C",X"F2",X"0C",X"32",X"0C",X"F2",X"3F",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0F",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"03",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"0C",X"00",X"0F",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0C",X"C0",X"0C",X"C0",X"0F",X"F0",X"00",X"C0",X"00",X"C0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"0C",X"00",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"0C",X"00",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"00",X"30",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"00",X"30",X"00",X"30",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"30",X"C2",X"30",X"C2",X"30",X"C2",X"3F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"0F",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"00",X"C2",X"3F",X"C2",X"30",X"02",X"3F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"00",X"C2",X"3F",X"C2",X"00",X"C2",X"3F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"33",X"02",X"33",X"02",X"3F",X"C2",X"03",X"02",X"03",X"02",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"30",X"02",X"3F",X"C2",X"00",X"C2",X"3F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"30",X"02",X"3F",X"C2",X"30",X"C2",X"3F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"00",X"C2",X"03",X"C2",X"03",X"02",X"03",X"02",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"30",X"C2",X"3F",X"C2",X"30",X"C2",X"3F",X"C2",X"AA",X"AA",
		X"AA",X"AA",X"00",X"02",X"3F",X"C2",X"30",X"C2",X"3F",X"C2",X"00",X"C2",X"00",X"C2",X"AA",X"AA",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",
		X"57",X"F0",X"15",X"7F",X"01",X"57",X"00",X"15",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"7F",X"00",X"57",X"F0",X"15",X"7F",X"01",X"57",X"00",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"FD",X"FF",X"55",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"3F",X"D5",X"F5",X"55",X"55",X"40",X"50",X"00",
		X"00",X"3F",X"0F",X"F5",X"FD",X"55",X"55",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D5",X"57",X"55",X"07",X"40",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"03",X"F7",X"FF",X"57",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"03",X"C3",X"03",X"C4",X"03",X"C4",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",
		X"57",X"F0",X"15",X"7F",X"01",X"57",X"00",X"15",X"00",X"01",X"00",X"00",X"00",X"FC",X"00",X"7C",
		X"00",X"3F",X"0F",X"F5",X"FD",X"55",X"55",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D5",X"54",X"55",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"3C",X"00",
		X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",
		X"03",X"C3",X"03",X"FF",X"03",X"C3",X"03",X"C4",X"03",X"C4",X"03",X"C4",X"03",X"C0",X"03",X"C3",
		X"C0",X"00",X"00",X"00",X"CF",X"CF",X"F7",X"D3",X"F3",X"D3",X"F3",X"D3",X"F3",X"C3",X"C3",X"CF",
		X"00",X"3C",X"00",X"3C",X"0F",X"FF",X"3C",X"3C",X"3C",X"7C",X"3C",X"7C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"F3",X"F3",X"C4",X"C4",X"F3",X"F3",X"F3",X"33",X"3F",X"3F",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"F3",X"FC",X"CF",X"5F",X"CF",X"0F",X"0F",X"FF",X"0F",X"50",X"4F",X"0F",
		X"00",X"00",X"0C",X"00",X"FC",X"3F",X"7C",X"F5",X"3C",X"F0",X"3C",X"7F",X"3C",X"17",X"3C",X"C3",
		X"00",X"00",X"00",X"00",X"C3",X"FC",X"CF",X"5F",X"4F",X"0F",X"0F",X"FF",X"CF",X"57",X"CF",X"0F",
		X"00",X"07",X"0C",X"C7",X"FF",X"C7",X"3D",X"C7",X"3C",X"47",X"3C",X"07",X"3C",X"07",X"3C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"7F",X"00",
		X"0F",X"FF",X"00",X"00",X"15",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"F3",X"44",X"04",X"01",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"5F",
		X"CF",X"FF",X"10",X"00",X"55",X"55",X"00",X"5F",X"05",X"FD",X"5F",X"D5",X"FD",X"50",X"D5",X"00",
		X"3D",X"3C",X"41",X"41",X"55",X"15",X"F5",X"00",X"7F",X"54",X"17",X"FD",X"05",X"5F",X"00",X"15",
		X"43",X"FC",X"10",X"01",X"05",X"54",X"00",X"00",X"00",X"00",X"50",X"00",X"F5",X"40",X"7F",X"D5",
		X"FF",X"FF",X"00",X"40",X"55",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FC",X"10",X"01",X"45",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"00",X"47",X"55",X"17",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0D",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"5F",X"05",X"FD",X"1F",X"D5",X"FD",X"50",X"D5",X"00",
		X"05",X"FD",X"5F",X"D5",X"FD",X"50",X"D5",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"01",X"57",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"FD",X"50",X"5F",X"F5",X"15",X"7F",X"00",X"55",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"D5",X"00",X"FF",X"54",X"57",X"FD",X"05",X"5F",X"00",X"15",
		X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"50",X"07",X"F5",X"47",X"7F",X"D7",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"01",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FA",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"55",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"AA",X"AF",X"EA",X"AF",X"EA",X"BF",X"EA",X"BF",X"FA",X"BF",X"FA",X"FF",X"FA",X"EF",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"55",X"52",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",
		X"40",X"44",X"10",X"10",X"04",X"40",X"04",X"10",X"04",X"40",X"FF",X"FF",X"55",X"55",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"EB",X"AE",X"EA",X"AF",X"EB",X"AF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"15",X"55",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"52",X"AA",X"02",X"AA",X"02",X"AA",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"55",X"55",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"AA",X"AF",X"EA",X"AF",X"EA",X"BF",X"FA",X"BF",X"FA",X"BF",X"FA",X"FF",X"FE",X"EF",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"D5",X"03",X"FD",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"50",X"00",X"D5",X"00",X"FD",X"50",X"FF",X"D5",X"FF",X"FD",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"D5",X"00",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",
		X"6B",X"EA",X"6B",X"EA",X"5B",X"EA",X"DB",X"EA",X"DB",X"EA",X"D7",X"EA",X"F7",X"EA",X"F7",X"EA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"2A",X"00",X"28",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"EB",X"AE",X"EA",X"AF",X"EB",X"AF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"6B",X"EA",
		X"FD",X"50",X"FF",X"D5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"50",X"00",X"D5",X"00",X"FD",X"54",X"FF",X"FF",X"FF",X"F7",X"FF",X"F7",
		X"00",X"2A",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"55",X"52",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A9",X"AA",X"BC",
		X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"7F",X"F7",X"75",X"C1",X"55",X"73",X"3F",X"0F",
		X"55",X"5A",X"55",X"56",X"FF",X"D6",X"FF",X"D6",X"FF",X"D5",X"05",X"DD",X"4D",X"5D",X"CC",X"1D",
		X"55",X"5A",X"55",X"56",X"FF",X"D6",X"FF",X"D6",X"FF",X"D5",X"C3",X"DD",X"F3",X"DD",X"CC",X"CD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"55",
		X"FF",X"FF",X"7F",X"FF",X"57",X"FF",X"55",X"7F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"57",X"FF",X"55",X"7F",
		X"FF",X"F7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FD",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"2A",
		X"AA",X"FF",X"A8",X"0F",X"AE",X"8F",X"AE",X"83",X"BA",X"A3",X"BA",X"A3",X"BA",X"A3",X"BA",X"A3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"3F",X"D0",X"FF",X"F4",X"00",X"00",X"00",X"00",
		X"C3",X"1F",X"F0",X"FF",X"FC",X"3F",X"3F",X"3F",X"3B",X"3F",X"EB",X"0F",X"AB",X"CD",X"AB",X"CD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"7F",X"FF",X"57",X"FF",X"55",X"7F",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"FD",X"57",X"FD",X"57",X"F5",X"57",X"F5",X"57",X"F5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",
		X"BA",X"A3",X"BA",X"A3",X"BA",X"A3",X"BA",X"A3",X"AE",X"83",X"AE",X"8F",X"AB",X"0F",X"AA",X"FF",
		X"FA",X"AA",X"FA",X"AE",X"FA",X"BF",X"FD",X"57",X"C9",X"57",X"F9",X"57",X"FB",X"55",X"FB",X"55",
		X"AB",X"CD",X"AB",X"CD",X"AB",X"C0",X"EB",X"0C",X"00",X"FC",X"C0",X"3C",X"C3",X"0C",X"4D",X"40",
		X"F5",X"EA",X"7D",X"EA",X"7D",X"EA",X"3D",X"6A",X"CF",X"6A",X"FF",X"6A",X"0F",X"5A",X"C3",X"DA",
		X"00",X"15",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"51",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",
		X"D5",X"6A",X"D5",X"AF",X"D5",X"AA",X"D6",X"BF",X"D6",X"AA",X"DA",X"FF",X"DA",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"FE",X"AA",X"AA",X"AA",X"FF",X"AA",X"AA",X"AA",X"FF",X"EA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A7",X"AA",X"A7",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FB",X"55",X"FB",X"95",X"FB",X"95",X"FB",X"95",X"BB",X"9F",X"BB",X"9F",X"BB",X"9F",X"AB",X"9F",
		X"54",X"3C",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"53",X"DA",X"55",X"56",X"55",X"56",X"55",X"5E",X"7F",X"7E",X"7F",X"7E",X"7F",X"7E",X"7F",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"55",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"15",X"55",X"15",X"55",X"00",X"00",X"00",X"00",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"0F",X"FF",X"0F",X"FF",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"F5",X"5F",X"F5",X"5F",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"5A",X"5D",X"5A",X"DD",X"5A",X"F5",X"5A",
		X"0A",X"A0",X"3E",X"A0",X"FE",X"81",X"FA",X"0A",X"E8",X"16",X"A0",X"56",X"81",X"56",X"00",X"02",
		X"AB",X"9F",X"6B",X"9F",X"6B",X"9F",X"6B",X"9F",X"5B",X"9F",X"5B",X"9F",X"5B",X"9F",X"5A",X"9F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"75",X"7D",X"55",X"75",X"A9",X"5A",X"55",X"65",X"7F",
		X"7F",X"7E",X"7F",X"7E",X"7F",X"7E",X"57",X"7E",X"55",X"7E",X"55",X"5E",X"55",X"5E",X"F5",X"56",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"0D",X"55",X"05",X"55",X"07",X"55",X"05",X"55",X"2A",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"5A",X"AA",X"5A",X"57",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"AA",X"5A",X"AA",X"AA",
		X"0F",X"C3",X"CF",X"F0",X"CF",X"FC",X"C3",X"FC",X"FB",X"FF",X"FA",X"FF",X"FA",X"BF",X"FA",X"AE",
		X"5A",X"9F",X"5A",X"9F",X"5A",X"9F",X"9A",X"9F",X"9A",X"9F",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"67",X"FF",X"97",X"FF",X"9F",X"F5",X"9F",X"D7",X"9F",X"DF",X"9F",X"D7",X"9F",X"F5",X"97",X"FF",
		X"FF",X"5A",X"FF",X"6A",X"FF",X"AA",X"FE",X"AA",X"FF",X"EA",X"FF",X"DA",X"FF",X"DA",X"FF",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A7",X"95",X"A5",X"95",X"AA",X"95",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",
		X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"00",X"7F",X"33",X"C3",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"01",X"11",
		X"00",X"01",X"00",X"55",X"05",X"55",X"1F",X"55",X"7D",X"55",X"FD",X"55",X"D5",X"55",X"F5",X"55",
		X"D5",X"55",X"F1",X"55",X"3C",X"15",X"0F",X"C1",X"03",X"FF",X"00",X"3F",X"00",X"05",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"50",X"03",X"40",X"0F",X"00",X"3C",X"00",X"F0",X"FF",X"C0",X"FC",X"00",X"40",X"00",X"00",X"00",
		X"03",X"80",X"03",X"00",X"00",X"00",X"0F",X"00",X"3C",X"00",X"BC",X"00",X"80",X"00",X"A0",X"00",
		X"B0",X"00",X"AC",X"00",X"2B",X"C0",X"0A",X"BC",X"02",X"AA",X"03",X"AA",X"03",X"80",X"03",X"80",
		X"03",X"80",X"03",X"80",X"FF",X"80",X"FF",X"F0",X"3F",X"FC",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"0F",X"FE",X"3F",X"FA",X"FF",X"E8",X"FE",X"A0",X"AA",X"80",X"AB",X"80",X"03",X"80",X"03",X"80",
		X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"FF",X"AA",X"FF",
		X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FB",X"FA",X"FE",X"FA",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"6B",X"EA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"AA",X"02",X"AA",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"B5",X"AA",X"B5",X"AA",X"BD",X"AA",X"AD",X"AA",X"AD",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"A5",X"55",X"65",X"55",X"65",X"55",X"96",X"65",X"22",X"20",
		X"00",X"08",X"55",X"00",X"55",X"40",X"69",X"50",X"59",X"54",X"59",X"55",X"A9",X"55",X"88",X"00",
		X"88",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"80",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"2A",X"80",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"22",X"20",X"A2",X"A8",X"00",X"00",X"00",X"00",X"50",X"00",X"01",X"40",X"00",X"14",X"00",X"01",
		X"2A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"03",X"01",X"33",X"01",X"30",X"16",X"55",X"5A",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"40",X"00",X"90",X"30",X"90",X"33",X"A5",X"03",X"A9",X"55",X"AA",X"AA",X"AA",X"AA",
		X"00",X"02",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"2A",X"02",X"AA",
		X"BB",X"B8",X"BB",X"B8",X"FB",X"F8",X"0A",X"A8",X"00",X"A8",X"00",X"28",X"00",X"08",X"00",X"00",
		X"0B",X"BB",X"0B",X"BB",X"0B",X"EB",X"0A",X"A8",X"0A",X"80",X"0A",X"00",X"08",X"00",X"00",X"00",
		X"54",X"00",X"84",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"84",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"0A",X"00",X"0B",X"C0",X"0B",X"B8",X"0B",X"BA",X"0B",X"EB",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"28",X"02",X"B8",X"0A",X"B8",X"2A",X"B8",X"BB",X"F8",
		X"02",X"A0",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"40",X"55",X"10",X"00",X"04",X"00",X"01",X"00",X"00",X"40",X"00",X"10",X"00",X"05",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"6A",X"80",X"0A",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"00",X"08",X"00",X"28",X"00",X"A8",X"00",X"28",X"00",
		X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F5",X"2A",X"D1",X"2A",X"85",X"00",X"D5",X"0A",X"F4",X"2A",X"80",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"04",X"00",
		X"50",X"00",X"54",X"50",X"55",X"05",X"50",X"50",X"14",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
