module gun(
input	clk,
input gun1up,
input gun1dw,
input gun2up,
input gun2dw,
output [2:0] gun1out,
output [2:0] gun2out
);

//0x06, 0x02, 0x00, 0x04, 0x05, 0x01, 0x03
wire [6:0]gun[6:0]gun = ()
endmodule 