library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_tile_bit0 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"27",X"77",X"77",X"77",X"77",X"27",X"0E",X"08",X"22",X"77",X"77",X"77",X"77",X"22",X"08",
		X"88",X"22",X"77",X"77",X"77",X"77",X"22",X"88",X"8E",X"27",X"77",X"77",X"77",X"77",X"27",X"8E",
		X"00",X"02",X"03",X"03",X"03",X"03",X"FF",X"7F",X"00",X"02",X"03",X"03",X"03",X"03",X"FF",X"7F",
		X"00",X"02",X"03",X"03",X"03",X"03",X"FF",X"7F",X"00",X"02",X"03",X"03",X"03",X"03",X"FF",X"7F",
		X"70",X"D8",X"88",X"48",X"90",X"88",X"D8",X"70",X"77",X"DD",X"88",X"4C",X"99",X"88",X"DD",X"77",
		X"77",X"DD",X"88",X"CC",X"99",X"88",X"DD",X"77",X"70",X"D8",X"88",X"C8",X"90",X"88",X"D8",X"70",
		X"00",X"01",X"1F",X"0F",X"FF",X"1F",X"E3",X"07",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"FC",X"F6",
		X"0F",X"CF",X"87",X"FF",X"E3",X"0F",X"1F",X"00",X"F6",X"FE",X"FC",X"FC",X"F0",X"E0",X"C0",X"00",
		X"00",X"01",X"1F",X"0F",X"FF",X"17",X"EF",X"0F",X"00",X"C0",X"F0",X"F0",X"F8",X"F8",X"FC",X"F6",
		X"07",X"C3",X"8F",X"FF",X"EF",X"0F",X"1F",X"00",X"F6",X"FE",X"FC",X"FC",X"F8",X"E0",X"80",X"00",
		X"00",X"0C",X"27",X"79",X"FC",X"00",X"C0",X"00",X"00",X"00",X"C0",X"E0",X"38",X"0C",X"04",X"04",
		X"00",X"9C",X"F8",X"E7",X"03",X"07",X"00",X"00",X"0C",X"1C",X"18",X"38",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"00",X"03",X"06",X"01",X"00",X"00",X"00",X"00",X"C0",X"E3",X"F9",X"E7",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"03",X"0F",X"01",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"30",X"08",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"0F",X"07",X"00",X"00",X"01",X"0F",X"06",X"18",X"FC",X"E4",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"7E",X"04",X"1E",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"06",X"07",X"2F",X"3F",X"7F",X"7F",X"00",X"00",X"08",X"8C",X"8E",X"DE",X"FE",X"FE",
		X"7F",X"FF",X"FF",X"F9",X"F0",X"70",X"20",X"00",X"FE",X"FE",X"FC",X"FE",X"7C",X"38",X"18",X"00",
		X"30",X"78",X"48",X"4D",X"40",X"60",X"20",X"00",X"00",X"08",X"04",X"04",X"08",X"10",X"10",X"08",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",X"00",X"01",X"01",X"7F",X"7F",X"21",X"01",X"00",X"00",
		X"31",X"79",X"59",X"4D",X"4F",X"67",X"23",X"00",X"46",X"6F",X"79",X"59",X"49",X"43",X"02",X"00",
		X"04",X"7F",X"7F",X"64",X"34",X"1C",X"0C",X"00",X"0E",X"5F",X"51",X"51",X"51",X"77",X"76",X"00",
		X"06",X"0F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"60",X"70",X"58",X"4F",X"47",X"40",X"40",X"00",
		X"36",X"4F",X"4D",X"5D",X"59",X"79",X"36",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"78",X"30",X"00",
		X"38",X"44",X"42",X"21",X"42",X"44",X"38",X"00",X"0D",X"26",X"77",X"59",X"4D",X"57",X"22",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"5A",X"99",X"BD",X"BD",X"99",X"42",X"3C",X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",X"00",
		X"36",X"7F",X"49",X"49",X"49",X"7F",X"7F",X"00",X"22",X"63",X"41",X"41",X"63",X"3E",X"1C",X"00",
		X"1C",X"3E",X"63",X"41",X"41",X"7F",X"7F",X"00",X"41",X"49",X"49",X"49",X"49",X"7F",X"7F",X"00",
		X"40",X"48",X"48",X"48",X"48",X"7F",X"7F",X"00",X"4F",X"4F",X"49",X"49",X"63",X"3E",X"1C",X"00",
		X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"7F",X"7F",X"41",X"00",X"00",X"00",
		X"7E",X"7F",X"01",X"01",X"01",X"03",X"02",X"00",X"41",X"63",X"37",X"1E",X"0C",X"7F",X"7F",X"00",
		X"01",X"01",X"01",X"01",X"01",X"7F",X"7F",X"00",X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",X"00",
		X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",X"00",
		X"30",X"78",X"48",X"48",X"48",X"7F",X"7F",X"00",X"3D",X"7F",X"46",X"45",X"41",X"7F",X"3E",X"00",
		X"39",X"7B",X"4E",X"44",X"44",X"7F",X"7F",X"00",X"26",X"6F",X"4D",X"59",X"59",X"7B",X"32",X"00",
		X"40",X"40",X"7F",X"7F",X"40",X"40",X"00",X"00",X"7E",X"7F",X"03",X"03",X"03",X"7F",X"7E",X"00",
		X"78",X"7C",X"06",X"03",X"06",X"7C",X"78",X"00",X"7C",X"7F",X"06",X"1C",X"06",X"7F",X"7C",X"00",
		X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"60",X"78",X"0F",X"0F",X"78",X"60",X"00",X"00",
		X"61",X"71",X"79",X"5D",X"4F",X"47",X"43",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"0F",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"E0",
		X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"0F",X"1F",X"1F",X"00",X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"1F",X"1F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"07",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"E0",X"10",X"E0",X"00",X"E0",X"10",
		X"03",X"00",X"00",X"04",X"04",X"07",X"00",X"00",X"E0",X"00",X"60",X"90",X"90",X"A0",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",
		X"03",X"00",X"02",X"05",X"05",X"02",X"00",X"00",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"07",X"02",X"00",X"C0",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"04",X"02",X"C0",X"20",X"C0",X"00",X"20",X"A0",X"A0",X"60",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"06",X"05",X"05",X"04",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"40",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"07",X"04",X"03",X"C0",X"20",X"C0",X"00",X"40",X"E0",X"40",X"C0",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"05",X"05",X"07",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"F0",X"E0",X"C1",X"83",X"83",X"80",X"80",X"00",X"00",X"00",X"08",X"1C",X"1F",X"1F",X"1F",
		X"80",X"CE",X"90",X"90",X"C0",X"F0",X"FF",X"DF",X"0F",X"0F",X"0E",X"06",X"06",X"04",X"00",X"00",
		X"00",X"00",X"06",X"06",X"07",X"0F",X"1F",X"1F",X"00",X"00",X"20",X"30",X"70",X"FC",X"FD",X"FF",
		X"0F",X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"FF",X"BF",X"3F",X"3E",X"3C",X"1C",X"18",X"00",
		X"0F",X"0E",X"0C",X"08",X"08",X"01",X"01",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"80",X"00",X"18",X"7E",X"C3",X"99",X"3C",X"66",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"7E",X"50",X"50",X"10",X"14",X"14",X"34",X"34",X"7E",X"02",X"02",X"00",X"78",X"78",X"7C",X"7C",
		X"34",X"3C",X"3C",X"18",X"00",X"42",X"42",X"7E",X"7C",X"7C",X"78",X"78",X"00",X"02",X"02",X"7E",
		X"7E",X"3C",X"3C",X"1C",X"1C",X"0C",X"0C",X"24",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"24",X"30",X"30",X"38",X"38",X"3C",X"3C",X"7E",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"7E",
		X"7E",X"3C",X"3C",X"3C",X"3C",X"2C",X"2C",X"2C",X"7E",X"4C",X"4C",X"04",X"04",X"30",X"30",X"30",
		X"2C",X"2C",X"2C",X"2C",X"00",X"00",X"00",X"7E",X"36",X"36",X"36",X"36",X"00",X"00",X"00",X"7E",
		X"AF",X"2E",X"2C",X"08",X"08",X"81",X"81",X"C3",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",
		X"A0",X"20",X"20",X"00",X"00",X"80",X"80",X"C0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"0F",X"00",X"38",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"00",X"00",X"00",X"81",X"83",X"83",X"A7",X"AF",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"00",X"00",X"00",X"80",X"80",X"80",X"A0",X"A0",X"AF",X"FF",X"00",X"00",X"00",X"00",X"00",X"AF",
		X"FA",X"FF",X"00",X"00",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FA",X"FA",X"FA",X"FB",X"FA",X"FA",X"FC",X"F8",X"E0",X"F0",X"F8",X"FC",X"FC",
		X"F8",X"FC",X"F8",X"90",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"C0",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",X"18",X"24",
		X"1E",X"21",X"1E",X"00",X"06",X"29",X"29",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"21",X"01",X"C1",X"83",X"03",X"07",X"07",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"C3",X"C0",X"C0",X"C0",X"C8",X"DE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AC",X"AC",X"AC",X"AE",X"AE",X"AE",X"AF",X"AE",X"AE",X"AC",X"B8",X"A0",X"B0",X"B8",X"AC",X"AC",
		X"A8",X"EC",X"E8",X"90",X"C0",X"E0",X"B0",X"B0",X"A0",X"C0",X"C0",X"A0",X"A0",X"C0",X"C0",X"C0",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",
		X"1E",X"00",X"19",X"25",X"25",X"13",X"00",X"00",X"18",X"24",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",
		X"1E",X"00",X"06",X"29",X"29",X"3A",X"00",X"00",X"18",X"24",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",
		X"1E",X"00",X"16",X"29",X"29",X"16",X"00",X"00",X"18",X"24",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",X"18",X"24",
		X"1E",X"21",X"1E",X"00",X"01",X"3F",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",X"18",X"24",
		X"1E",X"21",X"1E",X"00",X"19",X"25",X"25",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",X"18",X"24",
		X"1E",X"21",X"1E",X"00",X"36",X"29",X"29",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"74",X"54",X"5C",X"00",X"24",X"18",X"18",X"24",
		X"1E",X"21",X"1E",X"00",X"02",X"3F",X"22",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"00",X"00",X"0E",X"3F",X"1C",X"FF",X"0C",
		X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"3F",X"7F",X"07",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"04",X"02",X"02",X"02",X"01",X"FA",X"FA",X"FC",X"38",X"20",X"30",X"18",X"0C",X"FC",
		X"F8",X"FC",X"C8",X"90",X"C0",X"60",X"20",X"F0",X"E0",X"C0",X"40",X"20",X"20",X"40",X"40",X"C0",
		X"AC",X"FC",X"04",X"02",X"02",X"02",X"01",X"AE",X"AE",X"FC",X"38",X"20",X"30",X"18",X"0C",X"AC",
		X"A8",X"FC",X"C8",X"90",X"C0",X"60",X"30",X"B0",X"A0",X"C0",X"40",X"20",X"20",X"40",X"40",X"C0",
		X"00",X"F0",X"B8",X"8C",X"86",X"82",X"83",X"81",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"FF",
		X"83",X"82",X"86",X"8C",X"B8",X"E0",X"00",X"00",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"7F",X"3F",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"7F",X"76",X"37",X"03",X"00",X"FF",X"FF",X"FF",X"FE",X"18",X"F0",X"E0",X"00",
		X"00",X"03",X"03",X"13",X"30",X"23",X"13",X"30",X"00",X"00",X"20",X"30",X"10",X"20",X"30",X"10",
		X"23",X"13",X"33",X"30",X"07",X"0F",X"07",X"00",X"20",X"30",X"30",X"00",X"E0",X"B0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C7",X"00",X"00",X"00",X"00",X"70",X"0C",X"63",X"39",
		X"FF",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"BF",X"BF",X"7F",X"FC",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"01",X"07",X"03",X"00",X"03",X"07",X"7F",X"F0",X"C0",X"E0",X"00",
		X"0F",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"66",X"FC",X"05",X"1F",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",
		X"03",X"00",X"03",X"04",X"04",X"02",X"00",X"00",X"C0",X"00",X"20",X"A0",X"A0",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"4C",X"50",X"21",X"43",X"43",X"40",X"40",X"00",X"20",X"10",X"C8",X"80",X"00",X"08",X"10",
		X"43",X"24",X"44",X"43",X"34",X"4F",X"40",X"80",X"D0",X"20",X"20",X"C0",X"20",X"C0",X"00",X"00",
		X"20",X"4F",X"90",X"A1",X"43",X"43",X"40",X"40",X"00",X"C0",X"80",X"80",X"90",X"08",X"00",X"00",
		X"43",X"27",X"47",X"43",X"37",X"4F",X"40",X"20",X"C8",X"30",X"30",X"D0",X"20",X"E0",X"00",X"00",
		X"20",X"4F",X"90",X"A1",X"43",X"43",X"40",X"40",X"00",X"E0",X"10",X"C0",X"E0",X"60",X"10",X"10",
		X"43",X"24",X"44",X"43",X"34",X"4F",X"20",X"18",X"88",X"20",X"20",X"C8",X"30",X"E0",X"00",X"00",
		X"41",X"87",X"9B",X"A0",X"A7",X"48",X"48",X"27",X"C0",X"C0",X"10",X"00",X"80",X"40",X"40",X"90",
		X"27",X"48",X"48",X"A6",X"A0",X"9B",X"87",X"41",X"90",X"48",X"00",X"00",X"C8",X"D0",X"E0",X"80",
		X"11",X"27",X"5B",X"A0",X"A6",X"4E",X"4E",X"27",X"80",X"E0",X"D0",X"C8",X"00",X"00",X"48",X"90",
		X"27",X"4E",X"4E",X"A7",X"A0",X"5B",X"27",X"11",X"90",X"40",X"40",X"80",X"00",X"10",X"C0",X"C0",
		X"00",X"4C",X"50",X"21",X"43",X"43",X"40",X"40",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",
		X"43",X"24",X"44",X"43",X"34",X"4F",X"40",X"00",X"C0",X"20",X"20",X"C0",X"20",X"C0",X"00",X"00",
		X"00",X"4F",X"90",X"A1",X"43",X"43",X"40",X"40",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"43",X"27",X"47",X"43",X"37",X"4F",X"40",X"00",X"C0",X"20",X"20",X"C0",X"20",X"C0",X"00",X"00",
		X"00",X"4F",X"90",X"A1",X"43",X"43",X"40",X"40",X"00",X"00",X"00",X"C0",X"E0",X"60",X"00",X"00",
		X"43",X"24",X"44",X"43",X"34",X"4F",X"20",X"10",X"80",X"20",X"20",X"C0",X"20",X"C0",X"00",X"00",
		X"00",X"4C",X"90",X"A3",X"43",X"43",X"40",X"40",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"43",X"24",X"44",X"43",X"74",X"7F",X"77",X"77",X"C0",X"20",X"20",X"C0",X"20",X"D8",X"B8",X"B8",
		X"01",X"87",X"9B",X"A0",X"A7",X"48",X"48",X"27",X"C0",X"C0",X"80",X"00",X"80",X"40",X"40",X"80",
		X"27",X"48",X"48",X"A6",X"A0",X"9B",X"87",X"01",X"80",X"40",X"00",X"00",X"C0",X"C0",X"C0",X"80",
		X"01",X"47",X"9B",X"A0",X"A7",X"48",X"C8",X"E7",X"C0",X"C0",X"80",X"00",X"80",X"40",X"40",X"80",
		X"E7",X"C8",X"48",X"A7",X"A0",X"9B",X"47",X"01",X"80",X"40",X"40",X"80",X"00",X"00",X"C0",X"C0",
		X"01",X"27",X"5B",X"A0",X"A6",X"4E",X"4E",X"27",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"40",X"80",
		X"27",X"4E",X"4E",X"A7",X"A0",X"5B",X"27",X"01",X"80",X"40",X"40",X"80",X"00",X"00",X"C0",X"C0",
		X"01",X"27",X"5B",X"A0",X"A7",X"48",X"48",X"27",X"C0",X"C0",X"81",X"01",X"81",X"40",X"41",X"8F",
		X"27",X"48",X"48",X"A7",X"A0",X"5B",X"27",X"01",X"8F",X"41",X"40",X"81",X"01",X"01",X"C0",X"C0",
		X"00",X"48",X"50",X"21",X"43",X"43",X"40",X"40",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",
		X"40",X"2E",X"50",X"50",X"2E",X"50",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"48",X"90",X"A1",X"43",X"43",X"40",X"40",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"40",X"2E",X"58",X"58",X"2E",X"58",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"48",X"90",X"A1",X"43",X"43",X"40",X"40",X"00",X"00",X"00",X"C0",X"E0",X"60",X"00",X"00",
		X"40",X"2E",X"50",X"50",X"2E",X"50",X"2E",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"48",X"90",X"A3",X"47",X"46",X"40",X"40",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"40",X"2E",X"50",X"50",X"6E",X"70",X"7F",X"77",X"80",X"80",X"80",X"80",X"80",X"B8",X"B8",X"B8",
		X"01",X"83",X"9B",X"A0",X"A6",X"48",X"48",X"26",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"48",X"48",X"A6",X"A0",X"98",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",
		X"01",X"83",X"9B",X"A0",X"AE",X"50",X"D0",X"EE",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"D0",X"50",X"AE",X"A0",X"9B",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"01",X"23",X"58",X"A0",X"AE",X"50",X"50",X"2E",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"50",X"50",X"AE",X"A0",X"5B",X"23",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"01",X"23",X"5B",X"A0",X"AE",X"50",X"50",X"2E",X"C0",X"C0",X"01",X"01",X"01",X"00",X"01",X"07",
		X"2E",X"50",X"50",X"AE",X"A0",X"5B",X"23",X"01",X"07",X"01",X"00",X"01",X"01",X"01",X"C0",X"C0",
		X"00",X"40",X"40",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"0E",X"10",X"10",X"0E",X"50",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"81",X"03",X"03",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"0E",X"18",X"18",X"0E",X"58",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"81",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"60",X"00",X"00",
		X"00",X"0E",X"10",X"10",X"0E",X"50",X"2E",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"83",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"10",X"10",X"4E",X"70",X"7F",X"77",X"80",X"80",X"80",X"80",X"80",X"98",X"B8",X"B8",
		X"01",X"83",X"83",X"80",X"86",X"08",X"08",X"06",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"08",X"08",X"86",X"80",X"80",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",
		X"01",X"C3",X"83",X"80",X"8E",X"10",X"90",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"90",X"10",X"8E",X"80",X"83",X"C3",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"01",X"23",X"40",X"80",X"8E",X"10",X"10",X"0E",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"10",X"10",X"8E",X"80",X"43",X"23",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"01",X"23",X"43",X"80",X"8E",X"10",X"10",X"00",X"C0",X"C0",X"01",X"01",X"01",X"00",X"01",X"07",
		X"00",X"10",X"10",X"8E",X"80",X"43",X"23",X"01",X"07",X"01",X"00",X"01",X"01",X"01",X"C0",X"C0",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"77",X"77",X"F7",X"A3",X"88",X"DC",X"F7",X"63",X"B8",X"B8",X"BC",X"14",X"44",X"EC",X"BC",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"54",X"F7",X"A3",X"88",X"DC",X"F7",X"63",X"00",X"A8",X"BC",X"14",X"44",X"EC",X"BC",X"18",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"B8",X"B8",X"B8",X"B8",
		X"77",X"77",X"F7",X"A3",X"88",X"DC",X"F7",X"63",X"B8",X"B8",X"BC",X"14",X"44",X"EC",X"BC",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"F7",X"A3",X"88",X"DC",X"F7",X"63",X"B8",X"B8",X"BC",X"14",X"44",X"EC",X"BC",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"54",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"A8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"7C",X"E7",X"CF",X"67",X"30",X"67",X"CF",X"CF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"67",X"30",X"67",X"CF",X"E7",X"7C",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"7C",X"E6",X"CC",X"66",X"30",X"66",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"30",X"66",X"CC",X"E6",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"7C",X"E7",X"CF",X"67",X"30",X"67",X"CF",X"CF",X"00",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",
		X"67",X"30",X"67",X"CF",X"E7",X"7C",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"7C",X"E7",X"CF",X"67",X"30",X"67",X"CF",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"67",X"30",X"67",X"CF",X"E7",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"FC",X"FE",X"00",X"FE",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"00",X"FE",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"30",X"60",X"00",X"00",X"70",X"98",X"88",X"48",X"90",X"88",X"D8",X"70",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"FF",X"00",X"00",X"00",X"00",X"FF",X"C1",X"FD",X"C3",
		X"FF",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"D3",X"CB",X"C3",X"DF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"CD",
		X"1F",X"1F",X"1F",X"07",X"03",X"03",X"01",X"00",X"AD",X"9D",X"AD",X"CD",X"AD",X"9D",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"7C",X"78",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"01",X"01",X"00",X"00",X"01",X"03",X"07",X"C0",X"E0",X"E0",X"C0",X"00",X"C0",X"C0",X"00",
		X"00",X"06",X"03",X"03",X"03",X"07",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"06",X"06",X"06",X"07",X"03",X"00",X"00",X"00",X"20",X"30",X"30",X"20",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"01",X"01",X"01",X"03",X"0E",X"00",X"00",X"00",X"90",X"98",X"98",X"18",X"30",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E4",X"76",X"36",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"36",X"76",X"E4",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"20",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"20",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"01",X"00",X"07",X"03",X"03",X"06",X"1C",X"01",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"03",X"03",X"07",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"E0",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"07",X"0E",X"08",X"01",X"00",X"00",X"60",X"60",X"60",X"60",X"E0",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"18",X"38",X"70",X"60",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"30",X"30",X"70",X"00",
		X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"70",X"30",X"30",X"80",X"C0",X"C0",X"C0",
		X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"60",X"70",X"38",X"18",
		X"60",X"80",X"80",X"43",X"47",X"2F",X"17",X"13",X"00",X"00",X"00",X"C0",X"20",X"20",X"20",X"C0",
		X"13",X"17",X"2F",X"47",X"43",X"80",X"80",X"60",X"C0",X"20",X"20",X"20",X"C0",X"00",X"00",X"00",
		X"00",X"01",X"02",X"02",X"02",X"01",X"00",X"00",X"80",X"00",X"00",X"78",X"F4",X"F4",X"F4",X"78",
		X"00",X"00",X"01",X"02",X"02",X"02",X"01",X"00",X"78",X"F4",X"F4",X"F4",X"78",X"00",X"00",X"80",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"70",X"F8",X"FC",X"FC",X"FC",X"F8",X"70",X"F8",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"F8",X"70",X"00",X"00",X"00",
		X"0F",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"F8",X"FC",X"F8",
		X"01",X"01",X"03",X"07",X"0F",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"33",X"00",X"00",X"00",X"F8",X"FC",X"FE",X"FF",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3F",X"7F",X"7B",X"75",X"3F",X"1F",X"00",X"38",X"FC",X"FE",X"DE",X"EE",X"FC",X"F8",
		X"1F",X"3F",X"75",X"7B",X"7F",X"3F",X"1C",X"00",X"D8",X"FC",X"EE",X"DE",X"FE",X"FC",X"38",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"80",X"C0",X"71",X"10",
		X"10",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
