library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_samples is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_samples is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"76",X"78",X"77",X"78",X"88",X"76",X"68",X"9A",X"68",X"77",X"9A",X"65",X"85",X"67",X"97",X"89",
		X"76",X"69",X"58",X"88",X"57",X"67",X"8A",X"AB",X"CB",X"A8",X"54",X"52",X"48",X"A7",X"67",X"87",
		X"BA",X"8C",X"96",X"33",X"15",X"8C",X"AA",X"74",X"45",X"88",X"ED",X"B9",X"A0",X"01",X"68",X"EF",
		X"95",X"74",X"37",X"E9",X"8C",X"81",X"04",X"55",X"DF",X"A6",X"31",X"19",X"EF",X"CA",X"73",X"00",
		X"2A",X"EF",X"FA",X"00",X"58",X"FF",X"F8",X"32",X"00",X"39",X"FF",X"C4",X"00",X"8E",X"FF",X"D5",
		X"00",X"02",X"8F",X"FD",X"20",X"18",X"EF",X"FE",X"60",X"00",X"5D",X"FD",X"D3",X"00",X"6C",X"FF",
		X"E4",X"00",X"06",X"FF",X"DB",X"60",X"06",X"EF",X"DE",X"50",X"00",X"9F",X"FC",X"A4",X"00",X"7F",
		X"FB",X"A4",X"00",X"2C",X"FF",X"96",X"30",X"2C",X"FF",X"84",X"20",X"05",X"EF",X"B6",X"62",X"15",
		X"FF",X"D4",X"01",X"03",X"CF",X"F6",X"02",X"45",X"DF",X"F6",X"00",X"14",X"CF",X"F9",X"10",X"28",
		X"FF",X"D7",X"00",X"06",X"FF",X"B9",X"31",X"2A",X"FF",X"B5",X"10",X"05",X"FF",X"C7",X"57",X"9A",
		X"FF",X"D6",X"01",X"46",X"7B",X"B8",X"B7",X"AB",X"AA",X"63",X"42",X"55",X"43",X"4F",X"DD",X"F9",
		X"91",X"24",X"68",X"85",X"00",X"5B",X"FF",X"A8",X"00",X"07",X"DB",X"61",X"46",X"5C",X"FF",X"A0",
		X"02",X"7C",X"B8",X"43",X"66",X"9D",X"ED",X"40",X"28",X"B9",X"73",X"48",X"68",X"FF",X"B1",X"16",
		X"8A",X"B7",X"11",X"9F",X"A9",X"CD",X"50",X"39",X"DA",X"53",X"66",X"DA",X"96",X"88",X"25",X"7B",
		X"B3",X"06",X"DF",X"96",X"73",X"43",X"69",X"B9",X"51",X"7B",X"FF",X"84",X"00",X"37",X"EF",X"71",
		X"18",X"FF",X"CC",X"A2",X"00",X"6F",X"E7",X"15",X"7C",X"FD",X"B9",X"60",X"05",X"CD",X"72",X"69",
		X"ED",X"BA",X"66",X"01",X"8A",X"B6",X"18",X"9F",X"FA",X"72",X"23",X"37",X"88",X"82",X"8E",X"FF",
		X"73",X"41",X"22",X"9C",X"76",X"47",X"FF",X"F9",X"00",X"27",X"75",X"BD",X"51",X"5C",X"FB",X"61",
		X"34",X"54",X"6D",X"D5",X"39",X"CF",X"97",X"33",X"51",X"3A",X"FD",X"63",X"9D",X"F9",X"64",X"33",
		X"05",X"BF",X"B4",X"39",X"CE",X"B8",X"43",X"30",X"49",X"DC",X"74",X"69",X"EF",X"B6",X"23",X"31",
		X"8B",X"BA",X"76",X"5A",X"FE",X"A5",X"34",X"35",X"99",X"99",X"77",X"7A",X"BC",X"B6",X"64",X"46",
		X"57",X"78",X"BA",X"97",X"7A",X"A9",X"97",X"64",X"56",X"68",X"B9",X"85",X"59",X"9A",X"A7",X"73",
		X"57",X"7A",X"A7",X"66",X"88",X"6A",X"99",X"53",X"77",X"89",X"77",X"67",X"75",X"8B",X"B8",X"36",
		X"98",X"54",X"7A",X"98",X"55",X"7A",X"AA",X"89",X"74",X"35",X"BA",X"88",X"55",X"58",X"DD",X"B7",
		X"43",X"48",X"BA",X"96",X"53",X"4A",X"CC",X"95",X"43",X"4A",X"BB",X"64",X"56",X"8A",X"AA",X"56",
		X"55",X"78",X"85",X"67",X"98",X"99",X"85",X"47",X"AA",X"84",X"34",X"6A",X"AB",X"A6",X"34",X"8C",
		X"D8",X"31",X"35",X"AB",X"CB",X"63",X"47",X"BC",X"96",X"34",X"58",X"AA",X"A7",X"66",X"79",X"98",
		X"76",X"66",X"78",X"98",X"76",X"68",X"99",X"87",X"65",X"68",X"99",X"86",X"67",X"89",X"97",X"77",
		X"77",X"88",X"87",X"77",X"78",X"88",X"76",X"67",X"89",X"87",X"76",X"67",X"9A",X"96",X"45",X"7A",
		X"A8",X"86",X"56",X"8B",X"B8",X"55",X"57",X"9A",X"A7",X"44",X"69",X"BB",X"85",X"55",X"89",X"9A",
		X"86",X"45",X"8B",X"A7",X"55",X"77",X"99",X"A8",X"65",X"68",X"99",X"86",X"66",X"78",X"88",X"77",
		X"77",X"78",X"77",X"77",X"77",X"78",X"88",X"77",X"77",X"89",X"87",X"67",X"78",X"88",X"87",X"77",
		X"77",X"77",X"77",X"77",X"77",X"87",X"77",X"78",X"87",X"77",X"77",X"88",X"78",X"87",X"77",X"88",
		X"77",X"67",X"77",X"88",X"88",X"77",X"78",X"87",X"77",X"77",X"87",X"67",X"78",X"87",X"78",X"77",
		X"67",X"88",X"76",X"77",X"88",X"88",X"77",X"87",X"78",X"97",X"67",X"88",X"86",X"88",X"87",X"77",
		X"87",X"77",X"78",X"88",X"77",X"76",X"67",X"88",X"87",X"67",X"78",X"87",X"78",X"76",X"68",X"98",
		X"77",X"77",X"78",X"78",X"97",X"67",X"78",X"88",X"87",X"77",X"77",X"79",X"97",X"66",X"78",X"77",
		X"88",X"99",X"97",X"77",X"66",X"55",X"67",X"9C",X"CB",X"75",X"68",X"84",X"36",X"9B",X"74",X"5A",
		X"EE",X"83",X"37",X"95",X"25",X"9D",X"A4",X"37",X"DF",X"C6",X"13",X"69",X"62",X"6B",X"EB",X"31",
		X"5D",X"FD",X"50",X"37",X"95",X"29",X"EF",X"A0",X"02",X"9F",X"FD",X"72",X"21",X"33",X"7D",X"FF",
		X"A2",X"00",X"48",X"FF",X"FB",X"30",X"02",X"69",X"EF",X"FB",X"20",X"02",X"7D",X"FF",X"C5",X"00",
		X"03",X"9F",X"FF",X"B2",X"00",X"15",X"9F",X"FF",X"B2",X"00",X"38",X"CF",X"FF",X"90",X"00",X"16",
		X"CF",X"FE",X"60",X"00",X"38",X"BF",X"FF",X"90",X"00",X"26",X"CF",X"FF",X"71",X"00",X"4A",X"FF",
		X"FF",X"71",X"00",X"4B",X"FF",X"ED",X"50",X"00",X"5A",X"FF",X"FF",X"81",X"00",X"3A",X"FF",X"FF",
		X"90",X"00",X"5C",X"FD",X"CE",X"C3",X"00",X"28",X"EE",X"ED",X"D5",X"00",X"28",X"FF",X"DC",X"C5",
		X"00",X"05",X"EF",X"CC",X"E8",X"00",X"05",X"CF",X"DC",X"EA",X"20",X"04",X"BF",X"DB",X"CB",X"50",
		X"05",X"9D",X"DC",X"DD",X"60",X"01",X"8E",X"DA",X"AD",X"82",X"02",X"7E",X"EB",X"8B",X"92",X"00",
		X"6D",X"EC",X"9A",X"B5",X"00",X"7A",X"DB",X"9A",X"D6",X"00",X"5B",X"DA",X"89",X"C8",X"20",X"6A",
		X"DA",X"69",X"DB",X"40",X"18",X"EA",X"57",X"9C",X"61",X"38",X"C9",X"57",X"AE",X"82",X"05",X"AA",
		X"66",X"AC",X"B6",X"25",X"89",X"55",X"AE",X"C6",X"13",X"58",X"86",X"8B",X"DC",X"73",X"45",X"54",
		X"8B",X"FE",X"A3",X"10",X"38",X"B9",X"67",X"EF",X"A1",X"14",X"87",X"7A",X"FD",X"71",X"03",X"9A",
		X"74",X"7C",X"FB",X"40",X"56",X"54",X"AE",X"FB",X"50",X"26",X"A8",X"54",X"8D",X"FC",X"52",X"55",
		X"34",X"BF",X"E9",X"43",X"36",X"66",X"67",X"7A",X"DE",X"75",X"46",X"33",X"9C",X"DA",X"75",X"54",
		X"66",X"64",X"48",X"DF",X"C8",X"62",X"32",X"5A",X"CF",X"FA",X"20",X"15",X"34",X"6B",X"CD",X"DD",
		X"73",X"12",X"36",X"CF",X"FC",X"60",X"13",X"45",X"8C",X"B7",X"7C",X"F9",X"02",X"47",X"3A",X"DF",
		X"B8",X"40",X"35",X"85",X"9B",X"94",X"8A",X"C5",X"48",X"75",X"5A",X"8A",X"CC",X"61",X"55",X"65",
		X"CC",X"51",X"8C",X"CB",X"88",X"02",X"49",X"9C",X"FB",X"30",X"44",X"78",X"CB",X"54",X"3A",X"BC",
		X"89",X"75",X"34",X"A8",X"FA",X"73",X"36",X"37",X"7E",X"84",X"13",X"BD",X"FB",X"C3",X"23",X"1A",
		X"AF",X"C7",X"21",X"44",X"89",X"F9",X"81",X"2A",X"CE",X"B9",X"31",X"51",X"7C",X"FB",X"81",X"05",
		X"7B",X"BC",X"A5",X"00",X"4C",X"FF",X"D4",X"00",X"36",X"FF",X"FA",X"30",X"17",X"CC",X"EA",X"41",
		X"00",X"7F",X"FE",X"66",X"03",X"5F",X"FF",X"A4",X"10",X"6A",X"FC",X"D4",X"10",X"01",X"AF",X"FF",
		X"64",X"01",X"6E",X"FC",X"A3",X"10",X"88",X"EC",X"A1",X"32",X"14",X"AD",X"FE",X"81",X"51",X"8A",
		X"F9",X"78",X"52",X"59",X"6F",X"B8",X"35",X"03",X"67",X"EF",X"BC",X"34",X"2B",X"5C",X"8B",X"C8",
		X"11",X"56",X"FC",X"64",X"00",X"34",X"6D",X"FA",X"C3",X"34",X"64",X"CB",X"DD",X"71",X"04",X"BF",
		X"F6",X"82",X"02",X"27",X"EA",X"B7",X"A5",X"86",X"67",X"AB",X"DB",X"22",X"06",X"9F",X"FB",X"20",
		X"03",X"9C",X"C6",X"49",X"5F",X"7D",X"57",X"07",X"8D",X"B9",X"53",X"6C",X"CA",X"50",X"24",X"57",
		X"E9",X"37",X"99",X"F8",X"81",X"22",X"9F",X"FD",X"90",X"02",X"8F",X"E7",X"30",X"09",X"7C",X"B7",
		X"64",X"AC",X"F5",X"50",X"57",X"DD",X"BA",X"23",X"39",X"BE",X"87",X"01",X"49",X"8A",X"87",X"52",
		X"8E",X"FC",X"34",X"28",X"CA",X"F7",X"63",X"24",X"BC",X"D8",X"13",X"37",X"86",X"97",X"65",X"38",
		X"AD",X"CA",X"45",X"5B",X"B8",X"C2",X"A6",X"67",X"88",X"A5",X"57",X"69",X"64",X"85",X"A7",X"97",
		X"58",X"BA",X"F4",X"73",X"58",X"6A",X"B8",X"76",X"28",X"5D",X"C4",X"63",X"38",X"C9",X"87",X"74",
		X"56",X"7B",X"B8",X"B5",X"95",X"62",X"77",X"EC",X"C5",X"12",X"4A",X"AC",X"84",X"24",X"7B",X"C8",
		X"54",X"67",X"AA",X"A9",X"95",X"B6",X"94",X"67",X"79",X"8C",X"67",X"55",X"58",X"78",X"86",X"75",
		X"A8",X"69",X"87",X"96",X"77",X"58",X"4B",X"8D",X"58",X"46",X"78",X"BA",X"75",X"76",X"95",X"B6",
		X"66",X"69",X"88",X"95",X"67",X"97",X"76",X"67",X"87",X"89",X"77",X"35",X"A9",X"C6",X"64",X"37",
		X"7B",X"99",X"94",X"77",X"89",X"96",X"88",X"98",X"76",X"76",X"6A",X"9B",X"94",X"56",X"5A",X"97",
		X"86",X"66",X"7A",X"8A",X"85",X"75",X"7A",X"76",X"95",X"87",X"79",X"87",X"86",X"79",X"88",X"88",
		X"57",X"77",X"99",X"78",X"77",X"77",X"87",X"95",X"78",X"78",X"87",X"87",X"78",X"77",X"88",X"87",
		X"66",X"67",X"96",X"99",X"78",X"66",X"77",X"89",X"78",X"76",X"87",X"78",X"87",X"76",X"77",X"86",
		X"87",X"77",X"77",X"88",X"77",X"78",X"88",X"76",X"77",X"79",X"98",X"86",X"66",X"69",X"A8",X"86",
		X"77",X"79",X"88",X"76",X"78",X"98",X"76",X"76",X"88",X"88",X"76",X"77",X"89",X"77",X"65",X"88",
		X"88",X"77",X"86",X"88",X"87",X"76",X"68",X"88",X"87",X"77",X"78",X"88",X"77",X"87",X"89",X"87",
		X"76",X"88",X"89",X"77",X"67",X"89",X"88",X"77",X"77",X"88",X"87",X"77",X"77",X"88",X"78",X"67",
		X"77",X"88",X"88",X"67",X"76",X"88",X"87",X"77",X"87",X"78",X"78",X"87",X"87",X"77",X"77",X"78",
		X"88",X"77",X"76",X"78",X"87",X"77",X"88",X"78",X"67",X"78",X"88",X"77",X"77",X"78",X"77",X"87",
		X"88",X"78",X"67",X"87",X"87",X"78",X"77",X"88",X"78",X"76",X"77",X"78",X"87",X"87",X"77",X"77",
		X"78",X"87",X"77",X"77",X"87",X"88",X"77",X"77",X"87",X"88",X"87",X"77",X"87",X"77",X"78",X"77",
		X"77",X"77",X"88",X"78",X"77",X"77",X"88",X"77",X"78",X"87",X"77",X"78",X"77",X"87",X"77",X"78",
		X"87",X"77",X"78",X"78",X"88",X"77",X"87",X"88",X"78",X"77",X"77",X"78",X"88",X"87",X"66",X"77",
		X"88",X"87",X"77",X"78",X"88",X"77",X"77",X"79",X"67",X"68",X"88",X"87",X"78",X"88",X"97",X"97",
		X"67",X"76",X"77",X"77",X"67",X"78",X"87",X"46",X"69",X"87",X"56",X"78",X"89",X"86",X"66",X"67",
		X"76",X"77",X"76",X"77",X"67",X"87",X"78",X"98",X"7A",X"89",X"87",X"76",X"89",X"87",X"77",X"78",
		X"67",X"88",X"86",X"56",X"78",X"77",X"67",X"87",X"78",X"87",X"76",X"67",X"78",X"78",X"87",X"77",
		X"66",X"67",X"88",X"98",X"77",X"88",X"98",X"78",X"88",X"76",X"78",X"99",X"88",X"77",X"97",X"98",
		X"88",X"88",X"87",X"78",X"77",X"76",X"66",X"67",X"79",X"96",X"76",X"78",X"78",X"68",X"77",X"88",
		X"87",X"77",X"68",X"88",X"87",X"76",X"68",X"77",X"77",X"68",X"77",X"66",X"86",X"87",X"70",X"70",
		X"0F",X"FF",X"0F",X"0F",X"0F",X"FF",X"00",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"FF",X"0B",X"0F",
		X"0F",X"FF",X"00",X"0F",X"0F",X"F7",X"0F",X"0F",X"0F",X"F0",X"A0",X"07",X"7F",X"F0",X"F0",X"50",
		X"F8",X"F0",X"F0",X"81",X"FF",X"F0",X"F0",X"F0",X"FE",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",
		X"FD",X"F0",X"F0",X"F0",X"FF",X"F0",X"81",X"C1",X"FF",X"FC",X"00",X"0F",X"FF",X"F9",X"00",X"0F",
		X"FF",X"3F",X"03",X"0F",X"FF",X"E4",X"00",X"0F",X"9F",X"6D",X"06",X"0D",X"FF",X"F0",X"50",X"4D",
		X"DF",X"07",X"0F",X"0A",X"5F",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"0E",X"0F",X"FF",X"00",X"00",
		X"FF",X"F0",X"F0",X"B0",X"8F",X"FD",X"B0",X"00",X"FF",X"FF",X"F0",X"B0",X"FF",X"FF",X"F0",X"71",
		X"FF",X"F0",X"F0",X"B0",X"FF",X"FF",X"00",X"01",X"F1",X"F5",X"F0",X"F0",X"9E",X"1F",X"F9",X"0F",
		X"0F",X"FF",X"30",X"B0",X"FF",X"AF",X"9F",X"01",X"0F",X"F0",X"F0",X"F0",X"FD",X"F0",X"F0",X"F9",
		X"0F",X"F0",X"F0",X"F0",X"FF",X"FF",X"08",X"0F",X"FF",X"0F",X"00",X"F0",X"FF",X"EF",X"0F",X"0D",
		X"FB",X"F0",X"F0",X"FF",X"F4",X"F0",X"00",X"FF",X"F8",X"0B",X"0F",X"CF",X"06",X"F0",X"FE",X"9F",
		X"F2",X"0F",X"0F",X"F0",X"F0",X"CF",X"DF",X"0F",X"0B",X"F4",X"8F",X"FE",X"0F",X"0F",X"F0",X"20",
		X"0F",X"3F",X"00",X"F0",X"3E",X"FF",X"0F",X"00",X"F0",X"0F",X"0B",X"9F",X"F0",X"08",X"0F",X"0F",
		X"FF",X"30",X"F0",X"FF",X"00",X"60",X"FF",X"0A",X"FC",X"0F",X"0F",X"FF",X"0F",X"5F",X"50",X"FF",
		X"00",X"F0",X"F7",X"0F",X"6F",X"40",X"FF",X"0A",X"F0",X"F0",X"0F",X"0F",X"F0",X"FF",X"0F",X"30",
		X"F0",X"0F",X"04",X"F0",X"8F",X"0F",X"F0",X"F7",X"0F",X"B0",X"F0",X"0F",X"00",X"F2",X"0F",X"05",
		X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"FF",X"0F",X"F0",X"FF",X"0D",X"F0",X"3F",X"0F",X"F0",X"FF",
		X"81",X"FF",X"03",X"F0",X"0F",X"F0",X"FF",X"0F",X"F0",X"0F",X"E0",X"0F",X"00",X"F7",X"05",X"F3",
		X"0F",X"F0",X"FF",X"00",X"FF",X"00",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"FF",X"09",X"F8",
		X"0F",X"F7",X"0D",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"C0",X"0F",X"D0",X"FF",X"81",
		X"7F",X"E0",X"0F",X"B0",X"5F",X"90",X"FF",X"00",X"DF",X"00",X"FF",X"F0",X"FF",X"00",X"FF",X"00",
		X"FF",X"24",X"FB",X"04",X"FE",X"30",X"CF",X"06",X"F8",X"05",X"FF",X"91",X"FF",X"0F",X"F0",X"0F",
		X"F0",X"FF",X"F9",X"0F",X"E0",X"FF",X"00",X"FF",X"90",X"FF",X"00",X"F6",X"0F",X"F0",X"0F",X"D0",
		X"FF",X"00",X"F0",X"0F",X"F0",X"0F",X"0F",X"F0",X"0F",X"B0",X"FF",X"1F",X"00",X"F1",X"0F",X"F5",
		X"F0",X"0F",X"40",X"FF",X"FF",X"09",X"F0",X"65",X"00",X"00",X"00",X"CD",X"0F",X"FB",X"FF",X"0F",
		X"00",X"A3",X"90",X"03",X"50",X"00",X"CF",X"C0",X"0E",X"EB",X"00",X"FF",X"8F",X"FF",X"3C",X"FF",
		X"00",X"FF",X"00",X"FC",X"0F",X"F0",X"0F",X"CC",X"FD",X"08",X"E9",X"FB",X"02",X"C6",X"00",X"99",
		X"17",X"F4",X"01",X"D1",X"7E",X"EF",X"F0",X"7B",X"26",X"E9",X"FB",X"36",X"73",X"87",X"59",X"A5",
		X"89",X"CC",X"47",X"DA",X"9C",X"98",X"96",X"69",X"86",X"89",X"97",X"89",X"98",X"AB",X"AA",X"79",
		X"87",X"98",X"78",X"A9",X"99",X"89",X"88",X"99",X"98",X"68",X"87",X"79",X"88",X"88",X"70",X"70",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70",
		X"87",X"87",X"77",X"78",X"78",X"87",X"68",X"B9",X"56",X"6B",X"86",X"69",X"99",X"56",X"98",X"A4",
		X"79",X"97",X"47",X"9A",X"65",X"78",X"C6",X"84",X"97",X"77",X"6B",X"78",X"66",X"98",X"56",X"7A",
		X"96",X"66",X"7E",X"6A",X"08",X"A5",X"B2",X"C8",X"75",X"68",X"A9",X"56",X"79",X"86",X"88",X"76",
		X"98",X"B1",X"86",X"AA",X"39",X"5B",X"76",X"68",X"86",X"65",X"98",X"89",X"E6",X"60",X"6E",X"8B",
		X"1A",X"79",X"36",X"C9",X"90",X"68",X"B9",X"67",X"7F",X"28",X"19",X"F6",X"D0",X"C4",X"B5",X"6B",
		X"69",X"07",X"6D",X"A5",X"E5",X"C0",X"87",X"DD",X"09",X"0E",X"47",X"AB",X"81",X"14",X"FF",X"81",
		X"2F",X"B7",X"09",X"9E",X"51",X"76",X"F4",X"67",X"D8",X"00",X"8F",X"C3",X"5F",X"65",X"07",X"FB",
		X"B0",X"A7",X"D1",X"4E",X"A9",X"02",X"9F",X"C0",X"0A",X"F3",X"50",X"FF",X"49",X"0F",X"99",X"05",
		X"F7",X"71",X"7E",X"F5",X"2F",X"68",X"03",X"FF",X"B0",X"54",X"F3",X"5D",X"99",X"01",X"CF",X"B0",
		X"1F",X"E8",X"05",X"DF",X"71",X"57",X"F2",X"79",X"EB",X"02",X"7F",X"A6",X"B3",X"B0",X"7C",X"FF",
		X"05",X"3F",X"4B",X"A6",X"71",X"7A",X"F5",X"0B",X"BB",X"02",X"6F",X"94",X"36",X"E4",X"74",X"D6",
		X"22",X"8E",X"6A",X"F7",X"30",X"3F",X"FB",X"07",X"4F",X"25",X"BA",X"60",X"8E",X"E5",X"AC",X"B0",
		X"04",X"FF",X"60",X"3F",X"E8",X"18",X"43",X"4A",X"F7",X"C9",X"83",X"05",X"FC",X"C0",X"4B",X"FB",
		X"35",X"24",X"0D",X"DD",X"D9",X"30",X"14",X"FB",X"B0",X"38",X"BE",X"6A",X"01",X"1A",X"E9",X"FC",
		X"90",X"04",X"FF",X"81",X"28",X"AB",X"79",X"52",X"09",X"DB",X"F7",X"B0",X"11",X"FC",X"A1",X"0A",
		X"9F",X"25",X"24",X"99",X"C7",X"F3",X"B0",X"8A",X"CE",X"0B",X"0F",X"4D",X"41",X"30",X"EC",X"F9",
		X"64",X"04",X"4F",X"5C",X"06",X"99",X"D5",X"81",X"24",X"FF",X"DF",X"06",X"0B",X"DC",X"E0",X"90",
		X"F6",X"E5",X"01",X"0D",X"BF",X"F2",X"50",X"86",X"FA",X"44",X"0D",X"4F",X"48",X"00",X"3B",X"FF",
		X"84",X"03",X"8F",X"B7",X"33",X"B6",X"E6",X"90",X"14",X"CE",X"FE",X"50",X"05",X"FE",X"A0",X"69",
		X"89",X"8A",X"10",X"08",X"DF",X"F5",X"20",X"4F",X"DE",X"08",X"4C",X"77",X"A3",X"30",X"5B",X"FF",
		X"81",X"03",X"FD",X"D1",X"74",X"A8",X"88",X"36",X"08",X"8F",X"FA",X"20",X"3F",X"EE",X"09",X"3E",
		X"48",X"64",X"81",X"97",X"FF",X"C0",X"01",X"FF",X"C0",X"74",X"E4",X"88",X"66",X"06",X"9F",X"FC",
		X"00",X"1F",X"EB",X"16",X"7B",X"73",X"A5",X"60",X"5B",X"FF",X"C0",X"01",X"FE",X"B0",X"39",X"DB",
		X"26",X"58",X"02",X"8F",X"FC",X"00",X"0F",X"DC",X"06",X"6D",X"B3",X"65",X"90",X"36",X"FF",X"E4",
		X"00",X"CB",X"F0",X"92",X"E8",X"53",X"5B",X"35",X"2A",X"FF",X"D0",X"05",X"CF",X"87",X"0E",X"6D",
		X"16",X"3A",X"51",X"4E",X"FF",X"60",X"0B",X"DF",X"48",X"1D",X"88",X"43",X"A3",X"91",X"9F",X"FF",
		X"00",X"0E",X"FF",X"62",X"4A",X"85",X"64",X"92",X"85",X"9F",X"FF",X"01",X"0E",X"CF",X"90",X"46",
		X"E7",X"52",X"73",X"87",X"9A",X"FD",X"50",X"07",X"7F",X"96",X"06",X"CC",X"81",X"24",X"E9",X"53",
		X"DF",X"D4",X"00",X"9B",X"F5",X"61",X"BC",X"C2",X"04",X"AE",X"72",X"3C",X"FE",X"50",X"07",X"AF",
		X"69",X"3D",X"69",X"35",X"8B",X"B3",X"34",X"EF",X"BC",X"02",X"06",X"ED",X"F3",X"50",X"B7",X"F3",
		X"71",X"46",X"CD",X"8F",X"5D",X"02",X"17",X"FC",X"A0",X"53",X"FA",X"A0",X"03",X"EF",X"9A",X"29",
		X"AF",X"76",X"04",X"6D",X"DA",X"6A",X"88",X"64",X"71",X"A6",X"C4",X"69",X"BF",X"87",X"10",X"54",
		X"FB",X"C0",X"64",X"EB",X"65",X"04",X"9F",X"A6",X"54",X"BA",X"F2",X"71",X"87",X"EA",X"73",X"6C",
		X"8E",X"66",X"03",X"6C",X"D9",X"A1",X"68",X"9F",X"58",X"01",X"7E",X"E8",X"71",X"B8",X"E3",X"41",
		X"7A",X"9C",X"5A",X"59",X"7B",X"A3",X"90",X"95",X"E9",X"83",X"28",X"8E",X"79",X"04",X"3B",X"CB",
		X"94",X"43",X"9A",X"F5",X"90",X"87",X"E8",X"73",X"59",X"BF",X"8A",X"07",X"2A",X"7A",X"88",X"86",
		X"87",X"9D",X"59",X"06",X"4D",X"89",X"76",X"9A",X"C6",X"52",X"46",X"8B",X"8B",X"76",X"66",X"A7",
		X"A5",X"86",X"88",X"86",X"95",X"96",X"69",X"7D",X"86",X"25",X"79",X"97",X"76",X"87",X"79",X"98",
		X"83",X"97",X"A8",X"53",X"86",X"D6",X"88",X"8C",X"67",X"26",X"69",X"78",X"99",X"A4",X"75",X"8A",
		X"A5",X"75",X"B7",X"B5",X"84",X"96",X"8A",X"8A",X"48",X"38",X"7A",X"67",X"6A",X"8A",X"76",X"56",
		X"77",X"B8",X"95",X"58",X"7C",X"59",X"37",X"69",X"89",X"79",X"77",X"65",X"87",X"99",X"88",X"67",
		X"89",X"86",X"65",X"98",X"B7",X"95",X"67",X"78",X"97",X"77",X"67",X"49",X"89",X"85",X"65",X"98",
		X"C8",X"83",X"47",X"9B",X"77",X"67",X"9A",X"98",X"46",X"49",X"9A",X"95",X"75",X"A7",X"A5",X"75",
		X"78",X"88",X"77",X"68",X"79",X"78",X"67",X"58",X"7A",X"77",X"77",X"98",X"86",X"75",X"76",X"89",
		X"89",X"78",X"66",X"49",X"79",X"87",X"78",X"A9",X"85",X"55",X"88",X"98",X"89",X"88",X"67",X"69",
		X"79",X"56",X"68",X"B7",X"95",X"85",X"87",X"88",X"77",X"68",X"88",X"86",X"67",X"77",X"77",X"78",
		X"88",X"76",X"77",X"88",X"77",X"68",X"77",X"A7",X"96",X"76",X"98",X"87",X"67",X"78",X"77",X"78",
		X"87",X"77",X"87",X"87",X"77",X"78",X"87",X"86",X"88",X"97",X"76",X"67",X"79",X"88",X"76",X"78",
		X"98",X"76",X"77",X"97",X"87",X"77",X"78",X"88",X"67",X"69",X"88",X"77",X"77",X"77",X"78",X"78",
		X"78",X"77",X"77",X"88",X"87",X"88",X"87",X"77",X"77",X"87",X"87",X"86",X"97",X"87",X"86",X"76",
		X"88",X"98",X"76",X"67",X"89",X"87",X"67",X"78",X"78",X"78",X"77",X"77",X"77",X"88",X"87",X"87",
		X"87",X"76",X"78",X"99",X"87",X"66",X"88",X"97",X"76",X"77",X"89",X"97",X"66",X"79",X"98",X"66",
		X"78",X"97",X"76",X"78",X"98",X"77",X"67",X"78",X"89",X"87",X"66",X"78",X"88",X"77",X"77",X"88",
		X"87",X"76",X"77",X"89",X"88",X"67",X"78",X"88",X"87",X"66",X"78",X"98",X"76",X"66",X"88",X"87",
		X"77",X"77",X"88",X"88",X"67",X"68",X"89",X"87",X"67",X"78",X"87",X"78",X"88",X"77",X"78",X"77",
		X"77",X"77",X"88",X"88",X"77",X"77",X"77",X"88",X"88",X"77",X"77",X"88",X"87",X"77",X"77",X"88",
		X"88",X"67",X"78",X"87",X"76",X"77",X"88",X"78",X"77",X"77",X"88",X"87",X"67",X"88",X"87",X"77",
		X"88",X"87",X"77",X"78",X"77",X"77",X"87",X"77",X"77",X"87",X"77",X"77",X"87",X"87",X"87",X"78",
		X"78",X"77",X"77",X"78",X"88",X"77",X"77",X"87",X"77",X"77",X"77",X"88",X"87",X"77",X"77",X"88",
		X"87",X"77",X"78",X"88",X"77",X"78",X"88",X"87",X"77",X"78",X"88",X"77",X"77",X"77",X"88",X"87",
		X"77",X"78",X"77",X"77",X"88",X"87",X"67",X"78",X"87",X"78",X"77",X"77",X"88",X"77",X"77",X"88",
		X"87",X"77",X"78",X"78",X"87",X"76",X"77",X"88",X"77",X"77",X"88",X"87",X"77",X"78",X"88",X"77",
		X"77",X"77",X"88",X"87",X"77",X"88",X"77",X"77",X"87",X"77",X"78",X"88",X"77",X"78",X"87",X"77",
		X"78",X"87",X"78",X"87",X"77",X"77",X"88",X"77",X"77",X"88",X"87",X"77",X"77",X"78",X"87",X"77",
		X"77",X"87",X"87",X"77",X"78",X"88",X"87",X"77",X"78",X"78",X"77",X"78",X"78",X"87",X"87",X"87",
		X"78",X"87",X"78",X"88",X"87",X"77",X"88",X"88",X"78",X"77",X"87",X"77",X"78",X"78",X"87",X"77",
		X"77",X"78",X"77",X"78",X"78",X"77",X"87",X"88",X"89",X"77",X"78",X"88",X"77",X"87",X"87",X"77",
		X"67",X"77",X"87",X"87",X"88",X"87",X"77",X"78",X"88",X"77",X"87",X"86",X"78",X"77",X"77",X"68",
		X"88",X"87",X"87",X"78",X"76",X"87",X"78",X"67",X"77",X"97",X"89",X"78",X"76",X"87",X"79",X"67",
		X"77",X"87",X"77",X"77",X"76",X"88",X"77",X"77",X"88",X"87",X"88",X"88",X"87",X"78",X"67",X"88",
		X"67",X"97",X"58",X"67",X"95",X"7A",X"88",X"78",X"95",X"A8",X"76",X"77",X"88",X"97",X"78",X"78",
		X"86",X"78",X"67",X"77",X"97",X"57",X"87",X"67",X"A8",X"9A",X"67",X"87",X"98",X"93",X"8A",X"77",
		X"68",X"57",X"78",X"87",X"76",X"A7",X"59",X"68",X"77",X"A8",X"78",X"6A",X"64",X"79",X"67",X"66",
		X"86",X"88",X"97",X"48",X"58",X"A8",X"56",X"64",X"66",X"76",X"88",X"65",X"8A",X"79",X"66",X"85",
		X"66",X"6A",X"47",X"67",X"77",X"76",X"58",X"78",X"88",X"6A",X"97",X"6B",X"67",X"A5",X"87",X"69",
		X"58",X"55",X"86",X"A8",X"68",X"78",X"78",X"9A",X"85",X"96",X"58",X"5A",X"67",X"B5",X"97",X"69",
		X"67",X"66",X"68",X"87",X"A5",X"A5",X"88",X"2B",X"97",X"D6",X"8A",X"69",X"56",X"84",X"A9",X"68",
		X"68",X"76",X"99",X"7A",X"88",X"B7",X"87",X"8A",X"5A",X"56",X"A7",X"C5",X"9A",X"89",X"8A",X"7A",
		X"67",X"79",X"86",X"97",X"74",X"89",X"6A",X"7A",X"74",X"A7",X"85",X"8A",X"59",X"59",X"88",X"94",
		X"98",X"97",X"68",X"46",X"65",X"6A",X"76",X"A9",X"65",X"D7",X"8B",X"65",X"68",X"75",X"87",X"5A",
		X"39",X"87",X"99",X"AA",X"89",X"96",X"99",X"8A",X"86",X"66",X"76",X"9A",X"59",X"75",X"7A",X"78",
		X"98",X"74",X"B7",X"58",X"58",X"77",X"88",X"77",X"6B",X"69",X"96",X"88",X"87",X"86",X"69",X"86",
		X"99",X"98",X"B6",X"68",X"A7",X"88",X"86",X"A8",X"55",X"75",X"86",X"65",X"A4",X"7B",X"46",X"56",
		X"49",X"A4",X"AB",X"48",X"B6",X"88",X"95",X"78",X"68",X"94",X"89",X"96",X"8A",X"84",X"79",X"78",
		X"87",X"56",X"68",X"69",X"56",X"83",X"97",X"58",X"67",X"88",X"97",X"59",X"68",X"A5",X"59",X"65",
		X"67",X"84",X"A6",X"6B",X"67",X"97",X"68",X"89",X"87",X"96",X"86",X"5A",X"75",X"A5",X"69",X"49",
		X"95",X"86",X"59",X"57",X"94",X"97",X"69",X"69",X"A6",X"B8",X"66",X"6A",X"68",X"67",X"B5",X"99",
		X"69",X"77",X"85",X"A7",X"6A",X"66",X"85",X"85",X"67",X"86",X"87",X"59",X"76",X"97",X"49",X"47",
		X"78",X"A6",X"79",X"38",X"86",X"98",X"8B",X"67",X"86",X"77",X"57",X"69",X"75",X"B7",X"7B",X"79",
		X"A7",X"65",X"86",X"96",X"97",X"76",X"6B",X"48",X"83",X"89",X"5A",X"57",X"59",X"86",X"58",X"68",
		X"A4",X"A8",X"86",X"69",X"78",X"66",X"75",X"94",X"86",X"8A",X"59",X"98",X"75",X"97",X"77",X"76",
		X"95",X"6A",X"79",X"67",X"B5",X"78",X"7B",X"48",X"94",X"86",X"89",X"5A",X"88",X"68",X"77",X"96",
		X"87",X"88",X"79",X"87",X"68",X"78",X"86",X"96",X"89",X"5A",X"87",X"96",X"78",X"88",X"56",X"A5",
		X"68",X"5A",X"78",X"75",X"A6",X"89",X"79",X"79",X"68",X"79",X"5B",X"77",X"86",X"86",X"78",X"79",
		X"78",X"95",X"A5",X"A6",X"69",X"49",X"66",X"86",X"96",X"78",X"69",X"97",X"99",X"69",X"69",X"48",
		X"66",X"96",X"85",X"96",X"87",X"69",X"59",X"59",X"85",X"87",X"98",X"6A",X"85",X"97",X"70",X"70",
		X"88",X"88",X"77",X"8A",X"00",X"C0",X"FC",X"0C",X"F9",X"08",X"71",X"0F",X"90",X"FF",X"A8",X"FF",
		X"FA",X"F6",X"F8",X"09",X"00",X"FA",X"20",X"00",X"0B",X"69",X"95",X"F6",X"F0",X"F9",X"FF",X"F0",
		X"FA",X"DF",X"0A",X"FD",X"00",X"00",X"0C",X"FF",X"00",X"BF",X"7F",X"FF",X"FE",X"2F",X"07",X"5F",
		X"D0",X"00",X"D9",X"00",X"F0",X"F0",X"60",X"EF",X"FF",X"FF",X"FF",X"FE",X"F6",X"BB",X"81",X"00",
		X"48",X"07",X"D0",X"40",X"1F",X"FE",X"F9",X"F5",X"FF",X"FF",X"FF",X"C0",X"F2",X"95",X"30",X"00",
		X"00",X"AF",X"EF",X"F9",X"CF",X"FF",X"FF",X"FF",X"0F",X"19",X"0A",X"30",X"00",X"0F",X"C5",X"0A",
		X"5D",X"FF",X"FF",X"FF",X"00",X"F0",X"FF",X"90",X"00",X"B2",X"81",X"00",X"C5",X"FF",X"FF",X"FF",
		X"F0",X"AF",X"6F",X"D0",X"00",X"0B",X"F0",X"00",X"00",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"60",
		X"0A",X"00",X"09",X"00",X"00",X"0F",X"6F",X"FF",X"FF",X"FF",X"FF",X"FC",X"08",X"04",X"46",X"00",
		X"00",X"6F",X"F5",X"77",X"FD",X"FF",X"FF",X"85",X"FF",X"3F",X"B1",X"00",X"00",X"30",X"20",X"41",
		X"CF",X"FF",X"FF",X"14",X"FF",X"DF",X"B3",X"02",X"20",X"A0",X"00",X"00",X"4F",X"FF",X"FF",X"CF",
		X"F7",X"FC",X"00",X"08",X"C9",X"D0",X"00",X"00",X"2F",X"BF",X"FF",X"FF",X"FF",X"F4",X"00",X"00",
		X"2A",X"01",X"00",X"09",X"B4",X"0F",X"F6",X"FF",X"FF",X"FF",X"CC",X"00",X"89",X"00",X"00",X"67",
		X"50",X"9F",X"34",X"FF",X"FF",X"FF",X"FA",X"3F",X"FA",X"00",X"00",X"30",X"04",X"30",X"0F",X"FF",
		X"FF",X"FF",X"9B",X"FF",X"F1",X"21",X"00",X"00",X"00",X"00",X"6F",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"30",X"60",X"5C",X"3D",X"00",X"00",X"30",X"AA",X"FF",X"FF",X"FF",X"FC",X"06",X"10",X"23",X"26",
		X"00",X"39",X"53",X"A2",X"36",X"BF",X"FF",X"FF",X"FF",X"3A",X"40",X"00",X"00",X"84",X"89",X"C1",
		X"09",X"6F",X"FF",X"FF",X"FC",X"FF",X"F3",X"10",X"00",X"00",X"02",X"00",X"7C",X"FF",X"EF",X"FB",
		X"A8",X"FF",X"F8",X"62",X"75",X"03",X"00",X"00",X"5A",X"FF",X"FF",X"FC",X"CF",X"FC",X"45",X"07",
		X"68",X"C8",X"00",X"00",X"10",X"45",X"FF",X"FF",X"FF",X"FD",X"B7",X"05",X"0A",X"81",X"00",X"71",
		X"61",X"01",X"04",X"BF",X"FF",X"FF",X"FB",X"D7",X"98",X"00",X"00",X"13",X"68",X"20",X"05",X"CF",
		X"DD",X"FF",X"FF",X"FF",X"FA",X"00",X"00",X"00",X"00",X"00",X"1D",X"FF",X"FD",X"F7",X"CF",X"FF",
		X"EA",X"6A",X"62",X"60",X"00",X"00",X"07",X"8F",X"FF",X"FE",X"FF",X"FE",X"35",X"77",X"6C",X"E7",
		X"20",X"00",X"00",X"05",X"88",X"9F",X"FF",X"FF",X"C8",X"61",X"88",X"71",X"16",X"6B",X"30",X"00",
		X"00",X"9D",X"FF",X"FF",X"FF",X"AC",X"D4",X"00",X"00",X"28",X"88",X"30",X"16",X"D5",X"BD",X"FF",
		X"FF",X"FF",X"F9",X"61",X"00",X"00",X"20",X"00",X"7C",X"AC",X"BC",X"AC",X"BF",X"FF",X"FD",X"F9",
		X"68",X"64",X"00",X"00",X"12",X"7B",X"B9",X"BF",X"FF",X"FC",X"B9",X"B7",X"DC",X"99",X"43",X"00",
		X"00",X"32",X"02",X"9F",X"FF",X"FF",X"FB",X"67",X"B7",X"23",X"24",X"75",X"35",X"60",X"00",X"39",
		X"EF",X"FF",X"FF",X"FF",X"F8",X"10",X"00",X"41",X"46",X"61",X"36",X"37",X"79",X"AE",X"DE",X"FF",
		X"FF",X"C6",X"33",X"20",X"10",X"00",X"57",X"7A",X"AA",X"98",X"9B",X"FF",X"FF",X"FB",X"BB",X"A8",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70",
		X"77",X"77",X"76",X"67",X"77",X"78",X"88",X"99",X"98",X"88",X"87",X"76",X"66",X"67",X"77",X"88",
		X"88",X"88",X"87",X"77",X"76",X"66",X"67",X"78",X"89",X"99",X"99",X"88",X"77",X"66",X"66",X"77",
		X"88",X"88",X"88",X"88",X"77",X"76",X"66",X"66",X"78",X"89",X"99",X"99",X"88",X"77",X"66",X"66",
		X"77",X"77",X"88",X"88",X"87",X"77",X"66",X"66",X"67",X"88",X"99",X"99",X"88",X"87",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"87",X"77",X"77",X"77",
		X"77",X"77",X"78",X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"67",X"77",X"78",X"88",X"88",X"88",X"87",X"77",X"77",X"77",X"88",X"87",X"77",X"76",
		X"66",X"77",X"78",X"99",X"98",X"88",X"87",X"77",X"77",X"78",X"87",X"77",X"77",X"66",X"66",X"78",
		X"89",X"99",X"88",X"87",X"76",X"67",X"88",X"87",X"77",X"76",X"66",X"67",X"89",X"99",X"99",X"88",
		X"76",X"66",X"78",X"87",X"88",X"86",X"66",X"68",X"89",X"99",X"89",X"87",X"65",X"67",X"77",X"78",
		X"87",X"65",X"68",X"9A",X"99",X"9A",X"85",X"34",X"56",X"67",X"8B",X"A7",X"46",X"AB",X"A9",X"9B",
		X"B7",X"11",X"46",X"44",X"8B",X"C9",X"57",X"AC",X"A8",X"8A",X"96",X"24",X"77",X"46",X"9A",X"96",
		X"79",X"B9",X"78",X"A8",X"64",X"69",X"63",X"6A",X"97",X"58",X"BB",X"76",X"78",X"62",X"3A",X"A5",
		X"56",X"B8",X"48",X"CE",X"CA",X"66",X"60",X"05",X"9A",X"65",X"97",X"6C",X"CE",X"DA",X"56",X"61",
		X"38",X"A8",X"44",X"88",X"BC",X"CC",X"B4",X"25",X"44",X"8C",X"93",X"17",X"9A",X"BB",X"C8",X"12",
		X"59",X"8A",X"EA",X"30",X"7A",X"CB",X"BA",X"50",X"46",X"98",X"9C",X"72",X"39",X"BA",X"99",X"84",
		X"15",X"78",X"79",X"B7",X"37",X"CC",X"A8",X"A6",X"21",X"68",X"56",X"AB",X"64",X"AF",X"A8",X"8A",
		X"40",X"58",X"83",X"8B",X"84",X"8C",X"C7",X"7A",X"73",X"5A",X"C4",X"39",X"A5",X"5B",X"EA",X"26",
		X"76",X"4B",X"E9",X"13",X"85",X"29",X"EF",X"76",X"56",X"5A",X"FD",X"72",X"62",X"86",X"EE",X"83",
		X"42",X"65",X"87",X"73",X"55",X"98",X"C9",X"96",X"45",X"99",X"48",X"76",X"15",X"8F",X"7C",X"56",
		X"57",X"D6",X"78",X"84",X"37",X"FC",X"E7",X"85",X"7A",X"99",X"67",X"89",X"BC",X"7C",X"43",X"46",
		X"94",X"78",X"52",X"4C",X"D5",X"A8",X"47",X"7D",X"71",X"25",X"75",X"CF",X"B9",X"95",X"AB",X"83",
		X"48",X"78",X"DB",X"48",X"A3",X"6A",X"B9",X"01",X"44",X"5B",X"9B",X"4A",X"BA",X"E6",X"73",X"05",
		X"9F",X"D9",X"37",X"49",X"A4",X"60",X"27",X"5F",X"F8",X"83",X"39",X"87",X"34",X"74",X"9C",X"FA",
		X"8A",X"48",X"E8",X"83",X"92",X"6C",X"BB",X"9C",X"39",X"C9",X"52",X"72",X"5B",X"AD",X"7A",X"56",
		X"D4",X"A7",X"73",X"5A",X"8B",X"59",X"76",X"B3",X"84",X"24",X"88",X"77",X"84",X"8B",X"39",X"34",
		X"63",X"AB",X"A7",X"A3",X"8C",X"59",X"57",X"55",X"E8",X"C8",X"A8",X"7D",X"59",X"76",X"56",X"D6",
		X"98",X"46",X"87",X"76",X"86",X"5C",X"7A",X"63",X"A7",X"99",X"67",X"54",X"8B",X"AB",X"29",X"47",
		X"F8",X"C4",X"58",X"8C",X"E8",X"68",X"47",X"6A",X"81",X"46",X"98",X"93",X"72",X"4A",X"3A",X"93",
		X"77",X"C7",X"CB",X"24",X"B4",X"AA",X"9B",X"5B",X"D5",X"7B",X"61",X"9A",X"6B",X"77",X"58",X"6B",
		X"C3",X"47",X"5B",X"5D",X"C1",X"6A",X"88",X"D6",X"47",X"5A",X"A6",X"B6",X"53",X"89",X"CA",X"66",
		X"83",X"8C",X"7A",X"A7",X"58",X"76",X"86",X"68",X"88",X"87",X"76",X"68",X"78",X"77",X"78",X"7A",
		X"98",X"76",X"87",X"89",X"C5",X"89",X"57",X"C5",X"96",X"86",X"77",X"B8",X"96",X"37",X"89",X"5C",
		X"73",X"86",X"4A",X"85",X"A8",X"78",X"88",X"5B",X"48",X"86",X"96",X"99",X"A6",X"74",X"66",X"BA",
		X"59",X"67",X"9B",X"67",X"A5",X"4C",X"B5",X"A7",X"48",X"7B",X"9C",X"27",X"48",X"AD",X"76",X"55",
		X"A7",X"9B",X"63",X"46",X"7A",X"94",X"68",X"39",X"D5",X"77",X"54",X"9A",X"A8",X"A6",X"48",X"98",
		X"7A",X"76",X"76",X"A7",X"B7",X"75",X"A1",X"98",X"8A",X"85",X"4B",X"58",X"98",X"47",X"76",X"88",
		X"77",X"87",X"89",X"88",X"77",X"77",X"88",X"88",X"88",X"78",X"87",X"88",X"87",X"88",X"88",X"88",
		X"88",X"77",X"88",X"78",X"88",X"68",X"99",X"79",X"36",X"59",X"7D",X"A6",X"86",X"68",X"97",X"66",
		X"67",X"8A",X"8A",X"56",X"79",X"77",X"84",X"55",X"AA",X"A6",X"87",X"66",X"77",X"58",X"79",X"A9",
		X"75",X"96",X"97",X"89",X"85",X"9B",X"69",X"67",X"49",X"5A",X"57",X"57",X"88",X"B6",X"58",X"87",
		X"98",X"77",X"57",X"C8",X"87",X"63",X"86",X"9D",X"73",X"8B",X"6A",X"A6",X"39",X"57",X"C8",X"48",
		X"67",X"98",X"98",X"56",X"88",X"A9",X"29",X"87",X"8B",X"64",X"95",X"5C",X"82",X"69",X"6A",X"76",
		X"87",X"3C",X"B8",X"75",X"69",X"B7",X"98",X"46",X"97",X"CA",X"24",X"C6",X"C9",X"75",X"74",X"8B",
		X"98",X"38",X"69",X"6C",X"63",X"96",X"8E",X"72",X"59",X"6B",X"86",X"97",X"3D",X"C6",X"66",X"5A",
		X"96",X"96",X"28",X"6C",X"9A",X"45",X"78",X"D8",X"58",X"63",X"B7",X"98",X"56",X"B7",X"59",X"64",
		X"95",X"AA",X"64",X"89",X"7C",X"75",X"75",X"4D",X"98",X"66",X"7A",X"C6",X"89",X"68",X"A7",X"A8",
		X"58",X"C7",X"8A",X"57",X"93",X"C8",X"47",X"66",X"8C",X"38",X"83",X"88",X"68",X"63",X"6B",X"95",
		X"97",X"7A",X"4A",X"B6",X"58",X"A7",X"7B",X"66",X"93",X"8A",X"55",X"89",X"6A",X"69",X"A6",X"68",
		X"59",X"95",X"87",X"C5",X"6C",X"57",X"94",X"AA",X"55",X"B8",X"39",X"8A",X"B3",X"9A",X"45",X"8B",
		X"75",X"97",X"7B",X"38",X"B5",X"48",X"A7",X"96",X"5A",X"86",X"85",X"78",X"68",X"8A",X"66",X"B6",
		X"6A",X"58",X"86",X"69",X"A4",X"8B",X"7A",X"55",X"96",X"38",X"C9",X"29",X"B7",X"B3",X"7B",X"54",
		X"7C",X"86",X"67",X"AA",X"3B",X"75",X"77",X"89",X"95",X"5D",X"84",X"C4",X"78",X"48",X"CB",X"15",
		X"C8",X"B5",X"6C",X"53",X"8B",X"B2",X"89",X"6D",X"39",X"B3",X"38",X"9A",X"85",X"5A",X"94",X"A6",
		X"68",X"37",X"AA",X"53",X"D7",X"4B",X"48",X"94",X"6C",X"C2",X"6B",X"9A",X"47",X"B5",X"58",X"8A",
		X"57",X"77",X"96",X"88",X"77",X"78",X"87",X"77",X"77",X"77",X"77",X"77",X"77",X"87",X"78",X"78",
		X"77",X"87",X"68",X"98",X"77",X"78",X"96",X"88",X"77",X"78",X"88",X"77",X"88",X"78",X"77",X"77",
		X"78",X"87",X"78",X"87",X"67",X"88",X"57",X"99",X"66",X"96",X"97",X"5A",X"73",X"8A",X"A5",X"67",
		X"8B",X"37",X"B5",X"58",X"9A",X"69",X"48",X"C2",X"99",X"47",X"66",X"CB",X"23",X"B9",X"84",X"3D",
		X"91",X"7D",X"B2",X"8A",X"4C",X"44",X"D5",X"2B",X"A7",X"85",X"4B",X"95",X"76",X"98",X"36",X"AC",
		X"62",X"E7",X"5B",X"39",X"B1",X"5D",X"B1",X"69",X"9B",X"17",X"C7",X"25",X"BA",X"49",X"67",X"E1",
		X"6C",X"44",X"87",X"9B",X"33",X"CB",X"84",X"5D",X"82",X"48",X"D5",X"4D",X"59",X"92",X"CA",X"16",
		X"BB",X"37",X"86",X"D3",X"3D",X"72",X"9A",X"A4",X"95",X"7E",X"16",X"C4",X"58",X"69",X"B3",X"2D",
		X"A7",X"44",X"D9",X"15",X"9D",X"53",X"C8",X"89",X"4A",X"A2",X"69",X"C4",X"58",X"8C",X"53",X"B8",
		X"37",X"8C",X"57",X"67",X"D6",X"3B",X"72",X"89",X"98",X"72",X"BD",X"38",X"77",X"93",X"5B",X"C4",
		X"1C",X"A6",X"A4",X"AB",X"14",X"BE",X"23",X"B7",X"A8",X"1C",X"A0",X"79",X"E4",X"19",X"79",X"A1",
		X"BC",X"14",X"CC",X"46",X"78",X"D3",X"5C",X"75",X"58",X"D7",X"94",X"8F",X"35",X"C5",X"47",X"7C",
		X"79",X"36",X"F4",X"4A",X"75",X"77",X"B9",X"83",X"8E",X"46",X"86",X"74",X"59",X"C9",X"19",X"E4",
		X"98",X"48",X"54",X"9B",X"82",X"9D",X"58",X"75",X"85",X"58",X"B9",X"3A",X"D5",X"98",X"69",X"34",
		X"8C",X"92",X"AE",X"38",X"73",X"84",X"48",X"B9",X"29",X"F4",X"68",X"48",X"65",X"9A",X"A1",X"9F",
		X"48",X"86",X"A3",X"3A",X"E6",X"1A",X"D5",X"A7",X"4A",X"34",X"9C",X"91",X"9F",X"45",X"64",X"A5",
		X"6A",X"AA",X"26",X"F5",X"39",X"78",X"75",X"89",X"B3",X"7F",X"52",X"B7",X"68",X"57",X"AA",X"29",
		X"F3",X"49",X"57",X"85",X"7B",X"90",X"9F",X"37",X"84",X"97",X"49",X"9A",X"25",X"F6",X"18",X"87",
		X"87",X"A9",X"94",X"5E",X"A0",X"6B",X"57",X"7D",X"96",X"66",X"BA",X"06",X"B5",X"66",X"D8",X"58",
		X"89",X"C1",X"4D",X"52",X"8E",X"54",X"A7",X"8C",X"14",X"D4",X"47",X"E6",X"49",X"89",X"C1",X"5D",
		X"44",X"5D",X"A2",X"7D",X"67",X"53",X"D9",X"56",X"AC",X"36",X"E5",X"59",X"59",X"96",X"79",X"C4",
		X"5E",X"73",X"A6",X"68",X"76",X"7B",X"35",X"E6",X"3B",X"65",X"97",X"96",X"A6",X"4D",X"A1",X"99",
		X"58",X"8C",X"67",X"86",X"9B",X"26",X"B5",X"57",X"D8",X"38",X"85",X"86",X"4B",X"63",X"8E",X"82",
		X"9B",X"59",X"64",X"B6",X"38",X"E6",X"3A",X"96",X"A5",X"3C",X"53",X"AE",X"54",X"99",X"7A",X"44",
		X"B6",X"39",X"D6",X"59",X"89",X"A3",X"59",X"73",X"6C",X"A3",X"8D",X"54",X"97",X"78",X"67",X"AC",
		X"45",X"F7",X"29",X"87",X"74",X"6C",X"B1",X"8E",X"46",X"95",X"A6",X"29",X"C5",X"86",X"4E",X"52",
		X"A6",X"68",X"27",X"F6",X"1A",X"B6",X"96",X"4C",X"51",X"AD",X"57",X"96",X"9A",X"26",X"D3",X"49",
		X"79",X"B5",X"5E",X"61",X"B9",X"58",X"46",X"E8",X"1A",X"D3",X"7A",X"69",X"81",X"9F",X"44",X"A7",
		X"7A",X"26",X"D5",X"39",X"89",X"B4",X"7E",X"43",X"B9",X"57",X"48",X"D5",X"4A",X"77",X"A4",X"7B",
		X"63",X"77",X"C8",X"2A",X"B3",X"88",X"79",X"42",X"79",X"9A",X"36",X"D6",X"4A",X"A7",X"53",X"BD",
		X"78",X"66",X"C6",X"4B",X"95",X"34",X"CD",X"47",X"75",X"A7",X"3A",X"B2",X"38",X"BB",X"47",X"85",
		X"98",X"5C",X"72",X"67",X"BB",X"58",X"64",X"B9",X"68",X"64",X"55",X"A8",X"8A",X"26",X"C5",X"6A",
		X"55",X"55",X"8A",X"B4",X"4B",X"85",X"A7",X"69",X"35",X"9B",X"B4",X"8A",X"57",X"B4",X"88",X"46",
		X"68",X"99",X"93",X"6D",X"65",X"96",X"67",X"47",X"CC",X"33",X"C9",X"4A",X"67",X"B2",X"48",X"B8",
		X"5A",X"75",X"B5",X"5C",X"73",X"78",X"79",X"C5",X"8A",X"37",X"C4",X"6A",X"45",X"77",X"8D",X"53",
		X"98",X"79",X"57",X"A6",X"45",X"A8",X"A4",X"4A",X"94",X"A9",X"8A",X"43",X"7A",X"8B",X"76",X"A4",
		X"5D",X"86",X"B4",X"37",X"99",X"B5",X"66",X"58",X"96",X"99",X"44",X"6B",X"B7",X"5A",X"65",X"77",
		X"8A",X"63",X"67",X"78",X"8A",X"93",X"68",X"79",X"86",X"95",X"37",X"BA",X"77",X"96",X"48",X"99",
		X"95",X"37",X"88",X"89",X"A6",X"75",X"7A",X"A4",X"89",X"54",X"89",X"99",X"88",X"74",X"6A",X"A7",
		X"66",X"66",X"69",X"A8",X"87",X"76",X"6A",X"97",X"57",X"76",X"79",X"96",X"99",X"75",X"78",X"95",
		X"6A",X"74",X"6A",X"96",X"5B",X"C5",X"27",X"C8",X"37",X"C7",X"36",X"B9",X"45",X"BC",X"43",X"9B",
		X"64",X"6C",X"92",X"5B",X"A4",X"5A",X"C7",X"25",X"BA",X"35",X"AB",X"43",X"9C",X"63",X"8E",X"A2",
		X"4B",X"A4",X"38",X"D7",X"26",X"C7",X"37",X"BE",X"62",X"5B",X"83",X"7A",X"94",X"49",X"C8",X"26",
		X"AD",X"34",X"8B",X"85",X"79",X"B4",X"49",X"C6",X"46",X"9C",X"76",X"59",X"86",X"59",X"B6",X"47",
		X"A8",X"55",X"9A",X"A6",X"57",X"87",X"68",X"78",X"57",X"99",X"74",X"68",X"B9",X"75",X"79",X"75",
		X"79",X"66",X"8A",X"96",X"36",X"AB",X"A7",X"57",X"77",X"67",X"98",X"77",X"A9",X"43",X"7B",X"BB",
		X"75",X"56",X"87",X"76",X"98",X"57",X"97",X"56",X"7B",X"B9",X"64",X"79",X"74",X"8C",X"74",X"6A",
		X"85",X"47",X"99",X"C7",X"64",X"78",X"56",X"8C",X"65",X"7A",X"74",X"78",X"99",X"B7",X"55",X"79",
		X"66",X"9B",X"65",X"7B",X"84",X"66",X"9A",X"A8",X"55",X"67",X"57",X"AB",X"64",X"7B",X"74",X"69",
		X"87",X"9B",X"74",X"57",X"75",X"9B",X"94",X"68",X"86",X"79",X"86",X"79",X"A7",X"76",X"66",X"7A",
		X"A6",X"68",X"96",X"67",X"85",X"58",X"CB",X"54",X"67",X"87",X"87",X"87",X"77",X"98",X"77",X"78",
		X"78",X"AB",X"53",X"68",X"86",X"98",X"65",X"89",X"87",X"76",X"67",X"98",X"89",X"76",X"58",X"A7",
		X"66",X"97",X"67",X"98",X"67",X"88",X"65",X"8A",X"B6",X"69",X"76",X"48",X"A8",X"77",X"89",X"76",
		X"68",X"87",X"69",X"B9",X"56",X"77",X"76",X"A7",X"78",X"88",X"67",X"88",X"65",X"89",X"86",X"99",
		X"66",X"67",X"87",X"97",X"78",X"88",X"67",X"97",X"56",X"88",X"78",X"78",X"95",X"69",X"78",X"59",
		X"97",X"78",X"87",X"79",X"65",X"78",X"86",X"78",X"A8",X"56",X"88",X"77",X"98",X"67",X"88",X"78",
		X"86",X"68",X"87",X"78",X"87",X"79",X"77",X"88",X"85",X"78",X"88",X"78",X"86",X"68",X"70",X"70",
		X"88",X"89",X"89",X"99",X"87",X"67",X"89",X"AA",X"98",X"76",X"67",X"9A",X"98",X"76",X"78",X"AB",
		X"97",X"67",X"AB",X"97",X"79",X"BA",X"64",X"8B",X"86",X"7B",X"A3",X"5C",X"B5",X"4D",X"93",X"8F",
		X"66",X"E8",X"1A",X"81",X"7B",X"3C",X"F6",X"DF",X"6B",X"E2",X"77",X"06",X"50",X"98",X"7F",X"8C",
		X"F6",X"E9",X"0C",X"03",X"90",X"BA",X"9F",X"7D",X"F3",X"E4",X"59",X"08",X"35",X"F6",X"DF",X"4F",
		X"46",X"81",X"B0",X"9C",X"5F",X"5F",X"A9",X"91",X"B0",X"B1",X"BA",X"9D",X"7E",X"3C",X"09",X"0C",
		X"3F",X"6F",X"5E",X"1B",X"0B",X"3E",X"6D",X"7A",X"64",X"91",X"B5",X"F5",X"F3",X"B2",X"65",X"5C",
		X"7F",X"5E",X"27",X"56",X"B7",X"F4",X"E4",X"85",X"3C",X"4F",X"5E",X"59",X"74",X"93",X"E6",X"E8",
		X"99",X"1A",X"2D",X"6C",X"B7",X"A1",X"94",X"9B",X"7E",X"5A",X"83",X"94",X"CB",X"9D",X"48",X"62",
		X"C8",X"BE",X"48",X"53",X"C6",X"9D",X"48",X"82",X"A5",X"7F",X"79",X"B1",X"4B",X"6B",X"E5",X"6B",
		X"44",X"E9",X"6C",X"A3",X"6B",X"79",X"C8",X"26",X"B8",X"9D",X"93",X"6B",X"75",X"DC",X"44",X"9A",
		X"4C",X"E7",X"47",X"A8",X"7C",X"94",X"59",X"C7",X"8B",X"94",X"4A",X"D9",X"79",X"77",X"8A",X"BA",
		X"64",X"4C",X"F5",X"37",X"B7",X"99",X"89",X"57",X"A7",X"98",X"6B",X"A6",X"47",X"B3",X"EF",X"82",
		X"B6",X"78",X"99",X"89",X"88",X"87",X"88",X"78",X"78",X"88",X"88",X"98",X"88",X"88",X"88",X"89",
		X"87",X"78",X"98",X"87",X"88",X"97",X"78",X"89",X"98",X"89",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70",
		X"78",X"87",X"77",X"78",X"87",X"77",X"78",X"97",X"67",X"77",X"88",X"66",X"88",X"88",X"76",X"78",
		X"98",X"66",X"78",X"99",X"76",X"68",X"88",X"76",X"68",X"98",X"76",X"68",X"99",X"76",X"78",X"89",
		X"76",X"78",X"87",X"76",X"8A",X"86",X"67",X"78",X"88",X"75",X"78",X"77",X"98",X"77",X"77",X"88",
		X"78",X"86",X"88",X"67",X"98",X"67",X"77",X"88",X"A8",X"68",X"96",X"7A",X"75",X"77",X"78",X"99",
		X"77",X"88",X"68",X"97",X"56",X"77",X"8A",X"96",X"68",X"77",X"9A",X"86",X"67",X"78",X"A7",X"37",
		X"96",X"7B",X"85",X"67",X"78",X"BA",X"54",X"88",X"79",X"A7",X"66",X"77",X"8C",X"84",X"7A",X"78",
		X"B7",X"34",X"76",X"7D",X"92",X"6B",X"77",X"B8",X"24",X"87",X"7E",X"B1",X"4B",X"86",X"B9",X"13",
		X"98",X"7E",X"C1",X"4C",X"96",X"A9",X"13",X"A8",X"7E",X"B2",X"4B",X"97",X"B9",X"13",X"97",X"9C",
		X"51",X"59",X"9A",X"C7",X"26",X"98",X"CB",X"22",X"87",X"7E",X"C1",X"1A",X"87",X"FB",X"02",X"C7",
		X"6E",X"B0",X"2A",X"7A",X"E5",X"05",X"A7",X"AE",X"50",X"7A",X"7E",X"C1",X"0A",X"A6",X"CC",X"11",
		X"99",X"CE",X"60",X"7A",X"8B",X"D4",X"06",X"98",X"D9",X"01",X"89",X"9C",X"91",X"4A",X"8D",X"D3",
		X"08",X"A8",X"BB",X"21",X"88",X"BE",X"71",X"7A",X"8B",X"C4",X"18",X"8A",X"E8",X"03",X"97",X"AD",
		X"60",X"7B",X"9C",X"90",X"07",X"99",X"D8",X"05",X"C9",X"AA",X"10",X"7B",X"8C",X"A1",X"3A",X"AB",
		X"91",X"06",X"B9",X"BA",X"23",X"9A",X"B8",X"10",X"7B",X"AB",X"A3",X"38",X"AC",X"91",X"18",X"BA",
		X"B9",X"23",X"7A",X"CA",X"10",X"8A",X"9C",X"A1",X"38",X"9C",X"B1",X"09",X"C8",X"CB",X"12",X"88",
		X"CC",X"10",X"9E",X"8B",X"B1",X"17",X"8D",X"C3",X"08",X"E9",X"BB",X"11",X"68",X"DD",X"30",X"8E",
		X"9B",X"B1",X"06",X"7D",X"F4",X"07",X"FA",X"AA",X"10",X"68",X"EF",X"60",X"6D",X"BB",X"92",X"06",
		X"7F",X"F5",X"07",X"CA",X"DB",X"00",X"77",X"DF",X"60",X"5C",X"AB",X"B2",X"07",X"AC",X"F7",X"02",
		X"9A",X"BB",X"40",X"6C",X"CD",X"71",X"06",X"BA",X"B7",X"04",X"BC",X"C9",X"00",X"5C",X"9A",X"B2",
		X"19",X"BC",X"D3",X"06",X"D9",X"9C",X"40",X"69",X"CE",X"81",X"4D",X"BA",X"C4",X"04",X"BB",X"C9",
		X"21",X"8C",X"AB",X"60",X"3C",X"BB",X"A3",X"05",X"C8",X"99",X"11",X"B9",X"BF",X"60",X"6E",X"88",
		X"D4",X"07",X"B9",X"D9",X"02",X"AA",X"7C",X"90",X"4D",X"8A",X"F4",X"08",X"C5",X"AD",X"20",X"B9",
		X"8F",X"90",X"4A",X"79",X"E7",X"05",X"B5",X"CF",X"40",X"8A",X"7A",X"E5",X"07",X"98",X"CA",X"20",
		X"59",X"9B",X"B3",X"17",X"7B",X"F8",X"13",X"68",X"AD",X"A0",X"29",X"6C",X"F8",X"04",X"A7",X"AF",
		X"90",X"3A",X"6D",X"F6",X"04",X"B8",X"AF",X"60",X"48",X"8F",X"E4",X"04",X"BA",X"CE",X"40",X"38",
		X"BE",X"C5",X"04",X"DB",X"AC",X"50",X"2B",X"CB",X"C5",X"05",X"EA",X"8D",X"60",X"2D",X"AA",X"E7",
		X"06",X"EA",X"8D",X"71",X"2C",X"8B",X"E7",X"05",X"B9",X"AC",X"71",X"2A",X"8A",X"D8",X"00",X"6A",
		X"BA",X"93",X"27",X"BC",X"CA",X"30",X"3A",X"B9",X"A9",X"11",X"9B",X"AC",X"91",X"2B",X"EA",X"9A",
		X"20",X"8C",X"8A",X"A1",X"06",X"D9",X"6C",X"90",X"4C",X"89",X"C7",X"13",X"9A",X"78",X"C7",X"06",
		X"B8",X"AF",X"A2",X"4C",X"75",X"CD",X"20",X"79",X"7C",X"F8",X"15",X"A7",X"7D",X"B1",X"07",X"97",
		X"CD",X"61",X"5A",X"77",X"EB",X"11",X"77",X"7B",X"D7",X"27",X"95",X"7E",X"D3",X"05",X"86",X"BF",
		X"B5",X"47",X"79",X"DD",X"40",X"38",X"7B",X"FA",X"21",X"57",X"7A",X"E7",X"04",X"B8",X"8C",X"A2",
		X"04",X"87",X"8D",X"B2",X"29",X"74",X"AD",X"61",X"7A",X"47",X"FB",X"22",X"86",X"5C",X"F8",X"48",
		X"75",X"9C",X"B7",X"46",X"96",X"8D",X"93",X"37",X"54",X"AE",X"84",X"78",X"35",X"DB",X"56",X"94",
		X"4C",X"D7",X"68",X"54",X"7D",X"D6",X"78",X"35",X"BC",X"97",X"64",X"66",X"AA",X"76",X"55",X"56",
		X"99",X"78",X"86",X"46",X"BA",X"68",X"82",X"6B",X"A8",X"76",X"55",X"8A",X"97",X"88",X"44",X"AB",
		X"67",X"96",X"66",X"A9",X"77",X"85",X"59",X"97",X"89",X"85",X"68",X"97",X"79",X"73",X"8B",X"66",
		X"98",X"57",X"89",X"67",X"B6",X"4A",X"96",X"89",X"87",X"77",X"87",X"78",X"87",X"78",X"78",X"77",
		X"97",X"69",X"85",X"79",X"66",X"98",X"66",X"99",X"68",X"96",X"69",X"98",X"87",X"87",X"6A",X"96",
		X"78",X"76",X"8A",X"85",X"79",X"56",X"B9",X"56",X"97",X"78",X"97",X"58",X"96",X"89",X"76",X"79",
		X"87",X"78",X"76",X"88",X"77",X"78",X"77",X"98",X"76",X"88",X"78",X"76",X"77",X"88",X"78",X"87",
		X"68",X"A7",X"77",X"77",X"78",X"86",X"78",X"86",X"8A",X"66",X"86",X"78",X"98",X"77",X"78",X"88",
		X"97",X"67",X"77",X"78",X"97",X"68",X"78",X"98",X"86",X"77",X"68",X"98",X"76",X"87",X"7A",X"77",
		X"76",X"67",X"98",X"77",X"86",X"88",X"79",X"76",X"87",X"78",X"88",X"78",X"86",X"88",X"68",X"87",
		X"77",X"77",X"89",X"77",X"86",X"78",X"78",X"87",X"67",X"89",X"78",X"95",X"78",X"68",X"88",X"76",
		X"79",X"69",X"96",X"68",X"67",X"78",X"77",X"78",X"69",X"97",X"88",X"57",X"77",X"87",X"79",X"69",
		X"97",X"78",X"67",X"68",X"86",X"98",X"79",X"78",X"75",X"98",X"58",X"76",X"A6",X"9A",X"28",X"76",
		X"A7",X"77",X"49",X"99",X"95",X"68",X"5C",X"95",X"75",X"8B",X"98",X"45",X"87",X"C8",X"46",X"5A",
		X"B8",X"81",X"59",X"7C",X"84",X"65",X"E8",X"68",X"05",X"A8",X"A4",X"46",X"8F",X"A7",X"62",X"9B",
		X"C9",X"23",X"5A",X"D7",X"72",X"4B",X"9A",X"93",X"58",X"FB",X"56",X"25",X"CC",X"73",X"25",X"CB",
		X"65",X"15",X"BA",X"97",X"34",X"CF",X"B9",X"65",X"8C",X"D6",X"33",X"4F",X"94",X"60",X"6B",X"A7",
		X"32",X"4E",X"A4",X"71",X"4B",X"87",X"53",X"4D",X"C5",X"83",X"5C",X"AA",X"82",X"5C",X"D9",X"85",
		X"5A",X"CA",X"84",X"3B",X"FA",X"85",X"79",X"AD",X"64",X"47",X"FA",X"58",X"48",X"BC",X"73",X"45",
		X"FA",X"39",X"46",X"DA",X"65",X"35",X"F9",X"29",X"25",X"D9",X"64",X"24",X"F9",X"19",X"15",X"E7",
		X"67",X"15",X"F7",X"1A",X"06",X"F7",X"57",X"14",X"F8",X"19",X"05",X"F6",X"58",X"14",X"F8",X"19",
		X"05",X"F7",X"68",X"25",X"F9",X"18",X"15",X"F7",X"58",X"25",X"FA",X"08",X"14",X"F9",X"57",X"35",
		X"FB",X"16",X"24",X"DB",X"56",X"34",X"FC",X"25",X"23",X"BD",X"65",X"53",X"FF",X"24",X"44",X"AE",
		X"74",X"63",X"DF",X"33",X"53",X"AE",X"84",X"63",X"BF",X"43",X"73",X"8F",X"94",X"63",X"AF",X"51",
		X"83",X"7F",X"94",X"63",X"AF",X"61",X"75",X"7F",X"A3",X"63",X"8F",X"81",X"75",X"6F",X"A3",X"54",
		X"8F",X"91",X"76",X"5F",X"C2",X"63",X"6F",X"A0",X"86",X"5F",X"D2",X"54",X"6F",X"B0",X"77",X"5F",
		X"E2",X"55",X"4F",X"C0",X"78",X"5E",X"F3",X"45",X"3F",X"D0",X"78",X"4E",X"F3",X"35",X"3F",X"F0",
		X"68",X"3D",X"F3",X"25",X"1F",X"F1",X"57",X"3C",X"F4",X"15",X"1E",X"F2",X"25",X"39",X"F6",X"15",
		X"1C",X"F5",X"14",X"56",X"F9",X"15",X"39",X"F9",X"15",X"85",X"ED",X"23",X"56",X"FF",X"14",X"B4",
		X"CF",X"31",X"63",X"FF",X"21",X"93",X"9F",X"50",X"62",X"8F",X"71",X"55",X"4F",X"B0",X"55",X"5F",
		X"E0",X"5A",X"3D",X"F3",X"28",X"3E",X"F1",X"3A",X"39",X"F6",X"07",X"37",X"F6",X"06",X"53",X"FC",
		X"05",X"53",X"FE",X"05",X"B2",X"CF",X"43",X"82",X"DF",X"33",X"93",X"6F",X"81",X"73",X"6F",X"81",
		X"58",X"2F",X"E1",X"47",X"3F",X"F1",X"4D",X"19",X"F5",X"29",X"29",X"F5",X"18",X"33",X"FA",X"06",
		X"53",X"FC",X"05",X"90",X"DF",X"13",X"91",X"EF",X"23",X"B1",X"6F",X"71",X"84",X"4F",X"A0",X"67",
		X"1F",X"F1",X"48",X"2F",X"F1",X"4C",X"0A",X"F4",X"19",X"26",X"F7",X"06",X"43",X"FD",X"16",X"72",
		X"FF",X"15",X"B1",X"BF",X"42",X"91",X"7F",X"60",X"53",X"4F",X"C1",X"56",X"3F",X"F1",X"6A",X"1A",
		X"F5",X"29",X"27",X"F7",X"04",X"44",X"FD",X"15",X"53",X"FF",X"15",X"A1",X"BF",X"50",X"72",X"6F",
		X"A0",X"34",X"5F",X"E3",X"47",X"3F",X"F3",X"38",X"2B",X"F6",X"06",X"35",X"FD",X"03",X"75",X"FF",
		X"41",X"75",X"EF",X"51",X"33",X"9F",X"90",X"35",X"4F",X"F0",X"2A",X"6B",X"F6",X"07",X"76",X"FC",
		X"01",X"86",X"BF",X"40",X"86",X"CF",X"50",X"56",X"7F",X"A0",X"48",X"4F",X"F1",X"1B",X"68",X"F7",
		X"06",X"74",X"FF",X"02",X"B6",X"9F",X"60",X"77",X"7E",X"90",X"28",X"7B",X"E5",X"18",X"7A",X"F5",
		X"06",X"66",X"EC",X"02",X"A4",X"CF",X"50",X"B8",X"6F",X"B0",X"3A",X"3D",X"F3",X"0C",X"76",X"F9",
		X"07",X"A4",X"FD",X"01",X"A5",X"8F",X"60",X"96",X"6F",X"81",X"58",X"5D",X"E1",X"1B",X"49",X"F5",
		X"08",X"64",X"FC",X"03",X"B3",X"CF",X"40",X"A7",X"5F",X"B0",X"3A",X"2D",X"F4",X"0A",X"86",X"FB",
		X"03",X"A3",X"EF",X"31",X"B9",X"7F",X"B0",X"59",X"3E",X"F1",X"1B",X"89",X"F8",X"07",X"85",X"FD",
		X"03",X"96",X"BF",X"60",X"97",X"7F",X"B0",X"38",X"6B",X"F5",X"18",X"78",X"FA",X"02",X"87",X"AE",
		X"50",X"88",X"8E",X"A0",X"18",X"89",X"D6",X"08",X"89",X"EA",X"02",X"98",X"AE",X"40",X"87",X"7F",
		X"B0",X"2B",X"7A",X"F5",X"08",X"77",X"FB",X"03",X"A7",X"AF",X"50",X"78",X"7F",X"B0",X"2A",X"7A",
		X"E7",X"06",X"98",X"FC",X"12",X"A9",X"8D",X"81",X"39",X"7D",X"D2",X"1B",X"B7",X"C8",X"03",X"A7",
		X"BD",X"10",X"9A",X"8C",X"90",X"4A",X"7A",X"D4",X"06",X"97",X"AA",X"23",X"A8",X"8D",X"71",X"4A",
		X"89",X"C5",X"29",X"97",X"EC",X"13",X"B8",X"7D",X"81",X"69",X"6D",X"E2",X"2B",X"85",X"DA",X"15",
		X"96",X"BE",X"30",X"89",X"6C",X"B1",X"39",X"89",X"D8",X"03",X"A8",X"9D",X"61",X"6A",X"7D",X"E2",
		X"0B",X"A5",X"DB",X"03",X"B6",X"AF",X"40",X"9B",X"4B",X"D1",X"1B",X"87",X"F8",X"04",X"C6",X"7E",
		X"50",X"9D",X"5D",X"F1",X"0E",X"93",X"DA",X"04",X"E5",X"9F",X"30",X"BB",X"3C",X"D0",X"1D",X"75",
		X"E7",X"05",X"C6",X"8E",X"50",X"9B",X"4B",X"E2",X"1C",X"95",X"CB",X"03",X"C6",X"7E",X"60",X"7A",
		X"69",X"D5",X"1A",X"B5",X"CE",X"21",X"B9",X"5C",X"C0",X"3C",X"65",X"E8",X"05",X"B5",X"7F",X"60",
		X"AA",X"4C",X"F3",X"1C",X"84",X"DD",X"12",X"C6",X"5F",X"A0",X"4B",X"67",X"F8",X"08",X"B3",X"BF",
		X"40",X"A9",X"4D",X"D0",X"1B",X"55",X"FB",X"03",X"A5",X"8F",X"81",X"7A",X"3C",X"F4",X"09",X"84",
		X"CE",X"21",X"A6",X"5F",X"D1",X"29",X"78",X"EB",X"14",X"94",X"9F",X"60",X"49",X"7A",X"E7",X"06",
		X"95",X"DF",X"50",X"79",X"6B",X"D3",X"08",X"86",X"EE",X"20",X"AA",X"6D",X"D1",X"1A",X"66",X"EA",
		X"02",X"B8",X"6E",X"B0",X"3C",X"68",X"F7",X"04",X"A7",X"8E",X"81",X"59",X"6A",X"E6",X"06",X"96",
		X"9D",X"61",X"79",X"6B",X"E5",X"17",X"96",X"AE",X"50",X"79",X"5C",X"F4",X"19",X"95",X"CE",X"31",
		X"98",X"5D",X"E3",X"09",X"96",X"DE",X"21",X"97",X"5E",X"D1",X"0A",X"95",X"ED",X"11",X"B7",X"5F",
		X"C0",X"1B",X"86",X"EC",X"02",X"B7",X"7F",X"90",X"2B",X"76",X"FA",X"03",X"C6",X"8F",X"81",X"3B",
		X"67",X"F8",X"05",X"B5",X"AF",X"50",X"5A",X"5A",X"F5",X"07",X"A5",X"CF",X"30",X"79",X"5C",X"E3",
		X"08",X"95",X"DE",X"20",X"88",X"6C",X"C3",X"08",X"97",X"DD",X"30",X"79",X"6B",X"C4",X"17",X"96",
		X"CD",X"40",X"79",X"7A",X"D6",X"16",X"A7",X"BE",X"50",X"69",X"6A",X"E5",X"07",X"95",X"CF",X"50",
		X"67",X"7C",X"D5",X"17",X"76",X"CE",X"51",X"57",X"8C",X"D6",X"26",X"76",X"CD",X"72",X"47",X"9B",
		X"B8",X"34",X"77",X"9C",X"A3",X"39",X"98",X"BA",X"33",X"87",X"8D",X"B2",X"49",X"88",X"B9",X"33",
		X"88",X"8C",X"B3",X"48",X"88",X"A9",X"43",X"78",X"8B",X"B5",X"36",X"99",X"99",X"62",X"69",X"8B",
		X"B5",X"26",X"A9",X"99",X"62",X"69",X"9A",X"A6",X"14",X"AA",X"8A",X"72",X"5A",X"A9",X"B7",X"13",
		X"AB",X"8A",X"93",X"39",X"A9",X"BB",X"21",X"9A",X"8A",X"A4",X"27",X"98",X"BB",X"42",X"6A",X"99",
		X"96",X"24",X"AA",X"99",X"51",X"4A",X"C9",X"88",X"43",X"9C",X"99",X"83",X"18",X"D8",X"7A",X"61",
		X"7C",X"99",X"B6",X"26",X"C9",X"68",X"83",X"4A",X"A7",X"89",X"33",X"AC",X"66",X"A6",X"28",X"C8",
		X"8C",X"61",X"7C",X"76",X"A9",X"23",X"BA",X"79",X"92",X"29",X"C7",X"7B",X"61",X"7C",X"88",X"C7",
		X"17",X"C7",X"6B",X"92",X"4B",X"97",X"A8",X"13",X"AC",X"78",X"A5",X"17",X"C8",X"9C",X"72",X"7C",
		X"85",X"A9",X"34",X"B9",X"69",X"93",X"3A",X"C5",X"6C",X"71",X"8C",X"68",X"D8",X"26",X"B6",X"5B",
		X"A3",X"4A",X"86",X"BB",X"52",X"99",X"68",X"C8",X"35",X"97",X"8A",X"83",X"47",X"88",X"70",X"70",
		X"88",X"89",X"88",X"88",X"88",X"88",X"89",X"A8",X"54",X"8C",X"EC",X"63",X"36",X"9B",X"CC",X"B9",
		X"53",X"37",X"CE",X"C7",X"44",X"8B",X"CA",X"75",X"48",X"CB",X"53",X"2B",X"EF",X"E8",X"31",X"12",
		X"8E",X"FF",X"C4",X"00",X"7D",X"FF",X"63",X"35",X"78",X"AE",X"EE",X"93",X"10",X"5C",X"EE",X"C7",
		X"43",X"33",X"8E",X"FF",X"E6",X"10",X"06",X"CF",X"FD",X"63",X"22",X"5C",X"FF",X"F8",X"40",X"06",
		X"CF",X"FB",X"62",X"23",X"7C",X"FF",X"D6",X"20",X"29",X"DF",X"E9",X"43",X"34",X"9D",X"FE",X"B4",
		X"11",X"4A",X"CE",X"C7",X"33",X"49",X"CD",X"D9",X"43",X"36",X"BD",X"DB",X"64",X"35",X"AC",X"DB",
		X"74",X"46",X"9B",X"B9",X"76",X"67",X"9A",X"AA",X"86",X"66",X"8A",X"BA",X"86",X"57",X"9B",X"B9",
		X"76",X"67",X"89",X"BA",X"97",X"55",X"79",X"BB",X"96",X"67",X"89",X"99",X"99",X"87",X"77",X"89",
		X"99",X"77",X"78",X"88",X"89",X"99",X"97",X"76",X"79",X"9A",X"98",X"77",X"77",X"89",X"99",X"98",
		X"77",X"78",X"99",X"99",X"87",X"77",X"89",X"A9",X"97",X"77",X"89",X"99",X"98",X"77",X"78",X"99",
		X"98",X"77",X"78",X"89",X"88",X"88",X"88",X"88",X"99",X"87",X"77",X"89",X"99",X"98",X"77",X"78",
		X"99",X"99",X"87",X"77",X"89",X"99",X"87",X"78",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"77",
		X"88",X"88",X"88",X"88",X"87",X"88",X"99",X"87",X"77",X"88",X"99",X"88",X"88",X"87",X"88",X"99",
		X"88",X"88",X"98",X"88",X"88",X"98",X"87",X"88",X"99",X"88",X"78",X"88",X"88",X"88",X"88",X"78",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
