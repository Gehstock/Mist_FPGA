library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpa_13m is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpa_13m is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"00",X"E8",X"ED",X"56",X"3A",X"04",X"D0",X"A7",X"F2",X"00",X"33",X"CD",X"F4",X"05",
		X"CD",X"F2",X"06",X"CD",X"29",X"0D",X"C3",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",
		X"EB",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"D9",X"CD",X"6D",X"05",X"21",X"4E",X"E0",
		X"34",X"7E",X"23",X"E6",X"0F",X"20",X"01",X"34",X"23",X"35",X"23",X"35",X"3A",X"04",X"D0",X"A7",
		X"FA",X"93",X"00",X"21",X"4E",X"E0",X"34",X"01",X"03",X"00",X"21",X"4E",X"E0",X"35",X"10",X"FE",
		X"0D",X"20",X"FB",X"D9",X"08",X"FB",X"FB",X"C9",X"FB",X"CD",X"8A",X"0B",X"3E",X"01",X"32",X"4D",
		X"E0",X"32",X"0F",X"E5",X"3C",X"32",X"08",X"E5",X"C3",X"B7",X"0B",X"06",X"00",X"AF",X"32",X"4D",
		X"E0",X"21",X"46",X"E0",X"70",X"FB",X"CD",X"45",X"07",X"CD",X"8A",X"0B",X"C3",X"B7",X"0B",X"06",
		X"04",X"18",X"EA",X"CD",X"CB",X"05",X"3A",X"00",X"D0",X"2F",X"32",X"53",X"E0",X"CB",X"4F",X"28",
		X"15",X"3A",X"04",X"D0",X"CB",X"67",X"20",X"0E",X"21",X"46",X"E0",X"CB",X"4E",X"20",X"07",X"3A",
		X"00",X"D0",X"E6",X"01",X"20",X"F9",X"3A",X"04",X"D0",X"CB",X"5F",X"20",X"06",X"21",X"F3",X"E0",
		X"34",X"CB",X"46",X"FD",X"E5",X"DD",X"E5",X"CD",X"0E",X"04",X"3A",X"41",X"E0",X"A7",X"20",X"05",
		X"3E",X"02",X"32",X"48",X"E0",X"21",X"46",X"E0",X"46",X"CB",X"78",X"20",X"15",X"CB",X"48",X"20",
		X"1B",X"3A",X"48",X"E0",X"A7",X"20",X"1D",X"CB",X"50",X"20",X"11",X"3A",X"47",X"E0",X"A7",X"C2",
		X"8F",X"00",X"CB",X"40",X"28",X"06",X"CD",X"7A",X"04",X"CD",X"EC",X"01",X"DD",X"E1",X"FD",X"E1",
		X"D9",X"08",X"FB",X"C9",X"36",X"02",X"31",X"00",X"E8",X"FB",X"CD",X"29",X"0D",X"CD",X"33",X"05",
		X"28",X"FB",X"CD",X"38",X"0B",X"C3",X"B7",X"0B",X"31",X"00",X"E8",X"21",X"46",X"E0",X"35",X"FB",
		X"F2",X"68",X"00",X"CD",X"96",X"0B",X"AF",X"32",X"A6",X"E1",X"21",X"15",X"E5",X"35",X"28",X"1B",
		X"CD",X"D5",X"06",X"21",X"46",X"E0",X"CB",X"66",X"CA",X"B7",X"0B",X"CD",X"03",X"06",X"3A",X"15",
		X"E5",X"A7",X"C2",X"B7",X"0B",X"CD",X"03",X"06",X"C3",X"B7",X"0B",X"3E",X"1B",X"CD",X"75",X"0D",
		X"21",X"46",X"E0",X"CB",X"66",X"28",X"1F",X"21",X"ED",X"2A",X"CD",X"4E",X"03",X"3A",X"46",X"E0",
		X"1F",X"1F",X"1F",X"E6",X"01",X"3C",X"CD",X"BD",X"03",X"CD",X"03",X"06",X"CD",X"E4",X"05",X"3A",
		X"15",X"E5",X"A7",X"C2",X"B7",X"0B",X"21",X"02",X"2B",X"CD",X"4E",X"03",X"CD",X"1C",X"06",X"28",
		X"03",X"CD",X"03",X"06",X"CD",X"E8",X"05",X"CD",X"29",X"0D",X"21",X"2A",X"2A",X"CD",X"00",X"03",
		X"3E",X"11",X"A7",X"28",X"3D",X"3D",X"27",X"32",X"54",X"E0",X"11",X"33",X"82",X"0E",X"02",X"CD",
		X"AE",X"03",X"3E",X"40",X"32",X"50",X"E0",X"3A",X"50",X"E0",X"A7",X"3A",X"54",X"E0",X"28",X"E2",
		X"3A",X"48",X"E0",X"A7",X"20",X"0B",X"21",X"57",X"2C",X"CD",X"74",X"03",X"CD",X"27",X"05",X"18",
		X"E6",X"CD",X"33",X"05",X"28",X"E1",X"CD",X"DA",X"01",X"CD",X"DA",X"01",X"CD",X"BF",X"0C",X"C3",
		X"B7",X"0B",X"F3",X"AF",X"32",X"46",X"E0",X"C3",X"68",X"00",X"3A",X"40",X"E0",X"32",X"15",X"E5",
		X"21",X"00",X"00",X"22",X"00",X"E5",X"22",X"02",X"E5",X"C3",X"03",X"06",X"DD",X"21",X"00",X"E3",
		X"3E",X"20",X"32",X"E8",X"E0",X"DD",X"7E",X"00",X"3D",X"FA",X"00",X"02",X"21",X"0C",X"02",X"EF",
		X"11",X"10",X"00",X"DD",X"19",X"21",X"E8",X"E0",X"35",X"20",X"EA",X"C9",X"11",X"13",X"31",X"13",
		X"70",X"13",X"88",X"13",X"BC",X"13",X"C2",X"13",X"EB",X"13",X"21",X"14",X"09",X"18",X"E0",X"15",
		X"FA",X"15",X"2D",X"16",X"2D",X"16",X"49",X"16",X"5D",X"16",X"8F",X"16",X"3D",X"19",X"57",X"19",
		X"5E",X"19",X"D1",X"19",X"2F",X"1A",X"44",X"1A",X"92",X"1A",X"B9",X"1A",X"F0",X"1A",X"01",X"1B",
		X"27",X"1B",X"33",X"14",X"E0",X"18",X"AA",X"1E",X"28",X"1F",X"AC",X"20",X"C4",X"20",X"AA",X"1E",
		X"28",X"1F",X"00",X"20",X"1A",X"20",X"A4",X"1E",X"28",X"1F",X"4D",X"20",X"9C",X"20",X"23",X"1D",
		X"F3",X"1D",X"51",X"1E",X"9B",X"1E",X"9B",X"1C",X"BC",X"1C",X"14",X"1E",X"29",X"1E",X"CD",X"DC",
		X"0D",X"CD",X"0D",X"21",X"CD",X"3A",X"1B",X"CD",X"C7",X"1B",X"CD",X"A7",X"12",X"CD",X"E7",X"12",
		X"CD",X"DC",X"0D",X"3A",X"CF",X"E1",X"21",X"D0",X"E1",X"BE",X"28",X"E2",X"5F",X"16",X"E6",X"DD",
		X"21",X"00",X"00",X"DD",X"19",X"DD",X"4E",X"00",X"CB",X"21",X"20",X"11",X"21",X"CF",X"E1",X"BE",
		X"20",X"03",X"C6",X"04",X"77",X"DD",X"E5",X"C1",X"79",X"C6",X"04",X"18",X"D9",X"06",X"00",X"DD",
		X"70",X"00",X"DD",X"7E",X"01",X"21",X"A5",X"02",X"E5",X"21",X"D3",X"02",X"09",X"4E",X"23",X"66",
		X"69",X"E9",X"21",X"D0",X"E1",X"6E",X"26",X"E6",X"71",X"23",X"77",X"23",X"73",X"23",X"72",X"2C",
		X"7D",X"32",X"D0",X"E1",X"C9",X"22",X"06",X"FA",X"02",X"ED",X"02",X"22",X"03",X"2F",X"03",X"67",
		X"03",X"61",X"03",X"37",X"03",X"A6",X"0D",X"01",X"12",X"18",X"12",X"00",X"00",X"3A",X"4E",X"E0",
		X"DD",X"86",X"01",X"DD",X"77",X"01",X"DD",X"36",X"00",X"04",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"CD",X"DB",X"03",X"7E",X"06",X"12",X"FE",X"26",X"28",X"06",X"06",X"30",X"FE",X"27",X"20",X"0D",
		X"23",X"78",X"32",X"50",X"E0",X"3A",X"50",X"E0",X"A7",X"20",X"FA",X"18",X"E6",X"CD",X"C9",X"03",
		X"18",X"E1",X"3A",X"4E",X"E0",X"DD",X"BE",X"01",X"28",X"05",X"DD",X"36",X"00",X"04",X"C9",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"18",X"44",X"3A",X"50",X"E0",X"A7",X"20",X"0C",X"CD",X"2F",X"03",
		X"DD",X"35",X"01",X"C8",X"3E",X"04",X"32",X"50",X"E0",X"DD",X"36",X"00",X"07",X"C9",X"CD",X"DB",
		X"03",X"CD",X"C9",X"03",X"3E",X"03",X"32",X"50",X"E0",X"3A",X"50",X"E0",X"A7",X"20",X"FA",X"18",
		X"F0",X"3A",X"50",X"E0",X"A7",X"20",X"08",X"3E",X"04",X"32",X"50",X"E0",X"CD",X"FA",X"02",X"DD",
		X"36",X"00",X"08",X"C9",X"3A",X"4E",X"E0",X"CB",X"67",X"20",X"85",X"CD",X"DB",X"03",X"7E",X"23",
		X"FE",X"21",X"C8",X"FE",X"23",X"28",X"09",X"FE",X"22",X"28",X"F0",X"AF",X"12",X"13",X"18",X"EE",
		X"23",X"18",X"EB",X"7E",X"13",X"E6",X"0F",X"28",X"04",X"1B",X"CD",X"A6",X"03",X"2B",X"7E",X"1F",
		X"1F",X"1F",X"1F",X"CD",X"A7",X"03",X"7E",X"E6",X"0F",X"C6",X"30",X"12",X"13",X"C9",X"FD",X"21",
		X"00",X"04",X"FD",X"19",X"F5",X"1F",X"1F",X"1F",X"1F",X"CD",X"BD",X"03",X"F1",X"E6",X"0F",X"C6",
		X"30",X"12",X"FD",X"71",X"00",X"13",X"FD",X"23",X"C9",X"7E",X"23",X"FE",X"21",X"28",X"33",X"FE",
		X"23",X"28",X"12",X"FE",X"25",X"28",X"2D",X"FE",X"22",X"20",X"E6",X"5E",X"23",X"56",X"23",X"FD",
		X"21",X"00",X"04",X"FD",X"19",X"4E",X"23",X"3A",X"F9",X"E0",X"A7",X"C8",X"79",X"A7",X"C8",X"FE",
		X"03",X"38",X"0B",X"FE",X"06",X"28",X"03",X"FE",X"09",X"C0",X"C6",X"05",X"4F",X"C9",X"C6",X"0B",
		X"4F",X"C9",X"E1",X"C9",X"46",X"23",X"7E",X"23",X"CD",X"C1",X"03",X"10",X"FB",X"C9",X"21",X"3E",
		X"E0",X"11",X"41",X"E0",X"3A",X"00",X"D0",X"01",X"02",X"00",X"CD",X"34",X"04",X"21",X"3F",X"E0",
		X"13",X"3A",X"02",X"D0",X"1F",X"F6",X"04",X"0E",X"20",X"CD",X"34",X"04",X"3A",X"4C",X"E0",X"B0",
		X"32",X"01",X"D0",X"C9",X"1F",X"1F",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"E6",X"55",X"FE",
		X"54",X"28",X"0E",X"7E",X"E6",X"AA",X"C0",X"21",X"ED",X"E0",X"34",X"7E",X"E6",X"0F",X"C0",X"18",
		X"19",X"78",X"B1",X"47",X"3E",X"13",X"CD",X"7D",X"0D",X"1A",X"FE",X"01",X"28",X"11",X"FE",X"08",
		X"30",X"0B",X"21",X"47",X"E0",X"34",X"BE",X"C0",X"AF",X"77",X"3C",X"18",X"02",X"D6",X"08",X"21",
		X"48",X"E0",X"86",X"27",X"30",X"02",X"3E",X"99",X"77",X"C9",X"3A",X"46",X"E0",X"07",X"30",X"5B",
		X"11",X"01",X"D0",X"CB",X"67",X"28",X"07",X"3A",X"43",X"E0",X"3D",X"28",X"01",X"13",X"21",X"4A",
		X"E0",X"7E",X"23",X"77",X"2B",X"1A",X"2F",X"77",X"2B",X"E6",X"03",X"77",X"C9",X"3A",X"0B",X"E5",
		X"2A",X"F7",X"E0",X"BE",X"20",X"13",X"23",X"7E",X"54",X"5D",X"23",X"22",X"F7",X"E0",X"A7",X"28",
		X"04",X"FE",X"FF",X"20",X"D9",X"32",X"E0",X"E1",X"C9",X"21",X"4A",X"E0",X"3A",X"E0",X"E1",X"A7",
		X"28",X"13",X"3A",X"4E",X"E0",X"07",X"47",X"E6",X"01",X"3C",X"32",X"49",X"E0",X"78",X"E6",X"1E",
		X"20",X"03",X"36",X"20",X"C9",X"7E",X"36",X"FF",X"23",X"77",X"C9",X"21",X"4D",X"E0",X"3A",X"4E",
		X"E0",X"47",X"7E",X"A7",X"28",X"B7",X"FE",X"50",X"28",X"1D",X"CB",X"18",X"38",X"05",X"CB",X"18",
		X"38",X"01",X"34",X"0E",X"02",X"21",X"49",X"E0",X"FE",X"18",X"38",X"01",X"0D",X"71",X"23",X"36",
		X"00",X"FE",X"B0",X"D8",X"C3",X"7B",X"00",X"21",X"00",X"E3",X"7E",X"FE",X"04",X"20",X"0C",X"3A",
		X"09",X"E3",X"17",X"D8",X"36",X"08",X"0E",X"0A",X"C3",X"C2",X"02",X"FE",X"08",X"C8",X"21",X"4A",
		X"E0",X"36",X"20",X"23",X"36",X"00",X"C9",X"21",X"E2",X"2A",X"CD",X"00",X"03",X"3A",X"48",X"E0",
		X"C3",X"AE",X"03",X"21",X"D1",X"2A",X"CD",X"74",X"03",X"CD",X"27",X"05",X"21",X"86",X"2A",X"3A",
		X"48",X"E0",X"3D",X"28",X"03",X"21",X"97",X"2A",X"CD",X"00",X"03",X"3A",X"53",X"E0",X"E6",X"03",
		X"C8",X"1F",X"3A",X"48",X"E0",X"06",X"80",X"38",X"06",X"D6",X"01",X"27",X"C8",X"06",X"90",X"D6",
		X"01",X"27",X"F3",X"32",X"48",X"E0",X"78",X"32",X"46",X"E0",X"3C",X"FB",X"C9",X"21",X"00",X"E1",
		X"11",X"40",X"C8",X"01",X"40",X"00",X"ED",X"B0",X"1E",X"20",X"0E",X"20",X"ED",X"B0",X"1E",X"C0",
		X"0E",X"40",X"ED",X"B0",X"11",X"A0",X"C8",X"0E",X"20",X"ED",X"B0",X"0E",X"1C",X"7E",X"06",X"04",
		X"ED",X"79",X"0C",X"10",X"FB",X"23",X"3A",X"C3",X"E1",X"A7",X"28",X"2B",X"7E",X"E6",X"7F",X"01",
		X"40",X"00",X"CB",X"3F",X"30",X"01",X"04",X"20",X"F9",X"7E",X"07",X"E6",X"01",X"A8",X"5F",X"ED",
		X"A3",X"3A",X"00",X"88",X"E6",X"07",X"BB",X"C2",X"C3",X"00",X"0E",X"80",X"ED",X"A3",X"0E",X"60",
		X"ED",X"A3",X"0E",X"A0",X"ED",X"A3",X"7E",X"2F",X"D3",X"C0",X"C9",X"2A",X"DD",X"E1",X"7D",X"BC",
		X"C8",X"26",X"E0",X"7E",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"7D",X"3C",X"E6",X"07",
		X"32",X"DD",X"E1",X"C9",X"3E",X"40",X"18",X"02",X"3E",X"C0",X"32",X"50",X"E0",X"3A",X"50",X"E0",
		X"A7",X"20",X"FA",X"C9",X"21",X"00",X"E0",X"01",X"00",X"07",X"36",X"00",X"23",X"0B",X"78",X"B1",
		X"20",X"F8",X"C9",X"21",X"46",X"E0",X"7E",X"EE",X"08",X"77",X"21",X"00",X"E5",X"11",X"18",X"E5",
		X"06",X"18",X"1A",X"4F",X"7E",X"12",X"71",X"23",X"13",X"10",X"F7",X"C9",X"3A",X"46",X"E0",X"CB",
		X"5F",X"C9",X"4F",X"81",X"81",X"4F",X"06",X"00",X"21",X"0C",X"2A",X"09",X"3A",X"46",X"E0",X"A7",
		X"F0",X"11",X"00",X"E5",X"06",X"03",X"A7",X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"CD",
		X"AF",X"06",X"06",X"03",X"11",X"00",X"E5",X"21",X"08",X"E0",X"A7",X"1A",X"9E",X"23",X"13",X"10",
		X"FA",X"38",X"15",X"2A",X"00",X"E5",X"22",X"08",X"E0",X"3A",X"02",X"E5",X"32",X"0A",X"E0",X"3A",
		X"0E",X"E5",X"32",X"0B",X"E0",X"CD",X"85",X"06",X"11",X"84",X"80",X"CD",X"1C",X"06",X"28",X"03",
		X"11",X"A4",X"80",X"21",X"02",X"E5",X"0E",X"01",X"CD",X"E7",X"03",X"06",X"03",X"7E",X"CD",X"AE",
		X"03",X"2B",X"10",X"F9",X"C9",X"21",X"0B",X"E0",X"7E",X"0E",X"09",X"FE",X"1B",X"38",X"04",X"D6",
		X"1A",X"0E",X"06",X"C6",X"40",X"32",X"4A",X"80",X"3A",X"F9",X"E0",X"1F",X"79",X"30",X"02",X"C6",
		X"05",X"32",X"4A",X"84",X"11",X"43",X"80",X"0E",X"09",X"CD",X"E7",X"03",X"2B",X"18",X"CC",X"2A",
		X"01",X"E5",X"3A",X"45",X"E0",X"3D",X"F8",X"3D",X"28",X"01",X"24",X"CB",X"2C",X"25",X"3C",X"7C",
		X"20",X"05",X"A7",X"28",X"02",X"3E",X"FE",X"21",X"03",X"E5",X"BE",X"C0",X"7E",X"FE",X"03",X"C8",
		X"34",X"21",X"15",X"E5",X"34",X"3A",X"15",X"E5",X"3D",X"28",X"03",X"4F",X"3E",X"01",X"21",X"7C",
		X"80",X"CD",X"EC",X"06",X"CD",X"EC",X"06",X"28",X"03",X"79",X"C6",X"30",X"77",X"23",X"A7",X"C8",
		X"3C",X"C9",X"21",X"40",X"E0",X"3A",X"03",X"D0",X"47",X"3C",X"E6",X"03",X"20",X"02",X"3E",X"05",
		X"77",X"23",X"78",X"0F",X"0F",X"47",X"E6",X"03",X"32",X"45",X"E0",X"3A",X"04",X"D0",X"CB",X"57",
		X"78",X"28",X"1F",X"1F",X"1F",X"ED",X"44",X"E6",X"0F",X"CB",X"5F",X"28",X"01",X"3C",X"77",X"23",
		X"77",X"3A",X"04",X"D0",X"2F",X"1F",X"47",X"E6",X"01",X"23",X"77",X"78",X"1F",X"E6",X"01",X"23",
		X"77",X"C9",X"1F",X"1F",X"2F",X"47",X"3C",X"E6",X"03",X"77",X"78",X"1F",X"1F",X"E6",X"03",X"FE",
		X"02",X"DE",X"F5",X"18",X"DA",X"CD",X"29",X"0D",X"21",X"97",X"2C",X"CD",X"00",X"03",X"CD",X"27",
		X"05",X"21",X"57",X"2C",X"CD",X"4E",X"03",X"11",X"54",X"E0",X"01",X"20",X"00",X"3A",X"44",X"E0",
		X"A7",X"20",X"34",X"CD",X"9F",X"07",X"CD",X"E8",X"07",X"7E",X"FE",X"32",X"20",X"20",X"3E",X"53",
		X"32",X"5F",X"E0",X"32",X"68",X"E0",X"21",X"62",X"E0",X"7E",X"87",X"D6",X"30",X"FE",X"3A",X"38",
		X"06",X"D6",X"0A",X"77",X"2B",X"3E",X"31",X"77",X"21",X"54",X"E0",X"CD",X"4E",X"03",X"3A",X"47",
		X"E0",X"A7",X"20",X"FA",X"C3",X"E8",X"05",X"CD",X"D3",X"07",X"CD",X"DD",X"07",X"18",X"E9",X"21",
		X"67",X"2C",X"ED",X"B0",X"21",X"57",X"E0",X"3A",X"41",X"E0",X"11",X"08",X"00",X"FE",X"08",X"38",
		X"12",X"C6",X"28",X"77",X"19",X"36",X"53",X"23",X"23",X"23",X"36",X"31",X"11",X"06",X"00",X"19",
		X"36",X"00",X"C9",X"3D",X"C8",X"11",X"0B",X"00",X"19",X"C6",X"31",X"77",X"11",X"06",X"00",X"19",
		X"36",X"53",X"C9",X"21",X"7D",X"2C",X"ED",X"B0",X"21",X"5B",X"E0",X"18",X"CA",X"CD",X"E8",X"07",
		X"21",X"5B",X"E0",X"3A",X"42",X"E0",X"18",X"C2",X"21",X"54",X"E0",X"CD",X"4E",X"03",X"2A",X"54",
		X"E0",X"11",X"40",X"00",X"19",X"22",X"54",X"E0",X"21",X"57",X"E0",X"34",X"C9",X"21",X"77",X"E2",
		X"06",X"07",X"7E",X"A7",X"28",X"0B",X"2B",X"10",X"F9",X"C9",X"21",X"61",X"E2",X"06",X"12",X"18",
		X"F1",X"34",X"7D",X"D6",X"50",X"87",X"87",X"DD",X"77",X"01",X"C9",X"DD",X"7E",X"07",X"E6",X"F8",
		X"6F",X"26",X"20",X"29",X"29",X"DD",X"7E",X"03",X"1F",X"57",X"1F",X"1F",X"E6",X"1F",X"85",X"6F",
		X"C9",X"3A",X"00",X"E3",X"FE",X"06",X"30",X"7A",X"3A",X"E2",X"E1",X"DD",X"96",X"0F",X"ED",X"44",
		X"DD",X"77",X"03",X"FE",X"E0",X"38",X"6D",X"DD",X"4E",X"0B",X"0D",X"20",X"6B",X"FE",X"E8",X"30",
		X"67",X"E1",X"DD",X"36",X"00",X"00",X"DD",X"7E",X"0D",X"37",X"17",X"D8",X"37",X"17",X"21",X"18",
		X"2E",X"30",X"01",X"24",X"5F",X"16",X"00",X"19",X"46",X"DD",X"5E",X"01",X"16",X"E1",X"78",X"17",
		X"30",X"10",X"06",X"01",X"17",X"38",X"27",X"7B",X"FE",X"60",X"38",X"06",X"62",X"D6",X"5E",X"6F",
		X"36",X"00",X"FD",X"21",X"00",X"00",X"FD",X"19",X"7B",X"1F",X"1F",X"E6",X"3F",X"C6",X"50",X"6F",
		X"26",X"E2",X"11",X"04",X"00",X"FD",X"72",X"02",X"FD",X"19",X"10",X"F9",X"72",X"C9",X"CD",X"82",
		X"08",X"21",X"74",X"E1",X"01",X"00",X"18",X"71",X"23",X"10",X"FC",X"21",X"D1",X"E1",X"70",X"23",
		X"70",X"C9",X"E1",X"C9",X"DD",X"36",X"0B",X"01",X"DD",X"7E",X"0D",X"07",X"D8",X"17",X"21",X"18",
		X"2E",X"30",X"01",X"24",X"5F",X"16",X"00",X"19",X"DD",X"5E",X"01",X"16",X"E1",X"FD",X"21",X"00",
		X"00",X"FD",X"19",X"56",X"23",X"5E",X"23",X"4E",X"06",X"00",X"21",X"F5",X"08",X"09",X"4E",X"23",
		X"66",X"69",X"DD",X"4E",X"03",X"DD",X"7E",X"07",X"CD",X"ED",X"08",X"AF",X"E9",X"2F",X"47",X"3A",
		X"3C",X"E0",X"80",X"47",X"C9",X"69",X"09",X"5A",X"09",X"CF",X"09",X"CD",X"09",X"F5",X"0A",X"43",
		X"09",X"E2",X"0A",X"90",X"0A",X"56",X"0A",X"B7",X"0A",X"52",X"0A",X"9F",X"0A",X"C9",X"09",X"25",
		X"0B",X"76",X"09",X"97",X"09",X"BA",X"09",X"1E",X"0A",X"44",X"0A",X"34",X"09",X"25",X"09",X"1D",
		X"0B",X"B0",X"09",X"83",X"09",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"E6",X"1F",X"FE",X"0B",X"38",
		X"38",X"1C",X"18",X"35",X"3A",X"4E",X"E0",X"E6",X"03",X"28",X"01",X"14",X"CD",X"69",X"09",X"16",
		X"3B",X"18",X"1B",X"FD",X"21",X"A4",X"E1",X"FD",X"77",X"0A",X"FD",X"77",X"0E",X"FD",X"77",X"12",
		X"FD",X"77",X"16",X"CD",X"95",X"0A",X"3E",X"F8",X"80",X"47",X"CD",X"69",X"09",X"14",X"3E",X"10",
		X"81",X"4F",X"21",X"04",X"00",X"EB",X"FD",X"19",X"EB",X"DD",X"7E",X"0B",X"A7",X"79",X"20",X"35",
		X"C6",X"08",X"FE",X"20",X"38",X"35",X"FD",X"70",X"00",X"FD",X"73",X"01",X"FD",X"72",X"02",X"FD",
		X"71",X"03",X"C9",X"DD",X"7E",X"08",X"1E",X"07",X"CB",X"3F",X"CB",X"13",X"C6",X"7A",X"57",X"78",
		X"FE",X"80",X"D2",X"25",X"0B",X"18",X"DF",X"3E",X"08",X"80",X"47",X"FD",X"21",X"74",X"E1",X"79",
		X"FE",X"F8",X"D0",X"18",X"D1",X"C6",X"08",X"FE",X"F0",X"38",X"CB",X"FD",X"36",X"02",X"00",X"C9",
		X"3A",X"4E",X"E0",X"CB",X"57",X"28",X"BF",X"14",X"18",X"BC",X"3E",X"0E",X"80",X"60",X"47",X"2E",
		X"01",X"CD",X"E4",X"09",X"11",X"08",X"76",X"18",X"11",X"3E",X"0A",X"18",X"02",X"3E",X"05",X"80",
		X"60",X"47",X"2E",X"01",X"CD",X"E4",X"09",X"11",X"08",X"71",X"44",X"21",X"08",X"00",X"EB",X"FD",
		X"19",X"EB",X"2E",X"00",X"CD",X"69",X"09",X"FD",X"70",X"04",X"2D",X"20",X"29",X"3E",X"40",X"AB",
		X"FD",X"77",X"05",X"3E",X"08",X"FD",X"72",X"06",X"81",X"FD",X"77",X"07",X"C6",X"08",X"FE",X"F8",
		X"30",X"0A",X"FE",X"20",X"D0",X"DD",X"7E",X"0B",X"A7",X"28",X"06",X"C9",X"DD",X"7E",X"0B",X"A7",
		X"C8",X"FD",X"36",X"06",X"00",X"C9",X"14",X"FD",X"73",X"05",X"3E",X"10",X"18",X"D7",X"C5",X"D5",
		X"21",X"02",X"08",X"09",X"44",X"4D",X"79",X"C6",X"08",X"FE",X"D0",X"30",X"11",X"CD",X"83",X"09",
		X"11",X"04",X"00",X"FD",X"19",X"D1",X"C1",X"2E",X"00",X"FD",X"75",X"0A",X"18",X"A6",X"FD",X"36",
		X"02",X"00",X"18",X"EC",X"32",X"A6",X"E1",X"32",X"AA",X"E1",X"32",X"AE",X"E1",X"CD",X"95",X"0A",
		X"18",X"10",X"3E",X"18",X"18",X"02",X"3E",X"0D",X"FD",X"21",X"74",X"E1",X"80",X"47",X"3E",X"F8",
		X"81",X"4F",X"AF",X"CD",X"6F",X"0A",X"EB",X"11",X"08",X"00",X"FD",X"19",X"EB",X"3E",X"10",X"81",
		X"6F",X"FD",X"77",X"03",X"FD",X"77",X"07",X"FD",X"70",X"00",X"3E",X"F0",X"80",X"FD",X"77",X"04",
		X"FD",X"73",X"01",X"FD",X"73",X"05",X"FD",X"72",X"02",X"14",X"14",X"FD",X"72",X"06",X"15",X"C9",
		X"CD",X"95",X"0A",X"18",X"CD",X"3A",X"F9",X"E0",X"1F",X"D0",X"7B",X"F6",X"0C",X"5F",X"C9",X"FD",
		X"21",X"74",X"E1",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"0E",X"00",X"3E",X"18",X"80",X"47",X"AF",
		X"CD",X"6F",X"0A",X"FD",X"72",X"06",X"C9",X"3E",X"18",X"80",X"47",X"FD",X"21",X"74",X"E1",X"3E",
		X"F8",X"CD",X"CD",X"0A",X"21",X"0C",X"00",X"EB",X"FD",X"19",X"EB",X"3E",X"08",X"CD",X"6F",X"0A",
		X"FD",X"75",X"0B",X"D6",X"10",X"FD",X"77",X"08",X"FD",X"77",X"09",X"7A",X"C6",X"03",X"FD",X"77",
		X"0A",X"C9",X"FD",X"21",X"A4",X"E1",X"FD",X"77",X"06",X"CD",X"95",X"0A",X"21",X"08",X"F8",X"09",
		X"44",X"4D",X"C3",X"76",X"09",X"FD",X"21",X"A4",X"E1",X"FD",X"36",X"1A",X"00",X"CD",X"95",X"0A",
		X"3E",X"F8",X"CD",X"13",X"0B",X"3E",X"08",X"CD",X"0C",X"0B",X"3E",X"18",X"EB",X"11",X"08",X"00",
		X"FD",X"19",X"EB",X"CD",X"6F",X"0A",X"7A",X"C6",X"02",X"FD",X"77",X"06",X"C9",X"3A",X"4E",X"E0",
		X"CB",X"4F",X"28",X"01",X"1C",X"CD",X"76",X"09",X"DD",X"7E",X"01",X"FE",X"60",X"D8",X"EB",X"11",
		X"A0",X"FF",X"FD",X"19",X"EB",X"C3",X"76",X"09",X"CD",X"8E",X"0C",X"CD",X"BF",X"0C",X"3A",X"04",
		X"D0",X"CB",X"6F",X"C0",X"21",X"A9",X"2A",X"CD",X"00",X"03",X"3E",X"FF",X"32",X"51",X"E0",X"21",
		X"53",X"E0",X"7E",X"4E",X"A9",X"A1",X"1F",X"38",X"08",X"3A",X"51",X"E0",X"47",X"79",X"10",X"F3",
		X"C9",X"21",X"0E",X"E5",X"7E",X"3C",X"FE",X"34",X"30",X"E0",X"77",X"2A",X"16",X"E5",X"46",X"23",
		X"7E",X"E6",X"7F",X"23",X"FE",X"06",X"20",X"F6",X"78",X"32",X"0B",X"E5",X"22",X"16",X"E5",X"32",
		X"23",X"E5",X"22",X"2E",X"E5",X"CD",X"12",X"0D",X"18",X"C0",X"CD",X"B1",X"0C",X"21",X"94",X"26",
		X"22",X"16",X"E5",X"C3",X"BF",X"0C",X"2A",X"16",X"E5",X"2B",X"7E",X"2B",X"E6",X"7F",X"FE",X"06",
		X"20",X"F7",X"11",X"DC",X"E1",X"EB",X"7E",X"36",X"00",X"EB",X"A7",X"20",X"EC",X"7E",X"32",X"0B",
		X"E5",X"23",X"23",X"22",X"16",X"E5",X"C9",X"21",X"00",X"E1",X"01",X"00",X"04",X"CD",X"FA",X"05",
		X"DD",X"21",X"00",X"E3",X"DD",X"36",X"00",X"01",X"DD",X"36",X"10",X"09",X"DD",X"36",X"01",X"B0",
		X"DD",X"36",X"21",X"A0",X"DD",X"21",X"70",X"E3",X"3E",X"60",X"06",X"09",X"11",X"10",X"00",X"DD",
		X"77",X"01",X"DD",X"19",X"C6",X"04",X"10",X"F7",X"CD",X"96",X"0B",X"2B",X"46",X"3E",X"04",X"21",
		X"00",X"C0",X"05",X"F2",X"FA",X"0B",X"3E",X"07",X"26",X"A8",X"32",X"14",X"E5",X"22",X"06",X"E3",
		X"3E",X"02",X"32",X"08",X"E5",X"CD",X"8D",X"0D",X"3A",X"13",X"E5",X"3D",X"FE",X"05",X"CE",X"00",
		X"06",X"FB",X"1F",X"38",X"01",X"04",X"78",X"32",X"C5",X"E1",X"CD",X"81",X"29",X"A7",X"20",X"5F",
		X"21",X"0F",X"E5",X"CB",X"46",X"20",X"58",X"34",X"3A",X"10",X"E5",X"A7",X"28",X"58",X"21",X"5F",
		X"2A",X"CD",X"00",X"03",X"3A",X"10",X"E5",X"FE",X"04",X"38",X"02",X"3E",X"03",X"C6",X"30",X"32",
		X"56",X"81",X"3E",X"1C",X"CD",X"6F",X"0D",X"3E",X"40",X"32",X"0A",X"E3",X"0E",X"68",X"21",X"B6",
		X"30",X"46",X"CB",X"78",X"20",X"14",X"23",X"5E",X"23",X"7E",X"23",X"EB",X"26",X"83",X"71",X"26",
		X"87",X"70",X"0C",X"2C",X"BD",X"20",X"F5",X"EB",X"18",X"E7",X"3E",X"D3",X"21",X"D8",X"30",X"11",
		X"10",X"E2",X"46",X"CB",X"78",X"20",X"08",X"12",X"13",X"10",X"FC",X"3C",X"23",X"18",X"F3",X"21",
		X"46",X"E0",X"34",X"C3",X"6E",X"02",X"21",X"47",X"2A",X"CD",X"00",X"03",X"18",X"B4",X"AF",X"32",
		X"4D",X"E0",X"CD",X"95",X"0C",X"CD",X"03",X"06",X"21",X"00",X"E5",X"01",X"16",X"00",X"CD",X"FA",
		X"05",X"32",X"0F",X"E5",X"3A",X"40",X"E0",X"32",X"15",X"E5",X"21",X"62",X"21",X"22",X"16",X"E5",
		X"C9",X"21",X"DE",X"26",X"22",X"F7",X"E0",X"21",X"03",X"E5",X"01",X"11",X"00",X"18",X"DF",X"CD",
		X"29",X"0D",X"21",X"21",X"84",X"0E",X"06",X"3A",X"0E",X"E5",X"FE",X"1A",X"3E",X"00",X"38",X"01",
		X"3C",X"32",X"F9",X"E0",X"C5",X"0E",X"01",X"CD",X"E7",X"03",X"79",X"C1",X"06",X"1E",X"77",X"23",
		X"10",X"FC",X"23",X"23",X"0D",X"20",X"F5",X"21",X"0F",X"2B",X"CD",X"00",X"03",X"CD",X"68",X"06",
		X"CD",X"85",X"06",X"3A",X"46",X"E0",X"CB",X"67",X"28",X"0F",X"CD",X"03",X"06",X"CD",X"68",X"06",
		X"CD",X"03",X"06",X"21",X"72",X"2B",X"CD",X"00",X"03",X"CD",X"D5",X"06",X"CD",X"2C",X"21",X"CD",
		X"8A",X"29",X"3A",X"0E",X"E5",X"0E",X"02",X"FE",X"1A",X"38",X"04",X"D6",X"1A",X"0E",X"07",X"C6",
		X"40",X"32",X"52",X"80",X"79",X"32",X"52",X"84",X"C9",X"21",X"00",X"80",X"01",X"00",X"08",X"CD",
		X"FA",X"05",X"21",X"00",X"E1",X"01",X"C6",X"00",X"CD",X"FA",X"05",X"3A",X"43",X"E0",X"3D",X"28",
		X"09",X"21",X"46",X"E0",X"AF",X"CB",X"5E",X"28",X"01",X"3C",X"32",X"4C",X"E0",X"21",X"04",X"D0",
		X"AE",X"21",X"3C",X"E0",X"36",X"EF",X"16",X"FF",X"1F",X"30",X"03",X"14",X"36",X"F1",X"23",X"72",
		X"01",X"00",X"40",X"AF",X"ED",X"79",X"0C",X"10",X"FB",X"F3",X"CD",X"7D",X"0D",X"FB",X"C9",X"F3",
		X"CD",X"75",X"0D",X"FB",X"C9",X"E5",X"21",X"46",X"E0",X"CB",X"7E",X"E1",X"F0",X"E5",X"2A",X"DE",
		X"E1",X"26",X"E0",X"77",X"7D",X"3C",X"E6",X"07",X"32",X"DE",X"E1",X"E1",X"C9",X"CD",X"48",X"29",
		X"CD",X"C2",X"0C",X"06",X"20",X"C5",X"CD",X"06",X"11",X"21",X"E2",X"E1",X"7E",X"C6",X"08",X"77",
		X"C1",X"10",X"F2",X"C3",X"3B",X"0D",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"01",X"4A",X"30",X"81",
		X"4F",X"0A",X"4F",X"EB",X"11",X"20",X"00",X"7E",X"A7",X"20",X"03",X"19",X"18",X"F9",X"22",X"54",
		X"E0",X"0A",X"03",X"3D",X"C8",X"F2",X"CD",X"0D",X"3C",X"77",X"19",X"18",X"F4",X"3A",X"54",X"E0",
		X"3C",X"6F",X"E6",X"1F",X"20",X"E8",X"7D",X"D6",X"20",X"6F",X"18",X"E2",X"CD",X"5B",X"12",X"3A",
		X"E2",X"E1",X"21",X"09",X"E5",X"47",X"AE",X"E6",X"F8",X"C8",X"78",X"E6",X"F8",X"77",X"CD",X"06",
		X"11",X"3A",X"4D",X"E0",X"A7",X"C0",X"21",X"0B",X"E5",X"34",X"7E",X"5F",X"A7",X"28",X"07",X"E6",
		X"1F",X"20",X"03",X"CD",X"D6",X"29",X"7B",X"2A",X"16",X"E5",X"BE",X"20",X"0B",X"23",X"7E",X"E6",
		X"7F",X"32",X"D7",X"E1",X"23",X"22",X"16",X"E5",X"21",X"D7",X"E1",X"7E",X"3D",X"F8",X"36",X"00",
		X"FE",X"18",X"D2",X"45",X"0F",X"FE",X"17",X"28",X"26",X"D6",X"06",X"FA",X"8A",X"0E",X"D6",X"07",
		X"FA",X"F0",X"0E",X"87",X"87",X"87",X"5F",X"16",X"00",X"FD",X"21",X"00",X"10",X"FD",X"19",X"CD",
		X"93",X"0E",X"FD",X"7E",X"06",X"A7",X"28",X"03",X"CD",X"FD",X"07",X"DD",X"71",X"00",X"C9",X"3E",
		X"19",X"32",X"70",X"E3",X"C9",X"3E",X"01",X"32",X"DC",X"E1",X"2A",X"E4",X"E0",X"7D",X"E6",X"1F",
		X"F6",X"C0",X"6F",X"36",X"0A",X"01",X"20",X"00",X"5D",X"09",X"36",X"0B",X"7B",X"3D",X"E6",X"1F",
		X"F6",X"C0",X"6F",X"CD",X"81",X"29",X"C6",X"41",X"77",X"22",X"DA",X"E1",X"09",X"36",X"F2",X"01",
		X"E0",X"03",X"09",X"3A",X"F9",X"E0",X"C6",X"05",X"77",X"C9",X"3C",X"28",X"C8",X"C6",X"05",X"32",
		X"08",X"E5",X"C9",X"FD",X"7E",X"00",X"FE",X"02",X"28",X"1B",X"FE",X"07",X"38",X"1C",X"16",X"00",
		X"FD",X"5E",X"05",X"DD",X"21",X"70",X"E3",X"FD",X"46",X"04",X"DD",X"7E",X"00",X"A7",X"28",X"13",
		X"DD",X"19",X"10",X"F6",X"C9",X"21",X"D7",X"E1",X"36",X"11",X"11",X"F0",X"FF",X"DD",X"21",X"F0",
		X"E4",X"18",X"E4",X"FD",X"7E",X"00",X"DD",X"77",X"0C",X"FD",X"7E",X"01",X"DD",X"77",X"0D",X"3A",
		X"09",X"E5",X"D6",X"02",X"DD",X"77",X"0F",X"CD",X"3D",X"15",X"FD",X"86",X"03",X"DD",X"77",X"07",
		X"DD",X"36",X"0B",X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"0E",X"00",X"FD",X"4E",X"02",X"C9",
		X"3C",X"CA",X"40",X"0F",X"F5",X"FD",X"21",X"4E",X"10",X"CD",X"BA",X"0E",X"F1",X"C6",X"86",X"DD",
		X"77",X"0D",X"DD",X"71",X"00",X"21",X"4A",X"30",X"85",X"C6",X"80",X"6F",X"6E",X"FD",X"2A",X"E4",
		X"E0",X"11",X"20",X"00",X"7E",X"23",X"3D",X"F2",X"22",X"0F",X"3C",X"FD",X"77",X"00",X"FD",X"19",
		X"18",X"F2",X"C8",X"22",X"E6",X"E0",X"3D",X"28",X"11",X"FD",X"21",X"55",X"10",X"CD",X"9E",X"0E",
		X"DD",X"36",X"0A",X"00",X"DD",X"34",X"0E",X"DD",X"71",X"00",X"3E",X"0D",X"32",X"D7",X"E1",X"C9",
		X"2A",X"E6",X"E0",X"18",X"C8",X"D6",X"1F",X"FA",X"B7",X"0F",X"21",X"C5",X"E1",X"0E",X"FF",X"23",
		X"0C",X"D6",X"08",X"F2",X"4F",X"0F",X"C6",X"08",X"28",X"10",X"77",X"23",X"23",X"23",X"77",X"23",
		X"23",X"23",X"77",X"0D",X"F8",X"21",X"D6",X"E1",X"34",X"C9",X"77",X"FD",X"21",X"70",X"E3",X"11",
		X"10",X"00",X"06",X"19",X"0D",X"FA",X"A5",X"0F",X"FD",X"7E",X"00",X"D6",X"22",X"FE",X"06",X"30",
		X"19",X"6F",X"CB",X"4D",X"20",X"14",X"61",X"FD",X"7E",X"0D",X"FE",X"2A",X"20",X"01",X"24",X"25",
		X"20",X"08",X"CB",X"55",X"20",X"09",X"FD",X"36",X"00",X"24",X"FD",X"19",X"10",X"DA",X"C9",X"FD",
		X"36",X"0F",X"01",X"18",X"F5",X"FD",X"7E",X"00",X"D6",X"1E",X"FE",X"02",X"30",X"04",X"FD",X"36",
		X"00",X"24",X"FD",X"19",X"10",X"EF",X"C9",X"C6",X"08",X"FE",X"04",X"30",X"08",X"21",X"0B",X"E5",
		X"46",X"23",X"70",X"23",X"77",X"3A",X"D5",X"E1",X"A7",X"C8",X"5F",X"16",X"00",X"FD",X"21",X"FF",
		X"E3",X"FD",X"19",X"21",X"70",X"E3",X"1E",X"10",X"01",X"3A",X"05",X"7E",X"A7",X"CA",X"5D",X"10",
		X"19",X"10",X"F8",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
