library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_K1_High is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(3 downto 0)
);
end entity;

architecture prom of ROM_K1_High is
	type rom is array(0 to  2047) of std_logic_vector(3 downto 0);
	signal rom_data: rom := (
		X"3",X"4",X"4",X"A",X"1",X"1",X"F",X"C",X"C",X"5",X"5",X"5",X"1",X"1",X"0",X"3",
		X"4",X"4",X"A",X"1",X"1",X"B",X"4",X"5",X"5",X"6",X"6",X"1",X"1",X"0",X"4",X"4",
		X"4",X"A",X"1",X"0",X"4",X"4",X"5",X"5",X"6",X"6",X"1",X"1",X"0",X"4",X"4",X"4",
		X"A",X"1",X"0",X"3",X"4",X"5",X"5",X"6",X"6",X"1",X"0",X"0",X"4",X"4",X"4",X"A",
		X"0",X"0",X"3",X"4",X"5",X"6",X"6",X"F",X"9",X"0",X"0",X"4",X"4",X"4",X"A",X"0",
		X"0",X"3",X"3",X"5",X"6",X"6",X"B",X"A",X"0",X"0",X"4",X"4",X"4",X"A",X"0",X"0",
		X"3",X"3",X"4",X"C",X"C",X"C",X"2",X"0",X"0",X"4",X"4",X"4",X"A",X"0",X"0",X"2",
		X"2",X"3",X"2",X"2",X"2",X"1",X"0",X"0",X"4",X"4",X"4",X"A",X"0",X"0",X"2",X"2",
		X"2",X"2",X"2",X"2",X"1",X"0",X"0",X"4",X"4",X"4",X"A",X"0",X"0",X"2",X"2",X"2",
		X"2",X"2",X"1",X"1",X"0",X"0",X"4",X"4",X"4",X"A",X"0",X"0",X"2",X"2",X"2",X"2",
		X"1",X"1",X"1",X"0",X"F",X"5",X"4",X"4",X"A",X"0",X"7",X"9",X"2",X"2",X"2",X"1",
		X"1",X"1",X"0",X"B",X"5",X"4",X"4",X"A",X"0",X"7",X"D",X"C",X"C",X"C",X"C",X"C",
		X"C",X"C",X"5",X"5",X"4",X"4",X"3",X"3",X"4",X"C",X"C",X"8",X"4",X"4",X"4",X"4",
		X"8",X"8",X"4",X"4",X"4",X"3",X"3",X"C",X"3",X"3",X"3",X"9",X"4",X"4",X"F",X"3",
		X"3",X"C",X"9",X"5",X"2",X"F",X"2",X"3",X"3",X"3",X"D",X"4",X"4",X"B",X"2",X"3",
		X"3",X"D",X"5",X"2",X"A",X"2",X"3",X"3",X"3",X"3",X"8",X"8",X"2",X"2",X"3",X"3",
		X"4",X"9",X"2",X"2",X"2",X"2",X"3",X"3",X"3",X"3",X"2",X"2",X"2",X"3",X"3",X"4",
		X"E",X"2",X"2",X"1",X"2",X"2",X"2",X"2",X"2",X"2",X"1",X"1",X"3",X"3",X"4",X"E",
		X"2",X"1",X"1",X"2",X"2",X"3",X"2",X"2",X"1",X"1",X"C",X"9",X"3",X"4",X"5",X"E",
		X"1",X"1",X"1",X"9",X"2",X"2",X"2",X"1",X"F",X"7",X"E",X"3",X"4",X"5",X"E",X"1",
		X"1",X"F",X"D",X"2",X"2",X"1",X"1",X"B",X"0",X"2",X"4",X"4",X"5",X"A",X"1",X"1",
		X"B",X"1",X"9",X"1",X"1",X"F",X"7",X"0",X"2",X"4",X"4",X"5",X"A",X"1",X"0",X"6",
		X"6",X"D",X"1",X"1",X"B",X"7",X"0",X"2",X"4",X"4",X"5",X"A",X"0",X"0",X"6",X"6",
		X"1",X"8",X"C",X"0",X"7",X"0",X"2",X"4",X"4",X"5",X"A",X"0",X"0",X"6",X"6",X"0",
		X"0",X"0",X"0",X"4",X"4",X"E",X"5",X"5",X"5",X"A",X"0",X"0",X"A",X"5",X"0",X"0",
		X"0",X"0",X"4",X"4",X"B",X"5",X"5",X"5",X"A",X"0",X"7",X"E",X"4",X"4",X"4",X"4",
		X"4",X"4",X"8",X"5",X"5",X"5",X"5",X"A",X"0",X"7",X"7",X"4",X"4",X"4",X"4",X"3",
		X"8",X"4",X"5",X"5",X"5",X"5",X"A",X"0",X"7",X"7",X"9",X"4",X"4",X"4",X"8",X"5",
		X"5",X"5",X"5",X"5",X"5",X"A",X"0",X"7",X"7",X"D",X"8",X"8",X"C",X"5",X"5",X"5",
		X"5",X"5",X"5",X"5",X"4",X"2",X"3",X"C",X"C",X"C",X"C",X"9",X"3",X"3",X"C",X"C",
		X"C",X"C",X"5",X"4",X"3",X"C",X"4",X"4",X"4",X"4",X"D",X"5",X"F",X"3",X"3",X"4",
		X"4",X"9",X"4",X"F",X"3",X"2",X"2",X"3",X"4",X"5",X"9",X"B",X"1",X"2",X"3",X"3",
		X"D",X"4",X"B",X"2",X"2",X"2",X"3",X"3",X"5",X"E",X"2",X"1",X"2",X"3",X"4",X"5",
		X"3",X"2",X"1",X"2",X"2",X"2",X"3",X"5",X"E",X"1",X"1",X"2",X"3",X"4",X"5",X"E",
		X"2",X"1",X"2",X"2",X"2",X"4",X"4",X"E",X"1",X"0",X"1",X"3",X"4",X"4",X"A",X"1",
		X"1",X"4",X"6",X"8",X"4",X"4",X"E",X"0",X"0",X"0",X"3",X"4",X"5",X"A",X"1",X"2",
		X"4",X"E",X"0",X"4",X"5",X"E",X"0",X"1",X"0",X"3",X"4",X"4",X"A",X"1",X"2",X"3",
		X"D",X"F",X"5",X"5",X"E",X"0",X"1",X"7",X"3",X"4",X"4",X"A",X"0",X"0",X"3",X"4",
		X"B",X"5",X"5",X"E",X"1",X"7",X"7",X"3",X"4",X"4",X"A",X"0",X"0",X"2",X"3",X"4",
		X"4",X"6",X"B",X"1",X"0",X"7",X"3",X"4",X"4",X"A",X"0",X"0",X"2",X"3",X"4",X"4",
		X"F",X"1",X"0",X"0",X"7",X"3",X"4",X"4",X"A",X"0",X"0",X"2",X"3",X"3",X"3",X"B",
		X"1",X"0",X"0",X"7",X"4",X"4",X"4",X"A",X"0",X"0",X"9",X"2",X"3",X"2",X"1",X"2",
		X"1",X"1",X"7",X"4",X"4",X"4",X"A",X"0",X"7",X"D",X"1",X"2",X"2",X"1",X"2",X"1",
		X"1",X"E",X"5",X"5",X"4",X"A",X"0",X"7",X"7",X"9",X"1",X"1",X"1",X"1",X"1",X"7",
		X"B",X"5",X"6",X"4",X"A",X"0",X"7",X"7",X"D",X"0",X"0",X"0",X"0",X"0",X"F",X"5",
		X"5",X"5",X"4",X"A",X"0",X"7",X"7",X"7",X"C",X"C",X"C",X"C",X"C",X"B",X"5",X"5",
		X"5",X"5",X"3",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"9",X"3",X"C",X"C",X"C",X"C",
		X"9",X"F",X"3",X"3",X"3",X"3",X"3",X"3",X"4",X"D",X"F",X"3",X"3",X"3",X"4",X"D",
		X"A",X"2",X"2",X"2",X"2",X"3",X"3",X"4",X"5",X"A",X"2",X"3",X"3",X"4",X"5",X"A",
		X"2",X"2",X"2",X"2",X"3",X"3",X"4",X"4",X"A",X"2",X"2",X"3",X"4",X"5",X"A",X"2",
		X"2",X"2",X"2",X"2",X"3",X"4",X"4",X"A",X"2",X"2",X"3",X"4",X"6",X"A",X"1",X"1",
		X"8",X"8",X"8",X"3",X"4",X"4",X"A",X"1",X"1",X"3",X"4",X"4",X"A",X"1",X"0",X"6",
		X"D",X"0",X"3",X"4",X"4",X"A",X"1",X"1",X"A",X"4",X"5",X"A",X"1",X"7",X"7",X"6",
		X"8",X"4",X"4",X"5",X"A",X"1",X"0",X"A",X"4",X"5",X"A",X"0",X"0",X"7",X"6",X"E",
		X"3",X"4",X"5",X"A",X"1",X"0",X"A",X"4",X"5",X"D",X"0",X"7",X"7",X"7",X"E",X"3",
		X"4",X"6",X"A",X"0",X"0",X"A",X"4",X"5",X"1",X"9",X"0",X"7",X"7",X"E",X"3",X"3",
		X"F",X"A",X"0",X"0",X"A",X"4",X"5",X"3",X"C",X"C",X"7",X"7",X"E",X"3",X"3",X"D",
		X"B",X"0",X"0",X"A",X"4",X"5",X"F",X"3",X"2",X"0",X"7",X"E",X"3",X"3",X"3",X"1",
		X"0",X"0",X"A",X"4",X"5",X"A",X"3",X"1",X"0",X"7",X"E",X"2",X"2",X"2",X"1",X"0",
		X"0",X"A",X"4",X"5",X"A",X"2",X"1",X"0",X"0",X"E",X"2",X"2",X"1",X"1",X"0",X"0",
		X"A",X"4",X"5",X"A",X"1",X"1",X"0",X"0",X"C",X"2",X"2",X"1",X"1",X"0",X"7",X"B",
		X"5",X"5",X"A",X"1",X"1",X"0",X"F",X"7",X"9",X"1",X"1",X"0",X"0",X"F",X"5",X"5",
		X"5",X"A",X"1",X"0",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"C",X"B",X"5",X"5",X"5",
		X"8",X"0",X"A",X"0",X"A",X"0",X"9",X"9",X"0",X"0",X"C",X"9",X"9",X"0",X"0",X"C",
		X"9",X"9",X"0",X"0",X"C",X"9",X"9",X"0",X"0",X"8",X"8",X"E",X"D",X"E",X"9",X"5",
		X"0",X"0",X"9",X"0",X"0",X"D",X"2",X"C",X"9",X"5",X"0",X"0",X"9",X"0",X"0",X"D",
		X"1",X"C",X"9",X"5",X"0",X"0",X"9",X"0",X"0",X"D",X"1",X"C",X"9",X"5",X"0",X"0",
		X"9",X"0",X"0",X"D",X"0",X"8",X"8",X"E",X"D",X"D",X"C",X"D",X"B",X"F",X"3",X"A",
		X"0",X"8",X"0",X"0",X"A",X"0",X"A",X"0",X"C",X"0",X"F",X"2",X"1",X"2",X"9",X"0",
		X"8",X"4",X"8",X"6",X"8",X"D",X"F",X"C",X"D",X"F",X"F",X"0",X"8",X"4",X"8",X"6",
		X"8",X"D",X"F",X"C",X"D",X"F",X"8",X"4",X"8",X"6",X"8",X"D",X"F",X"C",X"D",X"F",
		X"F",X"D",X"8",X"0",X"F",X"F",X"A",X"0",X"A",X"0",X"A",X"0",X"2",X"3",X"3",X"A",
		X"0",X"8",X"C",X"8",X"C",X"8",X"B",X"A",X"2",X"8",X"B",X"A",X"0",X"B",X"B",X"1",
		X"6",X"C",X"8",X"C",X"C",X"D",X"F",X"E",X"B",X"C",X"D",X"F",X"A",X"C",X"D",X"0",
		X"E",X"C",X"A",X"C",X"C",X"0",X"9",X"E",X"4",X"B",X"3",X"A",X"C",X"1",X"6",X"7",
		X"8",X"B",X"0",X"A",X"2",X"8",X"B",X"0",X"2",X"D",X"3",X"8",X"B",X"A",X"0",X"9",
		X"6",X"9",X"6",X"C",X"C",X"1",X"F",X"2",X"D",X"3",X"4",X"B",X"F",X"E",X"A",X"0",
		X"9",X"6",X"9",X"6",X"C",X"C",X"1",X"F",X"3",X"E",X"A",X"0",X"1",X"A",X"0",X"4",
		X"2",X"F",X"3",X"B",X"B",X"1",X"6",X"3",X"1",X"5",X"3",X"B",X"4",X"3",X"8",X"C",
		X"B",X"4",X"3",X"8",X"C",X"A",X"0",X"9",X"C",X"6",X"5",X"4",X"5",X"2",X"9",X"6",
		X"5",X"2",X"C",X"C",X"1",X"D",X"2",X"8",X"6",X"0",X"4",X"8",X"4",X"9",X"4",X"D",
		X"A",X"D",X"C",X"5",X"D",X"1",X"A",X"E",X"C",X"A",X"D",X"0",X"B",X"B",X"0",X"0",
		X"C",X"4",X"9",X"3",X"4",X"E",X"3",X"7",X"D",X"A",X"F",X"9",X"A",X"0",X"9",X"0",
		X"C",X"3",X"F",X"A",X"5",X"8",X"D",X"A",X"A",X"8",X"E",X"A",X"0",X"A",X"C",X"9",
		X"A",X"9",X"9",X"B",X"C",X"3",X"9",X"A",X"C",X"C",X"1",X"F",X"A",X"0",X"4",X"C",
		X"A",X"D",X"0",X"2",X"0",X"4",X"4",X"8",X"3",X"A",X"0",X"B",X"A",X"1",X"6",X"8",
		X"B",X"A",X"0",X"8",X"4",X"B",X"0",X"1",X"0",X"A",X"1",X"2",X"B",X"D",X"0",X"0",
		X"2",X"B",X"D",X"2",X"A",X"6",X"D",X"1",X"A",X"0",X"8",X"4",X"B",X"0",X"1",X"0",
		X"B",X"A",X"2",X"6",X"0",X"1",X"D",X"0",X"A",X"1",X"2",X"B",X"D",X"0",X"0",X"2",
		X"B",X"F",X"0",X"A",X"4",X"8",X"B",X"A",X"8",X"3",X"A",X"0",X"B",X"9",X"A",X"2",
		X"0",X"1",X"3",X"1",X"A",X"C",X"D",X"1",X"B",X"A",X"0",X"1",X"1",X"A",X"0",X"0",
		X"3",X"0",X"A",X"F",X"9",X"1",X"7",X"9",X"9",X"9",X"A",X"B",X"3",X"A",X"9",X"A",
		X"2",X"9",X"3",X"B",X"2",X"4",X"8",X"2",X"3",X"C",X"B",X"C",X"C",X"F",X"D",X"0",
		X"F",X"E",X"A",X"6",X"4",X"9",X"0",X"F",X"E",X"B",X"E",X"4",X"F",X"0",X"A",X"B",
		X"0",X"4",X"8",X"B",X"2",X"D",X"3",X"C",X"C",X"3",X"0",X"4",X"5",X"3",X"6",X"A",
		X"6",X"A",X"6",X"4",X"A",X"0",X"B",X"0",X"3",X"8",X"4",X"B",X"0",X"3",X"0",X"8",
		X"D",X"F",X"9",X"B",X"6",X"0",X"0",X"0",X"A",X"0",X"B",X"A",X"2",X"F",X"9",X"A",
		X"C",X"C",X"1",X"F",X"A",X"0",X"8",X"A",X"8",X"8",X"B",X"A",X"3",X"F",X"A",X"0",
		X"1",X"0",X"C",X"F",X"B",X"0",X"9",X"3",X"C",X"0",X"B",X"2",X"B",X"A",X"3",X"F",
		X"A",X"0",X"1",X"0",X"C",X"F",X"9",X"2",X"B",X"0",X"C",X"0",X"B",X"1",X"B",X"A",
		X"3",X"0",X"B",X"A",X"0",X"1",X"1",X"B",X"C",X"D",X"0",X"A",X"2",X"9",X"C",X"B",
		X"C",X"0",X"D",X"0",X"A",X"2",X"9",X"C",X"0",X"8",X"8",X"1",X"B",X"C",X"C",X"D",
		X"B",X"6",X"B",X"A",X"3",X"0",X"A",X"8",X"9",X"9",X"A",X"0",X"9",X"A",X"9",X"8",
		X"9",X"D",X"9",X"D",X"9",X"2",X"A",X"C",X"9",X"A",X"9",X"9",X"9",X"8",X"B",X"C",
		X"3",X"9",X"A",X"2",X"1",X"3",X"6",X"A",X"0",X"2",X"6",X"3",X"2",X"9",X"3",X"C",
		X"C",X"1",X"F",X"6",X"A",X"B",X"1",X"0",X"A",X"C",X"D",X"0",X"A",X"6",X"2",X"0",
		X"D",X"2",X"B",X"E",X"4",X"F",X"2",X"B",X"A",X"3",X"2",X"9",X"6",X"B",X"2",X"3",
		X"1",X"D",X"E",X"D",X"E",X"B",X"A",X"0",X"8",X"9",X"A",X"A",X"B",X"0",X"8",X"8",
		X"B",X"2",X"6",X"3",X"9",X"6",X"4",X"D",X"3",X"A",X"B",X"2",X"1",X"D",X"F",X"B",
		X"A",X"3",X"0",X"9",X"6",X"6",X"E",X"0",X"D",X"0",X"A",X"0",X"8",X"D",X"B",X"E",
		X"C",X"0",X"9",X"1",X"B",X"A",X"3",X"0",X"E",X"D",X"E",X"D",X"C",X"1",X"9",X"0",
		X"A",X"1",X"9",X"E",X"4",X"F",X"3",X"0",X"C",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",
		X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"0",X"2",X"9",X"3",X"2",X"2",X"3",X"4",X"8",
		X"3",X"A",X"0",X"8",X"B",X"8",X"0",X"8",X"D",X"A",X"0",X"8",X"C",X"2",X"0",X"1",
		X"5",X"1",X"2",X"A",X"3",X"2",X"D",X"3",X"2",X"3",X"3",X"E",X"B",X"A",X"B",X"D",
		X"0",X"2",X"A",X"3",X"4",X"A",X"3",X"2",X"0",X"1",X"7",X"0",X"4",X"F",X"3",X"A",
		X"0",X"A",X"F",X"3",X"9",X"9",X"9",X"9",X"6",X"2",X"9",X"3",X"C",X"C",X"1",X"F",
		X"A",X"0",X"8",X"C",X"8",X"0",X"8",X"4",X"2",X"0",X"1",X"1",X"F",X"2",X"0",X"1",
		X"3",X"F",X"8",X"4",X"2",X"2",X"3",X"E",X"B",X"2",X"B",X"3",X"0",X"7",X"1",X"5",
		X"B",X"A",X"B",X"2",X"3",X"D",X"1",X"A",X"C",X"C",X"0",X"D",X"0",X"2",X"8",X"3");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
