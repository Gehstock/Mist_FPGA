library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"00",X"0F",X"00",X"F0",X"C0",X"00",X"22",X"00",X"32",X"C0",X"33",X"2C",X"33",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3F",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"F3",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"FF",X"00",X"FF",X"00",X"CC",X"00",X"BF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"22",X"00",X"22",X"00",X"32",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"00",X"CC",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"F3",X"33",X"FF",X"33",X"FF",X"E3",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"FF",X"CC",X"FF",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"33",X"CC",X"23",X"3C",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"E3",X"33",
		X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"FE",X"33",X"FE",X"EC",X"EE",X"C0",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"E3",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"FF",X"CC",X"FF",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"C3",X"33",X"3C",X"23",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"E3",X"33",
		X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"FE",X"33",X"EE",X"33",X"EE",X"CC",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"22",X"00",X"32",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"3C",X"03",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"CB",X"33",X"0C",X"33",X"00",X"32",X"00",X"C2",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"2C",X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"2C",X"22",X"C0",X"2C",X"00",
		X"2C",X"00",X"2C",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"FF",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"CF",X"00",X"0F",X"00",X"0B",X"00",X"BB",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",X"33",X"F3",X"33",X"F3",X"33",
		X"00",X"0C",X"00",X"CA",X"00",X"AF",X"00",X"CC",X"00",X"CC",X"CA",X"CC",X"CA",X"AC",X"0C",X"AB",
		X"AA",X"00",X"44",X"00",X"FF",X"00",X"FC",X"0C",X"FF",X"CA",X"AA",X"F4",X"AC",X"CF",X"CA",X"FF",
		X"C0",X"AB",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"AA",X"00",X"BB",X"00",X"CB",X"00",X"0B",
		X"CC",X"FF",X"CC",X"CF",X"BB",X"CC",X"BB",X"CB",X"BC",X"BC",X"BB",X"C0",X"0B",X"00",X"CC",X"00",
		X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"CC",X"33",X"00",X"33",X"00",X"C3",X"00",X"0C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"2C",X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"23",X"22",X"23",X"2C",X"C2",X"C0",X"C2",X"00",
		X"2C",X"00",X"2B",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0C",X"FF",X"0C",X"FF",X"00",X"CF",
		X"CC",X"00",X"CC",X"00",X"FF",X"00",X"CC",X"00",X"BC",X"F0",X"CC",X"FC",X"FF",X"CF",X"CF",X"CF",
		X"00",X"FF",X"CF",X"FF",X"CF",X"FF",X"CF",X"FF",X"00",X"FF",X"0C",X"FE",X"0C",X"EC",X"00",X"0C",
		X"CF",X"CF",X"CF",X"CF",X"EF",X"FE",X"CE",X"EE",X"CC",X"E0",X"CC",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"EE",X"00",X"EE",X"0C",X"EE",X"CE",X"EE",X"CC",X"EE",
		X"EE",X"00",X"EE",X"00",X"FF",X"C0",X"CF",X"EC",X"FF",X"ED",X"EC",X"ED",X"CC",X"FF",X"CC",X"CF",
		X"EC",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"CC",X"FF",X"00",X"FF",X"00",X"EE",X"00",X"DD",
		X"EE",X"FF",X"DE",X"DD",X"ED",X"DD",X"ED",X"DC",X"ED",X"C0",X"DD",X"00",X"CD",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"DF",X"00",X"FD",X"00",X"FF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"00",X"FF",X"00",X"FF",X"F0",X"FF",X"FD",
		X"00",X"CF",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"CC",X"FD",X"CF",X"FD",X"CF",X"FD",X"CF",X"FD",X"CF",X"FD",X"CF",X"FD",X"CF",X"FD",X"FC",X"FD",
		X"00",X"00",X"00",X"F0",X"00",X"FF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CF",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"99",X"FF",X"99",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"EF",X"FF",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"FF",X"00",X"FF",X"EE",X"FF",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"DD",X"0E",X"DD",X"00",X"DD",X"00",X"ED",
		X"FF",X"FC",X"0F",X"FC",X"00",X"FC",X"00",X"FC",X"D0",X"FC",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"00",X"CE",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"D0",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"FF",X"00",X"CF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"CF",X"00",X"FC",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"FF",X"FC",X"CF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FF",X"FC",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"0F",
		X"FF",X"FF",X"FF",X"FA",X"AA",X"AA",X"AA",X"AC",X"CC",X"CC",X"CC",X"CF",X"FF",X"FE",X"EE",X"EE",
		X"FF",X"AA",X"AA",X"AC",X"AA",X"CE",X"CC",X"FE",X"CC",X"CC",X"FF",X"00",X"CC",X"00",X"C0",X"00",
		X"ED",X"2A",X"22",X"2A",X"22",X"FF",X"FF",X"FE",X"FF",X"CC",X"CC",X"AA",X"AA",X"AA",X"CC",X"CC",
		X"FC",X"00",X"FA",X"00",X"CA",X"C0",X"CA",X"C0",X"AA",X"00",X"AC",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"1F",X"FF",X"E1",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"22",X"00",X"FF",X"EE",X"FF",X"EE",X"FF",X"11",
		X"CC",X"11",X"00",X"FE",X"00",X"FC",X"00",X"FB",X"00",X"BF",X"00",X"BB",X"00",X"CB",X"00",X"0C",
		X"11",X"DD",X"DD",X"CC",X"22",X"00",X"22",X"BC",X"FF",X"BB",X"2B",X"BC",X"BB",X"C0",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"0E",
		X"00",X"0F",X"00",X"F9",X"0F",X"8F",X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"CC",X"AA",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"EE",X"CC",X"CE",X"EE",X"0C",X"EE",X"AA",X"32",X"AA",X"F2",X"AA",X"CF",X"AA",X"AC",X"CC",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"05",X"FF",
		X"00",X"FF",X"00",X"33",X"00",X"33",X"FF",X"FF",X"FF",X"32",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C0",X"33",X"FF",X"33",X"FF",X"FF",X"22",X"22",X"EE",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"EE",X"00",X"EE",X"C0",X"FE",X"EE",X"FF",X"E5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"05",X"00",X"0E",X"00",X"0C",
		X"00",X"0E",X"00",X"F3",X"0F",X"3F",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"55",X"FF",X"EE",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"EE",X"0C",X"EE",X"00",X"32",X"BB",X"32",X"BB",X"E2",X"BB",X"FF",X"BB",X"B2",X"CC",X"BB",
		X"EE",X"00",X"33",X"C0",X"FF",X"EE",X"22",X"EE",X"FF",X"FE",X"FF",X"EF",X"FF",X"F5",X"55",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"EE",X"00",X"E5",X"00",X"5D",X"00",X"DC",X"00",
		X"EE",X"DD",X"EE",X"CE",X"22",X"BE",X"22",X"BF",X"22",X"FF",X"FF",X"EB",X"CC",X"BB",X"BB",X"BC",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",
		X"05",X"55",X"0C",X"55",X"00",X"EE",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"55",X"FF",X"55",X"55",X"EE",X"55",X"CE",X"EE",X"CC",X"EE",X"C0",X"EE",X"CF",X"32",
		X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"FC",X"32",X"FE",X"32",X"FF",X"E2",X"CC",X"FF",X"BB",X"CF",X"BB",X"BC",X"CC",X"BB",X"00",X"CC",
		X"FF",X"FF",X"FF",X"F5",X"55",X"55",X"55",X"5E",X"EE",X"ED",X"EE",X"DD",X"ED",X"2C",X"22",X"2F",
		X"EF",X"55",X"55",X"5D",X"55",X"CC",X"DD",X"00",X"CC",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"22",X"2B",X"22",X"2B",X"22",X"FF",X"FF",X"FE",X"FF",X"CC",X"CC",X"BB",X"BB",X"BB",X"CC",X"CC",
		X"FC",X"00",X"FB",X"00",X"CB",X"C0",X"CB",X"C0",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"0A",X"BB",X"0A",X"BA",X"0C",X"AF",X"00",X"FF",X"0A",X"FF",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"00",X"BB",X"AA",X"BB",X"AF",X"AA",X"AF",X"FA",X"AC",X"FA",
		X"0A",X"FF",X"0A",X"AA",X"0C",X"BA",X"00",X"CB",X"00",X"AA",X"00",X"AA",X"00",X"CA",X"00",X"0C",
		X"AA",X"FA",X"AA",X"AA",X"CA",X"44",X"AB",X"CC",X"AA",X"BC",X"AA",X"4B",X"AA",X"C4",X"AB",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"0A",X"BB",X"0A",X"BB",X"0C",X"AF",X"00",X"FF",X"0A",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"BB",X"AA",X"BB",X"AF",X"AA",X"AF",X"FA",X"AC",X"FA",
		X"0A",X"FF",X"0A",X"AA",X"0C",X"BA",X"00",X"CB",X"00",X"AA",X"00",X"AA",X"00",X"CA",X"00",X"AC",
		X"AA",X"FA",X"AA",X"AA",X"CA",X"44",X"CC",X"CC",X"AA",X"BC",X"AA",X"44",X"AA",X"C4",X"AB",X"0C",
		X"00",X"A0",X"0A",X"4A",X"A4",X"BA",X"AA",X"AA",X"CC",X"FF",X"0A",X"FF",X"AA",X"FF",X"AA",X"CC",
		X"00",X"AC",X"0A",X"4A",X"0A",X"BB",X"AA",X"BA",X"FF",X"AC",X"FF",X"AA",X"FF",X"AA",X"AC",X"AA",
		X"AA",X"AA",X"CB",X"AA",X"0C",X"BB",X"00",X"AA",X"0A",X"AA",X"0C",X"AA",X"00",X"CA",X"00",X"AA",
		X"AA",X"A4",X"AA",X"44",X"C4",X"CC",X"AB",X"4C",X"AA",X"44",X"AB",X"CC",X"B4",X"00",X"BB",X"00",
		X"00",X"00",X"00",X"A0",X"0A",X"4A",X"A4",X"BA",X"AA",X"AA",X"CC",X"FF",X"0A",X"FF",X"AA",X"FC",
		X"00",X"00",X"00",X"AC",X"0A",X"4A",X"0A",X"BB",X"AA",X"BA",X"FF",X"AC",X"FF",X"AA",X"CC",X"AA",
		X"AA",X"FC",X"AA",X"AA",X"CB",X"AA",X"0C",X"BB",X"00",X"AA",X"00",X"AA",X"0A",X"AA",X"0C",X"CA",
		X"AC",X"AA",X"AA",X"A4",X"AA",X"44",X"44",X"CC",X"AB",X"44",X"AA",X"4C",X"AB",X"C0",X"B4",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"0A",X"BB",X"0A",X"BA",X"0C",X"AF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"BB",X"AA",X"BB",X"AF",X"AA",X"AF",X"FA",
		X"0A",X"FF",X"0A",X"FF",X"0A",X"AA",X"0C",X"BA",X"00",X"AB",X"00",X"AA",X"00",X"CA",X"00",X"AC",
		X"AF",X"FA",X"AC",X"FA",X"AA",X"AA",X"CA",X"44",X"A4",X"BC",X"AA",X"B4",X"AA",X"C4",X"AA",X"B4",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"0A",X"BB",X"0A",X"BA",X"0C",X"AF",X"00",X"FF",X"0A",X"FF",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"00",X"BB",X"AA",X"BB",X"AF",X"AA",X"AF",X"FA",X"AF",X"FA",
		X"0A",X"FC",X"0A",X"AA",X"0C",X"BA",X"00",X"CB",X"00",X"AA",X"00",X"AA",X"00",X"CA",X"00",X"0A",
		X"AA",X"FA",X"AA",X"AA",X"CA",X"44",X"A4",X"CC",X"AA",X"BC",X"AA",X"44",X"AA",X"C4",X"AB",X"CC",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"0A",X"BB",X"0A",X"BA",X"0C",X"AA",X"00",X"AF",X"0A",X"AF",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"00",X"BB",X"AA",X"BB",X"FA",X"FA",X"FA",X"FF",X"FA",X"CF",
		X"0A",X"AF",X"0A",X"AA",X"0C",X"BA",X"00",X"CB",X"00",X"AA",X"00",X"AA",X"00",X"CA",X"00",X"CA",
		X"AA",X"FF",X"AA",X"AA",X"AC",X"44",X"BA",X"CC",X"AA",X"B4",X"AA",X"44",X"AA",X"CC",X"AB",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"44",X"0A",X"BA",X"0C",X"AA",X"0A",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"44",X"AA",X"BB",X"FA",X"FA",X"FA",X"FF",
		X"0A",X"AF",X"0A",X"AF",X"0C",X"BA",X"00",X"CB",X"00",X"AA",X"00",X"AA",X"00",X"AC",X"00",X"AC",
		X"FA",X"CF",X"AA",X"FF",X"AC",X"44",X"CC",X"CC",X"AA",X"B4",X"AA",X"44",X"AA",X"CC",X"AA",X"C0",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"0A",X"BA",X"0C",X"AF",X"00",X"FF",X"0A",X"FF",X"0A",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"44",X"AA",X"BB",X"AC",X"AA",X"AF",X"FA",X"4A",X"FF",X"CC",X"AA",
		X"0C",X"BA",X"00",X"CB",X"00",X"CA",X"00",X"AA",X"00",X"AA",X"00",X"CA",X"00",X"AC",X"00",X"C0",
		X"CC",X"44",X"44",X"CC",X"AB",X"C0",X"AA",X"B4",X"AA",X"4C",X"AA",X"C4",X"AB",X"44",X"CC",X"CC",
		X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FA",X"00",X"AC",X"0A",X"AC",X"0A",X"AA",X"0C",X"AA",
		X"00",X"00",X"00",X"00",X"AA",X"F0",X"CA",X"FF",X"CC",X"AB",X"CC",X"AB",X"CC",X"B4",X"AB",X"44",
		X"00",X"CB",X"00",X"AA",X"00",X"BA",X"00",X"BA",X"00",X"CA",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"BB",X"CB",X"AA",X"CB",X"AA",X"BB",X"AA",X"44",X"AA",X"CC",X"AB",X"00",X"CC",X"00",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AB",
		X"00",X"00",X"00",X"00",X"4B",X"00",X"CA",X"00",X"AC",X"BB",X"AA",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"AA",X"BA",X"CA",X"AA",X"0C",X"AA",X"0A",X"AA",X"AA",X"4A",X"CA",X"4B",X"0A",X"4C",X"0C",X"C0",
		X"BB",X"BC",X"AB",X"CB",X"AB",X"BC",X"AB",X"CA",X"B4",X"CA",X"B4",X"AA",X"CC",X"AA",X"BB",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"00",X"AC",X"00",X"AA",X"00",X"AB",
		X"00",X"00",X"00",X"00",X"4B",X"00",X"CA",X"00",X"AC",X"BB",X"AA",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"AA",X"BA",X"CA",X"AA",X"0C",X"AA",X"0A",X"AA",X"AA",X"4A",X"CA",X"4B",X"0A",X"4C",X"0C",X"CB",
		X"BB",X"BC",X"AB",X"CB",X"AB",X"BC",X"AB",X"CA",X"B4",X"CA",X"B4",X"AA",X"CC",X"AA",X"00",X"44",
		X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"AA",X"00",X"4B",X"0A",X"BB",X"00",X"AA",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"BB",X"AA",X"BB",X"AA",X"AB",X"FA",X"FA",
		X"0A",X"AF",X"0B",X"FF",X"0C",X"FF",X"00",X"BB",X"00",X"CA",X"00",X"AA",X"00",X"AA",X"00",X"CA",
		X"FA",X"FF",X"AA",X"CF",X"AC",X"44",X"CC",X"CC",X"AA",X"B4",X"AA",X"44",X"AA",X"C4",X"AB",X"0C",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FC",X"00",X"CC",X"0F",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FC",X"FF",X"FC",X"CF",X"FC",X"CF",
		X"0F",X"CC",X"0F",X"FF",X"00",X"EF",X"00",X"EE",X"0C",X"CC",X"0C",X"CC",X"00",X"CF",X"00",X"FF",
		X"FF",X"CF",X"FF",X"FF",X"CF",X"EE",X"FE",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"FC",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FC",X"00",X"CC",X"0F",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FC",X"FF",X"FC",X"CF",X"FC",X"CF",
		X"0F",X"CC",X"0F",X"FF",X"00",X"EF",X"00",X"EE",X"0C",X"CC",X"00",X"CC",X"00",X"CF",X"0C",X"CF",
		X"FF",X"CF",X"FF",X"FF",X"CF",X"EE",X"FE",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"FC",
		X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FC",X"00",X"CC",X"0F",X"CC",X"0F",X"CC",
		X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FC",X"FF",X"FC",X"CF",X"FC",X"CF",X"FF",X"CF",
		X"0F",X"FF",X"00",X"EF",X"00",X"EE",X"00",X"CC",X"0C",X"CC",X"00",X"CF",X"00",X"CF",X"0C",X"CC",
		X"FF",X"FF",X"CF",X"EE",X"CC",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",
		X"00",X"00",X"00",X"C0",X"0C",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"CC",X"0F",X"CC",X"FF",X"CB",
		X"00",X"00",X"00",X"C0",X"0C",X"CC",X"0C",X"CC",X"FF",X"CC",X"CC",X"F0",X"CC",X"FF",X"CB",X"FF",
		X"FF",X"CC",X"FF",X"FF",X"0E",X"FF",X"00",X"EE",X"0C",X"CF",X"CC",X"CF",X"00",X"FF",X"00",X"FF",
		X"FC",X"FF",X"FF",X"FE",X"FF",X"EE",X"CE",X"00",X"FF",X"CC",X"FF",X"CC",X"FF",X"C0",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FC",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FC",X"FF",X"FC",X"CF",
		X"0F",X"CC",X"0F",X"CC",X"0F",X"FF",X"00",X"EF",X"00",X"EE",X"00",X"CC",X"00",X"CC",X"00",X"CC",
		X"FB",X"CF",X"FF",X"CF",X"FF",X"FF",X"CF",X"EE",X"FE",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"C0",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FC",X"00",X"CC",X"0F",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FC",X"FF",X"FC",X"CF",X"FC",X"CF",
		X"0F",X"CC",X"0F",X"FF",X"00",X"EF",X"00",X"EE",X"00",X"CC",X"00",X"CC",X"00",X"CF",X"00",X"FF",
		X"FF",X"CF",X"FF",X"FF",X"CF",X"EE",X"CC",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"FC",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FF",X"00",X"FC",X"0F",X"FC",
		X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"CF",X"CF",X"CF",X"CC",X"CF",X"CC",
		X"0F",X"FC",X"0F",X"FF",X"00",X"CF",X"00",X"CE",X"00",X"CC",X"00",X"CC",X"00",X"CF",X"00",X"FF",
		X"FF",X"CC",X"FF",X"FF",X"FC",X"EE",X"CC",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"00",X"CF",X"00",X"FF",X"0F",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FF",X"FC",X"CF",X"CF",X"CF",X"CC",
		X"0F",X"FC",X"0F",X"FC",X"00",X"FF",X"00",X"EE",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"FC",
		X"CF",X"CC",X"FF",X"CC",X"FC",X"EE",X"EF",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"FC",
		X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CF",X"00",X"FC",X"00",X"CC",X"0F",X"CC",X"0F",X"CC",
		X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"CC",X"FC",X"FF",X"FC",X"CF",X"FC",X"CF",X"FF",X"CF",
		X"0F",X"FF",X"00",X"EF",X"0C",X"EE",X"00",X"CC",X"00",X"CC",X"00",X"CF",X"00",X"CF",X"0C",X"CC",
		X"CF",X"FF",X"CC",X"EE",X"EE",X"E0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CF",X"0C",X"FC",X"00",X"CC",X"0F",X"FF",X"0F",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"CC",X"FB",X"FF",X"FF",X"CF",X"CF",X"FF",X"CC",X"FF",
		X"0F",X"FF",X"00",X"EE",X"0C",X"EF",X"00",X"CF",X"00",X"FF",X"00",X"CF",X"0C",X"CC",X"00",X"00",
		X"CC",X"FF",X"FF",X"EE",X"FF",X"E0",X"FF",X"CC",X"FF",X"FF",X"FF",X"CC",X"FF",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"0F",X"FE",X"00",X"EF",X"0C",X"CC",X"00",X"CF",X"00",X"CF",X"00",X"CC",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"CC",X"FF",X"C0",X"FF",X"CC",X"CC",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FC",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"0F",X"FE",X"0C",X"EF",X"00",X"CC",X"00",X"CF",X"00",X"CF",X"00",X"CC",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"CC",X"FF",X"C0",X"CC",X"CC",X"CC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"FC",
		X"0C",X"FF",X"0F",X"FF",X"0F",X"FF",X"00",X"FC",X"0C",X"EE",X"0C",X"CC",X"0C",X"FF",X"00",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"FF",X"CC",X"FF",X"EC",X"FC",X"CC",X"CF",X"FF",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",
		X"00",X"EC",X"00",X"EE",X"00",X"EE",X"00",X"DE",X"00",X"ED",X"00",X"EE",X"00",X"EF",X"00",X"EF",
		X"CE",X"ED",X"CE",X"DD",X"CE",X"DC",X"DE",X"C0",X"ED",X"DC",X"FF",X"DD",X"FF",X"CD",X"FF",X"DC",
		X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"CE",X"00",X"CE",
		X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EC",X"ED",X"EC",X"ED",
		X"00",X"EE",X"00",X"EE",X"00",X"DE",X"0E",X"ED",X"00",X"EE",X"00",X"EF",X"00",X"EF",X"00",X"EE",
		X"EE",X"DD",X"EE",X"DC",X"EE",X"C0",X"DD",X"DC",X"FF",X"DD",X"FF",X"CC",X"FF",X"C0",X"FF",X"DC",
		X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"EC",X"00",X"EC",
		X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",X"CE",X"ED",
		X"00",X"EE",X"00",X"EE",X"00",X"DE",X"0E",X"ED",X"0C",X"EE",X"00",X"EF",X"00",X"EF",X"00",X"EE",
		X"CE",X"DD",X"CE",X"DC",X"DE",X"C0",X"ED",X"DD",X"FF",X"DC",X"FF",X"C0",X"FF",X"C0",X"FF",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"DE",X"00",X"ED",X"00",X"EE",X"0E",X"EF",X"0C",X"EF",
		X"CC",X"ED",X"CC",X"DD",X"CC",X"DC",X"DD",X"C0",X"EE",X"DD",X"FF",X"DC",X"FF",X"C0",X"FF",X"CD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"EE",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",
		X"00",X"EC",X"00",X"EC",X"00",X"EE",X"00",X"DE",X"00",X"ED",X"00",X"EE",X"00",X"EF",X"00",X"CF",
		X"EE",X"ED",X"CE",X"DD",X"CE",X"DC",X"DE",X"C0",X"ED",X"DC",X"FF",X"DD",X"FF",X"CD",X"FF",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",
		X"00",X"EC",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"CD",X"00",X"EE",X"00",X"EF",X"00",X"EF",
		X"CE",X"ED",X"CE",X"DD",X"CE",X"DC",X"DE",X"C0",X"ED",X"DC",X"FF",X"DD",X"FF",X"CD",X"FF",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"0E",X"EE",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"CE",X"00",X"CD",X"00",X"EE",X"00",X"EF",X"00",X"EF",
		X"CC",X"ED",X"CC",X"DD",X"CC",X"DC",X"DE",X"C0",X"ED",X"DC",X"FF",X"DD",X"FF",X"CD",X"FF",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"EE",X"DE",X"EE",X"DD",X"EE",X"DD",X"EE",X"ED",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"ED",X"00",X"EE",X"00",X"EE",X"00",X"CC",
		X"EE",X"ED",X"CC",X"DD",X"CC",X"DC",X"CC",X"C0",X"ED",X"DD",X"FF",X"DD",X"FF",X"CC",X"FF",X"DC",
		X"00",X"EC",X"00",X"DE",X"0E",X"DE",X"0E",X"EF",X"0E",X"CC",X"00",X"FF",X"00",X"EE",X"00",X"EE",
		X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EF",X"DD",X"EF",X"ED",X"CE",X"FD",X"CE",X"FF",X"CE",X"DD",
		X"00",X"EE",X"0E",X"DD",X"0C",X"EE",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"CE",X"00",X"0C",
		X"DE",X"DC",X"DD",X"CD",X"FF",X"DD",X"FF",X"DC",X"FF",X"C0",X"FF",X"DD",X"FF",X"CC",X"CC",X"00",
		X"00",X"0F",X"00",X"00",X"F0",X"EE",X"00",X"CF",X"0E",X"FE",X"0E",X"EE",X"00",X"EE",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"CE",X"DE",X"CC",X"ED",X"EE",X"ED",X"CC",X"ED",X"DD",X"ED",
		X"00",X"ED",X"00",X"DE",X"0E",X"EF",X"0C",X"EF",X"00",X"EF",X"00",X"EE",X"00",X"CE",X"00",X"0C",
		X"EE",X"DD",X"FF",X"DC",X"FF",X"CD",X"FF",X"DD",X"FF",X"CC",X"FF",X"DD",X"EE",X"CC",X"DC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"ED",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"CE",X"C0",X"EE",X"DC",X"EE",X"ED",X"DD",X"ED",X"EE",X"ED",
		X"00",X"DE",X"00",X"DF",X"0E",X"EF",X"0C",X"EF",X"00",X"EE",X"00",X"EE",X"00",X"CE",X"00",X"0C",
		X"FF",X"DD",X"FF",X"DC",X"FF",X"CD",X"FF",X"DC",X"FF",X"CD",X"EE",X"DD",X"EE",X"CC",X"DC",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"CE",X"C0",X"EE",X"DC",X"CE",X"ED",X"DD",X"ED",
		X"00",X"ED",X"00",X"DE",X"00",X"DF",X"00",X"EF",X"00",X"EE",X"00",X"EE",X"00",X"CE",X"00",X"0C",
		X"EE",X"ED",X"FF",X"DD",X"FF",X"DC",X"FF",X"CD",X"FF",X"DD",X"EE",X"DD",X"EE",X"CC",X"DC",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"EE",X"00",X"DE",X"0E",X"DE",X"0E",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"EE",X"DE",X"EE",X"DD",X"EE",X"DD",
		X"00",X"EE",X"00",X"EF",X"00",X"FC",X"0E",X"FE",X"0E",X"EE",X"0C",X"ED",X"00",X"EE",X"00",X"EF",
		X"EF",X"ED",X"FF",X"ED",X"FF",X"DD",X"CF",X"FC",X"CE",X"CD",X"ED",X"DD",X"FF",X"DC",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",X"0B",X"BC",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",
		X"BB",X"BB",X"BB",X"BB",X"0B",X"BC",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"CC",X"00",X"BB",
		X"CB",X"B4",X"FB",X"44",X"FC",X"44",X"CF",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FC",X"44",
		X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",X"0B",X"BC",X"BB",X"BB",
		X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",X"CB",X"B4",
		X"BB",X"BB",X"0B",X"BC",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"0B",X"CF",X"0C",X"CF",X"00",X"0C",
		X"FB",X"44",X"FC",X"44",X"CF",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"44",X"FF",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BC",X"0B",X"BC",X"BB",X"BB",
		X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",X"CB",X"B4",
		X"BB",X"BB",X"0B",X"BC",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"CF",X"00",X"CF",X"00",X"0C",
		X"FB",X"44",X"FC",X"44",X"CF",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"CC",X"FF",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BC",X"0B",X"BC",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",
		X"BB",X"BB",X"BB",X"BB",X"0B",X"BC",X"00",X"CF",X"00",X"FF",X"0B",X"FF",X"00",X"FF",X"00",X"CF",
		X"CB",X"B4",X"FB",X"44",X"FC",X"44",X"CF",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"BC",
		X"0B",X"BB",X"BB",X"BC",X"BB",X"BB",X"0B",X"CC",X"00",X"CF",X"00",X"FF",X"00",X"BF",X"00",X"BB",
		X"BB",X"B4",X"BB",X"B4",X"CB",X"44",X"FC",X"44",X"CC",X"CC",X"FF",X"44",X"FF",X"44",X"FF",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",X"0B",X"BC",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",
		X"BB",X"BB",X"BB",X"BB",X"0B",X"CC",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"CB",X"B4",X"FB",X"44",X"FC",X"44",X"CF",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FC",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",
		X"BB",X"BB",X"BB",X"BB",X"0B",X"CC",X"00",X"CB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"FF",
		X"CC",X"B4",X"FF",X"44",X"FF",X"44",X"CC",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FC",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"BB",X"B4",X"BB",X"B4",
		X"BB",X"BB",X"BB",X"BB",X"0B",X"BC",X"00",X"CF",X"00",X"FF",X"00",X"BF",X"00",X"BB",X"00",X"CB",
		X"CC",X"B4",X"FF",X"44",X"FF",X"44",X"CC",X"CC",X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FC",X"44",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"0B",X"FF",X"00",X"FF",X"0B",X"BB",X"0B",X"BB",X"BB",X"BF",
		X"00",X"00",X"BB",X"C0",X"BF",X"F0",X"BF",X"44",X"CB",X"44",X"FB",X"B4",X"FC",X"B4",X"CF",X"B4",
		X"BB",X"FF",X"0C",X"FF",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"0B",X"BF",X"0B",X"BF",X"00",X"BB",
		X"FF",X"44",X"FF",X"CC",X"FF",X"44",X"FF",X"44",X"FF",X"CC",X"FF",X"C0",X"FF",X"44",X"FF",X"44",
		X"00",X"00",X"00",X"00",X"00",X"CF",X"00",X"FB",X"0B",X"BF",X"00",X"FF",X"0B",X"FF",X"0B",X"FF",
		X"00",X"00",X"00",X"00",X"FB",X"00",X"FF",X"00",X"FF",X"44",X"FF",X"44",X"FF",X"F4",X"FF",X"FF",
		X"BB",X"FF",X"BB",X"FF",X"0B",X"FF",X"00",X"CF",X"00",X"FF",X"0B",X"BF",X"0B",X"BF",X"00",X"CC",
		X"FF",X"FF",X"FF",X"F4",X"FF",X"CC",X"FF",X"44",X"FF",X"44",X"FF",X"CC",X"FF",X"44",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"FC",
		X"0B",X"FF",X"BF",X"FF",X"BB",X"FF",X"CB",X"FF",X"0C",X"CF",X"0B",X"FF",X"0B",X"BF",X"0C",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"FF",X"44",X"FF",X"CC",X"FB",X"44",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"FC",X"FF",X"FF",
		X"0B",X"FF",X"BB",X"FF",X"BB",X"FF",X"CB",X"FF",X"0C",X"CF",X"00",X"FF",X"00",X"BF",X"00",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"FF",X"44",X"FF",X"44",X"FF",X"C4",X"FF",X"44",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"0B",X"BB",X"0C",X"BB",X"0B",X"FF",X"0B",X"CF",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"BF",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BB",X"FF",X"BB",X"BB",X"CB",X"CC",X"0C",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"BF",X"0B",X"CF",
		X"BF",X"FF",X"CB",X"4F",X"FC",X"44",X"CC",X"CC",X"FF",X"44",X"FF",X"44",X"FF",X"4C",X"FF",X"44",
		X"00",X"00",X"00",X"A0",X"AA",X"BA",X"A4",X"FF",X"CA",X"FF",X"0A",X"FC",X"AA",X"CF",X"AA",X"AA",
		X"00",X"00",X"00",X"AC",X"0A",X"BA",X"FF",X"BB",X"FF",X"AB",X"CC",X"AA",X"AF",X"FA",X"AA",X"AA",
		X"AA",X"AC",X"CB",X"AC",X"AA",X"BB",X"CA",X"AA",X"0C",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AC",
		X"CC",X"A4",X"CC",X"44",X"C4",X"C4",X"AB",X"44",X"AA",X"4C",X"AB",X"CC",X"B4",X"00",X"CB",X"00",
		X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CF",X"00",X"FC",X"00",X"CC",X"0F",X"CB",X"0F",X"CC",
		X"00",X"C0",X"0C",X"CC",X"0C",X"CC",X"FF",X"CC",X"FC",X"FF",X"FB",X"CF",X"FC",X"CF",X"FF",X"CF",
		X"0F",X"FF",X"00",X"EF",X"0C",X"EE",X"00",X"CC",X"00",X"CF",X"00",X"FF",X"0C",X"FF",X"00",X"CC",
		X"CF",X"FF",X"CC",X"EE",X"CC",X"E0",X"EE",X"CC",X"FF",X"CC",X"FF",X"FC",X"EF",X"F0",X"FF",X"CC",
		X"00",X"00",X"00",X"EC",X"00",X"DE",X"0E",X"EE",X"0E",X"EE",X"0E",X"CC",X"0C",X"CE",X"00",X"EE",
		X"00",X"00",X"00",X"EC",X"00",X"DE",X"EE",X"DD",X"EE",X"ED",X"EE",X"ED",X"CE",X"ED",X"CE",X"ED",
		X"00",X"EE",X"00",X"EE",X"0E",X"DE",X"0C",X"ED",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"EF",
		X"DD",X"DD",X"CE",X"DC",X"DE",X"C0",X"FF",X"DD",X"FF",X"DC",X"FF",X"C0",X"FF",X"C0",X"FF",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"0B",X"BB",X"0C",X"CC",X"0B",X"CB",X"0B",X"BB",X"BB",X"BC",
		X"00",X"00",X"B4",X"00",X"BB",X"C0",X"BB",X"44",X"BB",X"44",X"CB",X"44",X"FB",X"44",X"FC",X"44",
		X"BB",X"FF",X"CC",X"FF",X"0B",X"FF",X"0B",X"FF",X"0C",X"FF",X"0B",X"FF",X"0B",X"BF",X"0B",X"BB",
		X"CC",X"44",X"CE",X"EC",X"FF",X"C4",X"FF",X"E4",X"FF",X"EC",X"FF",X"E4",X"FF",X"C4",X"FF",X"44",
		X"00",X"03",X"00",X"3C",X"03",X"FF",X"03",X"CC",X"3C",X"CC",X"3C",X"CC",X"3C",X"CC",X"03",X"CC",
		X"30",X"00",X"C3",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"30",X"C4",X"20",X"CC",X"C2",X"CC",X"C2",
		X"03",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CF",X"CC",X"CC",X"CC",X"3C",X"C2",X"02",X"20",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"3C",X"00",X"FF",X"03",X"CA",X"03",X"CC",X"3C",X"CC",X"2C",X"CC",X"3C",X"CC",
		X"33",X"00",X"CC",X"00",X"CC",X"20",X"CC",X"C3",X"CC",X"CC",X"CC",X"FC",X"CC",X"CC",X"CC",X"CC",
		X"02",X"9C",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"CC",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"CC",X"03",X"FF",X"03",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"20",X"23",X"C3",X"CC",X"CC",X"CC",X"4C",X"CC",X"CC",X"5C",X"CC",
		X"3C",X"CC",X"3C",X"AC",X"3C",X"CC",X"3C",X"CC",X"03",X"CC",X"02",X"C9",X"00",X"CC",X"00",X"22",
		X"CC",X"C2",X"CC",X"C2",X"CC",X"20",X"CC",X"20",X"CC",X"00",X"CC",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"FF",X"FF",X"AA",X"FF",X"CA",X"AF",
		X"C0",X"00",X"AC",X"00",X"AC",X"00",X"AA",X"00",X"AA",X"00",X"AF",X"FF",X"FF",X"AA",X"FF",X"AA",
		X"0C",X"FF",X"00",X"FF",X"00",X"FA",X"00",X"AA",X"00",X"AA",X"00",X"AC",X"00",X"C0",X"00",X"00",
		X"AA",X"AC",X"AA",X"C0",X"FA",X"C0",X"FF",X"AC",X"CF",X"AC",X"0C",X"AC",X"00",X"C0",X"00",X"00",
		X"00",X"BB",X"00",X"FB",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0F",X"BF",
		X"00",X"00",X"00",X"BC",X"CF",X"BC",X"FF",X"BC",X"FB",X"C0",X"BB",X"C0",X"FF",X"C0",X"FF",X"BC",
		X"FF",X"BF",X"BB",X"BF",X"CC",X"FF",X"00",X"CF",X"00",X"0F",X"00",X"0F",X"00",X"0C",X"00",X"00",
		X"BF",X"FF",X"BB",X"FF",X"BB",X"BB",X"BB",X"CC",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AB",X"00",X"AA",X"BB",X"CA",X"BB",X"0A",X"AB",X"0C",X"AA",X"00",X"AA",
		X"AA",X"00",X"AB",X"00",X"AB",X"00",X"BB",X"00",X"BB",X"C0",X"BB",X"BB",X"AA",X"BB",X"BA",X"AA",
		X"00",X"AB",X"00",X"BB",X"0A",X"BB",X"0A",X"BC",X"0B",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"AA",X"AB",X"CC",X"AB",X"00",X"AA",X"C0",X"AA",X"C0",X"CA",X"C0",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"0C",X"00",X"0A",X"00",X"AF",X"00",X"CC",
		X"88",X"BB",X"CC",X"CC",X"99",X"0B",X"9C",X"77",X"C6",X"F7",X"6F",X"C7",X"66",X"CC",X"C5",X"F9",
		X"00",X"99",X"00",X"F9",X"00",X"99",X"06",X"88",X"6F",X"CC",X"66",X"C7",X"C5",X"C7",X"0C",X"0C",
		X"7C",X"99",X"3C",X"C8",X"CA",X"BC",X"CA",X"BC",X"CC",X"C3",X"3C",X"C3",X"3C",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"65",X"00",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"6F",X"00",X"61",X"00",X"66",X"00",X"06",X"00",X"00",
		X"00",X"00",X"60",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"55",X"00",X"55",X"00",X"5C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"6F",X"00",X"61",X"00",X"66",X"00",X"66",X"00",X"06",X"00",X"00",
		X"65",X"00",X"66",X"00",X"66",X"C0",X"66",X"C0",X"66",X"C0",X"65",X"C0",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",
		X"00",X"6F",X"00",X"F1",X"00",X"F1",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"05",
		X"66",X"00",X"66",X"C0",X"66",X"C0",X"65",X"C0",X"65",X"C0",X"55",X"C0",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",
		X"00",X"6F",X"00",X"6F",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"55",X"00",X"00",
		X"66",X"C0",X"66",X"5C",X"66",X"5C",X"66",X"5C",X"65",X"5C",X"55",X"C0",X"55",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"F1",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"66",X"C0",
		X"00",X"F1",X"00",X"16",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"55",X"00",X"05",
		X"66",X"5C",X"66",X"5C",X"66",X"5C",X"65",X"5C",X"55",X"5C",X"55",X"C0",X"55",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"66",X"5C",X"66",X"5C",
		X"00",X"11",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"55",X"00",X"00",
		X"66",X"55",X"66",X"55",X"66",X"55",X"66",X"55",X"66",X"5C",X"55",X"5C",X"55",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"F1",X"00",X"F1",X"06",X"16",
		X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"C0",X"66",X"5C",X"66",X"5C",X"66",X"55",
		X"06",X"16",X"06",X"66",X"06",X"66",X"06",X"66",X"00",X"66",X"00",X"66",X"00",X"55",X"00",X"05",
		X"66",X"55",X"66",X"55",X"66",X"55",X"65",X"55",X"55",X"5C",X"55",X"5C",X"55",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"00",X"FF",X"00",X"F1",X"00",X"F6",X"06",X"16",
		X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"66",X"5C",X"66",X"55",X"66",X"55",X"66",X"55",
		X"06",X"66",X"06",X"66",X"06",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"55",X"00",X"00",
		X"66",X"55",X"66",X"55",X"66",X"55",X"66",X"55",X"65",X"55",X"55",X"5C",X"55",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"06",X"00",X"F1",X"00",X"F1",X"06",X"16",X"06",X"66",X"6F",X"66",X"61",X"66",
		X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"5C",X"66",X"55",X"66",X"55",X"66",X"55",X"66",X"55",
		X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"66",X"05",X"66",X"00",X"55",X"00",X"55",X"00",X"05",
		X"66",X"55",X"66",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"5C",X"55",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"00",X"CB",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"CF",X"00",X"CF",X"00",X"CC",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"CC",X"00",X"CB",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"00",X"C1",X"00",X"C1",X"00",X"CC",X"00",X"CC",X"00",X"0C",X"00",X"00",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"B0",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"CF",X"00",X"F1",X"00",X"F1",X"00",X"C1",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"0C",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CB",X"00",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",
		X"00",X"CF",X"00",X"CF",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",
		X"CC",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"C0",X"CC",X"C0",X"CC",X"B0",X"CC",X"0B",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"CF",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"00",X"F1",X"00",X"C1",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"0C",
		X"CC",X"C0",X"CC",X"C0",X"CC",X"CB",X"CC",X"C0",X"CC",X"C0",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CF",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"BB",X"CC",X"B0",X"CC",X"C0",X"CC",X"C0",
		X"00",X"FC",X"00",X"1C",X"00",X"1C",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"C0",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"CF",X"00",X"F1",X"00",X"F1",X"0C",X"1C",
		X"00",X"00",X"00",X"B0",X"00",X"B0",X"CC",X"00",X"CC",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"CC",
		X"0C",X"1C",X"0C",X"CC",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"0C",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"C0",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CF",X"00",X"FF",X"00",X"F1",X"0C",X"F1",
		X"00",X"00",X"00",X"00",X"CC",X"B0",X"CC",X"B0",X"CC",X"C0",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"0C",X"1C",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"0C",X"00",X"CC",X"00",X"F1",X"0C",X"FC",X"0C",X"1C",X"CC",X"1C",X"CC",X"CC",
		X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CB",X"CC",X"BB",X"CC",X"BC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"0C",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"11",X"01",X"11",X"01",X"11",X"01",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"11",X"1C",X"11",X"1C",X"11",X"1C",X"11",X"1C",
		X"01",X"11",X"01",X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"1C",X"11",X"1C",X"1C",X"11",X"CC",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"65",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"CC",X"1C",X"C0",X"1C",X"C0",X"1C",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"C1",X"C1",X"01",X"C1",X"01",X"C1",X"01",
		X"1C",X"C0",X"1C",X"C0",X"CC",X"11",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"01",X"C1",X"01",X"C0",X"11",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"01",X"C1",X"01",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"C1",X"C1",X"C1",X"C1",
		X"01",X"C1",X"01",X"11",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"C1",X"11",X"11",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"0C",X"1C",X"11",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"0C",X"1C",X"01",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"1C",X"1C",
		X"00",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"1C",X"10",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"1C",X"1C",
		X"11",X"1C",X"0C",X"11",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"11",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"1C",X"1C",
		X"0C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"11",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"0C",X"1C",X"00",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1C",X"1C",X"1C",X"1C",
		X"00",X"1C",X"00",X"11",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"11",X"11",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BC",X"00",X"CC",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"22",X"0F",X"22",X"00",X"32",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"C0",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",X"23",X"22",X"23",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"00",X"F3",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"C0",X"33",X"22",X"33",X"33",X"33",X"33",X"33",X"33",
		X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"00",X"F3",X"00",X"FF",X"00",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"2C",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"32",X"C0",X"32",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B3",X"00",X"3F",X"00",X"FF",X"00",X"CF",X"00",X"0F",X"00",X"0F",X"00",X"0C",X"00",X"00",
		X"33",X"33",X"33",X"33",X"F3",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"E3",X"FF",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CC",X"FF",X"BB",X"BB",X"CB",X"BB",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"22",X"33",X"32",X"CC",X"32",X"CC",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"E3",X"33",X"EE",X"33",X"EE",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"00",X"2C",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"B3",X"0C",X"BF",X"00",X"CF",X"00",X"0F",X"00",X"0F",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"FE",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"E3",X"FF",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CC",X"FE",X"BB",X"BB",X"CB",X"BB",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"23",X"22",X"32",X"22",X"33",X"32",X"CC",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"E3",X"33",X"EE",X"33",X"EC",X"C3",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"00",X"2C",X"00",X"2C",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"03",X"33",X"33",X"C3",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"03",X"00",X"B3",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"23",X"C3",X"23",X"0C",X"C2",X"00",X"C2",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"22",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"32",X"CC",X"2C",X"00",X"C0",X"00",
		X"00",X"00",X"C0",X"00",X"BC",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3F",X"00",X"FF",X"00",X"F3",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"FF",X"00",X"FF",X"00",X"CF",X"00",X"BF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"3C",
		X"00",X"CA",X"00",X"A4",X"0C",X"FF",X"CA",X"FF",X"CA",X"CA",X"CA",X"CA",X"0C",X"CC",X"AA",X"CC",
		X"C0",X"00",X"AC",X"00",X"AC",X"00",X"FC",X"C0",X"AA",X"AC",X"AF",X"4A",X"AF",X"4A",X"AF",X"4A",
		X"CA",X"BC",X"AA",X"BB",X"AA",X"AB",X"AA",X"AA",X"AA",X"BB",X"CB",X"BC",X"BC",X"BC",X"C0",X"BB",
		X"AA",X"AA",X"CC",X"BC",X"CC",X"BC",X"BC",X"C0",X"BB",X"00",X"CC",X"00",X"B0",X"00",X"C0",X"00",
		X"00",X"33",X"00",X"33",X"03",X"CC",X"33",X"33",X"CC",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"C3",X"00",X"03",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"C3",X"33",X"0C",X"32",X"00",X"C2",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"22",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BC",X"32",X"C0",X"22",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"00",X"FF",X"0F",X"CC",X"0F",X"CC",X"CF",X"FC",X"C0",X"FF",X"CC",X"CC",
		X"C0",X"00",X"CC",X"00",X"C0",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"CC",X"CC",X"CC",X"CB",X"CC",
		X"CC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"CC",X"CE",X"C0",X"C0",X"00",X"CC",
		X"CC",X"C0",X"FC",X"E0",X"FF",X"E0",X"EF",X"00",X"EE",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"EE",X"00",X"EF",X"0C",X"EF",X"CC",X"EF",X"EC",X"EE",X"EC",X"EE",X"EE",X"EE",
		X"C0",X"00",X"CC",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"C0",X"CE",X"CC",X"CF",X"DD",X"EF",X"DD",
		X"EF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"CD",X"FD",X"CD",X"ED",X"CD",X"DC",
		X"EF",X"DD",X"EE",X"DD",X"DD",X"DD",X"DD",X"CC",X"CC",X"00",X"C0",X"00",X"DC",X"00",X"C0",X"00",
		X"DF",X"00",X"FF",X"00",X"FF",X"D0",X"CC",X"DD",X"CF",X"DF",X"CF",X"DF",X"CF",X"DF",X"CF",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"FD",X"00",X"FF",X"00",
		X"CF",X"DF",X"FC",X"DF",X"FF",X"DF",X"0F",X"DF",X"00",X"DF",X"00",X"DF",X"00",X"DF",X"00",X"EF",
		X"FF",X"F0",X"CF",X"F0",X"FC",X"F0",X"FC",X"F0",X"FC",X"F0",X"FC",X"F0",X"FC",X"F0",X"FC",X"F0",
		X"00",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"FF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"00",X"CF",X"00",X"CF",X"00",X"FF",X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"99",X"00",X"99",X"00",X"FF",X"EE",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"FF",X"00",X"FF",X"A0",
		X"00",X"EC",X"00",X"EC",X"00",X"EC",X"00",X"EC",X"DD",X"EC",X"ED",X"EC",X"CE",X"DD",X"0C",X"DD",
		X"CC",X"F0",X"FF",X"F0",X"FF",X"F0",X"0F",X"F0",X"00",X"F0",X"00",X"00",X"D0",X"00",X"DD",X"00",
		X"00",X"DD",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"0F",X"00",X"0C",X"F0",X"0C",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"F0",X"0C",X"F0",X"0F",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"FF",X"00",X"CC",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"CF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"CF",X"00",X"FC",X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FF",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"ED",X"DE",X"FE",
		X"AA",X"AC",X"AA",X"C0",X"CC",X"C0",X"CC",X"C0",X"FF",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FE",X"22",X"FF",X"2E",X"FD",X"FF",X"CD",X"EC",X"AA",X"CA",X"AA",X"AA",X"CC",X"CC",X"00",
		X"00",X"00",X"AC",X"00",X"AA",X"00",X"AA",X"00",X"AC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"32",X"FF",X"FF",X"FF",X"FF",X"11",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"EC",X"00",X"EE",X"C0",X"FE",X"E1",X"FF",X"1D",
		X"EE",X"11",X"CC",X"EE",X"00",X"32",X"0B",X"32",X"BB",X"FF",X"CB",X"B2",X"0C",X"BB",X"00",X"CC",
		X"11",X"CC",X"DE",X"00",X"CE",X"00",X"BF",X"00",X"FB",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"AA",X"00",X"CA",X"00",X"EC",
		X"00",X"FF",X"00",X"99",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"CA",X"AA",
		X"00",X"CE",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"AA",X"00",X"AA",X"00",X"CC",X"00",X"00",
		X"EC",X"CC",X"EE",X"EE",X"FC",X"EE",X"FA",X"32",X"FF",X"32",X"FC",X"FF",X"AA",X"CC",X"CA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"5F",X"FF",
		X"00",X"FF",X"FF",X"33",X"FF",X"33",X"33",X"FF",X"F3",X"32",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"33",X"C0",X"33",X"C0",X"FF",X"EE",X"22",X"EE",X"FE",X"FE",X"FF",X"FF",X"FF",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"EE",X"00",X"EE",X"C0",X"FE",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"5F",X"00",X"E5",X"00",X"CE",
		X"00",X"EE",X"00",X"33",X"FF",X"FF",X"FF",X"32",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"E5",X"55",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",
		X"EE",X"EE",X"CC",X"EE",X"FC",X"32",X"FC",X"32",X"FF",X"32",X"BE",X"FF",X"BB",X"32",X"CB",X"BB",
		X"EC",X"00",X"3F",X"00",X"F2",X"EC",X"2E",X"EE",X"FE",X"EE",X"FF",X"FE",X"FF",X"55",X"55",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"00",X"5C",X"00",X"DC",X"00",X"C0",X"00",
		X"EE",X"DC",X"DD",X"C0",X"22",X"CC",X"22",X"CB",X"2F",X"CB",X"FF",X"BB",X"CC",X"BB",X"BB",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"E5",X"55",X"CC",X"55",X"00",X"EE",X"00",X"CE",X"00",X"0E",X"00",X"0E",X"00",X"0E",
		X"FF",X"FF",X"5F",X"FF",X"55",X"55",X"E5",X"55",X"EE",X"EE",X"EE",X"EE",X"C3",X"EE",X"F3",X"32",
		X"00",X"FE",X"00",X"FF",X"00",X"CE",X"00",X"BE",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",
		X"C3",X"32",X"B3",X"32",X"FF",X"32",X"FF",X"FF",X"CC",X"FF",X"BB",X"CC",X"BB",X"BB",X"CC",X"CC",
		X"FF",X"FE",X"FF",X"55",X"55",X"55",X"55",X"ED",X"ED",X"DE",X"DE",X"CE",X"ED",X"0E",X"22",X"FE",
		X"55",X"50",X"55",X"C0",X"DD",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"FE",X"22",X"FF",X"2E",X"FE",X"FF",X"CE",X"EC",X"BB",X"CB",X"BB",X"BB",X"CC",X"CC",X"00",
		X"00",X"00",X"BC",X"00",X"BB",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"A4",X"A0",X"4B",X"A0",X"AB",X"AA",X"CA",X"FF",X"AA",X"FF",X"AA",X"CC",
		X"00",X"00",X"0A",X"C0",X"A4",X"AC",X"A4",X"BA",X"AA",X"AA",X"FF",X"CC",X"FF",X"AC",X"CF",X"A4",
		X"AA",X"CA",X"AA",X"AA",X"BB",X"AA",X"CC",X"BB",X"00",X"AA",X"0A",X"AA",X"AA",X"AA",X"CC",X"AA",
		X"CF",X"A4",X"AA",X"B4",X"AA",X"4C",X"BB",X"C0",X"BB",X"00",X"AB",X"C0",X"B4",X"BC",X"4C",X"C0",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"A4",X"A0",X"BB",X"AA",X"CA",X"FF",X"AA",X"FF",X"AA",X"CC",
		X"00",X"00",X"00",X"00",X"0A",X"C0",X"A4",X"AA",X"A4",X"BA",X"FF",X"CC",X"FF",X"AC",X"CF",X"A4",
		X"AA",X"CA",X"AA",X"AA",X"BB",X"AA",X"CC",X"BC",X"AA",X"AA",X"CA",X"AA",X"0C",X"AA",X"0A",X"AA",
		X"CF",X"A4",X"AA",X"44",X"AA",X"4C",X"44",X"C0",X"BB",X"00",X"AB",X"C0",X"B4",X"4C",X"4C",X"C0",
		X"AA",X"00",X"44",X"00",X"4B",X"00",X"BB",X"AA",X"AA",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"AA",
		X"AA",X"00",X"44",X"C0",X"4B",X"AC",X"AB",X"AC",X"FA",X"C0",X"FF",X"C0",X"FF",X"4C",X"CF",X"4C",
		X"AA",X"AA",X"BB",X"AC",X"CC",X"CC",X"AA",X"AA",X"AA",X"AA",X"CC",X"AA",X"00",X"AA",X"0A",X"CC",
		X"AA",X"4C",X"A4",X"C0",X"4C",X"00",X"BB",X"00",X"B4",X"C0",X"4C",X"00",X"C0",X"00",X"4C",X"00",
		X"00",X"00",X"AA",X"00",X"44",X"00",X"4B",X"00",X"BB",X"AA",X"AA",X"FA",X"AF",X"FA",X"AF",X"CA",
		X"00",X"00",X"AA",X"00",X"44",X"C0",X"4B",X"AC",X"AB",X"AC",X"FA",X"C0",X"FF",X"C0",X"FF",X"4C",
		X"AF",X"AA",X"AA",X"AA",X"BB",X"AC",X"CC",X"BA",X"0A",X"AA",X"AA",X"AA",X"AC",X"AA",X"C0",X"AA",
		X"FF",X"4C",X"AA",X"4C",X"A4",X"C0",X"4C",X"00",X"BB",X"C0",X"B4",X"00",X"4C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"44",X"A0",X"AB",X"AA",X"CA",X"FF",X"AA",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AC",X"A4",X"BA",X"AA",X"AA",X"FF",X"CC",X"FF",X"AC",
		X"AA",X"FF",X"AA",X"CC",X"AA",X"AA",X"BB",X"AA",X"CC",X"BB",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"FF",X"A4",X"CF",X"A4",X"AA",X"44",X"AA",X"4C",X"44",X"C0",X"BB",X"C0",X"AB",X"C0",X"BC",X"C0",
		X"00",X"00",X"0A",X"00",X"A4",X"A0",X"44",X"A0",X"AB",X"AA",X"CA",X"FF",X"AA",X"FF",X"AA",X"FF",
		X"00",X"00",X"0A",X"C0",X"A4",X"AC",X"A4",X"BA",X"AA",X"AA",X"FF",X"CC",X"FF",X"AC",X"FF",X"A4",
		X"AA",X"FA",X"AA",X"AA",X"BB",X"AA",X"AA",X"BB",X"CA",X"AA",X"0C",X"AA",X"00",X"AA",X"00",X"AA",
		X"FC",X"A4",X"AA",X"44",X"AA",X"4C",X"44",X"C0",X"BB",X"00",X"AB",X"C0",X"B4",X"4C",X"44",X"C0",
		X"00",X"00",X"0A",X"00",X"A4",X"A0",X"44",X"A0",X"AB",X"AA",X"CA",X"FF",X"AA",X"FF",X"AA",X"CC",
		X"00",X"00",X"0A",X"C0",X"A4",X"AC",X"A4",X"BA",X"AA",X"AA",X"FF",X"CC",X"FF",X"AC",X"FC",X"A4",
		X"AA",X"FC",X"AA",X"AA",X"BB",X"AA",X"CA",X"BB",X"0A",X"AA",X"0C",X"AA",X"00",X"AA",X"00",X"AA",
		X"AC",X"A4",X"AA",X"44",X"AA",X"4C",X"44",X"C0",X"BB",X"C0",X"AB",X"44",X"B4",X"4C",X"44",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"4C",X"A4",X"AA",X"44",X"AA",X"AA",X"FF",X"AA",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"C0",X"A4",X"AC",X"AA",X"BA",X"FF",X"AC",X"FF",X"A4",
		X"AA",X"CC",X"AA",X"FC",X"BB",X"AA",X"CC",X"BB",X"00",X"AA",X"0A",X"AA",X"0A",X"AA",X"0C",X"AA",
		X"FC",X"A4",X"AC",X"44",X"AA",X"4C",X"C4",X"C0",X"BB",X"4C",X"AB",X"C0",X"A4",X"00",X"B4",X"00",
		X"00",X"00",X"0A",X"00",X"A4",X"A0",X"BB",X"AA",X"AA",X"CC",X"AA",X"FF",X"AF",X"FA",X"AA",X"AC",
		X"00",X"00",X"0A",X"00",X"A4",X"A0",X"AA",X"4A",X"CF",X"AC",X"FF",X"AC",X"FF",X"A4",X"AA",X"44",
		X"BB",X"CC",X"CC",X"44",X"AA",X"AA",X"CA",X"AA",X"0C",X"AA",X"0A",X"AA",X"0A",X"AA",X"0C",X"CC",
		X"CA",X"4C",X"44",X"C0",X"BB",X"4C",X"BB",X"C0",X"AB",X"00",X"B4",X"C0",X"4C",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"FA",X"AF",X"AA",X"AA",X"AC",X"AA",X"CC",X"AA",X"CC",X"AA",X"AA",
		X"00",X"00",X"CF",X"00",X"FF",X"00",X"AA",X"4C",X"AC",X"4C",X"CC",X"44",X"CB",X"44",X"BB",X"4C",
		X"BB",X"AB",X"BB",X"AA",X"BB",X"AA",X"CB",X"AA",X"0C",X"AA",X"00",X"AA",X"00",X"CB",X"00",X"0C",
		X"B4",X"BC",X"B4",X"BC",X"BB",X"BC",X"AB",X"C0",X"B4",X"00",X"4C",X"00",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"0A",X"AC",X"AA",X"CA",X"AA",X"AB",X"AA",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"CB",X"BC",X"BB",X"BC",X"BB",X"C0",
		X"CA",X"AA",X"AC",X"AA",X"CA",X"AA",X"40",X"AA",X"40",X"AA",X"A4",X"BB",X"A4",X"CB",X"44",X"0C",
		X"CB",X"BB",X"4C",X"BC",X"44",X"C0",X"44",X"AC",X"4B",X"A4",X"4B",X"4C",X"CB",X"4C",X"0C",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"0A",X"CC",X"AA",X"AA",X"AA",X"AB",X"AA",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"CB",X"00",X"AC",X"B0",X"BB",X"B0",X"BB",X"C0",
		X"CA",X"AA",X"AC",X"AA",X"CA",X"AA",X"40",X"AA",X"40",X"AA",X"A4",X"BB",X"A4",X"CB",X"44",X"BC",
		X"CB",X"BB",X"4C",X"BC",X"44",X"C0",X"44",X"AC",X"4B",X"A4",X"4B",X"4C",X"CB",X"4C",X"0C",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AC",X"A4",X"AA",X"44",X"AA",X"A4",X"AA",X"AA",X"FF",
		X"10",X"00",X"00",X"00",X"00",X"01",X"AA",X"00",X"A4",X"A0",X"A4",X"BA",X"AA",X"BC",X"FF",X"A4",
		X"AA",X"FF",X"AA",X"CC",X"BA",X"AA",X"CC",X"BC",X"AA",X"AA",X"CA",X"AA",X"0C",X"AA",X"00",X"AA",
		X"FF",X"A4",X"AC",X"F4",X"AA",X"4C",X"C4",X"C0",X"AB",X"C0",X"AB",X"4C",X"B4",X"4C",X"BC",X"C0",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"CC",X"FF",X"CC",X"FF",X"BC",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"CC",X"00",X"CC",X"F0",X"BC",X"FE",
		X"FF",X"CF",X"FF",X"FF",X"EE",X"FF",X"00",X"EE",X"CC",X"FF",X"CC",X"FF",X"0C",X"FF",X"0C",X"FF",
		X"CC",X"FE",X"FF",X"EE",X"FF",X"E0",X"EE",X"00",X"FC",X"CC",X"FC",X"CC",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"CC",X"FF",X"CC",X"FF",X"BC",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"CC",X"00",X"CC",X"F0",X"BC",X"FE",
		X"FF",X"CF",X"FF",X"FF",X"EE",X"FF",X"00",X"EE",X"CC",X"FF",X"CC",X"FF",X"0C",X"FF",X"CC",X"FF",
		X"CC",X"FE",X"FF",X"EE",X"FF",X"E0",X"EE",X"00",X"FC",X"C0",X"FC",X"CC",X"FF",X"0C",X"FF",X"00",
		X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"CC",X"FF",X"CC",X"FF",X"BC",X"FF",X"CF",
		X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"CC",X"00",X"CC",X"F0",X"BC",X"FE",X"CC",X"FE",
		X"FF",X"FF",X"EE",X"FF",X"00",X"EC",X"CC",X"FF",X"CC",X"FF",X"0C",X"FF",X"0C",X"FF",X"CC",X"FF",
		X"FF",X"EE",X"FF",X"E0",X"EE",X"00",X"FC",X"C0",X"FC",X"CC",X"FF",X"00",X"FF",X"00",X"FC",X"CC",
		X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"FF",X"FF",X"CF",X"FC",X"CF",X"FC",X"CF",
		X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"C0",X"FC",X"C0",X"CF",X"00",X"CC",X"00",X"CC",X"E0",
		X"FC",X"FF",X"FF",X"FF",X"EE",X"FC",X"0E",X"CC",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",
		X"CC",X"E0",X"FF",X"E0",X"FE",X"00",X"EE",X"00",X"CC",X"00",X"CC",X"C0",X"FC",X"00",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"CC",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"CC",X"00",X"CC",X"F0",
		X"FF",X"BB",X"FF",X"BF",X"FF",X"FF",X"EE",X"FF",X"00",X"EE",X"0C",X"FF",X"0C",X"FF",X"00",X"CF",
		X"BC",X"FE",X"BC",X"FE",X"FF",X"EE",X"FF",X"E0",X"EE",X"00",X"FC",X"00",X"FC",X"00",X"CC",X"00",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"CC",X"FF",X"CC",X"FF",X"BC",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"CC",X"00",X"CC",X"F0",X"BC",X"FE",
		X"FF",X"CF",X"FF",X"FF",X"CC",X"FF",X"CC",X"EC",X"CC",X"FF",X"0C",X"FF",X"0C",X"FF",X"0C",X"FF",
		X"CC",X"FE",X"FF",X"EE",X"FF",X"E0",X"EE",X"00",X"FC",X"C0",X"FC",X"CC",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"CC",X"FF",X"CC",X"FF",X"CA",
		X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"CC",X"00",X"CC",X"F0",X"CA",X"FE",
		X"FF",X"CC",X"FF",X"FF",X"FC",X"FF",X"0C",X"EE",X"0C",X"FF",X"0C",X"FF",X"0C",X"FF",X"0C",X"FF",
		X"FC",X"FE",X"FF",X"EE",X"FF",X"E0",X"CE",X"00",X"FC",X"C0",X"FC",X"CC",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CF",X"CC",X"FF",X"FF",X"CC",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"C0",X"CC",X"F0",X"CC",X"FE",
		X"FF",X"CB",X"FF",X"CC",X"FF",X"FF",X"00",X"EE",X"0C",X"FF",X"0C",X"FF",X"0C",X"CF",X"0C",X"CF",
		X"CB",X"FE",X"FC",X"EE",X"FF",X"E0",X"EE",X"00",X"FC",X"00",X"FC",X"C0",X"FF",X"CC",X"FF",X"00",
		X"0C",X"00",X"CC",X"C0",X"CC",X"C0",X"CC",X"FF",X"0F",X"BC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CF",
		X"0C",X"00",X"CC",X"C0",X"CC",X"CC",X"FF",X"CC",X"BC",X"00",X"CC",X"F0",X"CC",X"FE",X"CC",X"FE",
		X"FF",X"FF",X"EE",X"FC",X"C0",X"EE",X"CC",X"FF",X"0C",X"FF",X"0C",X"FF",X"0C",X"FF",X"CC",X"FF",
		X"FF",X"EE",X"FF",X"E0",X"EE",X"CC",X"FC",X"C0",X"FC",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"CC",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"CC",X"FF",X"CF",X"CB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"FF",X"C0",X"CC",X"CC",X"FC",X"F0",X"FF",X"FE",X"FC",X"FE",
		X"FF",X"CC",X"EE",X"FF",X"C0",X"FF",X"CC",X"FF",X"0F",X"FF",X"CC",X"FF",X"CC",X"FF",X"00",X"0C",
		X"CF",X"EE",X"FE",X"E0",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"FF",X"C0",X"FC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FC",X"FF",X"CF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"CF",X"F0",X"FF",X"FE",
		X"FF",X"EE",X"FF",X"FF",X"EE",X"FF",X"CC",X"FF",X"00",X"FF",X"CC",X"FF",X"CC",X"FF",X"00",X"00",
		X"EF",X"FE",X"FE",X"EE",X"FF",X"E0",X"FC",X"CC",X"FF",X"00",X"FF",X"C0",X"FC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CF",X"00",X"FC",X"F0",X"FF",X"FE",
		X"FF",X"EE",X"FF",X"FF",X"EE",X"FF",X"CC",X"FF",X"00",X"FF",X"CC",X"FF",X"0C",X"FF",X"00",X"00",
		X"EF",X"FE",X"FE",X"EE",X"FF",X"EC",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"0C",X"FF",X"CC",X"CF",X"CC",X"CF",X"CC",X"FF",
		X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"FC",X"00",X"CC",X"C0",X"FC",X"CC",X"FF",X"CC",
		X"CF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CE",X"CB",X"CC",X"EF",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",
		X"FF",X"FE",X"FF",X"FE",X"CC",X"EE",X"FB",X"C0",X"EE",X"CC",X"FC",X"CC",X"CC",X"CC",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"EE",X"EC",X"EE",X"EC",X"CE",X"C0",
		X"EE",X"EC",X"EE",X"EC",X"0E",X"EC",X"00",X"ED",X"0E",X"DE",X"EE",X"FF",X"EC",X"FF",X"0E",X"FF",
		X"CE",X"C0",X"EE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"00",X"DD",X"C0",X"FD",X"C0",X"FD",X"00",
		X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",
		X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"EE",X"EC",X"EE",X"EC",X"EE",X"C0",X"EE",X"C0",
		X"EE",X"CC",X"0E",X"CC",X"00",X"DD",X"EE",X"EE",X"CE",X"FF",X"0C",X"FF",X"0E",X"FF",X"EE",X"FF",
		X"EE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"00",X"DD",X"C0",X"FD",X"D0",X"FD",X"C0",X"DD",X"00",
		X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",
		X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"EE",X"EC",X"EE",X"EC",X"CE",X"C0",X"CE",X"C0",
		X"EE",X"EC",X"0E",X"EC",X"00",X"ED",X"EE",X"DE",X"CE",X"FF",X"0C",X"FF",X"00",X"FF",X"EE",X"FF",
		X"EE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"D0",X"DD",X"C0",X"FD",X"00",X"FD",X"00",X"DD",X"C0",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"CE",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"EE",X"EC",X"EE",X"EC",X"EC",X"C0",
		X"EE",X"CE",X"EE",X"EE",X"0E",X"EE",X"00",X"EE",X"0E",X"DD",X"EE",X"FF",X"CC",X"FF",X"00",X"FF",
		X"EC",X"C0",X"EE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"D0",X"DD",X"C0",X"FD",X"00",X"FD",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"C0",X"ED",X"EE",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"CD",X"C0",X"ED",X"EC",X"EE",X"EC",X"EE",X"C0",
		X"EE",X"EE",X"EE",X"EC",X"0E",X"EC",X"00",X"ED",X"0E",X"DE",X"EE",X"FF",X"EC",X"FF",X"0E",X"FF",
		X"CE",X"C0",X"CE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"00",X"DD",X"C0",X"FD",X"C0",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"EE",X"EC",X"EE",X"EC",X"CE",X"C0",
		X"EE",X"EC",X"EE",X"EC",X"CE",X"EC",X"EC",X"ED",X"EE",X"DE",X"0E",X"FF",X"00",X"FF",X"0E",X"FF",
		X"CE",X"C0",X"EE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"00",X"DD",X"C0",X"FD",X"C0",X"FD",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"CE",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"EE",X"EC",X"EE",X"EC",X"EC",X"C0",
		X"EE",X"CE",X"EE",X"EE",X"EC",X"EE",X"0E",X"ED",X"0E",X"DE",X"0E",X"FF",X"00",X"FF",X"0E",X"FF",
		X"EC",X"C0",X"EE",X"C0",X"ED",X"00",X"DC",X"00",X"DD",X"00",X"DD",X"C0",X"FD",X"C0",X"FD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"C0",X"EC",X"EE",X"CD",X"EE",X"CE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"CD",X"C0",X"ED",X"EC",X"EE",X"EC",X"EE",X"C0",
		X"EE",X"CE",X"EE",X"CE",X"CE",X"EE",X"0C",X"ED",X"0E",X"DE",X"0E",X"CF",X"0C",X"EC",X"0E",X"EC",
		X"EC",X"C0",X"EC",X"C0",X"ED",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"D0",X"FD",X"C0",X"FD",X"00",
		X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"CE",X"FE",X"EE",X"FE",X"EF",X"EC",X"FF",X"EC",X"EE",X"EC",
		X"0E",X"00",X"EC",X"C0",X"CD",X"EC",X"FE",X"EC",X"CC",X"EC",X"FF",X"C0",X"EE",X"C0",X"EE",X"C0",
		X"0E",X"ED",X"E0",X"DD",X"EE",X"FF",X"CE",X"FF",X"0C",X"FF",X"EE",X"FF",X"CC",X"FF",X"00",X"CC",
		X"ED",X"00",X"DC",X"D0",X"DD",X"C0",X"FD",X"00",X"FD",X"00",X"FD",X"00",X"DC",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"ED",X"EC",X"DE",X"CC",X"EE",X"EE",X"EE",X"CC",X"EE",X"DD",
		X"F0",X"00",X"00",X"00",X"0E",X"0F",X"FC",X"00",X"EF",X"E0",X"EE",X"E0",X"EE",X"C0",X"EE",X"C0",
		X"EE",X"EE",X"0E",X"FF",X"E0",X"FF",X"CE",X"FF",X"0C",X"FF",X"EE",X"FF",X"CC",X"EE",X"00",X"CD",
		X"DE",X"C0",X"ED",X"00",X"FC",X"D0",X"FD",X"C0",X"FD",X"00",X"ED",X"00",X"EC",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"EC",X"0E",X"EE",X"EE",X"EE",X"EE",X"DD",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"ED",X"00",X"EE",X"00",X"EE",X"C0",X"EE",X"C0",X"DE",X"C0",
		X"EE",X"FF",X"0E",X"FF",X"E0",X"FF",X"CE",X"FF",X"EC",X"FF",X"EE",X"EE",X"CC",X"EE",X"00",X"CD",
		X"ED",X"C0",X"FD",X"00",X"FC",X"D0",X"FD",X"C0",X"ED",X"00",X"ED",X"00",X"EC",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"EC",X"0E",X"EE",X"EE",X"EC",X"EE",X"DD",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"ED",X"00",X"EE",X"00",X"EE",X"C0",X"EE",X"C0",
		X"EE",X"EE",X"EE",X"FF",X"0E",X"FF",X"E0",X"FF",X"EE",X"FF",X"EE",X"EE",X"CC",X"EE",X"00",X"CD",
		X"DE",X"C0",X"ED",X"C0",X"FD",X"00",X"FC",X"00",X"ED",X"00",X"ED",X"00",X"EC",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"C0",X"EC",X"EE",X"CD",X"EE",X"CE",X"EE",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"EE",X"00",X"CD",X"C0",X"ED",X"EC",X"EE",X"EC",
		X"EE",X"EE",X"EE",X"FE",X"EE",X"FF",X"CF",X"EC",X"EC",X"EC",X"EE",X"DE",X"CE",X"FF",X"0C",X"FF",
		X"FE",X"C0",X"FF",X"C0",X"CF",X"C0",X"FF",X"DC",X"DD",X"DC",X"DD",X"C0",X"DD",X"00",X"FD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"BB",X"4C",X"CB",X"4C",
		X"BB",X"BC",X"BB",X"BF",X"BB",X"CF",X"CC",X"FC",X"0B",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"CF",
		X"BB",X"44",X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"CC",X"C4",X"44",X"C4",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",
		X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"BB",X"4C",X"CB",X"4C",X"BB",X"44",
		X"BB",X"BF",X"BB",X"CF",X"CC",X"FC",X"0B",X"FF",X"BB",X"FF",X"BB",X"FF",X"CC",X"FF",X"00",X"FF",
		X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"FC",X"C4",X"FC",X"C4",X"FC",X"40",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",
		X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"CB",X"4C",X"CB",X"4C",X"BB",X"44",
		X"BB",X"BF",X"BB",X"CF",X"CC",X"FC",X"0B",X"FF",X"BB",X"FF",X"BB",X"FF",X"BC",X"FF",X"C0",X"FF",
		X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"FC",X"40",X"FC",X"C4",X"FC",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"CB",X"4C",X"CB",X"4C",
		X"BB",X"BC",X"BB",X"BF",X"BB",X"CF",X"CC",X"FC",X"0B",X"FF",X"BB",X"FF",X"BB",X"FF",X"CC",X"FF",
		X"BB",X"44",X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"40",X"FF",X"C4",X"FC",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BF",X"BB",X"CB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"BB",X"4C",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"BB",X"CF",X"CC",X"CC",X"BB",X"FF",X"BB",X"FF",X"0B",X"FF",
		X"BB",X"4C",X"CB",X"44",X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"C0",X"F4",X"C0",X"44",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"BB",X"4C",X"CB",X"4C",
		X"CB",X"BC",X"CC",X"BF",X"BB",X"CF",X"BB",X"FC",X"BB",X"FF",X"BB",X"FF",X"BB",X"FF",X"CB",X"FF",
		X"BB",X"44",X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"CC",X"C4",X"44",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"CF",X"BB",X"BB",X"BB",X"BB",X"CB",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"BB",X"4C",X"BC",X"4C",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"CC",X"0C",X"BF",X"BB",X"BC",X"BB",X"CC",X"BB",X"FF",X"CB",X"FF",
		X"BB",X"44",X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"CC",X"C4",X"44",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"CF",X"BB",X"BB",X"BB",X"BB",X"CB",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"B4",X"00",X"BB",X"4C",X"BB",X"C0",X"BB",X"4C",X"BC",X"4C",
		X"BB",X"CB",X"BB",X"BB",X"BB",X"CC",X"0C",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"FF",X"CB",X"FF",
		X"BC",X"44",X"BB",X"44",X"C4",X"4C",X"FC",X"C0",X"FF",X"00",X"FF",X"C0",X"CC",X"C4",X"44",X"C4",
		X"00",X"00",X"0C",X"BB",X"0F",X"FB",X"BB",X"FB",X"BB",X"BC",X"BB",X"BF",X"BB",X"CF",X"BB",X"FC",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"4C",X"FF",X"C0",X"BB",X"4C",X"BB",X"4C",X"FB",X"44",
		X"CB",X"FF",X"CC",X"FF",X"BB",X"FF",X"BB",X"FF",X"0C",X"FF",X"0C",X"FF",X"BB",X"FF",X"BB",X"FF",
		X"FF",X"C4",X"FF",X"CC",X"FC",X"C0",X"FF",X"C0",X"FF",X"C0",X"F4",X"4C",X"F4",X"4C",X"44",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"FF",X"BB",X"FF",X"BB",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FC",X"00",X"BF",X"00",X"FB",X"4C",X"FF",X"C0",X"FF",X"4C",X"FF",X"4C",
		X"FF",X"FF",X"BF",X"FF",X"CC",X"FF",X"BB",X"FF",X"BB",X"FF",X"0C",X"FF",X"BB",X"FF",X"CC",X"CB",
		X"FF",X"44",X"FF",X"44",X"FF",X"4C",X"FC",X"C0",X"FF",X"C0",X"FF",X"40",X"F4",X"4C",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BB",X"FF",X"BB",X"FF",X"CC",X"FF",X"BB",X"FF",X"CC",X"FF",
		X"FF",X"4C",X"FF",X"F4",X"FF",X"44",X"FF",X"4C",X"FC",X"C0",X"FF",X"4C",X"FF",X"4C",X"FC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BB",X"FF",X"BB",X"FF",X"BC",X"FF",X"BB",X"BF",X"CC",X"BB",
		X"FF",X"4C",X"FF",X"44",X"FF",X"44",X"FF",X"4C",X"FC",X"C0",X"FF",X"C0",X"FF",X"C0",X"FC",X"00",
		X"00",X"10",X"10",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"FB",X"FF",X"FB",
		X"10",X"00",X"00",X"10",X"C0",X"00",X"BB",X"00",X"FF",X"4C",X"CF",X"C0",X"FF",X"4C",X"FF",X"4C",
		X"FF",X"BB",X"BB",X"BC",X"BB",X"CF",X"CC",X"CC",X"0B",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"FF",
		X"FF",X"F4",X"BB",X"F4",X"C4",X"4C",X"FC",X"C0",X"FF",X"C0",X"F4",X"C0",X"44",X"04",X"C4",X"C4",
		X"00",X"00",X"AA",X"00",X"4B",X"00",X"BB",X"FA",X"AF",X"FA",X"AF",X"CA",X"FF",X"AA",X"AA",X"AC",
		X"00",X"00",X"AA",X"00",X"4B",X"AC",X"FB",X"AC",X"FF",X"C0",X"FF",X"C0",X"CF",X"4C",X"AA",X"4C",
		X"AA",X"CC",X"BB",X"CC",X"CB",X"CC",X"AA",X"AA",X"AA",X"AA",X"CC",X"AA",X"A0",X"AA",X"0A",X"CC",
		X"AA",X"4C",X"A4",X"C0",X"44",X"4C",X"BB",X"C0",X"B4",X"C0",X"4C",X"00",X"C4",X"00",X"4C",X"00",
		X"00",X"C0",X"0C",X"CC",X"CC",X"CC",X"CC",X"FF",X"0F",X"CC",X"FF",X"BB",X"FF",X"CC",X"FF",X"FF",
		X"CC",X"00",X"CC",X"00",X"CC",X"C0",X"FF",X"C0",X"CC",X"00",X"BC",X"F0",X"CB",X"FE",X"FC",X"FE",
		X"FF",X"FF",X"EE",X"CC",X"C0",X"EC",X"CC",X"FE",X"0C",X"FF",X"0C",X"FF",X"00",X"FF",X"CC",X"FF",
		X"FF",X"EE",X"CF",X"E0",X"EE",X"CC",X"FC",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"0C",X"FC",X"C0",
		X"00",X"00",X"0E",X"00",X"EC",X"C0",X"CD",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",X"EE",X"EC",
		X"00",X"00",X"0E",X"00",X"EC",X"C0",X"EE",X"EC",X"EE",X"EC",X"CC",X"EC",X"EC",X"C0",X"EE",X"C0",
		X"EE",X"DD",X"CE",X"EC",X"0C",X"ED",X"EE",X"FF",X"CE",X"FF",X"0C",X"FF",X"00",X"FF",X"E0",X"FF",
		X"EE",X"C0",X"ED",X"00",X"DC",X"D0",X"DD",X"C0",X"FD",X"00",X"FE",X"00",X"FE",X"00",X"FD",X"C0",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"BB",X"BF",X"BB",X"CF",
		X"00",X"00",X"C0",X"00",X"44",X"00",X"B4",X"4C",X"CC",X"C0",X"BC",X"4C",X"BB",X"4C",X"C4",X"44",
		X"CB",X"CC",X"CF",X"FC",X"BC",X"FF",X"BF",X"FF",X"CF",X"FF",X"0F",X"FF",X"BB",X"FF",X"BB",X"FF",
		X"EE",X"C4",X"FE",X"CC",X"FE",X"4C",X"FF",X"4C",X"FF",X"C0",X"FE",X"C0",X"F4",X"C0",X"44",X"C4",
		X"00",X"33",X"33",X"FC",X"CC",X"CC",X"CF",X"CC",X"CF",X"AC",X"AC",X"CC",X"CC",X"CC",X"C9",X"CC",
		X"00",X"00",X"20",X"00",X"C3",X"00",X"C2",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"5C",X"00",
		X"CC",X"5C",X"3C",X"CC",X"02",X"CC",X"00",X"CC",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"20",X"CC",X"20",X"CC",X"20",X"4C",X"20",X"CC",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"03",X"CC",X"3C",X"CC",X"CF",X"CF",X"CF",X"CC",X"FC",X"CC",X"CC",X"C5",X"AC",X"CC",
		X"00",X"00",X"23",X"00",X"CC",X"00",X"CC",X"00",X"5C",X"20",X"CC",X"C2",X"CC",X"C2",X"CC",X"42",
		X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3C",X"33",X"FF",X"CC",X"CC",X"CF",X"CC",
		X"00",X"00",X"00",X"00",X"23",X"00",X"CC",X"00",X"CC",X"20",X"CC",X"20",X"CF",X"20",X"CC",X"20",
		X"FC",X"CC",X"CC",X"FC",X"CC",X"C5",X"AC",X"CC",X"CC",X"CC",X"CC",X"CC",X"3C",X"CC",X"02",X"22",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"C2",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"FA",X"00",X"FA",X"00",X"FA",X"00",X"FA",X"FF",X"FA",X"FF",X"FA",X"AA",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"AC",X"FF",X"AC",X"AA",X"C0",
		X"AA",X"FF",X"CF",X"AF",X"0F",X"AF",X"FF",X"AC",X"FA",X"C0",X"FA",X"00",X"CC",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"FA",X"00",X"FF",X"00",X"CC",X"00",X"00",X"00",
		X"0F",X"C0",X"0F",X"BC",X"0F",X"BB",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"00",X"FB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"FB",X"00",X"FF",X"00",
		X"BB",X"FB",X"BB",X"FB",X"CC",X"FB",X"00",X"FB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",
		X"FF",X"BC",X"BF",X"BC",X"BB",X"BC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"BC",X"AA",X"BB",X"AA",X"AB",X"AA",X"AA",X"AB",X"AA",X"AA",X"CA",X"BA",
		X"BC",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",X"BB",X"00",X"BB",X"C0",X"AB",X"BB",X"AA",X"AB",
		X"AA",X"BA",X"AA",X"AA",X"AB",X"CA",X"BB",X"0A",X"BC",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AC",X"BC",X"C0",X"BC",X"00",X"BB",X"00",X"BB",X"00",X"AB",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"08",X"00",X"89",X"00",X"8C",X"00",X"99",X"00",X"CC",X"00",X"A0",X"00",X"AC",X"00",X"BC",
		X"00",X"40",X"99",X"B4",X"9C",X"4C",X"C0",X"C0",X"6C",X"3C",X"65",X"3C",X"65",X"CC",X"5C",X"8C",
		X"00",X"C7",X"09",X"8C",X"09",X"8C",X"6C",X"CC",X"65",X"77",X"55",X"F7",X"5C",X"73",X"C0",X"33",
		X"CC",X"8C",X"AA",X"8C",X"FA",X"C0",X"AB",X"00",X"BB",X"C0",X"CC",X"C0",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"FF",X"00",X"F6",X"00",X"66",X"00",X"66",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"5C",X"00",X"5C",X"00",X"5C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"F6",X"00",X"16",X"00",X"66",X"00",X"66",X"00",X"65",X"00",X"55",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"5C",X"00",X"5C",X"00",X"5C",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"F1",X"00",X"16",X"00",X"16",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"55",
		X"00",X"00",X"5C",X"00",X"65",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"5C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"16",X"06",X"16",X"06",X"66",X"06",X"66",X"06",X"66",X"06",X"66",X"00",X"65",X"00",X"55",
		X"5C",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"5C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",
		X"00",X"11",X"06",X"16",X"06",X"66",X"06",X"66",X"06",X"66",X"00",X"66",X"00",X"55",X"00",X"55",
		X"65",X"00",X"65",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"66",X"0F",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"65",X"00",
		X"6F",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"65",X"05",X"55",X"00",X"55",
		X"65",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"F6",X"06",X"16",X"06",X"16",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"66",X"06",X"66",X"00",X"55",X"00",X"55",
		X"66",X"C0",X"66",X"C0",X"65",X"C0",X"65",X"C0",X"55",X"00",X"55",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"66",X"66",X"66",X"6F",X"66",X"FF",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"65",X"00",X"65",X"00",X"65",X"C0",
		X"F1",X"66",X"61",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"65",X"06",X"55",X"00",X"55",
		X"65",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"00",X"55",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"16",X"06",X"66",X"6F",X"66",X"6F",X"66",X"61",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"66",X"00",X"66",X"C0",X"66",X"C0",X"66",X"5C",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"65",X"00",X"55",X"00",X"55",
		X"66",X"5C",X"65",X"5C",X"65",X"5C",X"55",X"C0",X"55",X"C0",X"55",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"66",X"06",X"66",X"6F",X"66",X"FF",X"66",X"FF",X"66",X"F1",X"66",X"16",X"66",
		X"00",X"00",X"00",X"00",X"55",X"00",X"65",X"00",X"65",X"C0",X"65",X"C0",X"65",X"5C",X"65",X"5C",
		X"16",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"55",X"55",X"55",X"05",X"55",X"00",X"55",
		X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"C0",X"55",X"C0",X"55",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",X"FC",X"00",X"CC",X"00",X"CC",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"00",X"FC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"00",X"FC",X"00",X"FC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",
		X"00",X"00",X"C0",X"00",X"CC",X"00",X"CC",X"00",X"CB",X"00",X"CC",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"0C",X"CC",X"0C",X"CC",X"0C",X"CC",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",
		X"C0",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"0C",X"1C",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",
		X"CC",X"00",X"CC",X"00",X"CC",X"B0",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"1C",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"CF",X"CC",X"CF",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"0C",X"1C",X"CC",X"CC",X"CF",X"CC",X"CF",X"CC",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"CF",X"CC",X"C1",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"00",X"CC",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"F1",X"0C",X"1C",X"CC",X"1C",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"00",X"BB",X"00",X"BC",X"00",X"CC",X"00",X"CC",X"C0",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"00",X"CC",X"00",X"CC",
		X"CC",X"C0",X"CC",X"C0",X"CC",X"C0",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"0C",X"CC",X"CC",X"CC",X"CF",X"CC",X"FF",X"CC",X"FF",X"CC",X"F1",X"CC",
		X"00",X"00",X"00",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"BB",X"BB",X"BB",X"BB",X"C0",
		X"1C",X"CC",X"1C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"00",X"CC",
		X"CC",X"C0",X"CC",X"C0",X"CC",X"C0",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",X"FC",X"00",X"CC",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"1C",X"CC",X"1C",X"C0",X"1C",X"C0",X"1C",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"C1",X"C1",X"01",X"C1",X"01",X"C1",X"01",
		X"1C",X"C0",X"1C",X"C0",X"1C",X"11",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"01",X"C1",X"01",X"C0",X"11",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"FF",X"00",X"F6",X"00",X"66",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"5C",X"00",X"5C",X"00",X"5C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"FF",X"00",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"5C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"1C",X"10",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"11",X"11",X"11",X"11",X"01",X"1C",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"11",X"CC",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"C1",X"C1",X"C1",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"C1",X"C0",X"C1",X"C0",
		X"C1",X"C1",X"C1",X"C1",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"C0",X"C1",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"CC",X"1C",X"10",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"CC",X"1C",X"10",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"CC",X"1C",X"10",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"1C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
