`define BUILD_DATE "190909"
`define BUILD_TIME "130142"
