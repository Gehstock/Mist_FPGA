library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"18",X"50",X"69",X"30",X"81",X"00",X"10",X"14",X"02",X"80",X"10",X"98",X"01",X"80",X"4C",
		X"C0",X"02",X"00",X"C4",X"40",X"22",X"00",X"88",X"00",X"12",X"92",X"82",X"60",X"12",X"03",X"00",
		X"00",X"20",X"82",X"00",X"00",X"00",X"A0",X"40",X"00",X"30",X"02",X"68",X"40",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"02",X"10",X"00",X"20",X"C3",X"9E",X"01",X"68",X"42",X"80",X"48",X"00",
		X"14",X"80",X"08",X"71",X"25",X"29",X"05",X"08",X"0D",X"05",X"00",X"11",X"70",X"80",X"45",X"03",
		X"4C",X"8E",X"04",X"4D",X"41",X"21",X"00",X"05",X"08",X"0D",X"89",X"01",X"85",X"03",X"25",X"00",
		X"20",X"01",X"28",X"21",X"40",X"00",X"C3",X"34",X"02",X"01",X"00",X"08",X"20",X"08",X"01",X"00",
		X"10",X"00",X"30",X"40",X"00",X"00",X"09",X"00",X"20",X"01",X"20",X"00",X"20",X"30",X"48",X"02",
		X"3A",X"27",X"60",X"3C",X"C3",X"9B",X"3B",X"21",X"88",X"00",X"46",X"45",X"9A",X"80",X"09",X"C0",
		X"82",X"96",X"42",X"81",X"00",X"83",X"8A",X"58",X"80",X"10",X"62",X"04",X"86",X"2A",X"C3",X"01",
		X"00",X"10",X"00",X"90",X"A0",X"00",X"10",X"50",X"22",X"10",X"50",X"00",X"60",X"00",X"02",X"80",
		X"10",X"00",X"1A",X"82",X"41",X"A0",X"0B",X"04",X"00",X"40",X"00",X"08",X"00",X"01",X"00",X"40",
		X"50",X"05",X"40",X"90",X"01",X"01",X"89",X"0C",X"0C",X"2B",X"04",X"40",X"0E",X"14",X"45",X"04",
		X"11",X"20",X"04",X"04",X"04",X"01",X"89",X"55",X"0C",X"02",X"29",X"40",X"83",X"D0",X"90",X"07",
		X"00",X"04",X"02",X"00",X"20",X"41",X"08",X"40",X"40",X"41",X"29",X"00",X"00",X"01",X"29",X"60",
		X"20",X"04",X"20",X"09",X"08",X"00",X"08",X"02",X"00",X"00",X"08",X"01",X"41",X"00",X"20",X"20",
		X"31",X"FF",X"67",X"ED",X"56",X"F3",X"3A",X"00",X"80",X"CD",X"6E",X"17",X"CD",X"D4",X"1A",X"CD",
		X"06",X"2B",X"CD",X"BA",X"1A",X"CD",X"55",X"17",X"CD",X"C6",X"02",X"31",X"FF",X"67",X"AF",X"32",
		X"00",X"A0",X"CD",X"BA",X"1A",X"CD",X"28",X"50",X"CD",X"07",X"26",X"06",X"03",X"C5",X"06",X"03",
		X"AF",X"CD",X"63",X"28",X"CD",X"30",X"50",X"3C",X"CD",X"63",X"28",X"CD",X"30",X"50",X"10",X"F0",
		X"21",X"02",X"90",X"CB",X"76",X"C1",X"CA",X"8C",X"01",X"05",X"20",X"E1",X"CD",X"38",X"50",X"CD",
		X"20",X"50",X"21",X"5F",X"60",X"CB",X"E6",X"21",X"F8",X"0E",X"22",X"D8",X"61",X"00",X"00",X"00",
		X"00",X"00",X"CD",X"36",X"1F",X"32",X"66",X"60",X"AF",X"32",X"67",X"60",X"32",X"65",X"60",X"32",
		X"6E",X"60",X"32",X"6F",X"60",X"C3",X"F7",X"03",X"21",X"1C",X"60",X"AF",X"77",X"21",X"21",X"60",
		X"77",X"CD",X"CD",X"3C",X"21",X"5F",X"60",X"CB",X"A6",X"C3",X"1B",X"01",X"3E",X"09",X"32",X"5E",
		X"60",X"C3",X"5F",X"03",X"C5",X"F5",X"06",X"1F",X"CD",X"28",X"05",X"F1",X"C1",X"C9",X"F5",X"E5",
		X"C5",X"3A",X"CD",X"61",X"FE",X"00",X"C2",X"2B",X"02",X"3A",X"5B",X"60",X"FE",X"00",X"C2",X"2B",
		X"02",X"3E",X"03",X"32",X"5B",X"60",X"3E",X"FF",X"21",X"03",X"90",X"ED",X"67",X"2F",X"21",X"E2",
		X"0B",X"CB",X"27",X"4F",X"06",X"00",X"09",X"D5",X"EB",X"CB",X"39",X"21",X"30",X"68",X"09",X"34",
		X"1A",X"BE",X"CA",X"D9",X"01",X"D1",X"C3",X"26",X"02",X"36",X"00",X"13",X"1A",X"D1",X"C3",X"FC",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"5E",X"60",X"86",
		X"77",X"47",X"3A",X"21",X"D3",X"FE",X"1D",X"20",X"08",X"78",X"FE",X"0A",X"30",X"03",X"32",X"61",
		X"D3",X"3A",X"5F",X"60",X"CB",X"47",X"20",X"0E",X"21",X"08",X"00",X"39",X"F9",X"01",X"5F",X"03",
		X"C5",X"21",X"FA",X"FF",X"39",X"F9",X"21",X"01",X"60",X"CB",X"E6",X"3A",X"00",X"80",X"FB",X"C1",
		X"E1",X"F1",X"ED",X"4D",X"F5",X"E5",X"C5",X"3A",X"CD",X"61",X"FE",X"00",X"C2",X"C1",X"02",X"3A",
		X"5B",X"60",X"FE",X"00",X"C2",X"C1",X"02",X"3E",X"03",X"32",X"5B",X"60",X"3E",X"FF",X"21",X"03",
		X"90",X"ED",X"6F",X"2F",X"21",X"E2",X"0B",X"CB",X"27",X"4F",X"06",X"00",X"09",X"D5",X"EB",X"CB",
		X"39",X"21",X"30",X"68",X"09",X"34",X"1A",X"BE",X"CA",X"6F",X"02",X"D1",X"C3",X"BC",X"02",X"36",
		X"00",X"13",X"1A",X"D1",X"C3",X"92",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"5E",X"60",X"86",X"77",X"47",X"3A",X"21",X"D3",X"FE",X"1D",X"20",X"08",X"78",
		X"FE",X"0A",X"30",X"03",X"32",X"61",X"D3",X"3A",X"5F",X"60",X"CB",X"47",X"20",X"0E",X"21",X"08",
		X"00",X"39",X"F9",X"01",X"5F",X"03",X"C5",X"21",X"FA",X"FF",X"39",X"F9",X"21",X"01",X"60",X"CB",
		X"E6",X"C1",X"E1",X"F1",X"ED",X"45",X"AF",X"32",X"5B",X"60",X"32",X"00",X"A0",X"32",X"C9",X"61",
		X"CD",X"40",X"50",X"32",X"CD",X"61",X"32",X"5E",X"60",X"C3",X"57",X"49",X"CD",X"F9",X"02",X"CD",
		X"0A",X"03",X"AF",X"21",X"68",X"60",X"77",X"23",X"77",X"23",X"77",X"21",X"00",X"60",X"06",X"1C",
		X"77",X"23",X"10",X"FC",X"CD",X"2F",X"03",X"FB",X"C9",X"06",X"09",X"21",X"73",X"60",X"AF",X"3C",
		X"77",X"AF",X"23",X"77",X"23",X"77",X"23",X"10",X"F6",X"C9",X"21",X"80",X"D3",X"06",X"09",X"C5",
		X"06",X"02",X"3E",X"FF",X"77",X"23",X"10",X"FC",X"DD",X"21",X"FC",X"2E",X"06",X"09",X"DD",X"7E",
		X"00",X"DD",X"23",X"77",X"23",X"10",X"F7",X"3E",X"FF",X"77",X"23",X"C1",X"10",X"E1",X"C9",X"06",
		X"32",X"AF",X"21",X"1C",X"60",X"77",X"23",X"10",X"FC",X"C9",X"F5",X"3A",X"5B",X"60",X"FE",X"00",
		X"28",X"04",X"3D",X"32",X"5B",X"60",X"3A",X"CD",X"61",X"FE",X"00",X"28",X"01",X"3D",X"32",X"CD",
		X"61",X"3A",X"00",X"90",X"CB",X"7F",X"20",X"05",X"3E",X"05",X"32",X"CD",X"61",X"F1",X"C9",X"21",
		X"5F",X"60",X"CB",X"C6",X"CB",X"A6",X"21",X"1C",X"60",X"AF",X"77",X"21",X"21",X"60",X"77",X"CD",
		X"CD",X"3C",X"AF",X"32",X"00",X"A0",X"CD",X"25",X"25",X"3E",X"01",X"32",X"E2",X"61",X"AF",X"32",
		X"C8",X"61",X"01",X"17",X"00",X"21",X"00",X"90",X"CB",X"6E",X"28",X"27",X"3A",X"5E",X"60",X"FE",
		X"02",X"38",X"04",X"CB",X"76",X"28",X"34",X"C5",X"CD",X"A5",X"1C",X"CD",X"E5",X"27",X"CD",X"55",
		X"27",X"CD",X"5A",X"2D",X"C1",X"0B",X"78",X"B1",X"20",X"DB",X"3A",X"C8",X"61",X"CD",X"63",X"28",
		X"2F",X"18",X"CC",X"3A",X"5F",X"60",X"CB",X"8F",X"32",X"5F",X"60",X"CD",X"36",X"1F",X"32",X"66",
		X"60",X"AF",X"32",X"67",X"60",X"21",X"5E",X"60",X"35",X"18",X"16",X"3A",X"5F",X"60",X"CB",X"CF",
		X"32",X"5F",X"60",X"CD",X"36",X"1F",X"32",X"66",X"60",X"32",X"67",X"60",X"C3",X"60",X"49",X"35",
		X"35",X"AF",X"C3",X"6C",X"49",X"21",X"68",X"60",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",
		X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"3E",X"FF",X"21",X"9D",X"60",X"06",X"06",X"77",X"23",
		X"10",X"FC",X"AF",X"32",X"9F",X"60",X"32",X"A2",X"60",X"21",X"1C",X"D6",X"22",X"63",X"60",X"21",
		X"5F",X"60",X"CB",X"96",X"CD",X"BA",X"1A",X"CD",X"E5",X"1B",X"AF",X"32",X"60",X"60",X"2F",X"32",
		X"62",X"60",X"3E",X"0C",X"32",X"61",X"60",X"CD",X"C6",X"1C",X"CD",X"44",X"21",X"CD",X"42",X"1D",
		X"CD",X"64",X"1D",X"CD",X"77",X"1D",X"CD",X"D1",X"1D",X"CD",X"8B",X"1E",X"06",X"06",X"3E",X"05",
		X"21",X"A1",X"D5",X"CD",X"7D",X"1E",X"CD",X"E0",X"1E",X"CD",X"26",X"28",X"06",X"05",X"3E",X"01",
		X"21",X"E1",X"D4",X"CD",X"7D",X"1E",X"21",X"E1",X"D0",X"36",X"2A",X"19",X"CD",X"44",X"1F",X"DD",
		X"21",X"1C",X"60",X"DD",X"36",X"00",X"82",X"DD",X"36",X"01",X"08",X"DD",X"36",X"02",X"0F",X"CD",
		X"7F",X"1F",X"DD",X"77",X"03",X"DD",X"70",X"04",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"DD",X"36",
		X"00",X"81",X"C3",X"D5",X"04",X"DD",X"21",X"70",X"60",X"ED",X"5F",X"0E",X"00",X"1F",X"CB",X"11",
		X"DD",X"71",X"00",X"ED",X"5F",X"E6",X"07",X"1F",X"CE",X"02",X"FE",X"05",X"20",X"0A",X"3A",X"E2",
		X"61",X"FE",X"00",X"3E",X"05",X"20",X"01",X"3C",X"DD",X"77",X"01",X"ED",X"5F",X"1F",X"E6",X"03",
		X"1F",X"CE",X"07",X"FE",X"08",X"20",X"1A",X"47",X"CD",X"36",X"1F",X"3C",X"4F",X"3A",X"65",X"60",
		X"FE",X"00",X"28",X"05",X"3A",X"67",X"60",X"18",X"03",X"3A",X"66",X"60",X"B9",X"78",X"38",X"01",
		X"3C",X"DD",X"77",X"02",X"C9",X"AF",X"32",X"C9",X"61",X"CD",X"CF",X"33",X"CD",X"77",X"1D",X"CD",
		X"85",X"04",X"CD",X"FE",X"28",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"3E",X"81",X"32",X"21",X"60",
		X"CD",X"F4",X"30",X"CD",X"1C",X"31",X"CD",X"54",X"31",X"CD",X"77",X"1D",X"CD",X"F4",X"1E",X"21",
		X"01",X"D1",X"CD",X"44",X"1F",X"21",X"1F",X"60",X"CD",X"7F",X"1F",X"77",X"23",X"70",X"CD",X"C7",
		X"1F",X"CD",X"8F",X"17",X"06",X"B4",X"CD",X"28",X"05",X"CD",X"C1",X"2A",X"AF",X"32",X"21",X"60",
		X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"18",X"19",X"21",X"01",X"90",X"CD",X"5A",X"2D",X"CB",X"7E",
		X"28",X"FC",X"CB",X"7E",X"20",X"FC",X"C5",X"CD",X"3A",X"03",X"CD",X"8F",X"17",X"C1",X"10",X"E8",
		X"C9",X"CD",X"44",X"21",X"CD",X"E3",X"33",X"CD",X"5C",X"21",X"CD",X"92",X"31",X"CD",X"DA",X"30",
		X"CD",X"CF",X"30",X"CD",X"44",X"31",X"3E",X"03",X"32",X"9B",X"61",X"CD",X"15",X"2B",X"CD",X"F4",
		X"30",X"CD",X"1C",X"31",X"CD",X"54",X"31",X"CD",X"F4",X"1E",X"21",X"01",X"D1",X"CD",X"44",X"1F",
		X"DD",X"21",X"1C",X"60",X"DD",X"36",X"00",X"82",X"DD",X"36",X"01",X"08",X"DD",X"36",X"02",X"0F",
		X"CD",X"7F",X"1F",X"DD",X"77",X"03",X"DD",X"70",X"04",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"DD",
		X"36",X"00",X"81",X"21",X"1C",X"D6",X"22",X"63",X"60",X"AF",X"32",X"60",X"60",X"2F",X"32",X"62",
		X"60",X"3E",X"0C",X"32",X"61",X"60",X"CD",X"C6",X"1C",X"CD",X"AE",X"05",X"18",X"23",X"11",X"05",
		X"00",X"21",X"2B",X"60",X"0E",X"00",X"7E",X"E6",X"03",X"28",X"08",X"19",X"0C",X"FE",X"04",X"20",
		X"F5",X"18",X"0D",X"CD",X"61",X"30",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"DD",X"36",X"00",X"81",
		X"C9",X"3A",X"65",X"60",X"FE",X"00",X"28",X"05",X"21",X"67",X"60",X"18",X"03",X"21",X"66",X"60",
		X"35",X"7E",X"F5",X"CD",X"77",X"1D",X"F1",X"DD",X"21",X"26",X"60",X"DD",X"36",X"00",X"42",X"DD",
		X"36",X"02",X"1F",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"C6",X"08",X"DD",X"77",X"01",
		X"DD",X"36",X"03",X"00",X"DD",X"36",X"04",X"00",X"C3",X"21",X"06",X"CD",X"C1",X"2A",X"AF",X"32",
		X"C9",X"61",X"CD",X"4C",X"1E",X"CD",X"44",X"21",X"CD",X"5C",X"21",X"CD",X"92",X"35",X"C3",X"56",
		X"05",X"21",X"00",X"60",X"CB",X"F6",X"21",X"27",X"60",X"AF",X"16",X"58",X"06",X"0F",X"10",X"06",
		X"2F",X"CD",X"4C",X"1E",X"06",X"0F",X"F5",X"C5",X"E5",X"D5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",
		X"D1",X"E1",X"C1",X"7E",X"BA",X"28",X"04",X"34",X"F1",X"18",X"E3",X"FE",X"56",X"28",X"0A",X"3E",
		X"82",X"32",X"26",X"60",X"23",X"16",X"56",X"18",X"EF",X"F1",X"3E",X"FF",X"CD",X"4C",X"1E",X"C3",
		X"30",X"07",X"CD",X"CF",X"33",X"21",X"66",X"60",X"3A",X"65",X"60",X"FE",X"00",X"28",X"03",X"21",
		X"67",X"60",X"34",X"34",X"E5",X"CD",X"85",X"04",X"E1",X"35",X"35",X"CD",X"FE",X"28",X"CD",X"C7",
		X"1F",X"CD",X"8F",X"17",X"3E",X"81",X"32",X"21",X"60",X"CD",X"F4",X"30",X"CD",X"1C",X"31",X"CD",
		X"54",X"31",X"CD",X"77",X"1D",X"CD",X"F4",X"1E",X"21",X"01",X"D1",X"CD",X"44",X"1F",X"21",X"1F",
		X"60",X"CD",X"7F",X"1F",X"77",X"23",X"70",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"06",X"B4",X"CD",
		X"28",X"05",X"CD",X"C1",X"2A",X"AF",X"32",X"21",X"60",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"CD",
		X"44",X"21",X"CD",X"E3",X"33",X"CD",X"5C",X"21",X"CD",X"92",X"31",X"CD",X"44",X"31",X"CD",X"54",
		X"31",X"CD",X"DA",X"30",X"CD",X"CF",X"30",X"CD",X"15",X"2B",X"AF",X"32",X"60",X"60",X"2F",X"32",
		X"62",X"60",X"3E",X"0C",X"32",X"61",X"60",X"CD",X"C6",X"1C",X"21",X"1C",X"D6",X"22",X"63",X"60",
		X"CD",X"F4",X"1E",X"21",X"01",X"D1",X"CD",X"44",X"1F",X"DD",X"21",X"1C",X"60",X"DD",X"36",X"00",
		X"82",X"DD",X"36",X"01",X"08",X"DD",X"36",X"02",X"0F",X"CD",X"7F",X"1F",X"DD",X"77",X"03",X"DD",
		X"70",X"04",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"DD",X"36",X"00",X"81",X"CD",X"AE",X"05",X"21",
		X"26",X"60",X"36",X"82",X"23",X"36",X"58",X"23",X"36",X"56",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",
		X"CD",X"E3",X"35",X"DD",X"21",X"B6",X"61",X"DD",X"36",X"00",X"60",X"DD",X"36",X"01",X"00",X"DD",
		X"36",X"02",X"00",X"DD",X"36",X"03",X"B4",X"AF",X"32",X"B5",X"61",X"32",X"B4",X"61",X"32",X"E1",
		X"61",X"21",X"CE",X"61",X"06",X"05",X"AF",X"77",X"23",X"10",X"FC",X"21",X"5F",X"60",X"CB",X"FE",
		X"21",X"96",X"61",X"36",X"58",X"23",X"36",X"56",X"23",X"36",X"08",X"3E",X"08",X"32",X"98",X"61",
		X"11",X"00",X"00",X"ED",X"53",X"99",X"61",X"21",X"5F",X"60",X"CB",X"B6",X"CD",X"FD",X"45",X"CD",
		X"3A",X"46",X"18",X"06",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"CD",X"5A",X"2D",X"21",X"5F",X"60",
		X"CB",X"66",X"20",X"08",X"21",X"02",X"90",X"CB",X"5E",X"CA",X"5E",X"09",X"CD",X"B1",X"39",X"CD",
		X"56",X"39",X"3A",X"E1",X"61",X"FE",X"00",X"20",X"03",X"CD",X"7E",X"40",X"CD",X"06",X"44",X"CD",
		X"FF",X"35",X"CD",X"99",X"3A",X"06",X"04",X"21",X"2B",X"60",X"11",X"05",X"00",X"CB",X"4E",X"C2",
		X"C8",X"07",X"19",X"10",X"F8",X"C3",X"EE",X"07",X"E5",X"23",X"23",X"3A",X"28",X"60",X"96",X"30",
		X"02",X"ED",X"44",X"FE",X"09",X"D2",X"EA",X"07",X"2B",X"3A",X"27",X"60",X"96",X"30",X"02",X"ED",
		X"44",X"FE",X"09",X"D2",X"EA",X"07",X"E1",X"C3",X"8B",X"08",X"E1",X"C3",X"C2",X"07",X"CD",X"B0",
		X"3C",X"E6",X"0F",X"FE",X"0F",X"20",X"1D",X"DD",X"21",X"21",X"60",X"DD",X"CB",X"00",X"4E",X"CA",
		X"14",X"08",X"DD",X"7E",X"01",X"DD",X"BE",X"06",X"C2",X"14",X"08",X"DD",X"7E",X"02",X"DD",X"BE",
		X"07",X"CA",X"98",X"08",X"3A",X"5F",X"60",X"CB",X"7F",X"20",X"30",X"3A",X"27",X"60",X"57",X"3A",
		X"28",X"60",X"5F",X"3A",X"26",X"60",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"02",
		X"28",X"0D",X"38",X"0F",X"FE",X"04",X"28",X"0E",X"7B",X"D6",X"04",X"5F",X"C3",X"6E",X"08",X"1D",
		X"C3",X"6E",X"08",X"14",X"14",X"14",X"14",X"14",X"C3",X"6E",X"08",X"3A",X"28",X"60",X"21",X"97",
		X"61",X"96",X"D2",X"57",X"08",X"ED",X"44",X"FE",X"05",X"D2",X"88",X"08",X"3A",X"27",X"60",X"2B",
		X"96",X"D2",X"66",X"08",X"ED",X"44",X"FE",X"05",X"D2",X"88",X"08",X"56",X"23",X"5E",X"CD",X"0A",
		X"3C",X"7E",X"FE",X"E5",X"CA",X"4A",X"09",X"FE",X"63",X"CA",X"EA",X"0A",X"FE",X"59",X"38",X"08",
		X"FE",X"62",X"DA",X"FE",X"09",X"CA",X"CC",X"09",X"C3",X"84",X"07",X"CB",X"86",X"CB",X"8E",X"CD",
		X"C7",X"1F",X"CD",X"8F",X"17",X"C3",X"F3",X"0A",X"21",X"21",X"60",X"CB",X"86",X"CB",X"8E",X"21",
		X"26",X"60",X"CB",X"8E",X"21",X"00",X"60",X"CB",X"CE",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"3E",
		X"05",X"32",X"E1",X"61",X"CD",X"26",X"1F",X"FE",X"13",X"38",X"02",X"3E",X"12",X"F5",X"3D",X"21",
		X"79",X"0C",X"06",X"00",X"4F",X"09",X"4E",X"3A",X"65",X"60",X"FE",X"00",X"20",X"06",X"DD",X"21",
		X"68",X"60",X"18",X"04",X"DD",X"21",X"6B",X"60",X"DD",X"7E",X"01",X"81",X"27",X"DD",X"77",X"01",
		X"DD",X"7E",X"00",X"88",X"27",X"DD",X"77",X"00",X"3A",X"65",X"60",X"FE",X"00",X"20",X"05",X"21",
		X"C4",X"D2",X"18",X"03",X"21",X"C3",X"D2",X"CD",X"06",X"1E",X"F1",X"11",X"00",X"04",X"3D",X"47",
		X"C6",X"C6",X"21",X"F0",X"D1",X"77",X"19",X"36",X"05",X"78",X"FE",X"06",X"38",X"04",X"3E",X"D9",
		X"18",X"02",X"3E",X"D8",X"21",X"10",X"D2",X"77",X"19",X"36",X"05",X"06",X"20",X"C5",X"CD",X"C7",
		X"1F",X"CD",X"8F",X"17",X"CD",X"5A",X"2D",X"C1",X"10",X"F3",X"21",X"F0",X"D1",X"36",X"32",X"11",
		X"00",X"04",X"19",X"36",X"00",X"21",X"10",X"D2",X"36",X"FF",X"19",X"36",X"00",X"21",X"5F",X"60",
		X"CB",X"F6",X"21",X"26",X"60",X"CB",X"CE",X"C3",X"84",X"07",X"3E",X"FF",X"77",X"1E",X"00",X"CD",
		X"2C",X"3C",X"21",X"00",X"60",X"CB",X"DE",X"21",X"A9",X"60",X"35",X"C2",X"84",X"07",X"CD",X"2F",
		X"3F",X"21",X"01",X"60",X"CB",X"CE",X"CD",X"2F",X"3F",X"21",X"9B",X"61",X"35",X"20",X"1E",X"3A",
		X"5F",X"60",X"CB",X"4F",X"28",X"17",X"3A",X"65",X"60",X"FE",X"00",X"28",X"09",X"3A",X"66",X"60",
		X"FE",X"00",X"28",X"09",X"18",X"16",X"3A",X"67",X"60",X"FE",X"00",X"20",X"0F",X"CD",X"CD",X"3C",
		X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"CD",X"54",X"40",X"C3",X"62",X"06",X"CD",X"99",X"3A",X"CD",
		X"F3",X"3C",X"CD",X"10",X"35",X"CD",X"CD",X"3C",X"21",X"26",X"60",X"CB",X"CE",X"CD",X"74",X"2C",
		X"06",X"80",X"CD",X"28",X"05",X"3A",X"65",X"60",X"2F",X"32",X"65",X"60",X"CD",X"CD",X"3F",X"21",
		X"5F",X"60",X"CB",X"56",X"CA",X"D5",X"04",X"CB",X"96",X"C3",X"0B",X"06",X"CD",X"E5",X"3F",X"CD",
		X"2B",X"3D",X"CD",X"9F",X"3D",X"CD",X"2C",X"3C",X"CD",X"BD",X"3D",X"7B",X"FE",X"01",X"20",X"1B",
		X"3A",X"65",X"60",X"FE",X"00",X"20",X"06",X"21",X"9F",X"60",X"34",X"18",X"04",X"21",X"A2",X"60",
		X"34",X"7E",X"FE",X"04",X"38",X"02",X"36",X"03",X"CD",X"54",X"31",X"C3",X"57",X"09",X"CD",X"E5",
		X"3F",X"CD",X"9F",X"3D",X"7B",X"FE",X"03",X"28",X"04",X"FE",X"02",X"20",X"04",X"7E",X"CD",X"5E",
		X"3E",X"D5",X"CD",X"2B",X"3D",X"D1",X"CD",X"2C",X"3C",X"CD",X"BD",X"3D",X"7B",X"FE",X"03",X"28",
		X"04",X"FE",X"02",X"20",X"12",X"CD",X"96",X"3E",X"7E",X"CB",X"BF",X"FE",X"00",X"28",X"0B",X"23",
		X"7E",X"E6",X"1F",X"FE",X"00",X"28",X"45",X"C3",X"57",X"09",X"AF",X"21",X"E2",X"61",X"BE",X"28",
		X"01",X"35",X"C3",X"89",X"49",X"21",X"00",X"60",X"CB",X"FE",X"06",X"00",X"48",X"04",X"CD",X"C2",
		X"0A",X"CD",X"10",X"50",X"06",X"00",X"0E",X"00",X"CD",X"FC",X"1B",X"3E",X"FF",X"08",X"21",X"9D",
		X"60",X"3A",X"65",X"60",X"FE",X"00",X"28",X"03",X"21",X"A0",X"60",X"08",X"77",X"21",X"01",X"60",
		X"CB",X"E6",X"21",X"5E",X"60",X"34",X"CD",X"26",X"28",X"C3",X"69",X"09",X"CD",X"2F",X"3F",X"21",
		X"00",X"60",X"CB",X"FE",X"06",X"01",X"48",X"CD",X"C2",X"0A",X"CD",X"08",X"50",X"06",X"00",X"0E",
		X"01",X"CD",X"FC",X"1B",X"3E",X"FF",X"08",X"21",X"9E",X"60",X"3A",X"65",X"60",X"FE",X"00",X"28",
		X"03",X"21",X"A1",X"60",X"08",X"77",X"21",X"01",X"60",X"CB",X"F6",X"3A",X"65",X"60",X"FE",X"00",
		X"20",X"06",X"21",X"66",X"60",X"34",X"18",X"04",X"21",X"67",X"60",X"34",X"CD",X"77",X"1D",X"C3",
		X"69",X"09",X"C5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"C1",X"3A",X"59",X"60",X"E6",X"0F",X"20",
		X"0C",X"78",X"FE",X"01",X"28",X"03",X"05",X"18",X"01",X"04",X"CD",X"FC",X"1B",X"3A",X"03",X"60",
		X"FE",X"00",X"20",X"DE",X"06",X"01",X"CD",X"FC",X"1B",X"C9",X"CD",X"E5",X"3F",X"CD",X"2B",X"3D",
		X"CD",X"05",X"40",X"21",X"01",X"60",X"CB",X"EE",X"CD",X"64",X"2D",X"CD",X"CD",X"3C",X"E5",X"21",
		X"5F",X"60",X"CB",X"66",X"E1",X"C2",X"78",X"01",X"3A",X"65",X"60",X"FE",X"00",X"20",X"13",X"3A",
		X"66",X"60",X"FE",X"00",X"20",X"1F",X"3A",X"67",X"60",X"FE",X"00",X"CA",X"96",X"0B",X"3E",X"01",
		X"18",X"37",X"3A",X"67",X"60",X"FE",X"00",X"20",X"0C",X"3A",X"66",X"60",X"FE",X"00",X"CA",X"96",
		X"0B",X"3E",X"02",X"18",X"24",X"3A",X"5F",X"60",X"CB",X"4F",X"28",X"17",X"3A",X"65",X"60",X"FE",
		X"00",X"20",X"09",X"3A",X"67",X"60",X"FE",X"00",X"20",X"24",X"18",X"07",X"3A",X"66",X"60",X"FE",
		X"00",X"20",X"1B",X"CD",X"99",X"3A",X"C3",X"93",X"05",X"F5",X"CD",X"99",X"3A",X"CD",X"F3",X"3C",
		X"CD",X"10",X"35",X"F1",X"CD",X"FC",X"2C",X"06",X"80",X"CD",X"28",X"05",X"18",X"09",X"CD",X"99",
		X"3A",X"CD",X"F3",X"3C",X"CD",X"10",X"35",X"CD",X"74",X"2C",X"06",X"80",X"CD",X"28",X"05",X"3A",
		X"65",X"60",X"2F",X"32",X"65",X"60",X"CD",X"CD",X"3F",X"21",X"5F",X"60",X"CB",X"56",X"C2",X"0B",
		X"06",X"CB",X"D6",X"C3",X"D5",X"04",X"CD",X"FC",X"2C",X"06",X"80",X"CD",X"28",X"05",X"21",X"1C",
		X"60",X"CB",X"86",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"CD",X"BA",X"1A",X"CD",X"00",X"50",X"3A",
		X"5E",X"60",X"FE",X"00",X"28",X"0A",X"21",X"02",X"90",X"CB",X"76",X"28",X"1D",X"C3",X"5F",X"03",
		X"21",X"02",X"90",X"CB",X"76",X"28",X"13",X"21",X"5F",X"60",X"CB",X"86",X"06",X"02",X"C5",X"06",
		X"B4",X"CD",X"28",X"05",X"C1",X"10",X"F7",X"C3",X"1B",X"01",X"3E",X"09",X"32",X"5E",X"60",X"C3",
		X"5F",X"03",X"01",X"01",X"01",X"02",X"01",X"03",X"01",X"04",X"01",X"05",X"02",X"01",X"02",X"03",
		X"03",X"01",X"03",X"02",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"D8",X"D0",X"DA",X"D0",X"9A",X"D1",X"DA",X"D1",X"14",X"D2",X"16",X"D2",X"18",X"D2",
		X"1A",X"D2",X"5A",X"D2",X"9A",X"D2",X"C6",X"D0",X"C8",X"D0",X"CA",X"D0",X"CC",X"D0",X"CE",X"D0",
		X"D0",X"D0",X"D2",X"D0",X"0A",X"D1",X"10",X"D1",X"12",X"D1",X"4A",X"D1",X"52",X"D1",X"86",X"D1",
		X"C6",X"D1",X"D0",X"D1",X"46",X"D2",X"50",X"D2",X"86",X"D2",X"CA",X"D2",X"D2",X"D2",X"0A",X"D3",
		X"10",X"D3",X"12",X"D3",X"46",X"D3",X"48",X"D3",X"4A",X"D3",X"4C",X"D3",X"4E",X"D3",X"50",X"D3",
		X"52",X"D3",X"08",X"06",X"07",X"07",X"9D",X"D4",X"97",X"06",X"BD",X"D5",X"75",X"05",X"9D",X"D6",
		X"86",X"4D",X"1C",X"19",X"0E",X"0C",X"12",X"0A",X"15",X"4D",X"4D",X"0E",X"21",X"1D",X"1B",X"0A",
		X"4D",X"4D",X"56",X"02",X"56",X"03",X"56",X"05",X"4D",X"10",X"15",X"20",X"25",X"30",X"35",X"40",
		X"45",X"50",X"55",X"60",X"65",X"70",X"75",X"80",X"85",X"90",X"95",X"18",X"30",X"60",X"48",X"78",
		X"90",X"A8",X"C0",X"10",X"11",X"1B",X"1C",X"10",X"1C",X"15",X"15",X"14",X"1A",X"15",X"16",X"19",
		X"14",X"10",X"14",X"12",X"14",X"62",X"70",X"88",X"A0",X"63",X"72",X"8C",X"A2",X"5E",X"66",X"74",
		X"9A",X"5B",X"64",X"74",X"94",X"59",X"64",X"74",X"90",X"5A",X"66",X"74",X"92",X"5C",X"64",X"74",
		X"96",X"5D",X"68",X"78",X"98",X"5C",X"6A",X"7C",X"96",X"5F",X"6C",X"80",X"9C",X"60",X"6E",X"84",
		X"9E",X"61",X"66",X"74",X"92",X"00",X"47",X"46",X"49",X"48",X"FF",X"4A",X"FF",X"00",X"41",X"39",
		X"00",X"40",X"42",X"43",X"00",X"44",X"45",X"01",X"39",X"01",X"35",X"36",X"37",X"01",X"FF",X"01",
		X"01",X"3D",X"01",X"40",X"3E",X"FF",X"01",X"3F",X"01",X"01",X"FC",X"06",X"F2",X"03",X"6D",X"06",
		X"C7",X"01",X"FC",X"03",X"6D",X"06",X"F2",X"06",X"C7",X"11",X"21",X"13",X"11",X"32",X"13",X"21",
		X"12",X"11",X"31",X"12",X"13",X"23",X"22",X"32",X"32",X"21",X"12",X"11",X"12",X"F5",X"D0",X"27",
		X"D1",X"2D",X"D1",X"39",X"D1",X"6F",X"D1",X"75",X"D1",X"A9",X"D1",X"AD",X"D1",X"B3",X"D1",X"B7",
		X"D1",X"69",X"D2",X"6D",X"D2",X"73",X"D2",X"77",X"D2",X"AF",X"D2",X"B5",X"D2",X"E7",X"D2",X"ED",
		X"D2",X"F9",X"D2",X"35",X"D3",X"32",X"3C",X"38",X"31",X"32",X"3B",X"38",X"33",X"33",X"3C",X"34",
		X"31",X"33",X"3B",X"34",X"33",X"20",X"01",X"13",X"12",X"20",X"11",X"33",X"33",X"12",X"10",X"FF",
		X"E5",X"5E",X"5B",X"59",X"5A",X"5C",X"5D",X"5C",X"5F",X"60",X"61",X"62",X"63",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"FF",X"0C",X"11",X"0A",X"17",X"10",X"0E",X"09",X"0A",X"2B",X"36",X"3A",X"3B",
		X"3C",X"3D",X"48",X"53",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"0D",X"10",X"11",X"18",X"1C",
		X"21",X"2C",X"31",X"3E",X"43",X"49",X"56",X"5A",X"61",X"64",X"65",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"70",X"AC",X"AE",X"EA",X"EE",X"AE",X"06",X"6D",X"C5",X"3E",X"95",X"C7",X"07",X"7D",X"BD",
		X"EF",X"EB",X"BF",X"07",X"D5",X"EF",X"BF",X"FE",X"EF",X"07",X"BD",X"97",X"AF",X"3F",X"3D",X"05",
		X"AD",X"AF",X"87",X"AF",X"AF",X"07",X"ED",X"C7",X"AF",X"6F",X"6D",X"05",X"D5",X"BF",X"EF",X"FB",
		X"BF",X"07",X"7D",X"ED",X"BF",X"BE",X"EF",X"07",X"3D",X"95",X"6B",X"C5",X"97",X"07",X"A9",X"AB",
		X"BA",X"BB",X"AB",X"03",X"77",X"07",X"DE",X"03",X"FD",X"05",X"DE",X"03",X"FE",X"03",X"AF",X"07",
		X"FD",X"05",X"DF",X"07",X"FF",X"07",X"DE",X"03",X"AF",X"07",X"E5",X"05",X"FF",X"07",X"FF",X"07",
		X"FE",X"07",X"DF",X"03",X"75",X"05",X"DF",X"03",X"FE",X"07",X"FF",X"07",X"BB",X"07",X"E5",X"05",
		X"01",X"02",X"03",X"05",X"03",X"06",X"09",X"15",X"08",X"16",X"24",X"40",X"DA",X"D0",X"10",X"D3",
		X"0A",X"D1",X"10",X"D1",X"12",X"D1",X"86",X"D1",X"9A",X"D1",X"DA",X"D1",X"1A",X"D2",X"5A",X"D2",
		X"86",X"D2",X"9A",X"D2",X"0A",X"D3",X"12",X"D3",X"C6",X"D0",X"C8",X"D0",X"CA",X"D0",X"CC",X"D0",
		X"CE",X"D0",X"D0",X"D0",X"D2",X"D0",X"D8",X"D0",X"D0",X"D1",X"14",X"D2",X"18",X"D2",X"50",X"D2",
		X"D2",X"D2",X"48",X"D3",X"4C",X"D3",X"4E",X"D3",X"FF",X"31",X"30",X"32",X"FF",X"31",X"31",X"FF",
		X"FF",X"FF",X"32",X"32",X"FF",X"FF",X"33",X"FF",X"10",X"0A",X"16",X"0E",X"FF",X"18",X"1F",X"0E",
		X"1B",X"01",X"1C",X"1D",X"FF",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"02",X"17",X"0D",X"FF",X"19",
		X"15",X"0A",X"22",X"0E",X"1B",X"AE",X"AB",X"A7",X"AB",X"AE",X"A7",X"AB",X"00",X"01",X"02",X"03",
		X"00",X"03",X"03",X"03",X"04",X"00",X"04",X"04",X"04",X"04",X"00",X"04",X"05",X"05",X"05",X"00",
		X"06",X"06",X"06",X"07",X"90",X"24",X"00",X"00",X"02",X"04",X"01",X"03",X"05",X"06",X"08",X"05",
		X"07",X"09",X"0A",X"0B",X"08",X"0C",X"0D",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"10",X"10",X"10",X"10",X"10",X"10",X"12",X"12",
		X"12",X"12",X"12",X"12",X"15",X"15",X"15",X"18",X"10",X"10",X"10",X"12",X"12",X"12",X"15",X"15",
		X"15",X"15",X"18",X"18",X"18",X"18",X"18",X"20",X"00",X"08",X"08",X"04",X"04",X"02",X"02",X"04",
		X"04",X"08",X"08",X"04",X"04",X"08",X"08",X"01",X"01",X"08",X"08",X"01",X"01",X"08",X"08",X"04",
		X"04",X"08",X"08",X"01",X"01",X"08",X"08",X"04",X"04",X"08",X"08",X"04",X"04",X"02",X"02",X"04",
		X"04",X"08",X"08",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"02",X"02",X"02",X"04",X"04",
		X"04",X"08",X"08",X"01",X"01",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"02",X"02",X"02",X"01",
		X"01",X"02",X"02",X"04",X"04",X"04",X"08",X"08",X"08",X"02",X"02",X"02",X"02",X"02",X"01",X"01",
		X"08",X"08",X"01",X"01",X"02",X"02",X"01",X"01",X"01",X"08",X"08",X"04",X"04",X"08",X"08",X"01",
		X"01",X"01",X"01",X"01",X"02",X"02",X"04",X"04",X"02",X"02",X"01",X"01",X"01",X"08",X"08",X"01",
		X"01",X"02",X"02",X"01",X"01",X"08",X"08",X"08",X"08",X"08",X"08",X"04",X"04",X"02",X"02",X"02",
		X"04",X"04",X"08",X"08",X"04",X"04",X"08",X"08",X"01",X"01",X"08",X"08",X"01",X"01",X"01",X"08",
		X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"01",
		X"01",X"01",X"08",X"08",X"08",X"04",X"04",X"08",X"08",X"01",X"01",X"02",X"02",X"01",X"01",X"08",
		X"08",X"08",X"08",X"FF",X"1C",X"D1",X"1E",X"D1",X"21",X"D1",X"23",X"D1",X"25",X"D1",X"28",X"D1",
		X"FF",X"D1",X"FF",X"1B",X"D1",X"1D",X"D1",X"1F",X"D1",X"20",X"D1",X"22",X"D1",X"24",X"D1",X"26",
		X"D1",X"27",X"D1",X"FF",X"D1",X"FF",X"27",X"D1",X"26",X"D1",X"24",X"D1",X"22",X"D1",X"20",X"D1",
		X"1F",X"D1",X"1D",X"D1",X"1B",X"D1",X"FF",X"D1",X"FF",X"1B",X"E2",X"1D",X"F1",X"1B",X"E2",X"1D",
		X"F1",X"27",X"D0",X"FF",X"C1",X"D1",X"41",X"D1",X"00",X"DF",X"FF",X"03",X"E1",X"0A",X"E2",X"FF",
		X"27",X"E0",X"29",X"D0",X"2B",X"D0",X"2C",X"E0",X"2C",X"D2",X"FF",X"EF",X"2E",X"A1",X"00",X"EF",
		X"2E",X"D1",X"00",X"EF",X"2E",X"D1",X"00",X"EF",X"2E",X"D1",X"00",X"EF",X"2E",X"A1",X"00",X"EF",
		X"2E",X"D1",X"00",X"EF",X"2E",X"D1",X"00",X"EF",X"2E",X"D1",X"00",X"EF",X"2E",X"A1",X"00",X"EF",
		X"FF",X"18",X"A2",X"18",X"E2",X"16",X"D2",X"16",X"E2",X"18",X"A2",X"18",X"E2",X"16",X"D2",X"16",
		X"E2",X"18",X"B2",X"1A",X"D2",X"1A",X"E2",X"1B",X"D2",X"1B",X"E2",X"1B",X"92",X"1A",X"C1",X"1A",
		X"E1",X"00",X"EF",X"1A",X"D1",X"1A",X"E1",X"18",X"D1",X"18",X"E1",X"1A",X"D1",X"1A",X"E1",X"1B",
		X"B1",X"1D",X"D1",X"1D",X"E1",X"1D",X"71",X"FF",X"14",X"A4",X"14",X"E4",X"13",X"D4",X"13",X"E4",
		X"14",X"A4",X"14",X"E4",X"13",X"D4",X"13",X"E4",X"14",X"B4",X"16",X"D4",X"16",X"E4",X"18",X"D4",
		X"18",X"E4",X"18",X"94",X"16",X"C4",X"16",X"E4",X"00",X"EF",X"16",X"D4",X"16",X"E4",X"15",X"D4",
		X"15",X"E4",X"16",X"D4",X"16",X"E4",X"18",X"B4",X"1A",X"D4",X"1A",X"E4",X"1A",X"74",X"FF",X"08",
		X"A4",X"00",X"EF",X"08",X"D4",X"00",X"EF",X"08",X"94",X"08",X"A4",X"00",X"EF",X"08",X"D4",X"00",
		X"EF",X"08",X"94",X"0A",X"A4",X"00",X"EF",X"0A",X"D4",X"00",X"EF",X"0A",X"94",X"0A",X"A4",X"00",
		X"EF",X"0A",X"D4",X"00",X"EF",X"0A",X"94",X"FF",X"08",X"A4",X"00",X"EF",X"08",X"D4",X"00",X"EF",
		X"08",X"94",X"08",X"A4",X"00",X"EF",X"08",X"D4",X"00",X"EF",X"08",X"94",X"0A",X"A4",X"00",X"EF",
		X"0A",X"D4",X"00",X"EF",X"0A",X"94",X"0A",X"A4",X"00",X"EF",X"0A",X"D4",X"00",X"EF",X"0A",X"94",
		X"FF",X"27",X"C1",X"1B",X"C1",X"1F",X"C1",X"22",X"C1",X"27",X"C1",X"2B",X"C1",X"27",X"C1",X"FF",
		X"0F",X"C1",X"16",X"C1",X"1B",X"C1",X"1F",X"C1",X"13",X"C1",X"22",X"C1",X"1F",X"C1",X"FF",X"22",
		X"C1",X"20",X"C1",X"1F",X"C1",X"1D",X"C1",X"1B",X"C1",X"1A",X"C1",X"1B",X"A1",X"FF",X"1F",X"C1",
		X"1D",X"0C",X"1B",X"0C",X"1A",X"C1",X"18",X"C1",X"16",X"C1",X"18",X"A1",X"FF",X"1B",X"D1",X"1D",
		X"D1",X"1F",X"D1",X"20",X"D1",X"22",X"D1",X"24",X"D1",X"26",X"D1",X"27",X"D1",X"FF",X"27",X"D1",
		X"26",X"D1",X"24",X"D1",X"22",X"D1",X"20",X"D1",X"1F",X"D1",X"1D",X"D1",X"1B",X"D1",X"FF",X"1F",
		X"92",X"1D",X"C2",X"1F",X"92",X"1D",X"C2",X"1B",X"D2",X"1B",X"E2",X"00",X"EF",X"1B",X"A2",X"1A",
		X"C2",X"18",X"92",X"18",X"D2",X"18",X"E2",X"00",X"EF",X"18",X"B2",X"18",X"E2",X"00",X"EF",X"18",
		X"A2",X"1B",X"C2",X"1F",X"A2",X"1D",X"C2",X"1D",X"42",X"FF",X"E1",X"00",X"03",X"A4",X"03",X"D4",
		X"03",X"E4",X"00",X"EF",X"03",X"D4",X"03",X"E4",X"00",X"EF",X"07",X"84",X"0C",X"A4",X"0C",X"D4",
		X"0C",X"E4",X"00",X"EF",X"0C",X"D4",X"0C",X"E4",X"00",X"EF",X"0C",X"84",X"FF",X"1B",X"81",X"18",
		X"A2",X"1B",X"D2",X"1B",X"E2",X"00",X"EF",X"1B",X"D2",X"1B",X"E2",X"00",X"EF",X"1B",X"D2",X"1B",
		X"E2",X"00",X"EF",X"1B",X"C2",X"18",X"C2",X"16",X"C2",X"18",X"C2",X"16",X"C2",X"13",X"D2",X"13",
		X"E2",X"00",X"EF",X"13",X"D2",X"13",X"E2",X"00",X"EF",X"13",X"82",X"11",X"B2",X"11",X"E2",X"00",
		X"EF",X"11",X"D2",X"11",X"E2",X"00",X"EF",X"11",X"D2",X"11",X"E2",X"00",X"EF",X"11",X"D2",X"11",
		X"E2",X"00",X"EF",X"11",X"B2",X"11",X"E2",X"00",X"EF",X"11",X"C2",X"16",X"D2",X"16",X"E2",X"00",
		X"EF",X"16",X"C2",X"18",X"C2",X"16",X"D2",X"16",X"E2",X"00",X"EF",X"16",X"82",X"FF",X"B1",X"18",
		X"08",X"A4",X"08",X"D4",X"08",X"E4",X"00",X"EF",X"08",X"D4",X"08",X"E4",X"00",X"EF",X"08",X"84",
		X"03",X"A4",X"03",X"D4",X"03",X"E4",X"00",X"EF",X"03",X"D4",X"03",X"E4",X"00",X"EF",X"03",X"84",
		X"05",X"A4",X"05",X"D4",X"05",X"E4",X"00",X"EF",X"05",X"D4",X"05",X"E4",X"00",X"EF",X"05",X"84",
		X"0A",X"A4",X"0A",X"D4",X"0A",X"E4",X"00",X"EF",X"0A",X"D4",X"0A",X"E4",X"00",X"EF",X"0A",X"84",
		X"FF",X"11",X"E1",X"1B",X"D0",X"00",X"CF",X"18",X"D0",X"00",X"CF",X"14",X"D0",X"00",X"CF",X"0F",
		X"D0",X"00",X"CF",X"11",X"B2",X"13",X"B1",X"14",X"B0",X"13",X"D0",X"11",X"D1",X"0F",X"D2",X"0E",
		X"D3",X"0C",X"D4",X"0A",X"D5",X"08",X"A0",X"24",X"C4",X"25",X"C2",X"24",X"C1",X"25",X"C2",X"24",
		X"C4",X"25",X"C8",X"24",X"C4",X"25",X"C2",X"24",X"C1",X"25",X"C2",X"24",X"C4",X"25",X"C8",X"24",
		X"C4",X"25",X"C2",X"24",X"C1",X"25",X"C2",X"24",X"C4",X"25",X"C8",X"FF",X"A1",X"14",X"A1",X"16",
		X"A1",X"18",X"C0",X"16",X"18",X"D0",X"00",X"CF",X"14",X"D0",X"00",X"CF",X"11",X"D0",X"00",X"CF",
		X"0C",X"D0",X"00",X"CF",X"0E",X"B2",X"0F",X"B1",X"11",X"B0",X"0F",X"D0",X"0E",X"D1",X"0C",X"D2",
		X"0A",X"D3",X"08",X"D4",X"07",X"D5",X"05",X"A0",X"27",X"C4",X"28",X"C2",X"27",X"C1",X"28",X"C2",
		X"27",X"C4",X"28",X"C8",X"27",X"C4",X"28",X"C2",X"27",X"C1",X"28",X"C2",X"27",X"C4",X"28",X"C8",
		X"27",X"C4",X"28",X"C2",X"27",X"C1",X"28",X"C2",X"27",X"C4",X"28",X"C8",X"FF",X"1F",X"A1",X"1D",
		X"C1",X"1D",X"41",X"FF",X"0E",X"17",X"F0",X"16",X"F0",X"15",X"F0",X"14",X"F0",X"16",X"F0",X"15",
		X"F0",X"14",X"F0",X"13",X"F0",X"15",X"F0",X"14",X"F0",X"13",X"F0",X"12",X"F0",X"14",X"F0",X"13",
		X"F0",X"12",X"F0",X"11",X"F0",X"13",X"F0",X"12",X"F0",X"11",X"F0",X"10",X"F0",X"12",X"F0",X"11",
		X"F0",X"10",X"F0",X"0F",X"F0",X"11",X"F0",X"10",X"F0",X"0F",X"F0",X"0E",X"F0",X"10",X"F0",X"0F",
		X"F0",X"0E",X"F0",X"0D",X"F0",X"0F",X"F0",X"0E",X"F0",X"0D",X"F0",X"0C",X"F0",X"0E",X"F0",X"0D",
		X"F0",X"0C",X"F0",X"0B",X"F0",X"FF",X"13",X"F0",X"12",X"F0",X"11",X"F0",X"10",X"F0",X"12",X"F0",
		X"11",X"F0",X"10",X"F0",X"0F",X"F0",X"11",X"F0",X"10",X"F0",X"0F",X"F0",X"0E",X"F0",X"10",X"F0",
		X"0F",X"F0",X"0E",X"F0",X"0D",X"F0",X"0F",X"F0",X"0E",X"F0",X"0D",X"F0",X"0C",X"F0",X"0E",X"F0",
		X"0D",X"F0",X"0C",X"F0",X"0B",X"F0",X"0D",X"F0",X"0C",X"F0",X"0B",X"F0",X"0A",X"F0",X"0C",X"F0",
		X"0B",X"F0",X"0A",X"F0",X"09",X"F0",X"0B",X"F0",X"0A",X"F0",X"09",X"F0",X"08",X"F0",X"0A",X"F0",
		X"09",X"F0",X"08",X"F0",X"07",X"F0",X"FF",X"20",X"D1",X"22",X"D1",X"24",X"D1",X"27",X"D1",X"29",
		X"D1",X"27",X"D1",X"24",X"D1",X"22",X"D1",X"20",X"D1",X"00",X"AF",X"1B",X"C0",X"00",X"CF",X"16",
		X"C1",X"00",X"CF",X"1B",X"C0",X"00",X"CF",X"16",X"C1",X"00",X"CF",X"1F",X"B0",X"1D",X"D1",X"1B",
		X"D0",X"1B",X"D0",X"1B",X"D0",X"16",X"D0",X"18",X"C1",X"1A",X"C1",X"1B",X"C1",X"1D",X"C1",X"1F",
		X"C0",X"00",X"CF",X"21",X"C0",X"00",X"CF",X"22",X"C0",X"00",X"9F",X"22",X"D0",X"24",X"D0",X"00",
		X"CF",X"24",X"D0",X"26",X"D0",X"00",X"CF",X"26",X"D0",X"27",X"D0",X"FF",X"15",X"E8",X"00",X"EF",
		X"15",X"B8",X"15",X"E8",X"00",X"EF",X"15",X"C8",X"18",X"A8",X"1B",X"D8",X"1B",X"E8",X"00",X"EF",
		X"1B",X"68",X"1A",X"68",X"FF",X"00",X"4F",X"00",X"4F",X"00",X"4F",X"00",X"4F",X"0F",X"68",X"0E",
		X"68",X"0C",X"68",X"0E",X"68",X"0F",X"88",X"0F",X"21",X"D1",X"23",X"D1",X"25",X"D1",X"28",X"D1",
		X"2A",X"D1",X"28",X"D1",X"25",X"D1",X"23",X"D1",X"21",X"D1",X"00",X"AF",X"0A",X"C0",X"00",X"CF",
		X"0F",X"C1",X"00",X"CF",X"0A",X"C0",X"00",X"CF",X"0F",X"C1",X"00",X"CF",X"16",X"B0",X"14",X"D1",
		X"13",X"D0",X"13",X"D0",X"13",X"D0",X"0F",X"D0",X"14",X"C1",X"11",X"C1",X"13",X"C1",X"14",X"C1",
		X"0F",X"C0",X"00",X"CF",X"11",X"C0",X"00",X"CF",X"16",X"C0",X"00",X"9F",X"16",X"D0",X"14",X"D0",
		X"00",X"CF",X"14",X"D0",X"11",X"D0",X"00",X"CF",X"11",X"D0",X"0F",X"D0",X"FF",X"00",X"EF",X"11",
		X"C8",X"0F",X"C8",X"11",X"C8",X"13",X"A8",X"14",X"C8",X"14",X"68",X"16",X"98",X"13",X"C8",X"17",
		X"98",X"13",X"D8",X"13",X"E8",X"00",X"EF",X"13",X"D8",X"13",X"E8",X"00",X"EF",X"13",X"A8",X"0F",
		X"88",X"11",X"C8",X"11",X"B8",X"11",X"E8",X"00",X"EF",X"00",X"F2",X"03",X"F2",X"06",X"F2",X"09",
		X"F2",X"0C",X"F2",X"0F",X"F2",X"12",X"F2",X"15",X"F2",X"18",X"F2",X"1B",X"F2",X"1E",X"F2",X"21",
		X"F2",X"24",X"F2",X"27",X"F2",X"2A",X"F2",X"FF",X"03",X"F2",X"06",X"F2",X"09",X"F2",X"0C",X"F2",
		X"0F",X"F2",X"12",X"F2",X"15",X"F2",X"18",X"F2",X"1B",X"F2",X"1E",X"F2",X"21",X"F2",X"24",X"F2",
		X"27",X"F2",X"2A",X"F2",X"2D",X"F2",X"FF",X"03",X"F0",X"04",X"F0",X"05",X"F0",X"06",X"F0",X"07",
		X"F0",X"08",X"F0",X"09",X"F0",X"0A",X"F0",X"0B",X"F0",X"0C",X"F0",X"0D",X"F0",X"0E",X"F0",X"09",
		X"F0",X"0A",X"F0",X"0B",X"F0",X"0C",X"F0",X"0D",X"F0",X"0E",X"F0",X"0F",X"F0",X"10",X"F0",X"11",
		X"F0",X"12",X"F0",X"13",X"F0",X"14",X"F0",X"0F",X"F0",X"10",X"F0",X"11",X"F0",X"12",X"F0",X"13",
		X"F0",X"14",X"F0",X"15",X"F0",X"16",X"F0",X"17",X"F0",X"18",X"F0",X"19",X"F0",X"1A",X"F0",X"15",
		X"F0",X"16",X"F0",X"17",X"F0",X"18",X"F0",X"19",X"F0",X"1A",X"F0",X"1B",X"F0",X"1C",X"F0",X"1D",
		X"F0",X"1E",X"F0",X"1F",X"F0",X"20",X"F0",X"1B",X"F0",X"1C",X"F0",X"1D",X"F0",X"1E",X"F0",X"1F",
		X"F0",X"20",X"F0",X"21",X"F0",X"22",X"F0",X"23",X"F0",X"24",X"F0",X"25",X"F0",X"26",X"F0",X"21",
		X"F0",X"22",X"F0",X"23",X"F0",X"24",X"F0",X"25",X"F0",X"26",X"F0",X"27",X"F0",X"28",X"F0",X"29",
		X"F0",X"2A",X"F0",X"2B",X"F0",X"2C",X"F0",X"27",X"F0",X"28",X"F0",X"29",X"F0",X"2A",X"F0",X"2B",
		X"F0",X"2C",X"F0",X"2D",X"F0",X"2E",X"F0",X"2F",X"F0",X"30",X"F0",X"31",X"F0",X"32",X"F0",X"FF",
		X"00",X"EF",X"FF",X"EF",X"03",X"D4",X"03",X"E4",X"00",X"EF",X"03",X"C4",X"05",X"C4",X"07",X"A4",
		X"08",X"A8",X"08",X"D8",X"08",X"E8",X"00",X"EF",X"08",X"D8",X"08",X"E8",X"00",X"EF",X"08",X"98",
		X"08",X"D8",X"08",X"E8",X"00",X"EF",X"08",X"A8",X"08",X"D8",X"08",X"E8",X"00",X"EF",X"08",X"D8",
		X"08",X"E8",X"00",X"EF",X"08",X"88",X"03",X"A8",X"03",X"D8",X"03",X"E8",X"00",X"EF",X"03",X"D8",
		X"03",X"E8",X"00",X"EF",X"03",X"98",X"03",X"D8",X"03",X"E8",X"00",X"EF",X"03",X"A8",X"03",X"D8",
		X"03",X"00",X"EF",X"FF",X"03",X"D8",X"03",X"E8",X"00",X"EF",X"03",X"88",X"08",X"A8",X"08",X"D8",
		X"08",X"E8",X"00",X"EF",X"08",X"D8",X"08",X"E8",X"00",X"EF",X"08",X"98",X"08",X"D8",X"08",X"E8",
		X"00",X"EF",X"08",X"A8",X"08",X"D8",X"08",X"E8",X"00",X"EF",X"08",X"D8",X"08",X"E8",X"00",X"EF",
		X"08",X"88",X"0A",X"A8",X"0A",X"D8",X"0A",X"E8",X"00",X"EF",X"0A",X"D8",X"0A",X"E8",X"00",X"EF",
		X"0A",X"98",X"0A",X"D8",X"0A",X"E8",X"00",X"EF",X"0A",X"A8",X"0A",X"D8",X"0A",X"E8",X"00",X"EF",
		X"0A",X"D8",X"03",X"A4",X"03",X"D4",X"03",X"E4",X"00",X"EF",X"03",X"D4",X"03",X"E4",X"00",X"EF",
		X"07",X"84",X"0C",X"A4",X"0C",X"D4",X"0C",X"E4",X"00",X"EF",X"0C",X"D4",X"0C",X"E4",X"00",X"EF",
		X"0C",X"84",X"05",X"B4",X"05",X"E4",X"00",X"EF",X"05",X"B4",X"05",X"E4",X"00",X"EF",X"05",X"D4",
		X"05",X"E4",X"00",X"EF",X"05",X"B4",X"05",X"E4",X"00",X"EF",X"05",X"C4",X"0A",X"B4",X"0A",X"E4",
		X"00",X"EF",X"0A",X"B4",X"0A",X"E4",X"00",X"EF",X"0A",X"B4",X"0A",X"E4",X"00",X"EF",X"0A",X"B4",
		X"0A",X"E4",X"00",X"EF",X"0A",X"D4",X"0A",X"E4",X"00",X"EF",X"0A",X"B4",X"0A",X"E4",X"00",X"EF",
		X"0A",X"D4",X"0A",X"E4",X"00",X"EF",X"0A",X"84",X"FF",X"E8",X"00",X"EF",X"0A",X"88",X"FF",X"27",
		X"E0",X"29",X"D0",X"2B",X"D0",X"2C",X"E0",X"2C",X"D2",X"FF",X"03",X"C1",X"05",X"C1",X"C1",X"A1",
		X"FF",X"18",X"B0",X"FF",X"04",X"D1",X"00",X"DF",X"04",X"D1",X"00",X"DF",X"04",X"D1",X"00",X"DF",
		X"00",X"B1",X"FF",X"1C",X"D1",X"00",X"DF",X"1C",X"D1",X"00",X"DF",X"1C",X"D1",X"00",X"DF",X"18",
		X"B1",X"FF",X"0A",X"B2",X"0C",X"B4",X"0A",X"B2",X"0C",X"B4",X"0A",X"C2",X"00",X"CF",X"0E",X"C4",
		X"00",X"CF",X"0F",X"B8",X"00",X"BF",X"0F",X"91",X"FF",X"00",X"5F",X"00",X"CF",X"13",X"91",X"FF",
		X"00",X"5F",X"00",X"CF",X"16",X"91",X"FF",X"00",X"DF",X"00",X"EF",X"03",X"B1",X"00",X"BF",X"13",
		X"D4",X"13",X"E4",X"00",X"DF",X"00",X"EF",X"13",X"D4",X"13",X"E4",X"00",X"DF",X"00",X"EF",X"0F",
		X"B4",X"00",X"BF",X"0A",X"D1",X"0A",X"E1",X"00",X"DF",X"00",X"EF",X"0A",X"D1",X"0A",X"E1",X"FF",
		X"00",X"DF",X"0F",X"C1",X"00",X"CF",X"1F",X"D4",X"00",X"DF",X"1F",X"D4",X"00",X"DF",X"1B",X"C4",
		X"00",X"CF",X"16",X"D1",X"00",X"DF",X"16",X"D1",X"FF",X"00",X"EF",X"1B",X"D1",X"00",X"DF",X"2B",
		X"E4",X"00",X"EF",X"2B",X"E4",X"00",X"EF",X"27",X"D4",X"00",X"DF",X"22",X"E1",X"00",X"EF",X"22",
		X"E1",X"FF",X"C5",X"47",X"3E",X"01",X"05",X"28",X"05",X"CB",X"27",X"C3",X"36",X"17",X"C1",X"C9",
		X"D5",X"F5",X"78",X"3D",X"5F",X"CB",X"27",X"83",X"DD",X"21",X"04",X"60",X"5F",X"16",X"00",X"DD",
		X"19",X"F1",X"D1",X"C9",X"C9",X"21",X"00",X"70",X"06",X"04",X"0E",X"00",X"C5",X"06",X"FF",X"3A",
		X"01",X"90",X"CB",X"77",X"20",X"F9",X"71",X"23",X"10",X"F5",X"C1",X"10",X"EF",X"C9",X"3E",X"9F",
		X"32",X"00",X"B0",X"32",X"00",X"C0",X"3E",X"BF",X"32",X"00",X"B0",X"32",X"00",X"C0",X"3E",X"DF",
		X"32",X"00",X"B0",X"32",X"00",X"C0",X"3E",X"FF",X"32",X"00",X"B0",X"32",X"00",X"C0",X"C9",X"21",
		X"5F",X"60",X"CB",X"66",X"CA",X"A1",X"17",X"21",X"00",X"60",X"AF",X"77",X"23",X"77",X"23",X"77",
		X"C9",X"DD",X"E5",X"21",X"00",X"60",X"7E",X"E6",X"FF",X"C2",X"E5",X"17",X"23",X"7E",X"E6",X"FF",
		X"C2",X"D0",X"17",X"23",X"7E",X"E6",X"FF",X"CA",X"BF",X"18",X"06",X"10",X"CB",X"1F",X"D2",X"C4",
		X"17",X"CD",X"FA",X"17",X"04",X"08",X"78",X"FE",X"18",X"CA",X"BF",X"18",X"08",X"C3",X"BC",X"17",
		X"06",X"08",X"CB",X"1F",X"D2",X"DA",X"17",X"CD",X"FA",X"17",X"04",X"08",X"78",X"FE",X"10",X"28",
		X"D2",X"08",X"C3",X"D2",X"17",X"06",X"00",X"CB",X"1F",X"D2",X"EF",X"17",X"CD",X"FA",X"17",X"04",
		X"08",X"78",X"FE",X"08",X"28",X"B6",X"08",X"C3",X"E7",X"17",X"C5",X"F5",X"E5",X"21",X"6D",X"1B",
		X"CB",X"20",X"48",X"06",X"00",X"09",X"46",X"23",X"4E",X"68",X"61",X"46",X"23",X"4F",X"78",X"E6",
		X"FF",X"CA",X"AF",X"18",X"79",X"5E",X"23",X"56",X"23",X"DD",X"21",X"03",X"60",X"1A",X"E6",X"C0",
		X"CA",X"46",X"18",X"DD",X"7E",X"00",X"CB",X"77",X"20",X"0C",X"ED",X"53",X"16",X"60",X"DD",X"CB",
		X"00",X"F6",X"05",X"C3",X"0D",X"18",X"05",X"CB",X"7F",X"20",X"D2",X"ED",X"53",X"19",X"60",X"DD",
		X"CB",X"00",X"FE",X"C3",X"0D",X"18",X"DD",X"7E",X"00",X"CB",X"47",X"C2",X"5A",X"18",X"ED",X"53",
		X"04",X"60",X"DD",X"CB",X"00",X"C6",X"05",X"C3",X"0D",X"18",X"CB",X"4F",X"C2",X"6B",X"18",X"ED",
		X"53",X"07",X"60",X"DD",X"CB",X"00",X"CE",X"05",X"C3",X"0D",X"18",X"CB",X"57",X"C2",X"7C",X"18",
		X"ED",X"53",X"0A",X"60",X"DD",X"CB",X"00",X"D6",X"05",X"C3",X"0D",X"18",X"CB",X"5F",X"C2",X"8D",
		X"18",X"ED",X"53",X"0D",X"60",X"DD",X"CB",X"00",X"DE",X"05",X"C3",X"0D",X"18",X"CB",X"67",X"C2",
		X"9E",X"18",X"ED",X"53",X"10",X"60",X"DD",X"CB",X"00",X"E6",X"05",X"C3",X"0D",X"18",X"05",X"CB",
		X"6F",X"C2",X"0D",X"18",X"ED",X"53",X"13",X"60",X"DD",X"CB",X"00",X"EE",X"C3",X"0D",X"18",X"E1",
		X"F1",X"C1",X"08",X"78",X"E6",X"07",X"3C",X"CD",X"32",X"17",X"2F",X"A6",X"77",X"08",X"C9",X"3A",
		X"03",X"60",X"06",X"06",X"DD",X"21",X"04",X"60",X"CB",X"3F",X"DA",X"DA",X"18",X"DD",X"23",X"DD",
		X"23",X"DD",X"23",X"05",X"CA",X"CF",X"19",X"C3",X"C8",X"18",X"08",X"DD",X"7E",X"02",X"FE",X"00",
		X"28",X"07",X"DD",X"35",X"02",X"08",X"C3",X"CD",X"18",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7E",
		X"FE",X"FF",X"C2",X"3E",X"19",X"3E",X"06",X"90",X"FE",X"03",X"38",X"14",X"D6",X"03",X"CB",X"27",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"F6",X"9F",X"32",X"00",X"C0",X"C3",X"1F",X"19",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"F6",X"9F",X"32",X"00",X"B0",X"3E",
		X"06",X"90",X"57",X"1E",X"01",X"7A",X"FE",X"00",X"28",X"06",X"15",X"CB",X"23",X"C3",X"25",X"19",
		X"7B",X"2F",X"5F",X"3A",X"03",X"60",X"A3",X"32",X"03",X"60",X"08",X"C3",X"CD",X"18",X"3E",X"06",
		X"90",X"FE",X"03",X"FA",X"9A",X"19",X"D6",X"03",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"CB",X"27",X"F6",X"80",X"4F",X"FD",X"21",X"07",X"1B",X"7E",X"E6",X"3F",X"CB",X"27",X"5F",X"16",
		X"00",X"FD",X"19",X"FD",X"7E",X"00",X"B1",X"32",X"00",X"C0",X"FD",X"7E",X"01",X"32",X"00",X"C0",
		X"23",X"3E",X"00",X"ED",X"67",X"B1",X"CB",X"E7",X"32",X"00",X"C0",X"3E",X"00",X"ED",X"6F",X"FD",
		X"21",X"F7",X"1A",X"23",X"DD",X"75",X"00",X"DD",X"74",X"01",X"5F",X"16",X"00",X"FD",X"19",X"FD",
		X"7E",X"00",X"3D",X"DD",X"77",X"02",X"08",X"C3",X"CD",X"18",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"CB",X"27",X"CB",X"27",X"F6",X"80",X"4F",X"FD",X"21",X"07",X"1B",X"7E",X"E6",X"3F",X"CB",X"27",
		X"5F",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"B1",X"32",X"00",X"B0",X"FD",X"7E",X"01",X"32",
		X"00",X"B0",X"23",X"AF",X"ED",X"67",X"B1",X"CB",X"E7",X"32",X"00",X"B0",X"C3",X"7B",X"19",X"CB",
		X"3F",X"38",X"0D",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"CB",X"3F",X"38",X"72",X"C3",X"B7",X"1A",
		X"08",X"DD",X"7E",X"02",X"FE",X"00",X"28",X"07",X"DD",X"35",X"02",X"08",X"C3",X"D3",X"19",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"7E",X"FE",X"FF",X"20",X"11",X"3E",X"FF",X"32",X"00",X"B0",X"3A",
		X"03",X"60",X"E6",X"BF",X"32",X"03",X"60",X"08",X"C3",X"D3",X"19",X"06",X"00",X"CB",X"3F",X"CB",
		X"10",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3D",X"CB",X"20",X"CB",X"20",
		X"B0",X"F6",X"E0",X"32",X"00",X"B0",X"23",X"3E",X"00",X"ED",X"67",X"F6",X"F0",X"32",X"00",X"B0",
		X"3E",X"00",X"ED",X"6F",X"FD",X"21",X"F7",X"1A",X"23",X"DD",X"75",X"00",X"DD",X"74",X"01",X"5F",
		X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"3D",X"DD",X"77",X"02",X"08",X"C3",X"D3",X"19",X"DD",
		X"7E",X"02",X"FE",X"00",X"28",X"06",X"DD",X"35",X"02",X"C3",X"B7",X"1A",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"7E",X"FE",X"FF",X"20",X"10",X"3E",X"FF",X"32",X"00",X"C0",X"3A",X"03",X"60",X"E6",
		X"7F",X"32",X"03",X"60",X"C3",X"B7",X"1A",X"06",X"00",X"CB",X"3F",X"CB",X"10",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3D",X"CB",X"20",X"CB",X"20",X"B0",X"F6",X"E0",X"32",
		X"00",X"C0",X"23",X"3E",X"00",X"ED",X"67",X"F6",X"F0",X"32",X"00",X"C0",X"3E",X"00",X"ED",X"6F",
		X"FD",X"21",X"F7",X"1A",X"23",X"DD",X"75",X"00",X"DD",X"74",X"01",X"5F",X"16",X"00",X"FD",X"19",
		X"FD",X"7E",X"00",X"3D",X"DD",X"77",X"02",X"DD",X"E1",X"C9",X"E5",X"F5",X"C5",X"21",X"80",X"D0",
		X"3E",X"FF",X"0E",X"18",X"23",X"06",X"1E",X"77",X"23",X"10",X"FC",X"23",X"0D",X"C2",X"C4",X"1A",
		X"C1",X"F1",X"E1",X"C9",X"3E",X"00",X"06",X"80",X"21",X"00",X"D0",X"77",X"23",X"10",X"FC",X"0E",
		X"00",X"06",X"18",X"77",X"11",X"20",X"00",X"19",X"10",X"F9",X"0C",X"0D",X"C2",X"F6",X"1A",X"0C",
		X"21",X"9F",X"D0",X"C3",X"E1",X"1A",X"C9",X"FF",X"E0",X"C0",X"A0",X"80",X"60",X"40",X"30",X"20",
		X"18",X"10",X"0C",X"08",X"04",X"02",X"01",X"08",X"3F",X"0F",X"3B",X"09",X"38",X"06",X"35",X"06",
		X"32",X"0A",X"2F",X"0E",X"2C",X"06",X"2A",X"00",X"28",X"0C",X"25",X"0A",X"23",X"0A",X"21",X"0C",
		X"1F",X"0F",X"1D",X"04",X"1C",X"0B",X"1A",X"03",X"19",X"0D",X"17",X"07",X"16",X"03",X"15",X"00",
		X"14",X"0E",X"12",X"0D",X"11",X"0D",X"10",X"0E",X"0F",X"00",X"0F",X"02",X"0E",X"06",X"0D",X"0A",
		X"0C",X"0E",X"0B",X"04",X"0B",X"0A",X"0A",X"00",X"0A",X"07",X"09",X"0F",X"08",X"07",X"08",X"0F",
		X"07",X"08",X"07",X"01",X"07",X"0B",X"06",X"05",X"06",X"0F",X"05",X"0A",X"05",X"05",X"05",X"00",
		X"05",X"0B",X"04",X"07",X"04",X"03",X"04",X"0F",X"03",X"0C",X"03",X"09",X"03",X"91",X"1B",X"D1",
		X"1B",X"D6",X"1B",X"9C",X"1B",X"9F",X"1B",X"DB",X"1B",X"A5",X"1B",X"AE",X"1B",X"AE",X"1B",X"B8",
		X"1B",X"BD",X"1B",X"C2",X"1B",X"A2",X"1B",X"C7",X"1B",X"99",X"1B",X"CC",X"1B",X"DE",X"1B",X"DE",
		X"1B",X"01",X"B4",X"0F",X"02",X"C3",X"0F",X"D6",X"0F",X"01",X"E9",X"0F",X"01",X"F4",X"0F",X"01",
		X"FB",X"0F",X"01",X"00",X"10",X"04",X"31",X"10",X"68",X"10",X"9F",X"10",X"C8",X"10",X"02",X"F1",
		X"10",X"00",X"11",X"02",X"0F",X"11",X"1E",X"11",X"02",X"2D",X"11",X"3E",X"11",X"02",X"4F",X"11",
		X"12",X"16",X"02",X"9F",X"11",X"00",X"12",X"02",X"43",X"12",X"94",X"12",X"02",X"E5",X"12",X"36",
		X"13",X"02",X"87",X"13",X"08",X"14",X"02",X"89",X"14",X"A8",X"14",X"01",X"C7",X"14",X"02",X"70",
		X"15",X"C1",X"15",X"19",X"17",X"06",X"03",X"0E",X"00",X"C5",X"06",X"00",X"CD",X"FC",X"1B",X"C1",
		X"10",X"02",X"18",X"04",X"0C",X"C5",X"18",X"F2",X"CD",X"6A",X"1C",X"C9",X"DD",X"21",X"55",X"0C",
		X"16",X"00",X"78",X"FE",X"02",X"20",X"02",X"1E",X"02",X"79",X"CB",X"27",X"CB",X"27",X"D5",X"16",
		X"00",X"5F",X"DD",X"19",X"D1",X"DD",X"5E",X"00",X"C5",X"DD",X"46",X"03",X"CB",X"38",X"CB",X"38",
		X"CB",X"38",X"CB",X"38",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"73",X"D5",X"11",X"20",X"00",X"19",
		X"D1",X"10",X"F7",X"CB",X"42",X"20",X"15",X"14",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"23",X"DD",
		X"46",X"03",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"18",X"DE",X"C1",X"78",X"FE",X"00",
		X"20",X"17",X"04",X"C5",X"01",X"20",X"00",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"09",X"DD",X"7E",
		X"03",X"E6",X"0F",X"47",X"1E",X"03",X"C3",X"2A",X"1C",X"C9",X"01",X"00",X"00",X"21",X"9E",X"D0",
		X"3E",X"4B",X"77",X"DD",X"21",X"52",X"0C",X"DD",X"09",X"DD",X"46",X"00",X"CD",X"9B",X"1C",X"0C",
		X"79",X"FE",X"03",X"20",X"EB",X"21",X"9D",X"D0",X"DD",X"21",X"61",X"0C",X"06",X"18",X"11",X"20",
		X"00",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"19",X"10",X"F7",X"C9",X"3C",X"11",X"20",X"00",X"19",
		X"77",X"19",X"10",X"FC",X"C9",X"23",X"CB",X"7E",X"28",X"FC",X"CB",X"7E",X"20",X"FC",X"E5",X"CD",
		X"3A",X"03",X"CD",X"8F",X"17",X"E1",X"CB",X"7E",X"28",X"FC",X"C9",X"C5",X"47",X"3E",X"01",X"10",
		X"02",X"C1",X"C9",X"07",X"18",X"F7",X"16",X"00",X"3A",X"62",X"60",X"FE",X"00",X"28",X"04",X"1E",
		X"06",X"18",X"02",X"1E",X"05",X"0E",X"00",X"06",X"0C",X"21",X"1C",X"D6",X"73",X"CD",X"24",X"1D",
		X"04",X"3E",X"17",X"B8",X"20",X"0A",X"0C",X"3E",X"04",X"B9",X"20",X"02",X"0E",X"00",X"06",X"00",
		X"3E",X"00",X"B9",X"20",X"05",X"3E",X"0C",X"B8",X"28",X"1E",X"3A",X"60",X"60",X"B9",X"20",X"15",
		X"3A",X"61",X"60",X"B8",X"20",X"0F",X"22",X"63",X"60",X"14",X"3A",X"62",X"60",X"FE",X"00",X"28",
		X"03",X"1D",X"18",X"01",X"1C",X"C3",X"DC",X"1C",X"AF",X"BA",X"20",X"07",X"3A",X"62",X"60",X"2F",
		X"32",X"62",X"60",X"C9",X"D5",X"CB",X"41",X"28",X"0A",X"CB",X"49",X"28",X"03",X"23",X"18",X"10",
		X"2B",X"18",X"0D",X"CB",X"49",X"28",X"05",X"11",X"E0",X"FF",X"18",X"03",X"11",X"20",X"00",X"19",
		X"D1",X"C9",X"3E",X"52",X"0E",X"00",X"21",X"9C",X"D0",X"08",X"3E",X"4E",X"06",X"16",X"77",X"CD",
		X"24",X"1D",X"08",X"77",X"CD",X"24",X"1D",X"10",X"FA",X"FE",X"55",X"28",X"06",X"3C",X"08",X"3C",
		X"0C",X"18",X"E9",X"C9",X"11",X"20",X"00",X"21",X"A3",X"D4",X"3E",X"01",X"06",X"0C",X"77",X"E5",
		X"23",X"77",X"E1",X"19",X"10",X"F8",X"C9",X"11",X"20",X"00",X"3A",X"65",X"60",X"FE",X"00",X"28",
		X"05",X"3A",X"67",X"60",X"18",X"03",X"3A",X"66",X"60",X"FE",X"07",X"38",X"02",X"3E",X"06",X"47",
		X"AF",X"08",X"3E",X"06",X"90",X"4F",X"C5",X"21",X"A3",X"D0",X"3E",X"E1",X"32",X"C8",X"61",X"AF",
		X"B8",X"3A",X"C8",X"61",X"28",X"08",X"77",X"3C",X"19",X"77",X"3D",X"19",X"10",X"F8",X"3E",X"FF",
		X"41",X"CB",X"20",X"32",X"C8",X"61",X"AF",X"B8",X"3A",X"C8",X"61",X"28",X"04",X"77",X"19",X"10",
		X"FC",X"08",X"FE",X"FF",X"28",X"0A",X"2F",X"08",X"21",X"A4",X"D0",X"3E",X"E3",X"C1",X"18",X"CC",
		X"C9",X"AF",X"CD",X"4C",X"1E",X"11",X"20",X"00",X"3A",X"5F",X"60",X"CB",X"4F",X"28",X"13",X"21",
		X"43",X"D2",X"36",X"02",X"19",X"36",X"17",X"19",X"C3",X"31",X"49",X"DD",X"21",X"6B",X"60",X"CD",
		X"06",X"1E",X"21",X"44",X"D2",X"36",X"01",X"19",X"36",X"1C",X"19",X"C3",X"3A",X"49",X"DD",X"21",
		X"68",X"60",X"CD",X"06",X"1E",X"C9",X"D5",X"C5",X"E5",X"06",X"03",X"21",X"DA",X"61",X"E5",X"DD",
		X"7E",X"00",X"4F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"77",X"23",X"79",X"E6",X"0F",
		X"77",X"DD",X"23",X"23",X"10",X"E9",X"E1",X"06",X"05",X"AF",X"BE",X"20",X"05",X"36",X"FF",X"23",
		X"10",X"F8",X"E1",X"DD",X"E5",X"DD",X"21",X"DA",X"61",X"11",X"20",X"00",X"06",X"06",X"DD",X"7E",
		X"00",X"77",X"DD",X"23",X"19",X"10",X"F7",X"DD",X"E1",X"C1",X"D1",X"C9",X"F5",X"C5",X"E5",X"FE",
		X"00",X"20",X"14",X"3E",X"03",X"21",X"44",X"D6",X"06",X"0A",X"CD",X"7D",X"1E",X"21",X"43",X"D6",
		X"06",X"0A",X"CD",X"7D",X"1E",X"18",X"12",X"3A",X"65",X"60",X"FE",X"00",X"20",X"07",X"21",X"44",
		X"D6",X"3E",X"04",X"18",X"EB",X"3E",X"04",X"18",X"E4",X"E1",X"C1",X"F1",X"C9",X"C5",X"D5",X"E5",
		X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"E1",X"D1",X"C1",X"C9",X"21",X"E2",X"D4",X"3E",X"07",
		X"06",X"03",X"CD",X"7D",X"1E",X"21",X"E2",X"D0",X"36",X"1D",X"11",X"20",X"00",X"19",X"36",X"18",
		X"19",X"36",X"19",X"19",X"4F",X"06",X"01",X"CD",X"BD",X"25",X"C9",X"FF",X"FF",X"2F",X"1E",X"17",
		X"12",X"1F",X"0E",X"1B",X"1C",X"0A",X"15",X"06",X"09",X"21",X"80",X"D3",X"DD",X"21",X"AB",X"1E",
		X"C5",X"06",X"0C",X"DD",X"7E",X"00",X"77",X"23",X"DD",X"23",X"10",X"F7",X"C1",X"10",X"ED",X"06",
		X"09",X"21",X"73",X"60",X"36",X"01",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"10",X"F5",X"C9",
		X"21",X"A1",X"D1",X"11",X"20",X"00",X"36",X"19",X"19",X"36",X"0A",X"19",X"36",X"1B",X"19",X"36",
		X"1D",X"19",X"18",X"06",X"21",X"21",X"D2",X"11",X"20",X"00",X"CD",X"26",X"1F",X"FE",X"00",X"28",
		X"24",X"FE",X"64",X"38",X"08",X"36",X"09",X"19",X"36",X"09",X"C3",X"25",X"1F",X"06",X"00",X"0E",
		X"0A",X"B9",X"38",X"04",X"91",X"04",X"18",X"F9",X"08",X"AF",X"B8",X"28",X"03",X"70",X"18",X"02",
		X"36",X"FF",X"19",X"08",X"77",X"C9",X"3A",X"65",X"60",X"CB",X"4F",X"28",X"05",X"3A",X"6F",X"60",
		X"18",X"03",X"3A",X"6E",X"60",X"C9",X"3A",X"02",X"90",X"CB",X"7F",X"28",X"04",X"3E",X"03",X"18",
		X"02",X"3E",X"05",X"C9",X"CD",X"26",X"1F",X"FE",X"00",X"20",X"04",X"36",X"FF",X"18",X"2F",X"3D",
		X"FE",X"12",X"38",X"02",X"3E",X"11",X"16",X"00",X"5F",X"FD",X"21",X"79",X"0C",X"FD",X"19",X"11",
		X"20",X"00",X"FD",X"7E",X"00",X"4F",X"E6",X"F0",X"28",X"0A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"77",X"19",X"79",X"E6",X"0F",X"77",X"19",X"36",X"00",X"19",X"36",X"00",X"C9",X"DD",
		X"E5",X"CD",X"26",X"1F",X"FE",X"00",X"28",X"07",X"3D",X"FE",X"12",X"38",X"02",X"3E",X"11",X"DD",
		X"21",X"93",X"0C",X"4F",X"06",X"00",X"DD",X"09",X"DD",X"46",X"00",X"0E",X"00",X"CB",X"27",X"CB",
		X"27",X"81",X"DD",X"E1",X"C9",X"DD",X"7E",X"01",X"FE",X"07",X"D2",X"AF",X"1F",X"3E",X"07",X"D6",
		X"07",X"5F",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"E6",X"0F",X"08",X"7B",X"FE",X"0B",
		X"DA",X"C5",X"1F",X"1E",X"0B",X"08",X"C9",X"DD",X"E5",X"CD",X"7D",X"44",X"CD",X"5A",X"2D",X"21",
		X"01",X"90",X"CB",X"7E",X"CA",X"D2",X"1F",X"21",X"59",X"60",X"34",X"7E",X"21",X"5A",X"60",X"E6",
		X"07",X"20",X"01",X"34",X"CD",X"3A",X"03",X"21",X"4E",X"60",X"AF",X"06",X"0B",X"77",X"23",X"10",
		X"FC",X"DD",X"21",X"1C",X"60",X"DD",X"7E",X"00",X"E6",X"03",X"C2",X"0C",X"20",X"04",X"3E",X"0A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
