library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity draw_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of draw_sp_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"0C",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"40",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"40",X"40",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"04",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",
		X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"44",X"44",X"44",X"00",
		X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"04",X"44",X"40",X"00",X"04",X"44",X"00",X"00",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"40",
		X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"40",X"44",X"44",
		X"04",X"00",X"44",X"44",X"04",X"00",X"44",X"44",X"04",X"00",X"44",X"44",X"04",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",
		X"44",X"00",X"04",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"04",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"40",X"44",X"44",X"44",X"40",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"04",X"44",X"44",X"40",X"04",X"44",X"44",X"40",X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",
		X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"40",X"44",X"00",
		X"04",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",
		X"44",X"00",X"04",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"04",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"04",X"44",X"00",X"44",
		X"04",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"00",
		X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",
		X"44",X"40",X"44",X"00",X"44",X"40",X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",
		X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",
		X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"00",X"44",X"04",X"44",X"04",X"44",X"04",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"40",X"00",X"00",X"44",X"40",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",
		X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",
		X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"40",
		X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"00",X"44",X"44",X"44",X"04",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",
		X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",
		X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"40",X"44",
		X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",
		X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",
		X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",
		X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",
		X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",X"44",X"04",X"40",X"44",
		X"44",X"04",X"40",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"40",
		X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"C0",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"0C",X"C0",X"CC",
		X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",
		X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",
		X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",
		X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",
		X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"C0",X"CC",
		X"CC",X"0C",X"C0",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"C0",
		X"CC",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"40",X"44",X"44",X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"40",X"44",X"44",
		X"44",X"40",X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",
		X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",
		X"44",X"40",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"40",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"40",X"04",X"44",X"04",X"44",X"00",X"44",
		X"04",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"04",X"00",X"44",X"44",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"C0",
		X"0C",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"C0",X"00",X"CC",
		X"CC",X"C0",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"C0",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"C0",X"CC",X"CC",X"CC",X"C0",X"0C",X"CC",X"0C",X"CC",X"00",X"CC",
		X"0C",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"0C",X"00",X"CC",X"CC",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"04",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"40",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"04",X"44",X"00",X"44",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",
		X"44",X"40",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"40",X"44",X"00",X"44",X"40",X"44",X"00",X"44",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"0C",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"C0",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"0C",X"CC",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"C0",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"C0",X"CC",X"00",X"CC",X"C0",X"CC",X"00",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"0C",X"CC",X"CC",X"00",X"0C",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"04",X"40",
		X"00",X"44",X"04",X"44",X"00",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",
		X"04",X"44",X"44",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"0C",X"C0",
		X"00",X"CC",X"0C",X"CC",X"00",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",
		X"0C",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",
		X"CC",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"60",X"00",X"CC",X"CC",X"C6",
		X"06",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"06",X"CC",
		X"CC",X"CC",X"06",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",
		X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",
		X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"06",X"CC",
		X"CC",X"CC",X"06",X"CC",X"CC",X"CC",X"6C",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",
		X"06",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"66",X"66",X"CC",X"00",X"00",X"06",X"CC",X"00",X"00",X"06",X"CC",
		X"00",X"00",X"06",X"CC",X"66",X"00",X"06",X"CC",X"CC",X"00",X"6C",X"CC",X"CC",X"00",X"6C",X"CC",
		X"CC",X"66",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C6",
		X"6C",X"CC",X"CC",X"60",X"06",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"60",X"00",X"CC",X"CC",X"C6",X"06",X"CC",X"CC",X"CC",
		X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",
		X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"06",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C6",
		X"00",X"CC",X"CC",X"66",X"06",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",
		X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"6C",X"CC",X"CC",X"CC",X"06",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C6",X"00",X"CC",X"CC",X"60",
		X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"C0",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"CC",
		X"CC",X"C0",X"CC",X"CC",X"CC",X"C0",X"CC",X"CC",X"CC",X"C0",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"0C",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C0",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"04",X"00",X"00",X"CC",X"04",X"00",X"40",
		X"C0",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"04",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"04",X"44",X"44",X"04",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"40",X"04",X"00",X"40",
		X"40",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"04",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"04",X"00",X"00",X"0C",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"04",X"04",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"04",X"04",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"04",X"44",X"44",X"04",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"40",X"04",X"00",X"40",
		X"40",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"04",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"04",X"44",X"44",X"04",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"40",X"04",X"00",X"40",
		X"40",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"04",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"04",X"00",X"44",X"40",X"44",
		X"04",X"44",X"44",X"44",X"00",X"44",X"40",X"4C",X"00",X"04",X"00",X"CC",X"40",X"04",X"00",X"CC",
		X"40",X"00",X"00",X"CC",X"44",X"00",X"04",X"CC",X"44",X"40",X"44",X"CC",X"44",X"00",X"44",X"CC",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"04",X"04",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"00",
		X"44",X"44",X"40",X"00",X"4C",X"CC",X"40",X"04",X"CC",X"CC",X"44",X"04",X"CC",X"CC",X"44",X"44",
		X"CC",X"CC",X"44",X"44",X"CC",X"4C",X"44",X"44",X"C4",X"44",X"C4",X"04",X"44",X"44",X"C4",X"04",
		X"44",X"44",X"CC",X"00",X"44",X"44",X"CC",X"00",X"44",X"44",X"CC",X"40",X"4C",X"44",X"CC",X"00",
		X"40",X"00",X"44",X"C4",X"40",X"04",X"4C",X"44",X"00",X"04",X"4C",X"44",X"00",X"44",X"CC",X"44",
		X"04",X"44",X"CC",X"44",X"00",X"44",X"CC",X"44",X"00",X"04",X"CC",X"44",X"40",X"04",X"CC",X"44",
		X"40",X"00",X"CC",X"44",X"44",X"04",X"CC",X"44",X"44",X"44",X"CC",X"44",X"44",X"44",X"CC",X"44",
		X"40",X"44",X"CC",X"44",X"40",X"44",X"C4",X"44",X"00",X"44",X"C4",X"44",X"04",X"44",X"44",X"44",
		X"00",X"4C",X"44",X"4C",X"00",X"4C",X"44",X"4C",X"40",X"4C",X"44",X"4C",X"40",X"4C",X"44",X"4C",
		X"44",X"CC",X"44",X"CC",X"44",X"CC",X"44",X"CC",X"44",X"CC",X"44",X"CC",X"40",X"CC",X"40",X"CC",
		X"40",X"CC",X"40",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"04",X"CC",X"00",X"CC",
		X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"40",X"CC",X"00",X"CC",X"40",X"CC",X"04",X"CC",
		X"CC",X"04",X"CC",X"00",X"CC",X"44",X"CC",X"04",X"CC",X"44",X"CC",X"04",X"CC",X"44",X"CC",X"44",
		X"CC",X"44",X"C4",X"44",X"CC",X"44",X"C4",X"44",X"CC",X"4C",X"44",X"04",X"C4",X"CC",X"44",X"04",
		X"C4",X"CC",X"44",X"00",X"44",X"CC",X"44",X"00",X"44",X"CC",X"44",X"40",X"44",X"CC",X"44",X"00",
		X"44",X"C4",X"40",X"00",X"44",X"44",X"00",X"04",X"4C",X"44",X"00",X"04",X"CC",X"44",X"00",X"44",
		X"CC",X"44",X"04",X"44",X"4C",X"44",X"00",X"44",X"44",X"44",X"00",X"04",X"44",X"44",X"40",X"04",
		X"44",X"44",X"40",X"00",X"04",X"44",X"44",X"00",X"00",X"C4",X"44",X"40",X"00",X"C4",X"44",X"00",
		X"00",X"C4",X"40",X"00",X"04",X"C4",X"40",X"04",X"44",X"C4",X"00",X"04",X"44",X"C4",X"00",X"44",
		X"44",X"C4",X"04",X"44",X"44",X"C4",X"00",X"44",X"C4",X"44",X"00",X"04",X"C4",X"44",X"40",X"04",
		X"40",X"CC",X"00",X"CC",X"44",X"CC",X"04",X"CC",X"44",X"CC",X"44",X"CC",X"44",X"CC",X"44",X"C4",
		X"40",X"4C",X"44",X"C4",X"40",X"4C",X"44",X"44",X"00",X"44",X"4C",X"44",X"00",X"44",X"CC",X"44",
		X"04",X"44",X"CC",X"44",X"00",X"44",X"CC",X"44",X"00",X"44",X"CC",X"44",X"40",X"44",X"44",X"40",
		X"40",X"04",X"44",X"40",X"44",X"04",X"44",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"44",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"04",X"44",X"44",X"04",X"00",X"44",X"40",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"40",
		X"40",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"04",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"4C",X"44",X"40",X"00",X"CC",X"44",X"44",X"00",X"CC",X"44",X"44",X"40",X"CC",X"44",X"44",X"00",
		X"44",X"40",X"40",X"00",X"44",X"00",X"40",X"04",X"44",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"04",X"04",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"04",X"04",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"04",X"44",X"44",X"04",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"40",X"04",X"00",X"40",
		X"40",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"00",X"04",X"44",
		X"40",X"00",X"00",X"40",X"40",X"04",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"04",X"44",X"44",X"04",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"40",X"04",X"00",X"40",
		X"40",X"00",X"00",X"40",X"44",X"00",X"04",X"44",X"44",X"40",X"44",X"44",X"C4",X"00",X"04",X"44",
		X"CC",X"00",X"00",X"40",X"CC",X"04",X"00",X"40",X"CC",X"CC",X"CC",X"CC",X"0C",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"04",X"04",X"00",X"00",X"04",X"44",X"40",X"00",X"44",
		X"44",X"44",X"04",X"44",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"04",X"04",X"00",X"40",X"04",
		X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"00",X"40",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"66",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"C6",X"66",X"00",X"CC",X"C6",
		X"00",X"00",X"CC",X"60",X"00",X"00",X"CC",X"60",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"06",X"CC",X"00",X"00",X"06",X"CC",X"00",X"00",X"6C",X"CC",X"00",
		X"00",X"6C",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"CC",X"00",X"00",X"CC",X"CC",X"60",X"00",X"CC",X"CC",X"C6",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"06",X"CC",X"66",X"CC",
		X"06",X"CC",X"00",X"CC",X"6C",X"CC",X"00",X"CC",X"6C",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"66",
		X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C6",X"66",X"00",
		X"CC",X"C6",X"CC",X"60",X"CC",X"C6",X"CC",X"C6",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"6C",X"CC",
		X"CC",X"CC",X"06",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C6",X"00",X"CC",
		X"CC",X"C6",X"00",X"CC",X"CC",X"C6",X"00",X"CC",X"CC",X"C6",X"00",X"CC",X"CC",X"C6",X"00",X"CC",
		X"CC",X"C6",X"00",X"CC",X"CC",X"C6",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",
		X"CC",X"CC",X"06",X"CC",X"6C",X"CC",X"6C",X"CC",X"6C",X"CC",X"CC",X"CC",X"06",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"C6",X"00",X"CC",X"CC",X"60",
		X"00",X"66",X"CC",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",
		X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",
		X"6C",X"CC",X"CC",X"C6",X"6C",X"CC",X"CC",X"C6",X"6C",X"C6",X"66",X"66",X"6C",X"C6",X"00",X"00",
		X"6C",X"C6",X"00",X"00",X"6C",X"C6",X"00",X"00",X"6C",X"C6",X"66",X"00",X"6C",X"C6",X"CC",X"60",
		X"6C",X"C6",X"CC",X"66",X"6C",X"CC",X"CC",X"C6",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",
		X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",
		X"06",X"66",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"6C",X"CC",X"00",X"00",X"6C",X"CC",X"00",X"00",X"6C",X"CC",X"66",X"00",X"6C",X"CC",
		X"CC",X"00",X"6C",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"66",X"CC",X"CC",
		X"CC",X"C6",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"C6",X"CC",X"CC",X"CC",X"66",X"CC",X"CC",X"CC",X"60",X"6C",X"CC",X"CC",X"00",
		X"66",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"06",X"CC",X"CC",X"00",X"06",X"CC",X"CC",
		X"00",X"6C",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",
		X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"06",X"CC",X"CC",X"CC",
		X"06",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",X"CC",X"6C",X"C6",X"CC",X"CC",X"CC",X"C6",X"CC",X"CC",
		X"CC",X"60",X"CC",X"CC",X"CC",X"60",X"CC",X"CC",X"CC",X"66",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"66",X"66",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
