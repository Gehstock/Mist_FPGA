library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MoonWar_speech_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MoonWar_speech_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"04",X"A0",X"05",X"40",X"05",X"C0",X"06",X"00",X"06",X"C0",X"07",X"20",X"07",X"A0",X"08",X"40",
		X"08",X"E0",X"09",X"C0",X"0A",X"40",X"0A",X"C0",X"0C",X"00",X"0C",X"E0",X"0D",X"80",X"0E",X"20",
		X"0E",X"60",X"0F",X"00",X"0F",X"E0",X"11",X"20",X"11",X"60",X"12",X"80",X"13",X"80",X"13",X"C0",
		X"14",X"40",X"15",X"A0",X"16",X"20",X"16",X"60",X"16",X"E0",X"17",X"60",X"17",X"C0",X"18",X"20",
		X"18",X"C0",X"19",X"E0",X"1A",X"00",X"1A",X"20",X"1A",X"40",X"1B",X"1F",X"1D",X"41",X"21",X"59",
		X"22",X"1C",X"22",X"9C",X"2A",X"41",X"2E",X"51",X"22",X"1D",X"22",X"9D",X"30",X"41",X"34",X"D1",
		X"36",X"41",X"3A",X"59",X"3A",X"78",X"3B",X"1F",X"3D",X"1D",X"3D",X"9D",X"45",X"49",X"45",X"6E",
		X"3B",X"9F",X"48",X"1C",X"48",X"1C",X"50",X"41",X"54",X"D9",X"55",X"41",X"59",X"51",X"5B",X"52",
		X"22",X"1D",X"22",X"9D",X"1B",X"1F",X"5D",X"41",X"5D",X"78",X"22",X"1C",X"22",X"9C",X"1B",X"1F",
		X"1B",X"1F",X"1B",X"7F",X"61",X"41",X"22",X"1D",X"22",X"1D",X"65",X"D0",X"1B",X"1F",X"67",X"40",
		X"22",X"1C",X"22",X"9C",X"1B",X"1F",X"1B",X"7F",X"6B",X"41",X"6F",X"D1",X"3B",X"1F",X"71",X"52",
		X"48",X"1C",X"48",X"1C",X"73",X"49",X"73",X"7C",X"79",X"1F",X"79",X"67",X"3B",X"1F",X"76",X"C9",
		X"3D",X"1C",X"3D",X"1C",X"7B",X"41",X"7F",X"51",X"7F",X"6F",X"22",X"1C",X"22",X"9C",X"1B",X"1F",
		X"1B",X"7E",X"81",X"40",X"22",X"1D",X"22",X"9D",X"22",X"1C",X"22",X"1C",X"85",X"41",X"89",X"51",
		X"48",X"9D",X"8F",X"1C",X"97",X"C1",X"8B",X"51",X"8D",X"50",X"8F",X"1C",X"8F",X"1D",X"8F",X"9C",
		X"79",X"1F",X"79",X"1F",X"79",X"7E",X"9B",X"41",X"9F",X"58",X"22",X"1D",X"22",X"9D",X"3B",X"1F",
		X"A0",X"52",X"A0",X"79",X"3B",X"1F",X"A2",X"51",X"A2",X"78",X"3B",X"1F",X"A4",X"51",X"A4",X"78",
		X"3B",X"9F",X"A6",X"49",X"5B",X"D2",X"1B",X"1F",X"A9",X"1E",X"AF",X"51",X"AF",X"78",X"79",X"1F",
		X"79",X"7F",X"B1",X"58",X"B1",X"78",X"3B",X"9F",X"79",X"1F",X"79",X"1F",X"79",X"7F",X"B2",X"4D",
		X"B2",X"66",X"3B",X"1F",X"B5",X"49",X"5B",X"D6",X"B8",X"41",X"BC",X"D1",X"BE",X"49",X"BE",X"7D",
		X"3B",X"1F",X"C1",X"D1",X"A9",X"1D",X"A9",X"1D",X"C3",X"4D",X"C3",X"78",X"1B",X"1F",X"C6",X"51",
		X"48",X"1C",X"48",X"1C",X"C8",X"41",X"C8",X"78",X"CC",X"9F",X"CE",X"41",X"D2",X"59",X"22",X"1D",
		X"22",X"9D",X"D3",X"41",X"D7",X"C9",X"DA",X"52",X"DC",X"59",X"DC",X"6E",X"3B",X"9F",X"3B",X"1F",
		X"3B",X"1F",X"3B",X"7E",X"DD",X"C1",X"48",X"1C",X"48",X"1C",X"E1",X"C1",X"E5",X"49",X"E5",X"67",
		X"3B",X"9F",X"3B",X"1F",X"3B",X"1F",X"3B",X"7E",X"E8",X"50",X"5B",X"D1",X"EA",X"51",X"EA",X"67",
		X"79",X"1F",X"79",X"1F",X"79",X"7F",X"EC",X"41",X"EC",X"75",X"79",X"1F",X"A9",X"9F",X"A9",X"FC",
		X"A9",X"F8",X"A9",X"F0",X"A9",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"99",X"72",X"63",X"69",X"99",X"99",X"99",X"97",X"72",X"5A",X"66",X"59",X"99",X"98",X"A6",X"65",
		X"E2",X"97",X"66",X"5D",X"99",X"69",X"99",X"99",X"8A",X"66",X"59",X"99",X"9D",X"75",X"99",X"98",
		X"76",X"68",X"96",X"66",X"65",X"99",X"9E",X"AA",X"69",X"9A",X"27",X"59",X"C5",X"95",X"AA",X"AD",
		X"29",X"9E",X"1A",X"67",X"61",X"64",X"7F",X"6F",X"2A",X"2A",X"1A",X"57",X"C5",X"94",X"7F",X"3F",
		X"29",X"A9",X"5E",X"1E",X"95",X"64",X"3F",X"6F",X"26",X"7A",X"1E",X"1A",X"D5",X"54",X"6F",X"6F",
		X"65",X"AA",X"1E",X"1A",X"D5",X"60",X"2F",X"AF",X"58",X"AD",X"5E",X"1A",X"D4",X"A0",X"3F",X"6F",
		X"95",X"7A",X"2A",X"57",X"95",X"E0",X"6A",X"AF",X"98",X"69",X"9E",X"62",X"59",X"D5",X"69",X"EE",
		X"97",X"5A",X"5D",X"75",X"D8",X"D7",X"5C",X"A3",X"35",X"CA",X"33",X"28",X"CA",X"35",X"CA",X"33",
		X"5A",X"28",X"9C",X"A5",X"D6",X"97",X"32",X"8D",X"72",X"8A",X"35",X"D6",X"96",X"8A",X"28",X"A5",
		X"72",X"97",X"5C",X"A3",X"32",X"8C",X"A5",X"A2",X"8C",X"A3",X"28",X"A2",X"8D",X"73",X"35",X"CA",
		X"5A",X"29",X"75",X"A2",X"97",X"28",X"CD",X"73",X"28",X"A3",X"33",X"5D",X"75",X"A5",X"D7",X"5C",
		X"69",X"68",X"CC",X"A3",X"35",X"D6",X"96",X"8A",X"35",X"CA",X"27",X"28",X"D6",X"97",X"5C",X"CA",
		X"29",X"75",X"D7",X"33",X"5C",X"CA",X"28",X"CA",X"33",X"28",X"D7",X"5C",X"A5",X"D7",X"5D",X"73",
		X"8D",X"75",X"CA",X"32",X"8A",X"5D",X"75",X"D6",X"97",X"5A",X"29",X"73",X"28",X"A2",X"8A",X"5A",
		X"28",X"D7",X"33",X"5A",X"5D",X"75",X"D6",X"8A",X"5D",X"68",X"A2",X"8A",X"5D",X"73",X"35",X"D7",
		X"29",X"8A",X"95",X"A9",X"67",X"98",X"7D",X"1F",X"69",X"5A",X"86",X"79",X"5E",X"65",X"AD",X"1F",
		X"78",X"2E",X"47",X"9A",X"1A",X"D1",X"B8",X"2F",X"B0",X"7D",X"0B",X"D0",X"BD",X"1A",X"A5",X"6A",
		X"8B",X"42",X"F0",X"2F",X"47",X"C2",X"F4",X"3F",X"8E",X"47",X"D4",X"3F",X"43",X"F4",X"B5",X"3F",
		X"9A",X"81",X"E0",X"BD",X"0A",X"F1",X"B5",X"2F",X"99",X"86",X"76",X"1A",X"1F",X"96",X"39",X"6F",
		X"8A",X"59",X"98",X"5E",X"67",X"99",X"6A",X"6B",X"89",X"A5",X"89",X"5A",X"A6",X"A1",X"A9",X"9E",
		X"98",X"69",X"5D",X"99",X"9A",X"79",X"6A",X"2A",X"89",X"D5",X"D5",X"E2",X"71",X"F8",X"69",X"7A",
		X"66",X"29",X"8A",X"65",X"9E",X"66",X"6D",X"1F",X"75",X"6A",X"1A",X"87",X"86",X"D4",X"F8",X"2E",
		X"67",X"61",X"A6",X"65",X"9E",X"82",X"F4",X"3F",X"A6",X"19",X"59",X"E9",X"0F",X"D6",X"75",X"6F",
		X"67",X"67",X"55",X"67",X"67",X"95",X"E9",X"6E",X"A2",X"62",X"65",X"9D",X"96",X"95",X"EA",X"7A",
		X"99",X"98",X"99",X"6A",X"26",X"56",X"AA",X"7A",X"A9",X"96",X"21",X"6A",X"27",X"61",X"AA",X"AA",
		X"A1",X"AA",X"95",X"45",X"AE",X"81",X"E6",X"BE",X"7A",X"15",X"AF",X"40",X"7A",X"A6",X"15",X"FF",
		X"A8",X"59",X"D9",X"D9",X"42",X"FD",X"41",X"FF",X"99",X"99",X"99",X"A6",X"05",X"FE",X"41",X"BE",
		X"66",X"66",X"62",X"66",X"66",X"76",X"9E",X"69",X"99",X"66",X"66",X"26",X"67",X"59",X"E9",X"AA",
		X"A5",X"99",X"66",X"66",X"59",X"99",X"AA",X"9D",X"6A",X"61",X"A6",X"3A",X"16",X"55",X"EA",X"7A",
		X"23",X"A6",X"71",X"7A",X"98",X"90",X"7E",X"7F",X"91",X"F5",X"7D",X"1F",X"56",X"90",X"7E",X"7F",
		X"C1",X"E5",X"BC",X"0B",X"97",X"90",X"7A",X"7F",X"D1",X"A1",X"BD",X"0F",X"87",X"90",X"6D",X"AF",
		X"99",X"85",X"AE",X"1A",X"47",X"E0",X"68",X"BF",X"86",X"A5",X"A8",X"7A",X"09",X"E2",X"65",X"7F",
		X"8A",X"63",X"66",X"87",X"63",X"5A",X"59",X"CA",X"5A",X"5A",X"29",X"69",X"8A",X"29",X"5E",X"29",
		X"68",X"A5",X"A5",X"A6",X"66",X"66",X"66",X"66",X"62",X"66",X"63",X"67",X"26",X"69",X"96",X"89",
		X"96",X"99",X"73",X"5A",X"63",X"5C",X"CC",X"CA",X"62",X"96",X"73",X"32",X"8C",X"D6",X"98",X"A6",
		X"29",X"8A",X"32",X"8C",X"A5",X"A5",X"CA",X"5C",X"A3",X"35",X"A2",X"8C",X"D6",X"76",X"27",X"5C",
		X"89",X"D6",X"75",X"A5",X"CC",X"A3",X"27",X"32",X"98",X"A6",X"28",X"CA",X"5A",X"35",X"9C",X"CD",
		X"73",X"35",X"A6",X"29",X"8A",X"65",X"CD",X"73",X"26",X"96",X"98",X"9D",X"89",X"D8",X"A3",X"27",
		X"8A",X"35",X"A5",X"A5",X"9C",X"D7",X"35",X"CD",X"69",X"67",X"62",X"97",X"32",X"97",X"5C",X"CA",
		X"33",X"5D",X"72",X"8C",X"9D",X"73",X"5A",X"35",X"A5",X"CC",X"D7",X"33",X"35",X"D6",X"8D",X"69",
		X"96",X"69",X"73",X"5C",X"D8",X"A5",X"CC",X"CC",X"A3",X"5A",X"33",X"32",X"8C",X"D8",X"9C",X"CD",
		X"73",X"59",X"D7",X"32",X"8C",X"CC",X"A5",X"9C",X"CA",X"33",X"33",X"28",X"CA",X"5C",X"D7",X"35",
		X"99",X"95",X"A9",X"AC",X"0B",X"C0",X"A5",X"FF",X"99",X"85",X"B9",X"6D",X"0B",X"C0",X"79",X"BF",
		X"96",X"59",X"F1",X"7D",X"0B",X"C0",X"79",X"BF",X"19",X"EA",X"95",X"99",X"8A",X"90",X"AD",X"AF",
		X"3A",X"89",X"95",X"79",X"66",X"15",X"BA",X"7F",X"9E",X"65",X"85",X"6A",X"66",X"55",X"AE",X"7B",
		X"98",X"A6",X"26",X"97",X"35",X"CD",X"89",X"D8",X"A2",X"8D",X"73",X"28",X"D7",X"35",X"A6",X"28",
		X"9C",X"D7",X"29",X"73",X"29",X"73",X"28",X"CD",X"8C",X"9D",X"68",X"A3",X"32",X"98",X"A3",X"5C",
		X"73",X"59",X"9D",X"8A",X"86",X"69",X"66",X"98",X"9D",X"8A",X"35",X"D7",X"63",X"28",X"CA",X"65",
		X"A3",X"62",X"75",X"A3",X"29",X"68",X"A5",X"D7",X"35",X"CA",X"32",X"8A",X"29",X"8A",X"65",X"CA",
		X"69",X"8C",X"9A",X"5C",X"A3",X"63",X"5A",X"5D",X"73",X"5C",X"D7",X"32",X"8A",X"35",X"9A",X"29",
		X"8A",X"35",X"C9",X"A3",X"32",X"8A",X"36",X"28",X"D7",X"32",X"8C",X"A3",X"5C",X"D7",X"35",X"D7",
		X"96",X"75",X"D6",X"8A",X"29",X"66",X"97",X"5C",X"D6",X"69",X"97",X"28",X"CC",X"A5",X"9D",X"67",
		X"5A",X"36",X"62",X"76",X"5A",X"27",X"5A",X"28",X"A5",X"D6",X"76",X"27",X"29",X"72",X"8C",X"D7",
		X"59",X"E6",X"76",X"19",X"D8",X"84",X"AE",X"EE",X"95",X"9A",X"A9",X"57",X"86",X"D0",X"3D",X"FF",
		X"A1",X"61",X"FD",X"4E",X"56",X"D0",X"79",X"FF",X"1F",X"81",X"E5",X"FD",X"02",X"E4",X"7C",X"7F",
		X"86",X"3B",X"80",X"FE",X"02",X"A4",X"BC",X"2F",X"79",X"4F",X"92",X"71",X"E8",X"1B",X"E0",X"3F",
		X"A5",X"6A",X"85",X"D5",X"F4",X"1F",X"D4",X"7F",X"67",X"A1",X"79",X"5A",X"84",X"7F",X"80",X"BF",
		X"39",X"D5",X"9D",X"6A",X"11",X"EF",X"50",X"BF",X"A6",X"26",X"65",X"D8",X"56",X"BA",X"05",X"FF",
		X"66",X"26",X"9A",X"26",X"5A",X"A1",X"B8",X"2B",X"75",X"67",X"66",X"66",X"57",X"E0",X"F8",X"2B",
		X"26",X"7A",X"55",X"9A",X"A6",X"51",X"7A",X"BE",X"95",X"5F",X"98",X"86",X"AA",X"54",X"69",X"FF",
		X"A0",X"6B",X"99",X"56",X"AA",X"54",X"69",X"FF",X"D4",X"6A",X"77",X"55",X"7B",X"60",X"5A",X"BF",
		X"A5",X"68",X"6B",X"95",X"1B",X"D0",X"66",X"BF",X"C4",X"B9",X"19",X"FD",X"03",X"E5",X"E4",X"7F",
		X"3D",X"46",X"BC",X"0B",X"C1",X"E1",X"B5",X"2F",X"D1",X"F4",X"2F",X"43",X"E1",X"A1",X"B5",X"2F",
		X"D0",X"F8",X"2F",X"43",X"D5",X"D5",X"F4",X"2F",X"76",X"26",X"98",X"6A",X"59",X"97",X"B4",X"3F",
		X"66",X"65",X"A6",X"68",X"99",X"A8",X"79",X"5F",X"66",X"65",X"A6",X"68",X"76",X"76",X"39",X"5F",
		X"66",X"65",X"A6",X"66",X"66",X"78",X"79",X"6A",X"66",X"65",X"A6",X"66",X"66",X"76",X"39",X"6A",
		X"A6",X"66",X"19",X"97",X"65",X"96",X"7A",X"AA",X"A9",X"66",X"1A",X"66",X"55",X"65",X"AF",X"6E",
		X"A9",X"69",X"5A",X"86",X"60",X"68",X"AF",X"6B",X"A9",X"69",X"5A",X"86",X"60",X"69",X"7F",X"6B",
		X"A9",X"69",X"8A",X"56",X"60",X"69",X"7F",X"6B",X"A9",X"67",X"59",X"C6",X"55",X"5D",X"7F",X"6B",
		X"9D",X"89",X"8A",X"62",X"55",X"99",X"EE",X"AA",X"A6",X"19",X"99",X"D8",X"98",X"67",X"7A",X"9A",
		X"99",X"99",X"89",X"89",X"A6",X"65",X"AA",X"7A",X"26",X"AA",X"61",X"86",X"A5",X"98",X"6A",X"AA",
		X"95",X"9D",X"A9",X"86",X"66",X"71",X"6A",X"6F",X"C5",X"94",X"BF",X"1D",X"42",X"F4",X"2A",X"7F",
		X"8A",X"90",X"BF",X"17",X"42",X"F4",X"2D",X"6F",X"83",X"E0",X"7F",X"5A",X"02",X"F4",X"3D",X"3F",
		X"61",X"B8",X"2F",X"57",X"42",X"F4",X"3D",X"3F",X"66",X"A9",X"1F",X"56",X"53",X"B4",X"79",X"7F",
		X"66",X"62",X"98",X"9D",X"6A",X"95",X"E9",X"2F",X"35",X"9D",X"66",X"67",X"67",X"95",X"A8",X"6F",
		X"95",X"9A",X"A6",X"19",X"6A",X"85",X"9A",X"AA",X"A1",X"5E",X"9E",X"55",X"99",X"A5",X"5E",X"2F",
		X"96",X"76",X"62",X"19",X"E7",X"65",X"67",X"AE",X"19",X"FD",X"59",X"0B",X"96",X"94",X"6E",X"7F",
		X"39",X"E9",X"58",X"5A",X"95",X"A0",X"7F",X"3F",X"7A",X"65",X"59",X"9A",X"95",X"61",X"7E",X"7B",
		X"66",X"36",X"66",X"59",X"D9",X"E5",X"78",X"7F",X"67",X"1A",X"89",X"D5",X"9A",X"A5",X"68",X"7F",
		X"39",X"6A",X"59",X"D5",X"95",X"F8",X"1E",X"3B",X"67",X"66",X"57",X"A1",X"95",X"B8",X"68",X"7F",
		X"89",X"99",X"9D",X"99",X"99",X"95",X"67",X"AF",X"95",X"99",X"F5",X"66",X"2A",X"90",X"6A",X"BF",
		X"95",X"D5",X"F9",X"59",X"5F",X"80",X"79",X"FF",X"86",X"63",X"E5",X"68",X"5B",X"90",X"79",X"FF",
		X"26",X"6A",X"98",X"D8",X"9A",X"50",X"B9",X"BF",X"76",X"75",X"99",X"76",X"26",X"16",X"AA",X"AE",
		X"99",X"89",X"99",X"D9",X"62",X"66",X"7A",X"77",X"99",X"98",X"99",X"D6",X"65",X"99",X"A9",X"E9",
		X"77",X"66",X"62",X"26",X"66",X"26",X"67",X"AA",X"98",X"9E",X"98",X"58",X"8D",X"A9",X"57",X"AE",
		X"99",X"99",X"D9",X"65",X"62",X"A9",X"86",X"AA",X"99",X"D8",X"89",X"D8",X"57",X"B6",X"15",X"BE",
		X"98",X"79",X"5A",X"96",X"66",X"A0",X"F8",X"2F",X"76",X"27",X"57",X"96",X"66",X"A0",X"F8",X"2F",
		X"A5",X"6A",X"1A",X"66",X"57",X"D0",X"F8",X"3B",X"95",X"E5",X"69",X"99",X"8E",X"85",X"F5",X"2F",
		X"99",X"A6",X"18",X"67",X"99",X"D6",X"39",X"E9",X"66",X"A6",X"25",X"5A",X"A5",X"D5",X"7A",X"7B",
		X"A0",X"6E",X"3E",X"03",X"83",X"F4",X"2E",X"3F",X"78",X"75",X"3F",X"57",X"42",X"F4",X"2D",X"7F",
		X"86",X"B4",X"3F",X"0F",X"02",X"F0",X"78",X"7F",X"5A",X"9A",X"A0",X"3F",X"03",X"D2",X"F0",X"3F",
		X"66",X"76",X"56",X"7A",X"16",X"A2",X"A5",X"3F",X"8A",X"75",X"59",X"E5",X"96",X"7A",X"64",X"7F",
		X"2B",X"55",X"9A",X"61",X"A5",X"7F",X"01",X"BF",X"3E",X"45",X"E7",X"61",X"85",X"EE",X"11",X"BF",
		X"79",X"86",X"9C",X"99",X"59",X"AA",X"51",X"FE",X"A6",X"26",X"66",X"66",X"16",X"AA",X"15",X"EE",
		X"8D",X"72",X"66",X"76",X"27",X"5D",X"97",X"5C",X"9D",X"75",X"99",X"E2",X"62",X"73",X"65",X"A2",
		X"8A",X"27",X"29",X"89",X"9A",X"5D",X"66",X"6A",X"25",X"9D",X"99",X"62",X"79",X"99",X"66",X"99",
		X"98",X"9D",X"87",X"86",X"A2",X"95",X"B8",X"2F",X"D1",X"F4",X"A8",X"79",X"1F",X"52",X"F0",X"3F",
		X"78",X"6A",X"17",X"99",X"87",X"D0",X"F5",X"2F",X"A1",X"E1",X"B4",X"7D",X"1B",X"82",X"B4",X"2F",
		X"78",X"2E",X"0E",X"8A",X"57",X"D0",X"FC",X"1F",X"C2",X"B4",X"2F",X"42",X"F0",X"B4",X"B8",X"2F",
		X"2A",X"A9",X"46",X"A9",X"46",X"E1",X"B5",X"3F",X"98",X"A8",X"A9",X"55",X"D6",X"A4",X"7D",X"6F",
		X"98",X"E6",X"26",X"1A",X"95",X"E4",X"7E",X"2B",X"A6",X"65",X"69",X"5E",X"56",X"62",X"AA",X"6A",
		X"A2",X"66",X"27",X"59",X"95",X"A6",X"7A",X"79",X"99",X"96",X"66",X"66",X"26",X"66",X"9E",X"9D",
		X"99",X"D6",X"61",X"69",X"9E",X"56",X"9A",X"A9",X"99",X"A2",X"29",X"89",X"86",X"B1",X"79",X"6F",
		X"96",X"A0",X"BC",X"0B",X"C1",X"F4",X"AC",X"2F",X"D4",X"AD",X"0B",X"C1",X"F4",X"A8",X"7D",X"1F",
		X"78",X"2F",X"07",X"D1",X"E5",X"A5",X"7C",X"1F",X"A5",X"3E",X"0B",X"57",X"57",X"D0",X"F8",X"2F",
		X"78",X"5E",X"1E",X"4A",X"C5",X"E5",X"B5",X"2F",X"89",X"99",X"89",X"9D",X"89",X"AA",X"65",X"AB",
		X"99",X"9D",X"56",X"99",X"85",X"F9",X"66",X"2F",X"95",X"ED",X"43",X"E5",X"90",X"FD",X"5D",X"6F",
		X"91",X"FA",X"94",X"3F",X"03",X"97",X"E0",X"7F",X"D0",X"FC",X"3D",X"0B",X"C0",X"E9",X"E1",X"3F",
		X"63",X"B0",X"3F",X"03",X"E0",X"7C",X"7D",X"2B",X"87",X"B4",X"2F",X"02",X"F0",X"A8",X"7D",X"2B",
		X"C4",X"BC",X"0F",X"52",X"E1",X"E1",X"B8",X"2F",X"A2",X"29",X"57",X"A1",X"9D",X"D5",X"B8",X"2F",
		X"A1",X"A6",X"1A",X"59",X"9A",X"95",X"F5",X"2F",X"96",X"72",X"36",X"1E",X"57",X"A2",X"A8",X"6E",
		X"66",X"62",X"76",X"66",X"23",X"A6",X"76",X"2E",X"66",X"66",X"27",X"63",X"5A",X"99",X"9C",X"7F",
		X"76",X"95",X"6B",X"52",X"66",X"79",X"C4",X"FF",X"6B",X"80",X"AF",X"50",X"6A",X"6A",X"81",X"FF",
		X"6B",X"80",X"EE",X"80",X"76",X"7A",X"55",X"BF",X"2B",X"C0",X"AE",X"50",X"9E",X"6A",X"55",X"BF",
		X"2F",X"80",X"7F",X"41",X"9A",X"A9",X"55",X"BF",X"3F",X"01",X"FA",X"12",X"1A",X"AE",X"41",X"BF",
		X"7E",X"05",X"E7",X"62",X"15",X"BE",X"01",X"FF",X"6A",X"95",X"5A",X"66",X"61",X"7F",X"50",X"BF",
		X"75",X"D7",X"5D",X"68",X"CC",X"CC",X"A2",X"8D",X"72",X"8C",X"CC",X"A3",X"29",X"72",X"8D",X"72",
		X"97",X"27",X"29",X"75",X"A2",X"8A",X"28",X"CD",X"75",X"A2",X"8D",X"72",X"8D",X"72",X"8C",X"A3",
		X"8A",X"33",X"28",X"D7",X"33",X"35",X"CC",X"D7",X"28",X"CC",X"CC",X"CC",X"CC",X"CA",X"35",X"9C",
		X"CA",X"5D",X"73",X"5C",X"CD",X"72",X"8D",X"73",X"5D",X"73",X"33",X"5D",X"73",X"28",X"A2",X"8A",
		X"8A",X"5C",X"CC",X"CC",X"CC",X"CD",X"73",X"32",X"8A",X"33",X"28",X"CC",X"CC",X"CC",X"CD",X"8C",
		X"CC",X"A3",X"35",X"CC",X"CA",X"27",X"5C",X"CA",X"5D",X"73",X"33",X"5C",X"A3",X"32",X"8C",X"A5",
		X"97",X"33",X"33",X"36",X"33",X"28",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"D8",X"CC",X"C9",
		X"D7",X"5C",X"CC",X"CC",X"D6",X"8C",X"CA",X"33",X"5C",X"A3",X"33",X"33",X"33",X"33",X"33",X"27",
		X"99",X"A2",X"76",X"16",X"57",X"A5",X"A9",X"AF",X"88",X"99",X"FD",X"46",X"07",X"E0",X"7E",X"6F",
		X"66",X"17",X"FC",X"18",X"47",X"E4",X"7D",X"7F",X"91",X"A7",X"BD",X"18",X"4E",X"D0",X"BC",X"6F",
		X"89",X"86",X"F9",X"1E",X"07",X"D0",X"A9",X"FF",X"85",X"D7",X"BC",X"28",X"0F",X"C0",X"B9",X"7F",
		X"86",X"57",X"F9",X"28",X"0F",X"D0",X"AC",X"7F",X"66",X"5A",X"AA",X"55",X"5A",X"94",X"5E",X"FE",
		X"66",X"A9",X"55",X"99",X"A9",X"55",X"AA",X"EE",X"2A",X"9D",X"56",X"95",X"A9",X"46",X"B6",X"BE",
		X"27",X"7A",X"55",X"96",X"7D",X"41",X"F7",X"BE",X"61",X"7F",X"1A",X"81",X"AD",X"45",X"A6",X"BF",
		X"66",X"39",X"6B",X"A0",X"1D",X"5B",X"C0",X"FF",X"A5",X"6A",X"86",X"65",X"9D",X"1B",X"D0",X"BF",
		X"66",X"A1",X"79",X"59",X"9D",X"4F",X"E0",X"7F",X"66",X"95",X"9D",X"86",X"A6",X"5A",X"B4",X"6F",
		X"66",X"62",X"68",X"6A",X"5A",X"A1",X"B8",X"2F",X"62",X"6A",X"55",X"DD",X"8A",X"67",X"A5",X"3F",
		X"A1",X"79",X"5A",X"5A",X"86",X"D4",X"F9",X"2B",X"69",X"5E",X"57",X"66",X"86",X"D4",X"BC",X"2B",
		X"69",X"5A",X"96",X"67",X"56",X"D4",X"BC",X"2B",X"69",X"5A",X"95",X"DA",X"56",X"D4",X"BC",X"2B",
		X"69",X"99",X"76",X"56",X"98",X"9A",X"A1",X"AF",X"D0",X"F8",X"7D",X"0B",X"C0",X"7A",X"E0",X"7F",
		X"C1",X"B5",X"B5",X"2F",X"40",X"B8",X"7D",X"2F",X"2B",X"12",X"F0",X"3F",X"05",X"DA",X"C4",X"BE",
		X"A5",X"96",X"66",X"1E",X"85",X"E9",X"A8",X"2F",X"E4",X"78",X"6C",X"0B",X"D0",X"BC",X"79",X"2F",
		X"D4",X"B8",X"3D",X"0B",X"C0",X"F8",X"A8",X"3F",X"B4",X"7D",X"0F",X"0A",X"C0",X"FC",X"79",X"2F",
		X"A1",X"6D",X"4A",X"D0",X"F8",X"78",X"AD",X"1F",X"75",X"7D",X"0B",X"C0",X"F8",X"79",X"7D",X"1F",
		X"66",X"A4",X"7E",X"03",X"F0",X"3D",X"B8",X"2F",X"38",X"5B",X"A8",X"0B",X"D0",X"7E",X"78",X"3F",
		X"35",X"7E",X"07",X"97",X"C0",X"BA",X"A0",X"BF",X"38",X"69",X"69",X"8A",X"57",X"E0",X"BC",X"2B",
		X"75",X"A3",X"28",X"C9",X"D7",X"59",X"D9",X"67",X"5D",X"69",X"75",X"D8",X"C7",X"97",X"5A",X"29",
		X"89",X"A5",X"A5",X"A6",X"26",X"97",X"5A",X"89",X"67",X"65",X"9D",X"96",X"69",X"89",X"A5",X"A2",
		X"67",X"5D",X"76",X"28",X"9E",X"22",X"98",X"CA",X"63",X"27",X"28",X"9A",X"65",X"A5",X"9A",X"66",
		X"63",X"28",X"9D",X"99",X"66",X"96",X"76",X"5A",X"27",X"59",X"D9",X"66",X"78",X"89",X"D6",X"75",
		X"96",X"98",X"9A",X"5D",X"8A",X"71",X"78",X"D8",X"CA",X"59",X"D9",X"69",X"98",X"99",X"D6",X"76",
		X"27",X"5D",X"8A",X"65",X"99",X"9D",X"6A",X"19",X"D8",X"D5",X"E6",X"5A",X"5D",X"69",X"75",X"99",
		X"96",X"66",X"76",X"59",X"D9",X"95",X"67",X"AE",X"C1",X"E1",X"BD",X"49",X"D7",X"94",X"3E",X"7F",
		X"D4",X"78",X"7F",X"07",X"92",X"B0",X"2E",X"6F",X"D4",X"75",X"AF",X"07",X"85",X"F0",X"2E",X"6F",
		X"6A",X"62",X"75",X"66",X"66",X"62",X"B4",X"3F",X"D0",X"FC",X"65",X"2F",X"02",X"E0",X"F8",X"3F",
		X"69",X"D5",X"9D",X"86",X"76",X"63",X"B4",X"3F",X"1F",X"47",X"F0",X"3F",X"03",X"97",X"D0",X"BF",
		X"82",X"F0",X"AC",X"3F",X"01",X"A7",X"A0",X"AF",X"57",X"D4",X"E5",X"BD",X"03",X"F0",X"68",X"BF",
		X"2B",X"42",X"F5",X"A8",X"0B",X"D4",X"5D",X"BF",X"2B",X"42",X"F5",X"A8",X"0B",X"D4",X"5D",X"BF",
		X"A5",X"6A",X"55",X"9A",X"85",X"B8",X"78",X"6F",X"96",X"79",X"59",X"9A",X"81",X"F5",X"E5",X"3F",
		X"89",X"E6",X"26",X"5A",X"81",X"F8",X"66",X"2F",X"67",X"A5",X"66",X"5E",X"12",X"B5",X"98",X"AE",
		X"5A",X"A5",X"5A",X"67",X"81",X"F8",X"78",X"6E",X"2A",X"1D",X"8A",X"96",X"63",X"A4",X"B8",X"2F",
		X"85",X"E6",X"A8",X"59",X"D9",X"D4",X"6D",X"7F",X"91",X"F4",X"BD",X"0F",X"56",X"D0",X"7D",X"AF",
		X"85",X"E5",X"F8",X"27",X"95",X"E0",X"3E",X"7F",X"56",X"A6",X"B5",X"27",X"95",X"E0",X"3E",X"7F",
		X"56",X"A6",X"B5",X"1E",X"89",X"A0",X"2F",X"3F",X"86",X"72",X"F0",X"79",X"2B",X"50",X"7D",X"EF",
		X"61",X"AA",X"D4",X"A8",X"3F",X"01",X"79",X"FF",X"D0",X"AE",X"75",X"65",X"3F",X"41",X"9D",X"FF",
		X"85",X"A9",X"AF",X"00",X"AF",X"06",X"85",X"FF",X"76",X"47",X"BE",X"40",X"AD",X"5E",X"55",X"BF",
		X"76",X"56",X"AA",X"55",X"96",X"79",X"55",X"FF",X"9C",X"89",X"A9",X"98",X"56",X"AA",X"15",X"EE",
		X"95",X"9A",X"61",X"67",X"A6",X"76",X"63",X"BA",X"79",X"85",X"9D",X"98",X"95",X"AE",X"91",X"BF",
		X"29",X"AA",X"80",X"F9",X"1A",X"1F",X"D0",X"BF",X"61",X"F8",X"A5",X"2F",X"00",X"F8",X"9C",X"AF",
		X"95",X"B8",X"78",X"2F",X"00",X"F9",X"78",X"7F",X"69",X"99",X"E9",X"0B",X"80",X"BD",X"69",X"3F",
		X"75",X"9C",X"5F",X"43",X"F0",X"A8",X"B5",X"2F",X"A1",X"6A",X"4A",X"D0",X"F8",X"69",X"B8",X"2F",
		X"69",X"5B",X"43",X"E0",X"E7",X"95",X"F8",X"2F",X"5E",X"53",X"D1",X"F4",X"7D",X"95",X"F8",X"2F",
		X"C5",X"62",X"BC",X"1D",X"5B",X"C0",X"5A",X"BF",X"D5",X"81",X"FD",X"78",X"0F",X"D0",X"A8",X"7F",
		X"2B",X"43",X"E0",X"FC",X"07",X"E5",X"58",X"EF",X"66",X"62",X"E4",X"7E",X"41",X"F8",X"78",X"2F",
		X"97",X"85",X"F8",X"0B",X"D0",X"F5",X"A8",X"2F",X"97",X"85",X"F8",X"0B",X"D0",X"F5",X"A8",X"2F",
		X"98",X"9A",X"A1",X"23",X"A9",X"99",X"66",X"AA",X"A6",X"19",X"D9",X"88",X"99",X"E9",X"55",X"EF",
		X"A6",X"56",X"69",X"98",X"88",X"EA",X"55",X"AF",X"79",X"85",X"A9",X"96",X"26",X"7A",X"55",X"AF",
		X"99",X"88",X"99",X"9A",X"66",X"66",X"3A",X"9E",X"99",X"89",X"66",X"66",X"99",X"99",X"9E",X"9E",
		X"A5",X"7A",X"1E",X"07",X"8A",X"A1",X"69",X"AA",X"3C",X"79",X"2B",X"47",X"42",X"F8",X"69",X"3F",
		X"35",X"BD",X"07",X"D6",X"90",X"BD",X"59",X"6F",X"92",X"BC",X"1D",X"8E",X"80",X"FC",X"2D",X"2F",
		X"91",X"FD",X"1A",X"8A",X"80",X"FC",X"2D",X"2F",X"69",X"A5",X"6A",X"57",X"52",X"F4",X"69",X"7F",
		X"97",X"5C",X"D9",X"67",X"83",X"9D",X"8D",X"78",X"67",X"59",X"9D",X"73",X"29",X"76",X"63",X"28",
		X"D8",X"99",X"A6",X"62",X"66",X"99",X"89",X"99",X"D6",X"66",X"99",X"72",X"8A",X"66",X"5A",X"66",
		X"66",X"63",X"A8",X"5E",X"81",X"E8",X"A5",X"6F",X"66",X"61",X"FC",X"0F",X"80",X"BC",X"78",X"3F",
		X"D0",X"F4",X"FD",X"0B",X"D0",X"3A",X"A5",X"6F",X"D0",X"BC",X"2E",X"0B",X"C0",X"6A",X"B0",X"7F",
		X"D0",X"BC",X"2E",X"0F",X"80",X"AA",X"A4",X"7F",X"C0",X"FC",X"65",X"7F",X"02",X"A0",X"F8",X"2F",
		X"82",X"F0",X"AC",X"3F",X"00",X"F9",X"A1",X"3F",X"82",X"F4",X"6E",X"1E",X"42",X"F0",X"78",X"AF",
		X"67",X"76",X"1A",X"66",X"16",X"A9",X"65",X"AF",X"87",X"98",X"65",X"E9",X"57",X"9E",X"85",X"EA",
		X"57",X"E0",X"7E",X"07",X"D4",X"F0",X"BC",X"1F",X"A1",X"A5",X"AD",X"0F",X"53",X"C2",X"F4",X"2F",
		X"D0",X"BC",X"68",X"2F",X"03",X"D4",X"F8",X"2F",X"D0",X"FC",X"2D",X"4B",X"50",X"FD",X"84",X"BF",
		X"66",X"98",X"67",X"69",X"57",X"E0",X"B8",X"2F",X"85",X"BE",X"03",X"E2",X"80",X"FD",X"19",X"7F",
		X"94",X"FD",X"4A",X"C5",X"D0",X"FD",X"0D",X"AF",X"89",X"98",X"E5",X"6A",X"1A",X"D1",X"B8",X"2F",
		X"67",X"56",X"A5",X"79",X"5A",X"D1",X"B8",X"2F",X"67",X"56",X"A1",X"A9",X"5A",X"D1",X"F5",X"2F",
		X"D1",X"F4",X"2F",X"42",X"F0",X"A8",X"B5",X"2F",X"A4",X"AD",X"0F",X"82",X"D6",X"A0",X"F5",X"2F",
		X"78",X"2F",X"43",X"E0",X"E5",X"E0",X"B8",X"2F",X"69",X"5E",X"56",X"99",X"97",X"A0",X"BC",X"2B",
		X"29",X"2F",X"0B",X"87",X"80",X"BE",X"03",X"F4",X"30",X"FD",X"1F",X"5B",X"00",X"BE",X"07",X"F0",
		X"84",X"FC",X"5E",X"2B",X"00",X"BF",X"03",X"F0",X"81",X"FC",X"5E",X"2E",X"00",X"BF",X"03",X"F0",
		X"91",X"F8",X"57",X"F4",X"74",X"3F",X"42",X"F6",X"91",X"EB",X"43",X"F4",X"E4",X"2F",X"03",X"F8",
		X"95",X"9E",X"45",X"AE",X"0B",X"8E",X"98",X"6F",X"8E",X"0E",X"47",X"2E",X"1A",X"A9",X"E5",X"3F",
		X"D2",X"83",X"D3",X"82",X"DA",X"1F",X"1F",X"C2",X"D5",X"83",X"87",X"83",X"DA",X"5B",X"8E",X"97",
		X"D2",X"91",X"CA",X"87",X"5E",X"A7",X"6A",X"39",X"C5",X"86",X"5A",X"62",X"9A",X"A7",X"6A",X"67",
		X"C5",X"95",X"66",X"9A",X"5A",X"7A",X"9D",X"99",X"C6",X"55",X"8A",X"67",X"5A",X"79",X"E9",X"69",
		X"DA",X"61",X"59",X"8D",X"D8",X"4E",X"1F",X"E9",X"DD",X"88",X"57",X"5A",X"59",X"4F",X"1F",X"E7",
		X"DD",X"86",X"17",X"66",X"59",X"4B",X"5F",X"DE",X"A6",X"A5",X"56",X"5A",X"57",X"4A",X"8F",X"DF",
		X"6A",X"9D",X"56",X"1A",X"8A",X"0A",X"1F",X"EA",X"96",X"8A",X"DD",X"07",X"6A",X"19",X"1F",X"F7",
		X"76",X"95",X"DF",X"50",X"7A",X"56",X"92",X"FF",X"3A",X"55",X"EA",X"16",X"56",X"AA",X"09",X"FF",
		X"A7",X"5A",X"52",X"C1",X"E5",X"9E",X"3D",X"2F",X"B4",X"7C",X"0F",X"81",X"B5",X"66",X"F4",X"3F",
		X"D2",X"9D",X"0F",X"C0",X"F4",X"F4",X"BC",X"3F",X"C3",X"D1",X"CB",X"03",X"E0",X"FC",X"2F",X"4A",
		X"C2",X"D2",X"5F",X"43",X"E0",X"BC",X"2F",X"0F",X"67",X"56",X"98",X"79",X"75",X"E5",X"DB",X"0F",
		X"1A",X"6E",X"07",X"E0",X"75",X"F4",X"3F",X"D0",X"0F",X"D0",X"EF",X"42",X"F0",X"35",X"B8",X"3F",
		X"5F",X"02",X"F6",X"0B",X"C0",X"A9",X"B8",X"3F",X"87",X"C1",X"6F",X"19",X"4B",X"C0",X"BE",X"D0",
		X"67",X"A5",X"66",X"1E",X"62",X"61",X"7E",X"2B",X"67",X"A1",X"75",X"6A",X"62",X"61",X"7E",X"3B",
		X"A5",X"E5",X"68",X"5E",X"56",X"62",X"7A",X"9E",X"A5",X"68",X"99",X"99",X"96",X"66",X"7A",X"9E",
		X"9D",X"99",X"59",X"99",X"98",X"98",X"AA",X"AA",X"27",X"7A",X"56",X"62",X"A1",X"74",X"7E",X"7B",
		X"62",X"6A",X"8A",X"86",X"A0",X"E4",X"2F",X"6F",X"95",X"6B",X"5A",X"82",X"E4",X"A4",X"2F",X"3F",
		X"95",X"7A",X"6A",X"46",X"E1",X"A0",X"2F",X"2F",X"C4",X"AA",X"6A",X"46",X"E1",X"A0",X"3E",X"3F",
		X"C4",X"7D",X"6E",X"06",X"D6",X"94",X"3E",X"3F",X"99",X"72",X"79",X"89",X"5A",X"A1",X"65",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
