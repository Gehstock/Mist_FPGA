library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"06",X"00",X"21",X"00",X"00",X"C3",X"10",X"08",X"31",X"FF",X"4B",X"26",X"50",X"36",X"00",X"CD",
		X"50",X"00",X"21",X"00",X"18",X"0E",X"03",X"CD",X"D0",X"01",X"CD",X"80",X"00",X"3A",X"A2",X"43",
		X"A7",X"CA",X"2D",X"00",X"CD",X"00",X"04",X"CD",X"00",X"27",X"C3",X"1A",X"00",X"3A",X"00",X"78",
		X"E6",X"40",X"CA",X"E0",X"03",X"CD",X"40",X"27",X"00",X"CD",X"60",X"17",X"A7",X"CA",X"46",X"00",
		X"CD",X"88",X"02",X"C3",X"1A",X"00",X"CD",X"E3",X"00",X"C3",X"1A",X"00",X"BF",X"E6",X"00",X"87",
		X"26",X"68",X"36",X"00",X"26",X"60",X"36",X"00",X"26",X"58",X"36",X"00",X"CD",X"6B",X"00",X"26",
		X"50",X"36",X"01",X"CD",X"6B",X"00",X"26",X"50",X"36",X"00",X"C9",X"21",X"F8",X"4B",X"3E",X"3F",
		X"36",X"00",X"2B",X"BC",X"C2",X"70",X"00",X"C9",X"CD",X"00",X"08",X"C3",X"BC",X"06",X"FF",X"FF",
		X"26",X"78",X"7E",X"E6",X"80",X"CA",X"80",X"00",X"7E",X"E6",X"80",X"C2",X"88",X"00",X"26",X"70",
		X"7E",X"21",X"A0",X"43",X"46",X"77",X"2C",X"70",X"2E",X"9B",X"CD",X"00",X"02",X"2E",X"8F",X"7E",
		X"FE",X"09",X"C8",X"D2",X"00",X"00",X"06",X"01",X"CD",X"BB",X"00",X"C8",X"2E",X"8F",X"34",X"7E",
		X"C6",X"20",X"32",X"42",X"41",X"C9",X"00",X"C9",X"00",X"C9",X"FF",X"21",X"A0",X"43",X"7E",X"2F",
		X"A0",X"2C",X"A6",X"C9",X"7E",X"E6",X"0F",X"F6",X"20",X"12",X"CD",X"10",X"02",X"05",X"C8",X"7E",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"F6",X"20",X"12",X"CD",X"10",X"02",X"2B",X"05",X"C2",X"C4",
		X"00",X"C9",X"FF",X"21",X"99",X"43",X"CD",X"00",X"02",X"01",X"01",X"00",X"CD",X"58",X"02",X"CA",
		X"E1",X"01",X"01",X"02",X"00",X"11",X"1F",X"01",X"CD",X"60",X"02",X"D2",X"96",X"01",X"01",X"20",
		X"01",X"CD",X"58",X"02",X"CA",X"88",X"06",X"0E",X"B0",X"CD",X"58",X"02",X"CA",X"E1",X"01",X"0E",
		X"C0",X"11",X"E0",X"01",X"CD",X"60",X"02",X"D2",X"0C",X"1B",X"01",X"00",X"02",X"11",X"C0",X"03",
		X"CD",X"60",X"02",X"D2",X"D0",X"1A",X"01",X"00",X"04",X"11",X"AF",X"04",X"CD",X"60",X"02",X"D2",
		X"C0",X"03",X"01",X"E6",X"04",X"11",X"FF",X"FF",X"CD",X"60",X"02",X"D2",X"B0",X"03",X"C9",X"FF",
		X"CD",X"A0",X"03",X"CD",X"80",X"00",X"CD",X"80",X"03",X"21",X"A3",X"43",X"36",X"02",X"2C",X"36",
		X"00",X"00",X"00",X"00",X"2E",X"B8",X"06",X"08",X"CD",X"D8",X"05",X"2E",X"BA",X"36",X"10",X"2E",
		X"BE",X"3A",X"00",X"78",X"E6",X"0C",X"07",X"07",X"C6",X"30",X"77",X"26",X"58",X"36",X"00",X"CD",
		X"80",X"00",X"C9",X"7E",X"E6",X"7F",X"06",X"CE",X"FE",X"1F",X"D8",X"06",X"FE",X"C8",X"06",X"AE",
		X"FE",X"5F",X"D8",X"06",X"FE",X"C8",X"06",X"CE",X"FE",X"7F",X"D8",X"06",X"FE",X"2D",X"7E",X"FE",
		X"09",X"C0",X"06",X"7E",X"C9",X"FF",X"7E",X"E6",X"1F",X"FE",X"06",X"D8",X"5F",X"7E",X"E6",X"E0",
		X"4F",X"2D",X"46",X"2E",X"A8",X"70",X"2C",X"71",X"01",X"60",X"18",X"CD",X"06",X"02",X"7E",X"2D",
		X"66",X"6F",X"7B",X"56",X"2C",X"5E",X"2D",X"4F",X"85",X"6F",X"79",X"D6",X"06",X"4F",X"CA",X"C8",
		X"01",X"CD",X"17",X"02",X"0D",X"C2",X"C1",X"01",X"7E",X"12",X"C3",X"40",X"17",X"C2",X"C0",X"01",
		X"56",X"2C",X"5E",X"7D",X"C6",X"05",X"6F",X"06",X"1A",X"CD",X"ED",X"01",X"0D",X"C2",X"D0",X"01",
		X"C9",X"CD",X"40",X"01",X"21",X"60",X"19",X"0E",X"03",X"C3",X"D0",X"01",X"FF",X"7E",X"12",X"23",
		X"CD",X"17",X"02",X"05",X"C2",X"ED",X"01",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"34",X"C0",X"2D",X"34",X"2C",X"C9",X"7E",X"81",X"77",X"2D",X"7E",X"88",X"77",X"2C",X"C9",X"FF",
		X"7B",X"C6",X"20",X"5F",X"D0",X"14",X"C9",X"7B",X"D6",X"20",X"5F",X"D0",X"15",X"C9",X"FF",X"FF",
		X"AF",X"7E",X"81",X"27",X"77",X"2D",X"7E",X"88",X"27",X"77",X"2D",X"7E",X"CE",X"00",X"27",X"77",
		X"2C",X"2C",X"C9",X"FF",X"FF",X"FF",X"37",X"3E",X"99",X"CE",X"00",X"91",X"86",X"27",X"77",X"2D",
		X"3E",X"99",X"CE",X"00",X"90",X"86",X"27",X"77",X"2D",X"3E",X"99",X"CE",X"00",X"86",X"27",X"77",
		X"2C",X"2C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"B9",X"C0",X"2D",X"7E",X"2C",X"B8",X"C9",
		X"CD",X"70",X"02",X"D8",X"CD",X"77",X"02",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"91",X"2D",X"7E",X"98",X"2C",X"C9",X"7B",X"96",X"2D",X"7A",X"9E",X"2C",X"C9",X"FF",X"FF",
		X"7D",X"B9",X"C0",X"7C",X"B8",X"C9",X"FF",X"FF",X"CD",X"40",X"01",X"21",X"C0",X"19",X"0E",X"02",
		X"CD",X"D0",X"01",X"0E",X"02",X"CD",X"60",X"17",X"FE",X"02",X"DA",X"A7",X"02",X"21",X"A0",X"1B",
		X"0E",X"01",X"CD",X"D0",X"01",X"0E",X"06",X"3A",X"00",X"70",X"2F",X"A1",X"C8",X"CD",X"CB",X"02",
		X"CD",X"F0",X"02",X"CD",X"2E",X"03",X"CD",X"50",X"03",X"CD",X"40",X"01",X"26",X"50",X"36",X"01",
		X"CD",X"40",X"01",X"26",X"50",X"36",X"00",X"C9",X"FF",X"FF",X"FF",X"0E",X"01",X"FE",X"02",X"CA",
		X"D4",X"02",X"0E",X"02",X"21",X"A2",X"43",X"71",X"3A",X"00",X"78",X"E6",X"10",X"CA",X"E3",X"02",
		X"79",X"07",X"4F",X"2E",X"8F",X"7E",X"91",X"77",X"C6",X"20",X"32",X"42",X"41",X"C9",X"FF",X"FF",
		X"11",X"83",X"43",X"21",X"8B",X"43",X"CD",X"14",X"03",X"D4",X"20",X"03",X"1E",X"87",X"2E",X"FF",
		X"CD",X"14",X"03",X"D4",X"20",X"03",X"2E",X"8B",X"11",X"41",X"41",X"06",X"06",X"CD",X"C4",X"00",
		X"C9",X"FF",X"FF",X"FF",X"1A",X"96",X"1D",X"2D",X"1A",X"9E",X"1D",X"2D",X"1A",X"9E",X"C9",X"FF",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"23",X"1A",X"77",X"C9",X"FF",X"FF",X"FF",X"21",X"80",
		X"43",X"36",X"00",X"23",X"7D",X"FE",X"88",X"C2",X"31",X"03",X"2E",X"83",X"11",X"61",X"42",X"06",
		X"06",X"CD",X"C4",X"00",X"2E",X"87",X"11",X"21",X"40",X"06",X"06",X"CD",X"C4",X"00",X"C9",X"FF",
		X"3A",X"00",X"78",X"E6",X"03",X"C6",X"03",X"47",X"21",X"90",X"43",X"70",X"2E",X"A2",X"7E",X"FE",
		X"01",X"CA",X"67",X"03",X"2E",X"91",X"70",X"2E",X"90",X"7E",X"F6",X"20",X"32",X"A2",X"42",X"2C",
		X"7E",X"F6",X"20",X"32",X"62",X"40",X"C9",X"21",X"8C",X"43",X"77",X"2C",X"77",X"C9",X"FF",X"FF",
		X"21",X"3F",X"43",X"11",X"1F",X"00",X"01",X"3F",X"03",X"72",X"2B",X"72",X"2B",X"7D",X"A3",X"B8",
		X"C2",X"89",X"03",X"72",X"2B",X"2B",X"2B",X"2B",X"7C",X"B9",X"C2",X"89",X"03",X"C9",X"FF",X"FF",
		X"21",X"3F",X"4B",X"11",X"47",X"00",X"72",X"2B",X"72",X"2B",X"7C",X"BB",X"C2",X"A6",X"03",X"C9",
		X"CD",X"73",X"01",X"21",X"A0",X"43",X"7E",X"E6",X"01",X"B0",X"77",X"C3",X"00",X"04",X"FF",X"FF",
		X"7E",X"0F",X"E6",X"1C",X"FE",X"10",X"DA",X"CC",X"03",X"2F",X"E6",X"0C",X"F6",X"20",X"6F",X"26",
		X"14",X"11",X"52",X"42",X"E5",X"CD",X"DC",X"07",X"E1",X"11",X"32",X"41",X"C3",X"DC",X"07",X"FF",
		X"3E",X"0F",X"21",X"8C",X"43",X"77",X"32",X"00",X"60",X"3E",X"8F",X"2C",X"77",X"32",X"00",X"68",
		X"3E",X"7F",X"30",X"C3",X"38",X"00",X"2E",X"BA",X"72",X"2C",X"73",X"C3",X"80",X"03",X"80",X"FF",
		X"21",X"0E",X"04",X"3A",X"A4",X"43",X"07",X"85",X"6F",X"7E",X"2C",X"6E",X"67",X"E9",X"04",X"30",
		X"04",X"AC",X"05",X"10",X"00",X"78",X"0A",X"EA",X"0B",X"60",X"24",X"00",X"05",X"D0",X"FF",X"FF",
		X"04",X"04",X"00",X"00",X"06",X"02",X"04",X"00",X"06",X"06",X"02",X"02",X"02",X"04",X"06",X"04",
		X"21",X"A4",X"43",X"36",X"01",X"2C",X"36",X"80",X"2E",X"A3",X"7E",X"36",X"00",X"FE",X"02",X"C8",
		X"77",X"2D",X"7E",X"FE",X"01",X"C8",X"2C",X"7E",X"A7",X"CA",X"A0",X"04",X"2E",X"90",X"7E",X"A7",
		X"C8",X"2E",X"A3",X"36",X"00",X"01",X"00",X"01",X"CD",X"60",X"04",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"21",X"00",X"50",X"11",X"20",X"43",X"70",X"1A",X"71",X"12",X"1C",X"7B",X"E6",X"03",X"C2",X"66",
		X"04",X"7B",X"E6",X"F0",X"D6",X"20",X"5F",X"D2",X"66",X"04",X"15",X"7A",X"FE",X"3F",X"C2",X"66",
		X"04",X"11",X"80",X"43",X"70",X"1A",X"71",X"12",X"1C",X"7B",X"FE",X"B8",X"C2",X"84",X"04",X"11",
		X"C0",X"4B",X"70",X"1A",X"71",X"12",X"1C",X"7B",X"FE",X"00",X"C2",X"92",X"04",X"C9",X"FF",X"FF",
		X"2E",X"A3",X"36",X"01",X"01",X"01",X"00",X"CD",X"60",X"04",X"C9",X"FF",X"21",X"A5",X"43",X"35",
		X"7E",X"2D",X"36",X"02",X"A7",X"C8",X"36",X"01",X"FE",X"7F",X"CA",X"F0",X"07",X"2E",X"9A",X"36",
		X"00",X"2C",X"36",X"00",X"E6",X"08",X"C2",X"E6",X"04",X"CD",X"08",X"05",X"00",X"21",X"A3",X"43",
		X"7E",X"A7",X"2E",X"83",X"11",X"61",X"42",X"CA",X"DF",X"04",X"2E",X"87",X"11",X"21",X"40",X"06",
		X"06",X"CD",X"C4",X"00",X"C9",X"FF",X"21",X"A3",X"43",X"7E",X"A7",X"11",X"61",X"42",X"CA",X"F4",
		X"04",X"11",X"21",X"40",X"06",X"06",X"CD",X"FB",X"04",X"C9",X"FF",X"3E",X"00",X"12",X"CD",X"10",
		X"02",X"05",X"C2",X"FB",X"04",X"C9",X"FF",X"FF",X"21",X"00",X"18",X"0E",X"01",X"C3",X"D0",X"01",
		X"21",X"A4",X"43",X"36",X"03",X"CD",X"EA",X"05",X"CD",X"80",X"05",X"CD",X"B8",X"05",X"3A",X"BB",
		X"43",X"A7",X"C8",X"C3",X"C4",X"32",X"FF",X"FF",X"FF",X"FF",X"21",X"38",X"05",X"11",X"C0",X"43",
		X"06",X"04",X"CD",X"E0",X"05",X"C3",X"A0",X"09",X"0C",X"10",X"64",X"D8",X"CD",X"42",X"05",X"C3",
		X"17",X"06",X"21",X"B0",X"43",X"56",X"2C",X"5E",X"21",X"40",X"1B",X"01",X"0B",X"04",X"C3",X"D6",
		X"0A",X"05",X"78",X"8E",X"23",X"47",X"7C",X"FE",X"40",X"C2",X"52",X"05",X"78",X"FE",X"40",X"CA",
		X"08",X"00",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"21",X"A2",X"43",X"7E",X"A7",X"C8",X"2E",X"B5",X"3A",X"83",X"43",X"E6",X"70",X"86",X"77",X"C9",
		X"21",X"B8",X"43",X"7E",X"E6",X"06",X"07",X"07",X"C6",X"98",X"6F",X"26",X"05",X"11",X"B0",X"43",
		X"06",X"08",X"CD",X"E0",X"05",X"C3",X"70",X"05",X"4B",X"3F",X"1D",X"D8",X"29",X"00",X"20",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"00",X"4A",X"46",X"1B",X"40",X"29",X"80",X"0C",X"00",
		X"4B",X"3F",X"1C",X"20",X"FF",X"FF",X"20",X"00",X"21",X"70",X"4B",X"06",X"08",X"36",X"04",X"2C",
		X"36",X"08",X"2C",X"36",X"80",X"2C",X"36",X"80",X"2C",X"05",X"C2",X"BD",X"05",X"C9",X"FF",X"FF",
		X"CD",X"F4",X"31",X"C3",X"BC",X"06",X"FF",X"FF",X"AF",X"77",X"23",X"05",X"C2",X"D9",X"05",X"C9",
		X"7E",X"12",X"23",X"13",X"05",X"C2",X"E0",X"05",X"C9",X"FF",X"21",X"C4",X"43",X"06",X"3C",X"CD",
		X"D8",X"05",X"21",X"50",X"43",X"06",X"30",X"CD",X"D8",X"05",X"2E",X"92",X"06",X"06",X"CD",X"D8",
		X"05",X"2E",X"9A",X"06",X"04",X"CD",X"D8",X"05",X"21",X"50",X"4B",X"06",X"9C",X"C3",X"D8",X"05",
		X"FF",X"FF",X"FF",X"FF",X"CD",X"50",X"06",X"AF",X"32",X"00",X"58",X"32",X"B9",X"43",X"21",X"B6",
		X"43",X"35",X"C0",X"2E",X"A4",X"36",X"02",X"2E",X"B8",X"7E",X"34",X"E6",X"0F",X"C0",X"11",X"3B",
		X"4A",X"01",X"0A",X"05",X"C5",X"D5",X"3E",X"00",X"12",X"13",X"05",X"C2",X"36",X"06",X"D1",X"C1",
		X"CD",X"17",X"02",X"0D",X"C2",X"34",X"06",X"C9",X"AF",X"2C",X"77",X"32",X"00",X"58",X"C9",X"FF",
		X"21",X"B0",X"43",X"56",X"2C",X"5E",X"2C",X"7E",X"2C",X"6E",X"67",X"7E",X"06",X"01",X"A7",X"C2",
		X"64",X"06",X"23",X"46",X"FE",X"3F",X"C2",X"6B",X"06",X"23",X"46",X"4F",X"23",X"79",X"12",X"CD",
		X"17",X"02",X"05",X"C2",X"6D",X"06",X"7A",X"FE",X"47",X"C2",X"5B",X"06",X"EB",X"21",X"B1",X"43",
		X"35",X"2C",X"72",X"2C",X"73",X"C9",X"47",X"20",X"01",X"06",X"02",X"11",X"F0",X"42",X"21",X"B0",
		X"06",X"CD",X"D6",X"0A",X"21",X"B0",X"43",X"36",X"4B",X"23",X"36",X"3A",X"23",X"36",X"16",X"23",
		X"36",X"40",X"3E",X"09",X"F5",X"CD",X"50",X"06",X"F1",X"3D",X"C2",X"A4",X"06",X"C9",X"FF",X"FF",
		X"60",X"70",X"61",X"00",X"C0",X"C8",X"C1",X"C9",X"A2",X"00",X"A3",X"00",X"21",X"B8",X"43",X"7E",
		X"07",X"E6",X"0C",X"47",X"FE",X"0C",X"CA",X"EA",X"06",X"2C",X"2C",X"7E",X"2C",X"86",X"3D",X"FE",
		X"03",X"DA",X"D6",X"06",X"3E",X"03",X"B0",X"C6",X"20",X"6F",X"26",X"04",X"46",X"3A",X"A3",X"43",
		X"E6",X"01",X"B0",X"32",X"00",X"50",X"C9",X"FF",X"CD",X"F4",X"7E",X"E6",X"10",X"0F",X"0F",X"0F",
		X"B0",X"47",X"2E",X"A4",X"7E",X"FE",X"07",X"C2",X"FB",X"06",X"04",X"78",X"C3",X"D7",X"06",X"FF",
		X"01",X"C0",X"43",X"11",X"E0",X"43",X"CD",X"18",X"07",X"79",X"C6",X"04",X"4F",X"C6",X"20",X"5F",
		X"50",X"FE",X"EC",X"C2",X"06",X"07",X"C9",X"C9",X"CD",X"20",X"07",X"C3",X"40",X"07",X"E6",X"EF",
		X"0A",X"67",X"E6",X"10",X"C8",X"7C",X"E6",X"EF",X"02",X"07",X"07",X"07",X"E6",X"07",X"C6",X"38",
		X"6F",X"26",X"07",X"6E",X"E9",X"6C",X"FF",X"8A",X"63",X"79",X"FF",X"9E",X"BE",X"FF",X"FF",X"FF",
		X"0A",X"67",X"E6",X"08",X"C8",X"7C",X"E6",X"07",X"67",X"0F",X"0F",X"0F",X"B4",X"F6",X"18",X"02",
		X"03",X"7C",X"C6",X"5B",X"6F",X"26",X"07",X"6E",X"E9",X"5E",X"0A",X"6D",X"88",X"FF",X"AA",X"D2",
		X"FF",X"FF",X"FF",X"EB",X"56",X"23",X"5E",X"2B",X"AF",X"12",X"EB",X"C9",X"EB",X"EB",X"23",X"23",
		X"56",X"23",X"5E",X"0A",X"12",X"0B",X"C9",X"12",X"23",X"EB",X"56",X"23",X"5E",X"2B",X"AF",X"12",
		X"CD",X"17",X"02",X"AF",X"12",X"EB",X"C9",X"23",X"EB",X"23",X"23",X"56",X"23",X"5E",X"0A",X"6F",
		X"26",X"14",X"7E",X"12",X"23",X"CD",X"17",X"02",X"7E",X"12",X"0B",X"C9",X"FF",X"EB",X"EB",X"56",
		X"23",X"5E",X"2B",X"AF",X"12",X"13",X"12",X"EB",X"C9",X"FF",X"EB",X"23",X"23",X"56",X"23",X"5E",
		X"0A",X"6F",X"26",X"14",X"7E",X"12",X"23",X"13",X"7E",X"12",X"0B",X"C9",X"23",X"13",X"EB",X"56",
		X"23",X"5E",X"2B",X"AF",X"12",X"13",X"12",X"CD",X"17",X"02",X"AF",X"12",X"1B",X"12",X"EB",X"C9",
		X"CD",X"4C",X"EB",X"23",X"23",X"56",X"23",X"5E",X"0A",X"6F",X"26",X"14",X"7E",X"12",X"23",X"13",
		X"7E",X"12",X"23",X"1B",X"CD",X"17",X"02",X"7E",X"12",X"23",X"13",X"7E",X"12",X"0B",X"C9",X"FF",
		X"3A",X"B9",X"43",X"32",X"00",X"58",X"CD",X"80",X"03",X"C3",X"2A",X"05",X"FF",X"FF",X"FF",X"FF",
		X"21",X"14",X"08",X"3A",X"B8",X"43",X"07",X"E6",X"1E",X"85",X"6F",X"7E",X"2C",X"6E",X"67",X"E9",
		X"C3",X"60",X"14",X"FF",X"06",X"14",X"08",X"34",X"22",X"80",X"34",X"00",X"05",X"3C",X"08",X"34",
		X"23",X"60",X"23",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"CD",X"76",X"08",X"CD",X"F0",X"0D",X"CD",X"AB",X"23",X"21",X"92",X"43",
		X"46",X"34",X"3A",X"BA",X"43",X"A7",X"CA",X"F6",X"21",X"FE",X"02",X"DC",X"58",X"0D",X"78",X"0F",
		X"DA",X"64",X"08",X"CD",X"50",X"0A",X"CD",X"00",X"30",X"CD",X"08",X"0F",X"CD",X"50",X"25",X"C3",
		X"40",X"0C",X"FF",X"FF",X"CD",X"1C",X"0D",X"CD",X"70",X"0D",X"CD",X"6C",X"0A",X"CD",X"78",X"0F",
		X"C3",X"80",X"20",X"FF",X"FF",X"FF",X"CD",X"00",X"07",X"CD",X"86",X"08",X"CD",X"A0",X"08",X"CD",
		X"A0",X"09",X"CD",X"7A",X"09",X"C9",X"21",X"EB",X"43",X"06",X"03",X"56",X"2B",X"5E",X"2B",X"72",
		X"2B",X"73",X"2B",X"05",X"C2",X"8B",X"08",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"E0",X"08",X"21",X"C4",X"43",X"CD",X"30",X"09",X"21",X"C8",X"43",X"3A",X"B8",X"43",X"E6",
		X"0F",X"FE",X"05",X"CA",X"30",X"09",X"7E",X"E6",X"08",X"C2",X"64",X"09",X"C9",X"FF",X"FF",X"FF",
		X"CD",X"50",X"0A",X"CD",X"00",X"30",X"CD",X"08",X"0F",X"CD",X"1C",X"0D",X"CD",X"70",X"0D",X"CD",
		X"6C",X"0A",X"3A",X"92",X"43",X"0F",X"DA",X"5C",X"08",X"C3",X"6D",X"08",X"CD",X"EA",X"08",X"CD",
		X"21",X"B8",X"43",X"7E",X"E6",X"0F",X"FE",X"06",X"D2",X"B0",X"22",X"2E",X"C2",X"CD",X"F8",X"08",
		X"01",X"00",X"16",X"C3",X"26",X"09",X"FF",X"FF",X"3A",X"A0",X"43",X"2F",X"E6",X"60",X"C8",X"E6",
		X"40",X"CA",X"0A",X"09",X"7E",X"FE",X"09",X"D8",X"35",X"C9",X"7E",X"FE",X"C0",X"D0",X"34",X"C9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"E6",X"07",X"81",X"4F",X"0A",X"2D",X"77",X"C9",X"FF",
		X"7E",X"E6",X"08",X"C2",X"64",X"09",X"EB",X"06",X"10",X"CD",X"BB",X"00",X"C8",X"7E",X"E6",X"EF",
		X"77",X"1A",X"F6",X"08",X"12",X"13",X"13",X"3A",X"C2",X"43",X"C6",X"04",X"12",X"13",X"3A",X"C3",
		X"43",X"D6",X"08",X"12",X"1B",X"EB",X"01",X"20",X"16",X"CD",X"26",X"09",X"3E",X"30",X"32",X"61",
		X"43",X"C9",X"FF",X"FF",X"2C",X"2C",X"2C",X"7E",X"D6",X"08",X"77",X"FE",X"1F",X"D0",X"2D",X"2D",
		X"2D",X"7E",X"E6",X"F7",X"77",X"C9",X"FF",X"FF",X"7E",X"E6",X"3A",X"C2",X"43",X"47",X"E6",X"07",
		X"07",X"21",X"38",X"0B",X"85",X"6F",X"78",X"96",X"32",X"9E",X"43",X"23",X"78",X"86",X"32",X"9F",
		X"43",X"C9",X"32",X"9F",X"43",X"C9",X"C6",X"00",X"11",X"65",X"41",X"06",X"04",X"C3",X"C4",X"00",
		X"01",X"C2",X"43",X"11",X"E2",X"43",X"CD",X"BA",X"09",X"0E",X"C6",X"1E",X"E6",X"CD",X"BA",X"09",
		X"0E",X"CA",X"1E",X"EA",X"C3",X"BA",X"09",X"FF",X"FF",X"FF",X"21",X"00",X"0A",X"0A",X"E6",X"F8",
		X"0F",X"0F",X"85",X"6F",X"7E",X"12",X"03",X"13",X"23",X"0A",X"E6",X"F8",X"0F",X"0F",X"0F",X"86",
		X"12",X"C9",X"FF",X"FF",X"3A",X"B8",X"43",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"3C",X"47",X"0E",
		X"00",X"16",X"05",X"3A",X"BC",X"43",X"0F",X"5F",X"D2",X"F0",X"09",X"78",X"81",X"27",X"47",X"4F",
		X"7B",X"15",X"C2",X"E6",X"09",X"21",X"DE",X"4B",X"71",X"2C",X"36",X"00",X"C3",X"98",X"09",X"00",
		X"43",X"20",X"43",X"00",X"42",X"E0",X"42",X"C0",X"42",X"A0",X"42",X"80",X"42",X"60",X"42",X"40",
		X"42",X"20",X"42",X"00",X"41",X"E0",X"41",X"C0",X"41",X"A0",X"41",X"80",X"41",X"60",X"41",X"40",
		X"41",X"20",X"41",X"00",X"40",X"E0",X"40",X"C0",X"40",X"A0",X"40",X"80",X"40",X"60",X"40",X"40",
		X"40",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"2C",X"2D",X"2E",X"2D",X"2E",X"2F",X"2F",X"30",X"31",X"32",X"31",X"30",X"31",X"2C",X"33",
		X"01",X"70",X"4B",X"11",X"B0",X"4B",X"C5",X"CD",X"18",X"07",X"C1",X"79",X"C6",X"04",X"4F",X"C6",
		X"40",X"5F",X"50",X"FE",X"D0",X"C2",X"56",X"0A",X"C9",X"FF",X"FF",X"FF",X"01",X"70",X"4B",X"11",
		X"B3",X"4B",X"C5",X"D5",X"0A",X"E6",X"18",X"CA",X"8A",X"0A",X"EB",X"56",X"2B",X"5E",X"2B",X"72",
		X"2B",X"73",X"EB",X"13",X"13",X"03",X"03",X"CD",X"BA",X"09",X"D1",X"C1",X"79",X"C6",X"04",X"4F",
		X"7B",X"C6",X"04",X"5F",X"FE",X"D3",X"C2",X"72",X"0A",X"C9",X"FF",X"FF",X"21",X"DB",X"4B",X"01",
		X"D4",X"4B",X"0A",X"FE",X"48",X"C2",X"E6",X"0E",X"36",X"04",X"EB",X"13",X"0B",X"CD",X"BA",X"09",
		X"1B",X"3E",X"49",X"12",X"3A",X"D2",X"4B",X"32",X"62",X"43",X"C9",X"FF",X"21",X"DD",X"4B",X"5E",
		X"2D",X"56",X"2D",X"1A",X"C6",X"14",X"86",X"6F",X"26",X"0A",X"7E",X"12",X"3A",X"DB",X"4B",X"A7",
		X"C2",X"90",X"0E",X"C9",X"FF",X"FF",X"D5",X"C5",X"7E",X"12",X"23",X"13",X"05",X"C2",X"D8",X"0A",
		X"C1",X"D1",X"CD",X"17",X"02",X"0D",X"C2",X"D6",X"0A",X"C9",X"21",X"E2",X"43",X"56",X"2C",X"5E",
		X"2E",X"A5",X"35",X"7E",X"CA",X"15",X"0B",X"FE",X"1F",X"DA",X"80",X"03",X"CA",X"A0",X"0B",X"D6",
		X"20",X"C3",X"B8",X"0B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"2D",X"36",X"05",X"2D",X"7E",X"C6",X"90",X"6F",X"7E",X"A7",X"C8",
		X"35",X"E5",X"CD",X"67",X"03",X"E1",X"7E",X"A7",X"C8",X"2E",X"A4",X"36",X"00",X"C9",X"FF",X"FF",
		X"FF",X"F0",X"E0",X"B0",X"C0",X"D0",X"C0",X"B0",X"00",X"08",X"01",X"09",X"01",X"09",X"02",X"0A",
		X"02",X"0A",X"01",X"09",X"01",X"09",X"00",X"08",X"2E",X"BA",X"36",X"21",X"B8",X"43",X"7E",X"FE",
		X"10",X"D8",X"78",X"87",X"27",X"47",X"7E",X"FE",X"30",X"D8",X"78",X"87",X"27",X"47",X"C9",X"FF",
		X"21",X"A5",X"43",X"34",X"7E",X"FE",X"40",X"CA",X"A0",X"03",X"21",X"00",X"1A",X"0E",X"01",X"FE",
		X"80",X"C2",X"95",X"0B",X"21",X"A4",X"43",X"36",X"00",X"2E",X"90",X"7E",X"2C",X"B6",X"C0",X"AF",
		X"2E",X"98",X"77",X"2C",X"77",X"2E",X"A2",X"77",X"2C",X"7E",X"A7",X"C8",X"36",X"00",X"01",X"00",
		X"01",X"CD",X"60",X"04",X"C9",X"CD",X"D0",X"01",X"CD",X"E4",X"01",X"C3",X"88",X"16",X"FF",X"FF",
		X"21",X"B8",X"43",X"7E",X"E6",X"0E",X"C8",X"FE",X"04",X"DA",X"AD",X"0B",X"35",X"2C",X"AF",X"77",
		X"32",X"00",X"58",X"C3",X"A0",X"03",X"FF",X"FF",X"0F",X"DA",X"78",X"0F",X"E6",X"7E",X"C6",X"A0",
		X"6F",X"26",X"2A",X"7E",X"23",X"6E",X"67",X"FE",X"17",X"CA",X"DC",X"0B",X"01",X"1F",X"00",X"EB",
		X"09",X"EB",X"01",X"04",X"03",X"C3",X"D6",X"0A",X"FF",X"FF",X"FF",X"FF",X"01",X"5D",X"00",X"EB",
		X"09",X"EB",X"01",X"08",X"06",X"CD",X"EE",X"0B",X"CD",X"EE",X"0B",X"C3",X"D6",X"0A",X"7A",X"FE",
		X"43",X"C0",X"7B",X"FE",X"40",X"D8",X"D6",X"20",X"5F",X"7D",X"80",X"6F",X"0D",X"C9",X"FF",X"FE",
		X"7E",X"D6",X"03",X"BA",X"D0",X"C6",X"05",X"BA",X"D8",X"23",X"7E",X"2B",X"D6",X"08",X"BB",X"D0",
		X"C6",X"10",X"BB",X"D8",X"2B",X"7E",X"23",X"11",X"08",X"39",X"FE",X"30",X"DA",X"2A",X"0C",X"11",
		X"03",X"53",X"FE",X"C0",X"DA",X"2A",X"0C",X"11",X"15",X"1F",X"3A",X"BA",X"43",X"FE",X"02",X"D2",
		X"A4",X"0E",X"3A",X"B8",X"43",X"E6",X"70",X"C6",X"10",X"83",X"5F",X"16",X"1A",X"C3",X"A4",X"0E",
		X"21",X"FF",X"43",X"06",X"05",X"CD",X"8B",X"08",X"CD",X"56",X"0C",X"CD",X"6B",X"0C",X"CD",X"D8",
		X"0C",X"C9",X"FF",X"FF",X"FF",X"FF",X"21",X"CC",X"43",X"E5",X"CD",X"84",X"0C",X"E1",X"7D",X"C6",
		X"04",X"6F",X"FE",X"E0",X"C2",X"59",X"0C",X"C9",X"FF",X"FF",X"FF",X"01",X"CE",X"43",X"11",X"EE",
		X"43",X"CD",X"BA",X"09",X"03",X"03",X"03",X"13",X"13",X"13",X"79",X"FE",X"E2",X"C2",X"71",X"0C",
		X"C9",X"FF",X"FF",X"FF",X"7E",X"E6",X"08",X"C8",X"00",X"00",X"2C",X"7E",X"EE",X"04",X"77",X"2C",
		X"2C",X"7E",X"C6",X"04",X"77",X"FE",X"F9",X"D2",X"6E",X"09",X"2D",X"47",X"CD",X"B4",X"0C",X"78",
		X"FE",X"B0",X"D8",X"C3",X"00",X"20",X"4E",X"0A",X"EB",X"2C",X"FE",X"E8",X"D2",X"6E",X"09",X"C9",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"DC",X"D8",X"FE",X"E9",X"D0",X"3A",X"9F",X"43",X"BE",X"D8",X"3A",
		X"9E",X"43",X"BE",X"D0",X"3E",X"04",X"32",X"A4",X"43",X"3E",X"60",X"32",X"A5",X"43",X"3E",X"FF",
		X"32",X"63",X"43",X"C9",X"FF",X"FF",X"FF",X"FF",X"01",X"CC",X"43",X"11",X"EC",X"43",X"C5",X"CD",
		X"18",X"07",X"C1",X"79",X"C6",X"04",X"4F",X"C6",X"20",X"5F",X"50",X"A7",X"C2",X"DE",X"0C",X"C9",
		X"21",X"DC",X"4B",X"36",X"49",X"2C",X"36",X"A9",X"21",X"9D",X"43",X"3A",X"DE",X"4B",X"77",X"2E",
		X"A4",X"36",X"06",X"2C",X"36",X"60",X"2E",X"63",X"36",X"FF",X"2E",X"B8",X"34",X"E1",X"E1",X"C9",
		X"CD",X"80",X"00",X"CD",X"A0",X"03",X"E1",X"E1",X"C9",X"FF",X"FF",X"FF",X"01",X"70",X"4B",X"21",
		X"50",X"4B",X"CD",X"30",X"0D",X"0C",X"0C",X"2C",X"3E",X"90",X"B9",X"C2",X"22",X"0D",X"C9",X"FF",
		X"56",X"23",X"0A",X"03",X"03",X"E6",X"08",X"C8",X"5E",X"EB",X"7E",X"07",X"C6",X"00",X"6F",X"26",
		X"17",X"0A",X"86",X"02",X"03",X"23",X"0A",X"86",X"02",X"EB",X"57",X"0B",X"0A",X"B2",X"E6",X"07",
		X"C0",X"34",X"C0",X"2D",X"34",X"2C",X"C9",X"EB",X"2E",X"94",X"78",X"0F",X"DA",X"61",X"0D",X"36",
		X"01",X"7E",X"A7",X"C8",X"2E",X"B8",X"7E",X"E6",X"F0",X"C8",X"E1",X"C3",X"C0",X"08",X"FF",X"FF",
		X"01",X"70",X"4B",X"21",X"50",X"4B",X"CD",X"86",X"0D",X"79",X"C6",X"04",X"4F",X"3E",X"90",X"B9",
		X"C2",X"76",X"0D",X"C9",X"FF",X"FF",X"56",X"23",X"5E",X"23",X"0A",X"E6",X"08",X"C8",X"EB",X"7E",
		X"A7",X"CA",X"D8",X"0D",X"07",X"C6",X"C0",X"6F",X"26",X"16",X"03",X"03",X"03",X"7E",X"23",X"0F",
		X"DA",X"B4",X"0D",X"0F",X"DA",X"C6",X"0D",X"0A",X"0F",X"E6",X"03",X"86",X"0B",X"C3",X"CC",X"0D",
		X"0F",X"E6",X"03",X"86",X"0A",X"0F",X"E6",X"03",X"86",X"67",X"0B",X"0A",X"07",X"E6",X"0C",X"84",
		X"C3",X"CC",X"0D",X"E6",X"04",X"84",X"0B",X"0A",X"0F",X"E6",X"03",X"86",X"6F",X"26",X"16",X"7E",
		X"0B",X"02",X"0B",X"EB",X"C9",X"7E",X"0B",X"02",X"0A",X"E6",X"F7",X"02",X"EB",X"C9",X"1B",X"1B",
		X"3A",X"94",X"43",X"12",X"67",X"13",X"36",X"00",X"C9",X"12",X"6F",X"13",X"7E",X"C9",X"FF",X"FF",
		X"01",X"C4",X"43",X"21",X"E6",X"43",X"CD",X"04",X"0E",X"01",X"C8",X"43",X"21",X"EA",X"43",X"CD",
		X"04",X"0E",X"C9",X"CC",X"0A",X"E6",X"08",X"C8",X"7E",X"C6",X"08",X"57",X"2C",X"5E",X"1A",X"D6",
		X"2C",X"FE",X"12",X"CA",X"3C",X"0E",X"DA",X"50",X"0E",X"2D",X"56",X"1A",X"FE",X"60",X"D8",X"FE",
		X"D0",X"D0",X"E6",X"07",X"07",X"07",X"C6",X"C0",X"6F",X"26",X"2A",X"03",X"03",X"0A",X"E6",X"07",
		X"BE",X"D0",X"23",X"BE",X"D8",X"C3",X"70",X"0E",X"FF",X"FF",X"FF",X"FF",X"AF",X"12",X"0A",X"E6",
		X"F7",X"02",X"2D",X"56",X"3E",X"FF",X"32",X"66",X"43",X"06",X"88",X"C3",X"2D",X"20",X"23",X"3E",
		X"FE",X"03",X"C2",X"3E",X"0E",X"E5",X"7B",X"D6",X"69",X"07",X"07",X"07",X"6F",X"26",X"3E",X"7E",
		X"21",X"BC",X"43",X"B6",X"77",X"E1",X"FE",X"1F",X"CA",X"F8",X"0C",X"C3",X"3E",X"0E",X"FF",X"FF",
		X"23",X"0A",X"E6",X"F8",X"86",X"57",X"03",X"0A",X"E6",X"F8",X"5F",X"21",X"70",X"4B",X"7E",X"23",
		X"23",X"E6",X"08",X"C4",X"00",X"0C",X"23",X"23",X"3E",X"90",X"BD",X"C2",X"7E",X"0E",X"C9",X"FF",
		X"3A",X"92",X"43",X"E6",X"0C",X"0F",X"0F",X"C6",X"48",X"6F",X"26",X"0A",X"7E",X"32",X"A6",X"49",
		X"C9",X"02",X"0C",X"00",X"2B",X"2B",X"0B",X"0B",X"0B",X"0A",X"E6",X"F7",X"02",X"7E",X"E6",X"F7",
		X"77",X"7D",X"C6",X"42",X"6F",X"46",X"23",X"4E",X"21",X"70",X"43",X"7E",X"E6",X"1F",X"CA",X"D5",
		X"0E",X"2E",X"74",X"7E",X"E6",X"1F",X"CA",X"D5",X"0E",X"2E",X"78",X"7E",X"E6",X"1F",X"CA",X"D5",
		X"0E",X"2E",X"7C",X"00",X"00",X"72",X"2C",X"73",X"2C",X"70",X"2C",X"71",X"CD",X"F0",X"0E",X"00",
		X"2E",X"BA",X"35",X"E1",X"E1",X"E9",X"36",X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2E",X"64",X"7B",X"FE",X"10",X"DA",X"FA",X"0E",X"2E",X"69",X"36",X"FF",X"C9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"E2",X"43",X"56",X"2C",X"5E",X"01",X"02",
		X"02",X"CD",X"56",X"0F",X"C8",X"00",X"00",X"21",X"9E",X"43",X"7E",X"D6",X"0A",X"47",X"2C",X"4E",
		X"21",X"70",X"4B",X"7E",X"2C",X"2C",X"E6",X"08",X"C4",X"38",X"0F",X"2C",X"2C",X"3E",X"90",X"BD",
		X"C2",X"23",X"0F",X"C9",X"FF",X"FF",X"FF",X"FF",X"2C",X"7E",X"2D",X"FE",X"D4",X"D8",X"FE",X"E7",
		X"D0",X"7E",X"B9",X"D0",X"B8",X"D8",X"CD",X"C4",X"0C",X"11",X"05",X"39",X"2B",X"2B",X"C3",X"AD",
		X"0E",X"AD",X"0E",X"FF",X"FF",X"FF",X"C5",X"D5",X"1A",X"FE",X"60",X"DA",X"63",X"0F",X"FE",X"D0",
		X"DA",X"72",X"0F",X"13",X"05",X"C2",X"58",X"0F",X"D1",X"C1",X"CD",X"17",X"02",X"0D",X"C2",X"56",
		X"0F",X"C9",X"D1",X"C1",X"C9",X"E2",X"56",X"2C",X"21",X"70",X"43",X"CD",X"C0",X"2F",X"21",X"74",
		X"43",X"CD",X"C0",X"2F",X"21",X"78",X"43",X"CD",X"C0",X"2F",X"21",X"7C",X"43",X"C3",X"C0",X"2F",
		X"7E",X"E6",X"1F",X"C8",X"35",X"7E",X"E6",X"FE",X"2C",X"2C",X"56",X"2C",X"5E",X"6F",X"26",X"2A",
		X"7E",X"2C",X"4E",X"6F",X"26",X"15",X"06",X"00",X"EB",X"09",X"EB",X"3E",X"A0",X"91",X"0F",X"4F",
		X"06",X"35",X"C5",X"01",X"08",X"00",X"C3",X"BC",X"0F",X"C3",X"AD",X"0E",X"7A",X"FE",X"43",X"C2",
		X"E9",X"0F",X"7B",X"FE",X"40",X"DA",X"E9",X"0F",X"D6",X"20",X"5F",X"2C",X"2C",X"41",X"FE",X"40",
		X"DA",X"E9",X"0F",X"D6",X"20",X"5F",X"2C",X"2C",X"78",X"81",X"47",X"7B",X"FE",X"40",X"DA",X"E9",
		X"0F",X"D6",X"20",X"5F",X"2C",X"2C",X"78",X"81",X"47",X"E3",X"7D",X"80",X"6F",X"E3",X"01",X"DF",
		X"FF",X"EB",X"C9",X"00",X"C3",X"40",X"35",X"68",X"3E",X"05",X"32",X"96",X"43",X"C3",X"A4",X"0E",
		X"05",X"1A",X"1A",X"1B",X"1C",X"1C",X"1D",X"1E",X"1E",X"1F",X"10",X"10",X"11",X"12",X"12",X"13",
		X"14",X"15",X"16",X"16",X"17",X"17",X"17",X"17",X"16",X"0F",X"0F",X"12",X"12",X"11",X"11",X"11",
		X"11",X"00",X"FF",X"FF",X"05",X"1D",X"1E",X"1F",X"10",X"10",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",
		X"19",X"18",X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"10",X"10",X"11",X"12",X"12",X"13",
		X"0F",X"0F",X"15",X"16",X"16",X"16",X"17",X"17",X"17",X"17",X"00",X"FF",X"05",X"1C",X"1C",X"1C",
		X"1D",X"1D",X"1E",X"1E",X"1E",X"1E",X"1F",X"1F",X"10",X"10",X"10",X"10",X"11",X"12",X"12",X"13",
		X"0F",X"0F",X"0F",X"14",X"15",X"15",X"15",X"16",X"16",X"16",X"16",X"17",X"17",X"17",X"17",X"17",
		X"17",X"00",X"FF",X"FF",X"05",X"1C",X"1C",X"1C",X"1C",X"1D",X"1E",X"1E",X"1F",X"10",X"10",X"10",
		X"10",X"10",X"11",X"12",X"12",X"13",X"14",X"14",X"14",X"14",X"15",X"16",X"16",X"17",X"18",X"18",
		X"18",X"18",X"19",X"1A",X"1B",X"1C",X"1C",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"10",X"11",
		X"12",X"13",X"14",X"14",X"0F",X"06",X"00",X"FF",X"05",X"1C",X"1C",X"1D",X"1E",X"1E",X"1F",X"10",
		X"10",X"11",X"12",X"13",X"14",X"14",X"14",X"14",X"04",X"02",X"02",X"02",X"02",X"03",X"1C",X"1C",
		X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"11",X"12",X"12",X"13",X"14",X"14",X"06",X"00",X"FF",
		X"05",X"1F",X"1F",X"1E",X"1E",X"1E",X"1D",X"1C",X"1C",X"1C",X"1C",X"1B",X"1A",X"19",X"18",X"18",
		X"17",X"16",X"15",X"14",X"0F",X"06",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"09",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"FF",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"05",X"1C",X"1B",X"1A",X"1A",X"19",X"18",X"18",X"18",X"17",X"16",X"16",X"15",
		X"0F",X"0F",X"0F",X"13",X"13",X"12",X"12",X"12",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"00",X"FF",X"FF",X"05",X"1C",X"1C",X"1B",X"1A",X"1A",X"19",X"18",X"19",X"1A",X"1B",X"1C",
		X"1D",X"1E",X"1F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"17",X"16",X"16",X"15",
		X"14",X"14",X"14",X"13",X"13",X"12",X"12",X"12",X"12",X"11",X"11",X"11",X"00",X"FF",X"05",X"1D",
		X"1D",X"1D",X"1D",X"1C",X"1C",X"1B",X"1A",X"19",X"18",X"18",X"18",X"18",X"17",X"16",X"15",X"14",
		X"14",X"13",X"13",X"13",X"13",X"0F",X"04",X"02",X"02",X"02",X"02",X"03",X"1C",X"1B",X"1B",X"1B",
		X"1B",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"10",X"10",X"11",X"12",X"13",X"14",X"14",X"15",
		X"15",X"15",X"15",X"06",X"00",X"FF",X"05",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"1A",
		X"1A",X"19",X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"15",X"14",X"14",X"14",X"13",X"13",X"12",
		X"12",X"11",X"10",X"1F",X"1E",X"1E",X"1D",X"1D",X"1C",X"1C",X"1C",X"1B",X"1B",X"1A",X"1A",X"19",
		X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"15",X"14",X"14",X"0F",X"0F",X"0F",X"0F",X"06",X"00",
		X"FF",X"FF",X"05",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1A",X"1A",X"1A",X"19",X"18",X"18",
		X"18",X"18",X"18",X"17",X"16",X"16",X"16",X"15",X"0F",X"0F",X"0F",X"14",X"13",X"13",X"12",X"12",
		X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"05",X"1C",X"1C",X"1C",X"1C",X"1B",
		X"1B",X"1A",X"1A",X"19",X"18",X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"14",X"14",X"0F",X"0F",
		X"0F",X"0F",X"04",X"01",X"01",X"01",X"01",X"01",X"03",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"11",
		X"12",X"13",X"14",X"14",X"06",X"00",X"FF",X"FF",X"05",X"19",X"19",X"1A",X"1A",X"1A",X"1B",X"1B",
		X"1C",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"10",X"11",X"12",X"13",X"14",X"0F",X"06",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0A",X"09",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"00",X"FF",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"05",X"1C",X"1D",
		X"1E",X"1E",X"1F",X"10",X"10",X"10",X"10",X"11",X"12",X"12",X"13",X"0F",X"0F",X"0F",X"14",X"15",
		X"16",X"16",X"16",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"00",X"FF",X"FF",
		X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"16",X"15",X"14",X"14",X"14",X"13",X"12",
		X"12",X"11",X"10",X"10",X"10",X"1F",X"1E",X"1D",X"1C",X"1C",X"1C",X"1B",X"1A",X"19",X"18",X"17",
		X"16",X"0F",X"0F",X"13",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"10",X"10",X"1F",X"1F",
		X"00",X"FF",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"16",X"16",X"16",X"15",X"14",X"14",X"13",
		X"12",X"12",X"11",X"10",X"10",X"1F",X"1E",X"1E",X"1D",X"1C",X"1C",X"1B",X"1A",X"1A",X"19",X"18",
		X"18",X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"0F",X"0F",X"0F",X"13",X"12",X"12",X"11",X"11",
		X"11",X"11",X"10",X"10",X"10",X"10",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"FF",X"FF",X"FF",
		X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"16",X"16",X"17",X"18",X"18",X"18",X"19",X"1A",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"10",X"11",X"12",X"12",X"13",X"0F",X"0F",X"0F",X"0F",X"15",
		X"16",X"16",X"17",X"18",X"18",X"18",X"19",X"19",X"19",X"19",X"19",X"19",X"00",X"FF",X"15",X"15",
		X"16",X"16",X"16",X"16",X"17",X"17",X"18",X"18",X"18",X"18",X"19",X"1A",X"1B",X"1B",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"13",X"13",X"12",X"12",X"11",X"10",X"10",X"10",X"10",X"1F",X"1E",X"1D",X"0F",
		X"0F",X"0F",X"0F",X"15",X"16",X"16",X"17",X"17",X"18",X"18",X"18",X"19",X"19",X"1A",X"19",X"18",
		X"17",X"17",X"00",X"FF",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"17",X"18",
		X"19",X"1A",X"1B",X"05",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"09",X"09",X"09",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"00",X"17",X"17",X"00",X"FF",X"FF",X"17",X"17",X"17",X"17",X"16",X"16",X"16",X"15",
		X"14",X"13",X"12",X"11",X"10",X"1F",X"1E",X"1D",X"1C",X"1B",X"19",X"17",X"15",X"13",X"13",X"14",
		X"14",X"14",X"14",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"1C",X"1D",X"1E",X"1F",X"1F",
		X"00",X"FF",X"15",X"15",X"15",X"15",X"15",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1D",X"1D",
		X"1D",X"1E",X"1F",X"10",X"11",X"13",X"14",X"14",X"15",X"15",X"15",X"15",X"0F",X"0F",X"04",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"1B",X"1B",X"19",X"19",X"19",X"19",X"00",X"FF",
		X"17",X"17",X"17",X"17",X"17",X"16",X"15",X"14",X"14",X"14",X"13",X"12",X"11",X"10",X"10",X"1F",
		X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"18",X"17",X"17",X"16",X"16",X"15",X"15",X"0F",X"0F",
		X"0F",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"FF",X"FF",
		X"30",X"40",X"31",X"41",X"00",X"42",X"33",X"43",X"00",X"44",X"35",X"45",X"00",X"46",X"37",X"47",
		X"38",X"48",X"00",X"49",X"3A",X"4A",X"00",X"4B",X"3C",X"4C",X"00",X"4D",X"3E",X"4E",X"3F",X"4F",
		X"C0",X"C8",X"C1",X"C9",X"C2",X"CA",X"C3",X"CB",X"C4",X"CC",X"C5",X"CD",X"C6",X"00",X"C7",X"CF",
		X"60",X"76",X"61",X"00",X"68",X"93",X"69",X"00",X"80",X"94",X"81",X"71",X"88",X"96",X"89",X"91",
		X"60",X"70",X"61",X"00",X"68",X"70",X"69",X"00",X"80",X"70",X"81",X"00",X"88",X"79",X"89",X"99",
		X"A0",X"00",X"A1",X"00",X"A2",X"00",X"A3",X"00",X"A4",X"00",X"A5",X"00",X"A6",X"00",X"A7",X"00",
		X"C3",X"F1",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"60",X"70",X"61",X"00",X"68",X"78",X"69",X"00",X"80",X"90",X"81",X"00",X"88",X"98",X"89",X"99",
		X"62",X"72",X"63",X"73",X"6A",X"7A",X"6B",X"7B",X"82",X"92",X"83",X"00",X"8A",X"9A",X"8B",X"9B",
		X"64",X"74",X"65",X"75",X"6C",X"7C",X"6D",X"7D",X"84",X"00",X"85",X"95",X"8C",X"9C",X"8D",X"9D",
		X"66",X"00",X"67",X"77",X"6E",X"00",X"6F",X"7F",X"86",X"00",X"87",X"97",X"8E",X"9E",X"8F",X"9F",
		X"B0",X"00",X"B1",X"00",X"A0",X"00",X"A1",X"00",X"A8",X"B8",X"A9",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"A2",X"00",X"A3",X"00",X"FF",X"FF",X"FF",X"FF",X"AA",X"BA",X"AB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"A4",X"00",X"A5",X"00",X"AC",X"BC",X"AD",X"BD",X"B2",X"B4",X"B3",X"B5",
		X"FF",X"FF",X"FF",X"FF",X"A6",X"00",X"A7",X"00",X"FF",X"FF",X"FF",X"FF",X"AE",X"BE",X"AF",X"BF",
		X"D6",X"DD",X"E9",X"EC",X"E3",X"F3",X"E1",X"F1",X"E4",X"F4",X"EB",X"EE",X"D8",X"EF",X"DF",X"DD",
		X"E0",X"F0",X"E1",X"DA",X"E9",X"DA",X"EA",X"F1",X"E2",X"F2",X"DE",X"DC",X"00",X"00",X"D6",X"FF",
		X"E9",X"EC",X"EA",X"ED",X"EB",X"EE",X"D8",X"EF",X"00",X"00",X"DF",X"DD",X"E0",X"F0",X"E1",X"F1",
		X"E2",X"F2",X"DE",X"DC",X"00",X"00",X"D6",X"D9",X"D7",X"DA",X"D8",X"DB",X"00",X"00",X"D0",X"D3",
		X"D1",X"D4",X"D2",X"D5",X"DF",X"FF",X"FE",X"FC",X"DE",X"FE",X"DC",X"B6",X"FF",X"CE",X"7E",X"FF",
		X"00",X"DD",X"DF",X"FF",X"00",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D6",X"D9",X"FF",X"E9",X"F9",X"EC",X"EB",X"FB",X"EE",X"D8",X"DB",X"EF",X"00",X"FE",X"DD",X"00",
		X"E0",X"F0",X"FF",X"E2",X"F2",X"00",X"DC",X"00",X"00",X"00",X"FF",X"00",X"D0",X"D3",X"DF",X"D2",
		X"D5",X"00",X"00",X"DC",X"00",X"00",X"00",X"00",X"D6",X"D9",X"00",X"D8",X"DB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DF",X"DD",X"00",X"DE",X"DC",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"D0",X"F6",X"DE",X"D1",X"F7",X"F5",X"D2",X"F8",X"DF",X"00",X"D0",X"D3",X"FF",X"D1",X"D4",X"00",
		X"D2",X"D5",X"00",X"D6",X"D9",X"DF",X"D7",X"DA",X"00",X"D8",X"DB",X"00",X"DF",X"DD",X"00",X"DE",
		X"FC",X"00",X"DD",X"DC",X"00",X"00",X"DE",X"00",X"DC",X"FE",X"00",X"00",X"DF",X"00",X"54",X"55",
		X"56",X"57",X"58",X"00",X"59",X"5A",X"53",X"5C",X"5D",X"00",X"54",X"59",X"5B",X"57",X"5C",X"00",
		X"55",X"5A",X"53",X"58",X"5D",X"00",X"00",X"54",X"00",X"53",X"57",X"00",X"00",X"56",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"14",X"18",X"1C",X"00",X"04",X"08",X"0C",X"20",X"24",X"28",X"2C",X"30",X"34",X"38",X"3C",
		X"80",X"84",X"88",X"8C",X"90",X"94",X"98",X"9C",X"A0",X"A4",X"A8",X"AC",X"B0",X"B4",X"B8",X"BC",
		X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"40",X"44",X"48",X"4C",X"50",X"54",X"58",X"5C",
		X"C0",X"C4",X"C8",X"FF",X"FF",X"D4",X"FF",X"DC",X"FF",X"E4",X"E8",X"EC",X"FF",X"F4",X"FF",X"FC",
		X"00",X"02",X"6F",X"00",X"02",X"7E",X"7F",X"00",X"13",X"00",X"05",X"7C",X"7D",X"00",X"13",X"39",
		X"3A",X"2C",X"2C",X"2C",X"2C",X"2C",X"3B",X"3C",X"00",X"11",X"00",X"02",X"3D",X"36",X"37",X"38",
		X"3D",X"00",X"13",X"00",X"02",X"60",X"33",X"34",X"35",X"60",X"00",X"13",X"00",X"04",X"32",X"00",
		X"15",X"00",X"03",X"DC",X"DD",X"A9",X"AA",X"DE",X"F4",X"00",X"11",X"FB",X"9C",X"FE",X"00",X"02",
		X"A7",X"A8",X"00",X"13",X"00",X"1A",X"00",X"1A",X"AF",X"21",X"86",X"19",X"06",X"06",X"CD",X"B0",
		X"16",X"21",X"F8",X"1A",X"06",X"08",X"CD",X"B0",X"16",X"21",X"95",X"0B",X"06",X"09",X"CD",X"B0",
		X"16",X"C6",X"6B",X"4F",X"11",X"F1",X"37",X"19",X"7E",X"81",X"77",X"C9",X"32",X"23",X"41",X"C9",
		X"86",X"23",X"05",X"C2",X"B0",X"16",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"02",X"08",X"02",X"08",X"04",X"0C",X"04",X"0C",X"04",X"28",X"04",X"28",X"02",X"2C",
		X"01",X"30",X"01",X"30",X"01",X"30",X"01",X"30",X"02",X"2C",X"01",X"30",X"01",X"30",X"01",X"10",
		X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",
		X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",
		X"FF",X"FF",X"01",X"00",X"FF",X"00",X"00",X"FF",X"00",X"01",X"00",X"FF",X"00",X"01",X"02",X"00",
		X"04",X"02",X"02",X"02",X"FE",X"02",X"FC",X"02",X"FE",X"00",X"FC",X"FE",X"04",X"FE",X"00",X"01",
		X"02",X"00",X"02",X"01",X"02",X"02",X"01",X"02",X"00",X"02",X"FF",X"02",X"FE",X"02",X"FE",X"01",
		X"FE",X"00",X"FE",X"FF",X"FE",X"FE",X"FF",X"FE",X"00",X"FE",X"01",X"FE",X"02",X"FE",X"02",X"FF",
		X"47",X"3A",X"00",X"78",X"E6",X"10",X"C8",X"EB",X"7A",X"FE",X"18",X"C0",X"7B",X"FE",X"95",X"36",
		X"22",X"C8",X"FE",X"9C",X"36",X"0E",X"C8",X"FE",X"B5",X"36",X"24",X"C8",X"70",X"C9",X"FE",X"FF",
		X"3A",X"00",X"78",X"E6",X"10",X"3A",X"8F",X"43",X"C8",X"0F",X"E6",X"0F",X"C9",X"FF",X"FF",X"FF",
		X"00",X"00",X"FE",X"DC",X"00",X"00",X"00",X"D6",X"D9",X"E5",X"DD",X"00",X"DD",X"E9",X"F9",X"E7",
		X"EC",X"DE",X"FE",X"E3",X"FA",X"ED",X"F3",X"DF",X"00",X"E4",X"EA",X"F9",X"F4",X"FF",X"DD",X"EB",
		X"FB",X"E8",X"EE",X"00",X"00",X"D8",X"DB",X"E6",X"EF",X"DC",X"00",X"00",X"FD",X"DE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"DD",X"00",X"00",X"00",X"00",X"E0",X"E7",
		X"F0",X"CE",X"00",X"FF",X"E1",X"F9",X"DA",X"00",X"00",X"00",X"EA",X"FA",X"F1",X"DC",X"00",X"DD",
		X"E2",X"E8",X"F2",X"DF",X"00",X"00",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D6",X"D9",X"FF",X"00",X"00",X"00",X"E9",X"F9",
		X"EC",X"00",X"00",X"00",X"EB",X"FB",X"EE",X"00",X"00",X"00",X"D8",X"DB",X"EF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"20",X"FF",X"FF",X"FF",X"FF",X"10",X"15",X"0E",X"0B",X"14",X"05",X"21",X"00",X"00",X"00",
		X"12",X"05",X"0B",X"0F",X"12",X"04",X"00",X"00",X"00",X"10",X"15",X"0E",X"0B",X"14",X"05",X"22",
		X"43",X"21",X"FF",X"FF",X"FF",X"FF",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"00",
		X"43",X"22",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"2A",X"20",X"00",X"00",X"00",X"00",X"00",
		X"07",X"05",X"0C",X"04",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"2A",X"20",X"00",X"00",X"00",
		X"43",X"25",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"02",X"09",X"14",X"14",X"05",X"00",X"07",
		X"05",X"0C",X"04",X"00",X"05",X"09",X"0E",X"17",X"05",X"12",X"06",X"05",X"0E",X"00",X"00",X"00",
		X"43",X"27",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"1F",X"00",X"21",X"13",X"10",X"09",X"05",
		X"0C",X"05",X"12",X"00",X"00",X"21",X"0D",X"15",X"05",X"0E",X"1A",X"05",X"00",X"00",X"1F",X"00",
		X"43",X"29",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"1F",X"00",X"22",X"13",X"10",X"09",X"05",
		X"0C",X"05",X"12",X"00",X"00",X"22",X"0D",X"15",X"05",X"0E",X"1A",X"05",X"0E",X"00",X"1F",X"00",
		X"43",X"2D",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"10",X"15",X"0E",X"0B",X"14",X"05",X"14",
		X"01",X"02",X"0C",X"0C",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"30",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"23",X"20",X"00",X"28",X"20",X"00",X"21",X"25",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"20",X"00",X"21",X"20",X"20",X"2B",X"24",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"37",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"2B",X"29",X"26",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"3A",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"20",X"20",X"2B",X"26",X"20",X"20",X"00",X"25",X"20",X"20",X"2B",X"24",X"20",X"20",X"20",
		X"43",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",
		X"00",X"00",X"21",X"29",X"28",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"3D",X"21",X"00",X"21",X"00",X"16",X"0E",X"09",X"16",X"05",X"12",X"13",X"01",X"0C",X"00",
		X"16",X"09",X"04",X"05",X"0F",X"00",X"13",X"10",X"09",X"05",X"0C",X"00",X"07",X"0D",X"02",X"08",
		X"43",X"3E",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"28",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"2C",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"15",X"12",X"00",
		X"13",X"10",X"09",X"05",X"0C",X"05",X"12",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"28",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"10",
		X"09",X"05",X"0C",X"05",X"0E",X"04",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"00",X"00",X"00",X"00",X"00",X"65",X"65",X"00",
		X"00",X"00",X"00",X"00",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"00",X"00",X"65",
		X"00",X"00",X"00",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"00",X"00",X"65",X"00",X"00",X"00",X"65",X"65",X"65",X"65",X"00",X"00",X"00",X"65",
		X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"65",X"65",
		X"65",X"65",X"65",X"65",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"65",X"00",X"00",X"00",X"00",X"00",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",
		X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"00",
		X"00",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"43",X"0A",X"20",X"03",X"42",X"8A",X"35",X"03",X"42",X"0A",X"4A",X"03",X"41",X"8A",X"5F",X"01",
		X"41",X"4A",X"66",X"03",X"40",X"CA",X"7B",X"03",X"40",X"4A",X"90",X"04",X"FF",X"FF",X"FF",X"FF",
		X"21",X"E8",X"4B",X"35",X"CA",X"F8",X"1A",X"7E",X"2C",X"6E",X"26",X"1A",X"56",X"2C",X"5E",X"2C",
		X"46",X"2C",X"4E",X"FE",X"20",X"C2",X"B8",X"0B",X"21",X"1E",X"08",X"19",X"EB",X"26",X"1A",X"68",
		X"06",X"07",X"C3",X"D6",X"0A",X"6C",X"00",X"6C",X"34",X"2C",X"7E",X"FE",X"C8",X"CA",X"00",X"1C",
		X"C6",X"04",X"77",X"2D",X"36",X"40",X"C3",X"80",X"03",X"C3",X"E4",X"01",X"CD",X"00",X"04",X"21",
		X"E8",X"4B",X"36",X"40",X"2C",X"36",X"B0",X"21",X"A4",X"43",X"7E",X"FE",X"03",X"C8",X"36",X"02",
		X"2E",X"BA",X"36",X"01",X"C9",X"FF",X"00",X"CD",X"BC",X"06",X"C3",X"2E",X"06",X"06",X"CF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CA",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"3A",X"00",X"60",X"3D",X"2C",
		X"00",X"33",X"36",X"2C",X"30",X"34",X"37",X"2C",X"00",X"35",X"38",X"2C",X"00",X"60",X"3D",X"2C",
		X"00",X"00",X"00",X"3B",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"32",X"00",X"36",X"39",X"36",X"39",X"00",X"32",X"34",X"00",X"3B",X"3D",X"3B",X"3D",X"00",X"34",
		X"43",X"2C",X"32",X"32",X"32",X"32",X"00",X"00",X"00",X"00",X"00",X"0E",X"05",X"15",X"05",X"12",
		X"00",X"01",X"0E",X"07",X"12",X"09",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"2C",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"10",X"09",X"05",
		X"0C",X"05",X"12",X"00",X"21",X"00",X"0F",X"04",X"05",X"12",X"00",X"22",X"00",X"00",X"00",X"00",
		X"43",X"29",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"03",X"08",X"14",X"15",X"0E",X"07",X"00",
		X"00",X"0E",X"05",X"15",X"05",X"12",X"00",X"01",X"15",X"06",X"14",X"12",X"01",X"07",X"00",X"00",
		X"43",X"2C",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"1A",X"09",X"05",X"0C",X"01",X"0E",X"06",X"0C",
		X"15",X"07",X"00",X"1A",X"15",X"12",X"00",X"00",X"02",X"01",X"13",X"09",X"13",X"00",X"00",X"00",
		X"CD",X"46",X"01",X"CD",X"27",X"1B",X"CD",X"E4",X"01",X"11",X"5D",X"26",X"19",X"11",X"20",X"00",
		X"3E",X"F4",X"06",X"1A",X"86",X"19",X"05",X"C2",X"14",X"1C",X"1E",X"24",X"19",X"86",X"77",X"C9",
		X"3F",X"04",X"87",X"3F",X"10",X"8F",X"3F",X"04",X"00",X"04",X"86",X"00",X"10",X"8E",X"00",X"04",
		X"3F",X"04",X"85",X"3F",X"10",X"8D",X"3F",X"04",X"00",X"04",X"84",X"00",X"10",X"8C",X"00",X"04",
		X"3F",X"05",X"87",X"3F",X"0E",X"8F",X"3F",X"05",X"00",X"05",X"86",X"00",X"0E",X"8E",X"00",X"05",
		X"3F",X"05",X"85",X"3F",X"0E",X"8D",X"3F",X"05",X"00",X"05",X"84",X"00",X"0E",X"8C",X"00",X"05",
		X"3F",X"06",X"87",X"3F",X"0C",X"8F",X"3F",X"06",X"00",X"06",X"86",X"00",X"0C",X"8E",X"00",X"06",
		X"83",X"3F",X"05",X"85",X"3F",X"0C",X"8D",X"3F",X"05",X"8B",X"82",X"00",X"05",X"84",X"00",X"0C",
		X"8C",X"00",X"05",X"8A",X"3F",X"01",X"83",X"3F",X"05",X"87",X"3F",X"0A",X"8F",X"3F",X"05",X"8B",
		X"3F",X"01",X"00",X"01",X"82",X"00",X"05",X"86",X"00",X"0A",X"8E",X"00",X"05",X"8A",X"00",X"01",
		X"3F",X"02",X"83",X"3F",X"04",X"85",X"3F",X"0A",X"8D",X"3F",X"04",X"8B",X"3F",X"02",X"00",X"02",
		X"82",X"00",X"04",X"84",X"00",X"0A",X"8C",X"00",X"04",X"8A",X"00",X"02",X"3F",X"03",X"83",X"3F",
		X"04",X"87",X"3F",X"08",X"8F",X"3F",X"04",X"8B",X"3F",X"03",X"00",X"03",X"82",X"00",X"04",X"86",
		X"00",X"08",X"8E",X"00",X"04",X"8A",X"00",X"03",X"3F",X"04",X"83",X"3F",X"03",X"85",X"3F",X"08",
		X"8D",X"3F",X"03",X"8B",X"3F",X"04",X"00",X"04",X"82",X"00",X"03",X"84",X"00",X"08",X"8C",X"00",
		X"03",X"8A",X"00",X"04",X"3F",X"05",X"83",X"3F",X"03",X"87",X"3F",X"06",X"8F",X"3F",X"03",X"8B",
		X"3F",X"05",X"00",X"05",X"82",X"00",X"03",X"86",X"00",X"06",X"8E",X"00",X"03",X"8A",X"00",X"05",
		X"3F",X"06",X"83",X"3F",X"02",X"85",X"3F",X"06",X"8D",X"3F",X"02",X"8B",X"3F",X"06",X"80",X"00",
		X"05",X"82",X"00",X"02",X"84",X"00",X"06",X"8C",X"00",X"02",X"8A",X"00",X"05",X"88",X"78",X"81",
		X"3F",X"05",X"83",X"3F",X"02",X"87",X"3F",X"04",X"8F",X"3F",X"02",X"8B",X"3F",X"05",X"89",X"78",
		X"00",X"01",X"79",X"80",X"00",X"04",X"82",X"00",X"02",X"86",X"00",X"04",X"8E",X"00",X"02",X"8A",
		X"00",X"04",X"88",X"79",X"00",X"01",X"00",X"02",X"7A",X"81",X"3F",X"04",X"83",X"3F",X"01",X"85",
		X"3F",X"04",X"8D",X"3F",X"01",X"8B",X"3F",X"04",X"89",X"7A",X"00",X"02",X"00",X"03",X"7B",X"80",
		X"00",X"03",X"82",X"00",X"01",X"84",X"00",X"04",X"8C",X"00",X"01",X"8A",X"00",X"03",X"88",X"7B",
		X"00",X"03",X"00",X"04",X"78",X"81",X"3F",X"03",X"83",X"3F",X"01",X"87",X"3F",X"02",X"8F",X"3F",
		X"01",X"8B",X"3F",X"03",X"89",X"78",X"00",X"04",X"00",X"05",X"79",X"80",X"00",X"02",X"82",X"00",
		X"01",X"86",X"00",X"02",X"8E",X"00",X"01",X"8A",X"00",X"02",X"88",X"79",X"00",X"05",X"00",X"06",
		X"7A",X"81",X"3F",X"02",X"83",X"85",X"3F",X"02",X"8D",X"8B",X"3F",X"02",X"89",X"7A",X"00",X"06",
		X"00",X"07",X"7B",X"80",X"00",X"01",X"82",X"84",X"00",X"02",X"8C",X"8A",X"00",X"01",X"88",X"7B",
		X"00",X"04",X"00",X"01",X"00",X"01",X"00",X"01",X"6E",X"6C",X"6B",X"00",X"05",X"78",X"81",X"3F",
		X"01",X"83",X"87",X"8F",X"8B",X"3F",X"01",X"89",X"78",X"00",X"05",X"5F",X"65",X"67",X"6E",X"6C",
		X"6B",X"00",X"06",X"79",X"80",X"82",X"86",X"8E",X"8A",X"88",X"79",X"00",X"06",X"5F",X"65",X"67",
		X"6E",X"6C",X"6B",X"00",X"07",X"7A",X"81",X"83",X"8B",X"89",X"7A",X"00",X"07",X"5F",X"65",X"67",
		X"6D",X"6C",X"6B",X"00",X"08",X"7B",X"7E",X"7F",X"7B",X"00",X"08",X"5E",X"65",X"67",X"6D",X"6C",
		X"6A",X"00",X"09",X"7C",X"7D",X"00",X"09",X"5E",X"65",X"67",X"6D",X"6C",X"6A",X"00",X"02",X"42",
		X"43",X"00",X"0B",X"52",X"52",X"52",X"52",X"00",X"02",X"64",X"66",X"6D",X"69",X"00",X"01",X"42",
		X"43",X"40",X"41",X"00",X"0B",X"51",X"51",X"51",X"51",X"4E",X"4F",X"63",X"63",X"00",X"01",X"69",
		X"00",X"01",X"40",X"41",X"00",X"0F",X"4E",X"4F",X"4C",X"4D",X"60",X"60",X"00",X"01",X"68",X"00",
		X"03",X"50",X"50",X"50",X"50",X"50",X"50",X"00",X"09",X"4C",X"4D",X"00",X"04",X"00",X"01",X"63",
		X"00",X"18",X"00",X"18",X"00",X"01",X"00",X"01",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",
		X"26",X"25",X"24",X"23",X"22",X"21",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"26",X"25",
		X"24",X"23",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"0C",X"19",X"19",X"19",X"07",
		X"04",X"00",X"09",X"00",X"0C",X"19",X"19",X"15",X"16",X"17",X"19",X"00",X"08",X"00",X"0C",X"19",
		X"07",X"05",X"06",X"19",X"19",X"19",X"00",X"07",X"00",X"0C",X"19",X"03",X"17",X"19",X"19",X"19",
		X"19",X"19",X"00",X"06",X"00",X"0D",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"00",X"05",
		X"00",X"0D",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"00",X"04",X"00",X"0E",X"19",
		X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"00",X"03",X"00",X"0F",X"19",X"19",X"19",X"19",
		X"19",X"07",X"04",X"19",X"19",X"00",X"02",X"00",X"10",X"19",X"19",X"19",X"15",X"16",X"17",X"19",
		X"19",X"19",X"00",X"02",X"00",X"04",X"07",X"04",X"00",X"0B",X"19",X"07",X"05",X"06",X"19",X"00",
		X"01",X"19",X"19",X"00",X"01",X"00",X"03",X"15",X"16",X"17",X"00",X"0C",X"03",X"17",X"19",X"19",
		X"19",X"19",X"19",X"00",X"01",X"00",X"02",X"07",X"05",X"06",X"00",X"0E",X"19",X"19",X"19",X"19",
		X"19",X"19",X"00",X"01",X"00",X"02",X"03",X"17",X"00",X"10",X"19",X"19",X"19",X"19",X"19",X"00",
		X"01",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"10",X"4A",X"25",X"38",X"10",X"4A",X"A7",
		X"48",X"10",X"48",X"E9",X"58",X"10",X"49",X"CB",X"68",X"10",X"4A",X"4D",X"78",X"10",X"49",X"4F",
		X"00",X"00",X"49",X"60",X"10",X"00",X"4A",X"02",X"20",X"00",X"49",X"04",X"30",X"00",X"49",X"A6",
		X"40",X"00",X"48",X"A8",X"50",X"00",X"4A",X"4A",X"60",X"00",X"49",X"6C",X"70",X"00",X"48",X"6E",
		X"80",X"00",X"4A",X"F0",X"90",X"00",X"49",X"D2",X"A0",X"00",X"48",X"F4",X"B0",X"00",X"4A",X"76",
		X"58",X"20",X"48",X"EB",X"70",X"20",X"4A",X"2E",X"80",X"20",X"49",X"50",X"88",X"20",X"4A",X"91",
		X"C0",X"20",X"49",X"78",X"D0",X"20",X"48",X"BA",X"48",X"40",X"49",X"C9",X"C8",X"40",X"4A",X"19",
		X"00",X"10",X"49",X"A0",X"10",X"10",X"49",X"22",X"20",X"10",X"4A",X"04",X"30",X"10",X"4A",X"66",
		X"40",X"10",X"48",X"E8",X"50",X"10",X"49",X"CA",X"60",X"10",X"4A",X"4C",X"70",X"10",X"49",X"4E",
		X"80",X"10",X"48",X"70",X"90",X"10",X"49",X"92",X"A0",X"10",X"4A",X"B4",X"B0",X"10",X"49",X"36",
		X"60",X"10",X"48",X"CC",X"68",X"10",X"4A",X"ED",X"78",X"10",X"4A",X"0F",X"90",X"10",X"48",X"D2",
		X"30",X"30",X"49",X"66",X"98",X"30",X"4A",X"33",X"B8",X"30",X"49",X"D7",X"C0",X"30",X"4A",X"F8",
		X"7E",X"E6",X"02",X"C8",X"54",X"7D",X"C6",X"20",X"5F",X"1A",X"C6",X"08",X"47",X"13",X"1A",X"4F",
		X"0A",X"FE",X"40",X"D8",X"FE",X"6F",X"D0",X"78",X"D6",X"08",X"57",X"59",X"2B",X"2B",X"7E",X"E6",
		X"F7",X"77",X"0A",X"FE",X"50",X"DA",X"40",X"20",X"3E",X"00",X"02",X"06",X"88",X"21",X"90",X"4B",
		X"0E",X"0F",X"CD",X"68",X"20",X"70",X"2C",X"2C",X"72",X"2C",X"73",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"E6",X"03",X"FE",X"02",X"C2",X"58",X"20",X"21",X"A0",X"4B",X"0E",X"FF",X"CD",X"68",X"20",X"36",
		X"80",X"2C",X"2C",X"70",X"2C",X"73",X"C9",X"FF",X"3E",X"00",X"02",X"06",X"6B",X"C3",X"2D",X"20",
		X"CD",X"76",X"08",X"C3",X"BC",X"33",X"FF",X"FF",X"7E",X"A1",X"C8",X"2C",X"2C",X"2C",X"2C",X"7E",
		X"A1",X"C8",X"2C",X"2C",X"2C",X"2C",X"7E",X"A1",X"C8",X"2C",X"2C",X"2C",X"2C",X"C9",X"FF",X"FF",
		X"3A",X"92",X"43",X"0F",X"0F",X"DA",X"9C",X"20",X"21",X"90",X"4B",X"E5",X"CD",X"B0",X"20",X"E1",
		X"7D",X"C6",X"04",X"6F",X"FE",X"A0",X"C2",X"89",X"20",X"C9",X"FF",X"FF",X"21",X"A0",X"4B",X"E5",
		X"CD",X"D4",X"20",X"E1",X"7D",X"C6",X"04",X"6F",X"FE",X"B0",X"C2",X"9F",X"20",X"C9",X"FF",X"FF",
		X"7E",X"E6",X"0F",X"C8",X"35",X"7E",X"2C",X"2C",X"56",X"2C",X"5E",X"6F",X"26",X"2A",X"6E",X"26",
		X"15",X"01",X"1E",X"00",X"EB",X"09",X"C3",X"26",X"21",X"21",X"C5",X"01",X"0C",X"00",X"C3",X"BC",
		X"0F",X"FF",X"FF",X"FF",X"7E",X"A7",X"C8",X"35",X"7E",X"2C",X"2C",X"56",X"2C",X"5E",X"E6",X"07",
		X"C6",X"F8",X"6F",X"26",X"20",X"6E",X"26",X"15",X"1B",X"1B",X"EB",X"01",X"DE",X"FF",X"C3",X"0C",
		X"21",X"C3",X"98",X"2A",X"FF",X"FF",X"FF",X"FF",X"56",X"EB",X"E5",X"DF",X"D9",X"D3",X"CD",X"FF",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"1A",X"77",X"13",X"23",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"23",
		X"1A",X"77",X"13",X"09",X"C9",X"D0",X"01",X"DE",X"FF",X"7C",X"FE",X"43",X"C2",X"00",X"21",X"7D",
		X"FE",X"40",X"DA",X"00",X"21",X"D6",X"20",X"6F",X"1C",X"1C",X"1C",X"FE",X"40",X"DA",X"0C",X"21",
		X"D6",X"20",X"6F",X"1C",X"1C",X"1C",X"C3",X"18",X"21",X"90",X"21",X"C3",X"A5",X"21",X"F0",X"F9",
		X"21",X"B8",X"43",X"7E",X"E6",X"04",X"C0",X"00",X"00",X"2E",X"92",X"7E",X"21",X"92",X"43",X"7E",
		X"FE",X"C0",X"D2",X"84",X"21",X"E6",X"04",X"47",X"7E",X"0F",X"0F",X"0F",X"4F",X"E6",X"18",X"C6",
		X"30",X"80",X"6F",X"26",X"22",X"56",X"23",X"5E",X"23",X"79",X"E6",X"07",X"86",X"6F",X"26",X"22",
		X"7E",X"12",X"C9",X"FF",X"0F",X"0F",X"0F",X"4F",X"7E",X"E6",X"04",X"C6",X"48",X"6F",X"26",X"22",
		X"56",X"23",X"5E",X"23",X"79",X"E6",X"07",X"86",X"6F",X"26",X"22",X"6E",X"EB",X"7E",X"23",X"A6",
		X"01",X"DF",X"FF",X"09",X"A6",X"23",X"A6",X"E6",X"F0",X"FE",X"40",X"C0",X"01",X"1F",X"00",X"09",
		X"EB",X"3E",X"08",X"32",X"62",X"43",X"E5",X"CD",X"C0",X"21",X"E1",X"C3",X"DC",X"07",X"22",X"CD",
		X"7D",X"FE",X"70",X"C0",X"21",X"C2",X"43",X"7E",X"FE",X"50",X"D0",X"2E",X"C8",X"7E",X"E6",X"08",
		X"C0",X"7E",X"F6",X"08",X"77",X"23",X"36",X"57",X"23",X"01",X"B8",X"1F",X"7B",X"FE",X"D8",X"CA",
		X"E5",X"21",X"01",X"C0",X"2F",X"70",X"23",X"71",X"2E",X"EA",X"36",X"00",X"2C",X"36",X"00",X"C9",
		X"0F",X"0F",X"C6",X"3A",X"5F",X"16",X"78",X"0F",X"D2",X"04",X"22",X"CD",X"40",X"0C",X"CD",X"78",
		X"0F",X"CD",X"80",X"20",X"21",X"94",X"43",X"34",X"7E",X"FE",X"60",X"D8",X"2E",X"A4",X"36",X"02",
		X"2E",X"60",X"36",X"FF",X"2E",X"B8",X"E5",X"E5",X"7E",X"E6",X"0E",X"FE",X"04",X"CA",X"F0",X"0C",
		X"E1",X"E1",X"34",X"FE",X"00",X"CA",X"74",X"22",X"2E",X"BA",X"36",X"10",X"C3",X"80",X"03",X"FF",
		X"4A",X"A9",X"50",X"00",X"48",X"6E",X"50",X"00",X"48",X"38",X"58",X"00",X"48",X"18",X"58",X"00",
		X"49",X"44",X"50",X"00",X"49",X"F2",X"50",X"00",X"4A",X"D8",X"60",X"00",X"4A",X"99",X"60",X"00",
		X"29",X"2A",X"2B",X"2A",X"2B",X"2A",X"29",X"28",X"61",X"62",X"61",X"60",X"61",X"62",X"61",X"60",
		X"6C",X"70",X"6C",X"68",X"6C",X"70",X"6C",X"68",X"40",X"42",X"41",X"43",X"44",X"46",X"45",X"47",
		X"48",X"4A",X"49",X"4B",X"2E",X"BB",X"36",X"08",X"2C",X"36",X"00",X"C3",X"80",X"03",X"03",X"15",
		X"21",X"B9",X"43",X"7E",X"0F",X"0F",X"0F",X"E6",X"1F",X"C6",X"20",X"5F",X"16",X"4B",X"3E",X"00",
		X"12",X"CD",X"17",X"02",X"7A",X"FE",X"47",X"C2",X"8E",X"22",X"CD",X"60",X"20",X"21",X"9B",X"43",
		X"7E",X"0F",X"D8",X"2E",X"B9",X"35",X"7E",X"32",X"00",X"58",X"C0",X"2D",X"34",X"C3",X"80",X"03",
		X"CD",X"C0",X"22",X"CD",X"E6",X"22",X"01",X"00",X"16",X"21",X"C2",X"43",X"C3",X"26",X"09",X"FF",
		X"21",X"9C",X"43",X"3A",X"A0",X"43",X"2F",X"E6",X"60",X"CA",X"D6",X"22",X"34",X"E6",X"40",X"C8",
		X"35",X"35",X"C9",X"FF",X"FF",X"FF",X"3A",X"9B",X"43",X"0F",X"00",X"D0",X"7E",X"35",X"A7",X"F0",
		X"34",X"34",X"C9",X"FF",X"FF",X"FF",X"21",X"9C",X"43",X"7E",X"A7",X"F2",X"0B",X"23",X"2F",X"3C",
		X"FE",X"7C",X"DA",X"F9",X"22",X"3E",X"7C",X"36",X"84",X"CD",X"26",X"23",X"21",X"C2",X"43",X"7E",
		X"91",X"77",X"FE",X"08",X"D0",X"36",X"08",X"C3",X"21",X"23",X"FF",X"FE",X"7C",X"DA",X"13",X"23",
		X"3E",X"7C",X"77",X"CD",X"26",X"23",X"21",X"C2",X"43",X"7E",X"81",X"77",X"FE",X"C1",X"D8",X"36",
		X"C0",X"2E",X"9C",X"36",X"00",X"C9",X"0F",X"0F",X"0F",X"4F",X"E6",X"07",X"C6",X"50",X"5F",X"16",
		X"23",X"1A",X"47",X"79",X"0F",X"0F",X"0F",X"E6",X"01",X"4F",X"3A",X"9B",X"43",X"E6",X"07",X"C6",
		X"58",X"5F",X"16",X"23",X"1A",X"A0",X"C8",X"0C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"FE",X"E0",X"D0",X"A9",X"D4",X"E0",X"F8",X"80",
		X"21",X"C0",X"1B",X"0E",X"02",X"CD",X"D0",X"01",X"CD",X"76",X"08",X"21",X"B9",X"43",X"3E",X"FF",
		X"77",X"32",X"00",X"58",X"2E",X"94",X"34",X"7E",X"FE",X"01",X"C2",X"81",X"23",X"2E",X"67",X"36",
		X"FF",X"FE",X"C0",X"C0",X"2E",X"B8",X"34",X"C3",X"80",X"03",X"36",X"00",X"2D",X"7E",X"FE",X"5E",
		X"CD",X"F8",X"24",X"CD",X"A0",X"24",X"CD",X"60",X"20",X"CD",X"78",X"0F",X"CD",X"F0",X"32",X"CD",
		X"A8",X"31",X"C3",X"76",X"32",X"FF",X"FF",X"FF",X"CD",X"76",X"08",X"21",X"B8",X"43",X"7E",X"E6",
		X"04",X"47",X"2E",X"92",X"7E",X"E6",X"03",X"B0",X"07",X"C6",X"C4",X"6F",X"26",X"23",X"7E",X"2C",
		X"6E",X"67",X"E9",X"FF",X"21",X"5C",X"24",X"30",X"24",X"3C",X"24",X"48",X"0A",X"9C",X"0A",X"BC",
		X"09",X"D4",X"37",X"D0",X"FF",X"FF",X"21",X"B8",X"43",X"7E",X"E6",X"0F",X"FE",X"01",X"CA",X"98",
		X"3A",X"FE",X"03",X"CA",X"98",X"3A",X"FE",X"05",X"CA",X"D0",X"3A",X"FE",X"07",X"CA",X"D0",X"3A",
		X"FE",X"09",X"D8",X"FE",X"0B",X"DA",X"02",X"3B",X"CD",X"02",X"3B",X"FF",X"98",X"3F",X"FF",X"FF",
		X"00",X"00",X"00",X"21",X"DC",X"4B",X"7E",X"D6",X"08",X"57",X"2C",X"5E",X"21",X"BA",X"43",X"36",
		X"10",X"2E",X"A4",X"36",X"02",X"2C",X"35",X"7E",X"C8",X"2D",X"36",X"06",X"FE",X"1E",X"D8",X"CA",
		X"80",X"03",X"FE",X"1F",X"CA",X"A0",X"03",X"D6",X"20",X"CD",X"B8",X"0B",X"C3",X"D4",X"09",X"7E",
		X"21",X"70",X"4B",X"CD",X"54",X"24",X"2E",X"74",X"C3",X"54",X"24",X"FF",X"21",X"78",X"4B",X"CD",
		X"54",X"24",X"2E",X"7C",X"C3",X"54",X"24",X"FF",X"21",X"80",X"4B",X"CD",X"54",X"24",X"2E",X"84",
		X"C3",X"54",X"24",X"FF",X"7E",X"E6",X"08",X"C8",X"2C",X"7E",X"FE",X"28",X"D0",X"7D",X"C6",X"41",
		X"6F",X"7E",X"C6",X"08",X"57",X"2C",X"7E",X"C6",X"02",X"5F",X"1A",X"A7",X"C0",X"3E",X"3E",X"12",
		X"C9",X"00",X"1C",X"C3",X"D6",X"0A",X"78",X"81",X"CD",X"95",X"24",X"2E",X"D3",X"77",X"21",X"BB",
		X"43",X"3E",X"08",X"96",X"07",X"2E",X"9A",X"86",X"07",X"47",X"2E",X"6F",X"7E",X"E6",X"1E",X"80",
		X"32",X"D1",X"4B",X"C9",X"1F",X"80",X"0D",X"C8",X"80",X"0D",X"C8",X"80",X"0D",X"C8",X"87",X"C9",
		X"21",X"95",X"43",X"7E",X"A7",X"C0",X"2E",X"B9",X"7E",X"A7",X"C2",X"B1",X"24",X"2E",X"95",X"36",
		X"FF",X"47",X"2E",X"B8",X"7E",X"E6",X"F0",X"4F",X"21",X"60",X"1F",X"E5",X"CD",X"CD",X"24",X"E1",
		X"7D",X"C6",X"04",X"6F",X"FE",X"00",X"C2",X"BB",X"24",X"C9",X"FF",X"FF",X"FF",X"7E",X"B8",X"C0",
		X"2C",X"7E",X"A9",X"E6",X"10",X"C0",X"79",X"BE",X"D8",X"2C",X"56",X"2C",X"5E",X"7D",X"E6",X"04",
		X"C6",X"EC",X"6F",X"26",X"24",X"CD",X"DC",X"07",X"03",X"C9",X"FF",X"FF",X"70",X"72",X"71",X"73",
		X"74",X"76",X"75",X"77",X"FF",X"FF",X"FF",X"FF",X"CD",X"1A",X"25",X"79",X"A7",X"C8",X"21",X"B9",
		X"43",X"7E",X"91",X"77",X"32",X"00",X"58",X"E6",X"07",X"C0",X"CD",X"50",X"06",X"21",X"B1",X"43",
		X"7E",X"FE",X"1F",X"C0",X"36",X"3F",X"C9",X"FF",X"FF",X"FF",X"21",X"95",X"43",X"7E",X"2F",X"E6",
		X"04",X"4F",X"2E",X"B9",X"7E",X"E6",X"C0",X"07",X"07",X"81",X"07",X"07",X"07",X"C3",X"26",X"23",
		X"3A",X"00",X"70",X"2F",X"E6",X"10",X"0F",X"0F",X"0F",X"00",X"81",X"07",X"07",X"07",X"4F",X"FE",
		X"40",X"DA",X"26",X"23",X"0E",X"40",X"C3",X"26",X"23",X"5E",X"5F",X"06",X"04",X"C3",X"C4",X"00",
		X"21",X"BA",X"43",X"3E",X"20",X"96",X"0F",X"E6",X"0F",X"57",X"2E",X"9F",X"86",X"4F",X"2D",X"7E",
		X"D6",X"0A",X"92",X"FE",X"E0",X"DA",X"69",X"25",X"AF",X"47",X"2E",X"9A",X"7E",X"82",X"FE",X"40",
		X"DA",X"75",X"25",X"3E",X"40",X"C6",X"88",X"57",X"2E",X"92",X"7E",X"E6",X"06",X"07",X"C6",X"70",
		X"6F",X"26",X"4B",X"E5",X"CD",X"94",X"25",X"E1",X"7D",X"C6",X"10",X"6F",X"E5",X"CD",X"94",X"25",
		X"E1",X"C9",X"FF",X"FF",X"7E",X"E6",X"08",X"C8",X"2C",X"2C",X"7E",X"B8",X"D8",X"B9",X"D0",X"2D",
		X"7E",X"FE",X"30",X"7A",X"D2",X"A9",X"25",X"C6",X"20",X"2C",X"2C",X"BE",X"D8",X"4E",X"2D",X"46",
		X"C3",X"B7",X"25",X"00",X"4F",X"2D",X"46",X"3A",X"B8",X"43",X"16",X"03",X"FE",X"10",X"DA",X"CA",
		X"25",X"16",X"04",X"FE",X"20",X"DA",X"CA",X"25",X"16",X"05",X"21",X"CC",X"43",X"7E",X"E6",X"08",
		X"CA",X"E0",X"25",X"7D",X"C6",X"04",X"6F",X"15",X"C2",X"CD",X"25",X"E1",X"E1",X"C9",X"FF",X"FF",
		X"78",X"C6",X"04",X"47",X"79",X"C6",X"0C",X"4F",X"36",X"08",X"2C",X"78",X"0F",X"E6",X"03",X"57",
		X"79",X"E6",X"04",X"82",X"C6",X"58",X"77",X"2C",X"70",X"2C",X"71",X"E1",X"E1",X"C9",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"3A",X"B9",X"43",X"2F",X"0F",X"0F",X"0F",X"E6",X"1F",X"21",X"D2",
		X"4B",X"77",X"2C",X"3A",X"D1",X"4B",X"BE",X"DA",X"50",X"26",X"3A",X"D5",X"4B",X"57",X"E6",X"03",
		X"5F",X"3A",X"9B",X"43",X"07",X"07",X"E6",X"0C",X"83",X"C6",X"D0",X"6F",X"26",X"3E",X"7A",X"0F",
		X"0F",X"E6",X"07",X"86",X"57",X"3A",X"B9",X"43",X"92",X"32",X"B9",X"43",X"32",X"00",X"58",X"3A",
		X"9B",X"43",X"0F",X"D2",X"D0",X"26",X"CD",X"68",X"26",X"C3",X"AA",X"26",X"C2",X"3A",X"26",X"3A",
		X"2C",X"3A",X"9B",X"43",X"07",X"07",X"E6",X"0C",X"86",X"C6",X"D0",X"6F",X"26",X"3E",X"3A",X"B9",
		X"43",X"86",X"C3",X"39",X"26",X"D2",X"AE",X"26",X"3A",X"6E",X"43",X"C6",X"02",X"47",X"3A",X"9A",
		X"43",X"57",X"0F",X"0F",X"E6",X"0F",X"80",X"47",X"21",X"BB",X"43",X"3E",X"08",X"96",X"0F",X"E6",
		X"03",X"80",X"47",X"5E",X"00",X"3A",X"D6",X"4B",X"C6",X"E0",X"6F",X"26",X"3E",X"78",X"BE",X"DA",
		X"93",X"26",X"46",X"7A",X"E6",X"F8",X"80",X"47",X"7B",X"FE",X"04",X"D2",X"A4",X"26",X"2F",X"00",
		X"E6",X"03",X"80",X"47",X"78",X"32",X"D5",X"4B",X"C9",X"58",X"21",X"D3",X"4B",X"7E",X"35",X"A7",
		X"C0",X"34",X"2E",X"D6",X"7E",X"FE",X"0C",X"D0",X"FE",X"08",X"D8",X"2C",X"96",X"07",X"47",X"3A",
		X"6F",X"43",X"E6",X"03",X"2E",X"D4",X"77",X"2F",X"E6",X"03",X"3C",X"4F",X"C3",X"76",X"24",X"C9",
		X"21",X"A8",X"4B",X"01",X"00",X"08",X"11",X"00",X"80",X"7E",X"A7",X"CA",X"E5",X"26",X"7A",X"07",
		X"D2",X"E4",X"26",X"51",X"59",X"0C",X"7D",X"90",X"6F",X"FE",X"68",X"C2",X"D9",X"26",X"3A",X"D2",
		X"4B",X"82",X"83",X"E6",X"1F",X"32",X"D6",X"4B",X"7B",X"92",X"32",X"D7",X"4B",X"C9",X"FF",X"FF",
		X"21",X"A2",X"43",X"7E",X"A7",X"C8",X"2C",X"7E",X"E6",X"01",X"07",X"07",X"C6",X"83",X"6F",X"3E",
		X"FF",X"32",X"97",X"43",X"11",X"70",X"43",X"CD",X"48",X"27",X"1C",X"1C",X"1C",X"7B",X"FE",X"80",
		X"C2",X"17",X"27",X"1E",X"9D",X"3A",X"A4",X"43",X"FE",X"06",X"DA",X"39",X"27",X"1A",X"47",X"0E",
		X"00",X"CD",X"20",X"02",X"AF",X"12",X"32",X"97",X"43",X"3A",X"97",X"43",X"A7",X"CC",X"68",X"27",
		X"CD",X"A8",X"27",X"C3",X"43",X"3B",X"FF",X"FF",X"1A",X"1C",X"E6",X"1F",X"FE",X"01",X"C0",X"1A",
		X"A7",X"C8",X"0F",X"0F",X"0F",X"0F",X"47",X"E6",X"F0",X"4F",X"78",X"E6",X"0F",X"47",X"CD",X"20",
		X"02",X"AF",X"12",X"32",X"97",X"43",X"C9",X"FF",X"E5",X"11",X"61",X"42",X"06",X"06",X"3A",X"A3",
		X"43",X"A7",X"CA",X"78",X"27",X"11",X"21",X"40",X"CD",X"C4",X"00",X"E1",X"11",X"BD",X"43",X"EB",
		X"7E",X"2C",X"B6",X"C8",X"2C",X"EB",X"CD",X"14",X"03",X"D0",X"3A",X"A3",X"43",X"C6",X"90",X"6F",
		X"34",X"CD",X"67",X"03",X"3E",X"FF",X"32",X"6A",X"43",X"2E",X"BE",X"7E",X"36",X"00",X"0F",X"0F",
		X"0F",X"0F",X"2D",X"77",X"C9",X"FF",X"FF",X"FF",X"21",X"8C",X"43",X"7E",X"32",X"00",X"60",X"2C",
		X"7E",X"32",X"00",X"68",X"36",X"0F",X"2D",X"36",X"0F",X"C9",X"C9",X"FF",X"FF",X"21",X"63",X"43",
		X"7E",X"A7",X"C8",X"FE",X"40",X"DA",X"CA",X"27",X"36",X"40",X"35",X"2E",X"8C",X"36",X"8F",X"E1",
		X"C9",X"FF",X"21",X"61",X"43",X"06",X"7F",X"7E",X"A7",X"CA",X"E2",X"27",X"06",X"FF",X"3D",X"E6",
		X"02",X"77",X"78",X"30",X"C9",X"E9",X"CD",X"7C",X"3D",X"CD",X"98",X"3D",X"78",X"A7",X"C8",X"21",
		X"8D",X"43",X"36",X"2F",X"79",X"A7",X"C8",X"0F",X"E6",X"06",X"F6",X"20",X"77",X"C9",X"C9",X"FF",
		X"10",X"24",X"10",X"00",X"10",X"24",X"10",X"4C",X"10",X"74",X"10",X"A8",X"10",X"74",X"10",X"A8",
		X"10",X"D0",X"10",X"FC",X"10",X"D0",X"10",X"FC",X"10",X"D0",X"10",X"FC",X"10",X"D0",X"10",X"FC",
		X"11",X"C2",X"11",X"24",X"11",X"C2",X"11",X"24",X"11",X"4E",X"11",X"86",X"11",X"4E",X"11",X"EA",
		X"11",X"86",X"12",X"18",X"12",X"46",X"12",X"18",X"12",X"46",X"12",X"18",X"12",X"46",X"12",X"18",
		X"2D",X"12",X"2C",X"00",X"2D",X"12",X"2C",X"00",X"2C",X"D4",X"2D",X"5C",X"2C",X"D4",X"2C",X"36",
		X"2D",X"32",X"2C",X"64",X"2C",X"A8",X"2D",X"32",X"2C",X"A8",X"2C",X"64",X"2C",X"A8",X"2D",X"32",
		X"12",X"70",X"13",X"78",X"12",X"70",X"13",X"78",X"12",X"A2",X"12",X"E0",X"13",X"A2",X"13",X"0E",
		X"13",X"A2",X"13",X"D0",X"13",X"0E",X"13",X"44",X"13",X"0E",X"13",X"D0",X"13",X"44",X"13",X"0E",
		X"2E",X"AE",X"2E",X"74",X"2E",X"AE",X"2E",X"56",X"2E",X"74",X"2E",X"8C",X"2E",X"EC",X"2E",X"8C",
		X"2E",X"74",X"2E",X"8C",X"2E",X"EC",X"2E",X"8C",X"2E",X"EC",X"2E",X"8C",X"2E",X"EC",X"2E",X"8C",
		X"2D",X"E8",X"2D",X"8A",X"2D",X"E8",X"2D",X"AC",X"2E",X"28",X"2D",X"C4",X"2E",X"28",X"2D",X"C4",
		X"2D",X"AC",X"2D",X"C4",X"2E",X"28",X"2D",X"C4",X"2E",X"28",X"2D",X"C4",X"2E",X"28",X"2D",X"C4",
		X"2C",X"00",X"2C",X"D4",X"2C",X"00",X"2F",X"6A",X"2F",X"94",X"2C",X"D4",X"2F",X"6A",X"2C",X"36",
		X"2F",X"94",X"2C",X"64",X"2C",X"A8",X"2C",X"64",X"2C",X"A8",X"2F",X"94",X"2C",X"64",X"2C",X"A8",
		X"12",X"70",X"12",X"A2",X"12",X"70",X"12",X"A2",X"2F",X"42",X"13",X"0E",X"12",X"E0",X"2F",X"1C",
		X"13",X"0E",X"2F",X"1C",X"2F",X"42",X"13",X"44",X"13",X"44",X"2F",X"1C",X"2F",X"42",X"13",X"44",
		X"41",X"30",X"00",X"18",X"31",X"28",X"C8",X"18",X"51",X"40",X"10",X"A0",X"13",X"20",X"C8",X"A0",
		X"41",X"40",X"C8",X"28",X"61",X"40",X"00",X"28",X"12",X"20",X"60",X"A0",X"61",X"50",X"40",X"A0",
		X"61",X"38",X"28",X"28",X"51",X"30",X"C8",X"38",X"13",X"20",X"00",X"18",X"15",X"40",X"00",X"A0",
		X"61",X"50",X"C8",X"A0",X"41",X"20",X"28",X"28",X"31",X"20",X"A0",X"A0",X"13",X"20",X"C8",X"18",
		X"13",X"04",X"00",X"18",X"51",X"30",X"08",X"18",X"13",X"04",X"C8",X"18",X"31",X"20",X"B8",X"18",
		X"13",X"30",X"80",X"A0",X"51",X"28",X"C8",X"38",X"61",X"40",X"28",X"28",X"13",X"08",X"00",X"A0",
		X"51",X"40",X"00",X"A0",X"13",X"08",X"70",X"A0",X"51",X"40",X"C8",X"A0",X"32",X"30",X"C8",X"18",
		X"22",X"20",X"00",X"18",X"31",X"30",X"00",X"28",X"51",X"40",X"B8",X"A0",X"31",X"20",X"28",X"A0",
		X"11",X"10",X"50",X"48",X"13",X"30",X"00",X"18",X"41",X"40",X"68",X"48",X"12",X"10",X"C8",X"18",
		X"21",X"30",X"70",X"48",X"21",X"20",X"C8",X"38",X"31",X"30",X"60",X"48",X"11",X"10",X"00",X"28",
		X"21",X"20",X"58",X"48",X"21",X"30",X"00",X"28",X"31",X"30",X"70",X"48",X"21",X"20",X"C8",X"28",
		X"31",X"20",X"50",X"48",X"13",X"30",X"C8",X"18",X"21",X"20",X"68",X"48",X"21",X"40",X"00",X"18",
		X"31",X"30",X"58",X"48",X"31",X"20",X"00",X"38",X"21",X"20",X"60",X"48",X"31",X"30",X"C8",X"38",
		X"31",X"20",X"50",X"48",X"31",X"30",X"C8",X"28",X"21",X"20",X"58",X"48",X"31",X"30",X"00",X"38",
		X"41",X"40",X"70",X"48",X"41",X"38",X"00",X"18",X"11",X"10",X"68",X"48",X"41",X"40",X"C8",X"18",
		X"21",X"30",X"60",X"48",X"41",X"20",X"C8",X"18",X"31",X"30",X"70",X"48",X"13",X"20",X"00",X"18",
		X"F2",X"20",X"50",X"20",X"4A",X"20",X"44",X"20",X"34",X"40",X"2A",X"40",X"1C",X"60",X"0E",X"60",
		X"00",X"60",X"1C",X"60",X"00",X"60",X"0E",X"60",X"2A",X"40",X"3E",X"20",X"34",X"40",X"3E",X"20",
		X"F2",X"20",X"50",X"20",X"4A",X"20",X"44",X"20",X"34",X"40",X"2A",X"40",X"1C",X"60",X"0E",X"60",
		X"1C",X"60",X"2A",X"40",X"3E",X"20",X"34",X"40",X"3E",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"20",X"50",X"20",X"4A",X"20",X"44",X"20",X"34",X"40",X"2A",X"40",X"1C",X"60",X"2A",X"40",
		X"34",X"40",X"3E",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"C4",X"BB",X"B2",X"A9",X"A0",X"B2",X"A9",X"A0",X"B2",X"A9",X"A0",X"00",X"00",X"00",X"00",
		X"F2",X"C4",X"BB",X"B2",X"BB",X"B2",X"A9",X"A0",X"A9",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"C4",X"BB",X"C4",X"B2",X"BB",X"A9",X"B2",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"56",X"EB",X"E5",X"D9",X"D3",X"CD",X"E5",X"EB",X"C3",X"98",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"15",X"90",X"15",X"84",X"15",X"6C",X"17",X"CA",X"15",X"6C",X"17",X"CA",X"17",X"A0",X"17",X"70",
		X"17",X"A0",X"17",X"70",X"17",X"CA",X"17",X"70",X"17",X"A0",X"17",X"CA",X"15",X"6C",X"15",X"78",
		X"08",X"00",X"00",X"FF",X"02",X"00",X"F8",X"FF",X"08",X"02",X"02",X"FF",X"04",X"00",X"FA",X"FF",
		X"08",X"04",X"04",X"FF",X"06",X"00",X"FC",X"FF",X"08",X"06",X"06",X"FF",X"08",X"00",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"03",X"02",X"02",X"02",X"02",X"03",X"FF",
		X"03",X"02",X"02",X"01",X"01",X"02",X"02",X"03",X"03",X"02",X"01",X"00",X"00",X"01",X"02",X"03",
		X"03",X"02",X"01",X"00",X"00",X"01",X"02",X"03",X"03",X"02",X"02",X"01",X"01",X"02",X"02",X"03",
		X"FF",X"03",X"02",X"02",X"02",X"02",X"03",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"FF",X"FF",X"01",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"01",X"03",X"03",X"03",X"03",X"01",X"FF",
		X"01",X"03",X"03",X"00",X"00",X"03",X"03",X"01",X"01",X"03",X"00",X"02",X"02",X"00",X"03",X"01",
		X"01",X"03",X"00",X"02",X"02",X"00",X"03",X"01",X"01",X"03",X"03",X"00",X"00",X"03",X"03",X"01",
		X"FF",X"01",X"03",X"03",X"03",X"03",X"01",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"FF",X"FF",
		X"A0",X"42",X"04",X"00",X"AB",X"42",X"88",X"40",X"B6",X"41",X"88",X"00",X"A0",X"42",X"0C",X"40",
		X"AB",X"42",X"46",X"00",X"B6",X"41",X"C6",X"40",X"A0",X"42",X"4A",X"00",X"A9",X"41",X"CA",X"40",
		X"1B",X"1C",X"2E",X"2D",X"2E",X"2D",X"1C",X"1B",X"00",X"00",X"00",X"CE",X"B9",X"CE",X"B9",X"B7",
		X"B6",X"B7",X"B6",X"00",X"00",X"00",X"FC",X"FD",X"FE",X"FF",X"FC",X"FD",X"FE",X"FF",X"00",X"00",
		X"38",X"10",X"48",X"E7",X"48",X"20",X"48",X"49",X"68",X"30",X"4A",X"8D",X"C0",X"40",X"4A",X"98",
		X"B0",X"50",X"49",X"76",X"90",X"60",X"48",X"72",X"50",X"70",X"49",X"6A",X"28",X"00",X"49",X"E5",
		X"08",X"10",X"49",X"41",X"55",X"20",X"4A",X"0B",X"88",X"30",X"49",X"71",X"A8",X"40",X"4A",X"F5",
		X"D0",X"50",X"48",X"77",X"78",X"60",X"48",X"6F",X"28",X"70",X"48",X"84",X"10",X"00",X"4A",X"FE",
		X"12",X"12",X"11",X"10",X"1F",X"1E",X"1F",X"10",X"10",X"11",X"12",X"13",X"14",X"14",X"15",X"16",
		X"17",X"18",X"18",X"19",X"1A",X"1B",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"11",X"12",X"13",
		X"14",X"0F",X"0F",X"0F",X"0F",X"15",X"16",X"17",X"18",X"17",X"16",X"15",X"15",X"16",X"17",X"18",
		X"18",X"19",X"19",X"19",X"00",X"FF",X"13",X"13",X"13",X"14",X"14",X"15",X"15",X"14",X"14",X"13",
		X"12",X"11",X"11",X"10",X"1F",X"1E",X"1E",X"1D",X"1C",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",
		X"15",X"0F",X"0F",X"13",X"12",X"12",X"11",X"11",X"11",X"11",X"10",X"10",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"00",X"FF",X"FF",X"13",X"13",X"13",X"12",X"12",X"12",X"11",X"10",X"10",X"10",X"10",X"1F",
		X"1E",X"1D",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"11",X"12",X"13",X"14",X"14",X"15",X"16",X"17",
		X"18",X"19",X"1A",X"1B",X"1C",X"1C",X"1B",X"1A",X"19",X"18",X"18",X"18",X"18",X"18",X"17",X"16",
		X"15",X"0F",X"0F",X"0F",X"0F",X"13",X"13",X"12",X"12",X"12",X"12",X"11",X"11",X"11",X"11",X"10",
		X"10",X"10",X"1F",X"1F",X"1F",X"00",X"FF",X"FF",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"11",X"13",X"14",X"15",X"17",X"18",X"17",X"16",X"15",X"0F",X"06",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"13",X"12",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"00",X"FF",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0E",X"0E",X"05",
		X"1C",X"1B",X"1A",X"19",X"18",X"18",X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"14",X"13",X"12",
		X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"12",X"13",X"0F",X"06",X"0A",X"0A",X"0B",X"0B",
		X"0B",X"0B",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0C",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"11",X"11",X"12",X"12",X"13",X"13",X"14",X"14",X"14",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"1C",X"1B",X"1A",X"1A",X"19",X"19",X"00",
		X"FF",X"FF",X"11",X"11",X"12",X"12",X"13",X"13",X"14",X"15",X"17",X"18",X"19",X"1B",X"1C",X"1D",
		X"1F",X"10",X"11",X"11",X"12",X"12",X"13",X"13",X"14",X"14",X"0F",X"0F",X"04",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"03",X"1C",X"1D",X"1E",X"1F",X"1F",X"00",X"FF",X"13",X"13",X"13",X"13",
		X"13",X"13",X"12",X"11",X"10",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",
		X"14",X"14",X"14",X"13",X"13",X"0F",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"1C",X"1D",X"1E",X"1F",X"1F",X"1F",X"1F",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"09",X"0A",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"FF",X"FF",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0A",X"09",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"00",X"FF",X"FF",X"1C",X"1C",X"1D",X"1E",X"1F",X"10",X"10",X"11",X"12",X"12",X"13",X"0F",
		X"06",X"0B",X"0B",X"0B",X"0A",X"09",X"08",X"08",X"09",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"FF",X"FF",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"18",X"18",X"18",X"19",X"1A",X"1A",X"1B",X"1C",X"1C",X"1C",X"1D",X"1E",X"1E",X"1F",X"10",X"10",
		X"10",X"10",X"11",X"12",X"12",X"13",X"14",X"14",X"14",X"14",X"15",X"15",X"16",X"16",X"17",X"18",
		X"18",X"18",X"19",X"1A",X"1A",X"0F",X"0F",X"0F",X"13",X"12",X"11",X"10",X"10",X"1F",X"1E",X"0F",
		X"0F",X"16",X"17",X"17",X"17",X"17",X"00",X"FF",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"18",X"18",X"18",X"19",X"1A",X"1B",X"1C",X"1C",X"1C",X"1D",X"1E",X"1E",X"1F",X"10",X"10",X"10",
		X"11",X"12",X"12",X"13",X"0F",X"0F",X"0F",X"15",X"15",X"16",X"16",X"16",X"17",X"17",X"17",X"17",
		X"17",X"17",X"17",X"17",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"06",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0A",X"09",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"00",X"FF",X"FF",X"08",X"08",X"08",X"08",X"08",X"09",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0A",X"09",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"FF",X"FF",X"1C",X"1B",X"1A",X"19",
		X"18",X"18",X"17",X"16",X"15",X"0F",X"06",X"08",X"08",X"08",X"09",X"0A",X"0B",X"0B",X"0A",X"09",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"FF",X"FF",X"16",X"15",
		X"14",X"14",X"13",X"12",X"11",X"10",X"1F",X"1E",X"1E",X"1D",X"1C",X"1C",X"1C",X"1B",X"1A",X"1A",
		X"19",X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"14",X"14",X"14",X"14",X"13",X"12",X"12",X"11",
		X"11",X"10",X"10",X"10",X"1F",X"1E",X"1D",X"0F",X"0F",X"0F",X"15",X"16",X"17",X"18",X"18",X"18",
		X"19",X"1A",X"0F",X"0F",X"0F",X"13",X"12",X"12",X"11",X"11",X"00",X"FF",X"16",X"15",X"14",X"14",
		X"13",X"12",X"11",X"10",X"10",X"1F",X"1E",X"1D",X"1C",X"1C",X"1C",X"1C",X"1B",X"1A",X"1A",X"19",
		X"18",X"18",X"18",X"18",X"17",X"16",X"16",X"15",X"14",X"14",X"14",X"13",X"13",X"12",X"12",X"12",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"FF",X"15",X"15",X"15",X"15",
		X"15",X"15",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1D",X"1E",X"1F",X"10",X"11",X"12",X"12",
		X"13",X"0F",X"0F",X"0F",X"06",X"0B",X"0B",X"0B",X"0B",X"0D",X"0D",X"0D",X"0B",X"0B",X"0B",X"0B",
		X"00",X"FF",X"0B",X"0B",X"0D",X"0D",X"0B",X"0D",X"0B",X"0D",X"0B",X"0B",X"0A",X"0A",X"0A",X"09",
		X"09",X"09",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"0A",X"0B",X"0B",X"0D",X"0D",
		X"0B",X"0B",X"0D",X"0D",X"0B",X"0B",X"0D",X"00",X"FF",X"FF",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"12",X"11",X"10",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",
		X"14",X"0F",X"0F",X"0F",X"0F",X"0F",X"06",X"09",X"08",X"08",X"0E",X"0E",X"0E",X"08",X"08",X"0E",
		X"0E",X"00",X"FF",X"FF",X"11",X"10",X"1F",X"10",X"11",X"10",X"1F",X"10",X"11",X"10",X"1F",X"10",
		X"11",X"11",X"12",X"0F",X"06",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0A",
		X"09",X"08",X"08",X"08",X"0E",X"0E",X"0E",X"0E",X"08",X"08",X"08",X"0E",X"0E",X"00",X"FF",X"FF",
		X"7E",X"E6",X"1F",X"C8",X"35",X"7E",X"CA",X"EC",X"2F",X"E6",X"E7",X"C2",X"95",X"0F",X"2C",X"46",
		X"2C",X"56",X"2C",X"5E",X"7B",X"E6",X"1F",X"FE",X"04",X"D8",X"1D",X"21",X"E0",X"FF",X"19",X"36",
		X"20",X"21",X"E2",X"4B",X"70",X"06",X"02",X"C3",X"C4",X"00",X"FF",X"FF",X"2C",X"2C",X"2C",X"7E",
		X"E6",X"1F",X"FE",X"04",X"D8",X"35",X"2D",X"2D",X"2D",X"7E",X"C3",X"96",X"0F",X"FF",X"FF",X"FF",
		X"21",X"93",X"43",X"7E",X"34",X"07",X"E6",X"06",X"C6",X"16",X"6F",X"26",X"30",X"7E",X"23",X"6E",
		X"67",X"E9",X"FF",X"FF",X"FF",X"FF",X"30",X"20",X"30",X"A0",X"31",X"94",X"31",X"40",X"FF",X"FF",
		X"21",X"D0",X"4B",X"7E",X"A7",X"C0",X"23",X"23",X"7E",X"A7",X"CA",X"3F",X"30",X"35",X"7E",X"E6",
		X"03",X"C0",X"2D",X"7E",X"E6",X"F0",X"C8",X"7E",X"D6",X"10",X"77",X"2D",X"36",X"01",X"C9",X"3E",
		X"FF",X"32",X"D9",X"4B",X"11",X"D1",X"4B",X"21",X"B4",X"43",X"7E",X"2C",X"6E",X"67",X"06",X"04",
		X"CD",X"E0",X"05",X"7D",X"E6",X"7F",X"C2",X"5D",X"30",X"7D",X"C6",X"80",X"6F",X"7D",X"32",X"B5",
		X"43",X"CD",X"78",X"30",X"0F",X"E6",X"3F",X"4F",X"21",X"D2",X"4B",X"7E",X"91",X"36",X"03",X"D8",
		X"FE",X"04",X"D8",X"77",X"C9",X"FF",X"FF",X"FF",X"21",X"B8",X"43",X"7E",X"0F",X"0F",X"E6",X"1C",
		X"4F",X"2C",X"2C",X"3E",X"10",X"96",X"81",X"4F",X"2E",X"9A",X"7E",X"0F",X"E6",X"7F",X"FE",X"20",
		X"DA",X"95",X"30",X"3E",X"1F",X"81",X"4F",X"C9",X"C3",X"8B",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"D0",X"4B",X"7E",X"FE",X"01",X"C0",X"21",X"70",X"4B",X"01",X"08",X"00",X"7E",X"E6",X"08",
		X"CA",X"B4",X"30",X"04",X"2C",X"2C",X"2C",X"2C",X"0D",X"C2",X"AD",X"30",X"21",X"E4",X"4B",X"70",
		X"21",X"D0",X"4B",X"36",X"00",X"3A",X"BA",X"43",X"90",X"C8",X"36",X"02",X"2C",X"47",X"7E",X"E6",
		X"0F",X"2E",X"D7",X"77",X"B8",X"D8",X"70",X"C9",X"4B",X"7E",X"FE",X"02",X"C0",X"34",X"2E",X"D3",
		X"3A",X"C2",X"43",X"96",X"16",X"00",X"D2",X"ED",X"30",X"2F",X"3C",X"16",X"20",X"47",X"0F",X"0F",
		X"0F",X"E6",X"1F",X"5F",X"CD",X"78",X"30",X"0F",X"00",X"E6",X"3F",X"4F",X"78",X"E6",X"0F",X"91",
		X"D2",X"05",X"31",X"3E",X"00",X"83",X"FE",X"20",X"DA",X"0D",X"31",X"3E",X"1F",X"E6",X"1E",X"B2",
		X"47",X"21",X"D4",X"4B",X"7E",X"FE",X"40",X"3E",X"00",X"D2",X"1E",X"31",X"3E",X"40",X"B0",X"47",
		X"3A",X"B8",X"43",X"E6",X"0F",X"FE",X"01",X"3E",X"00",X"CA",X"2E",X"31",X"3E",X"80",X"B0",X"5F",
		X"16",X"28",X"2E",X"D5",X"1A",X"77",X"2C",X"1C",X"1A",X"77",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"D0",X"4B",X"7E",X"FE",X"03",X"C0",X"36",X"00",X"11",X"70",X"4B",X"01",X"50",X"4B",X"3A",
		X"D3",X"4B",X"32",X"D8",X"4B",X"1A",X"E6",X"08",X"CA",X"6C",X"31",X"13",X"13",X"13",X"13",X"03",
		X"03",X"00",X"00",X"7B",X"FE",X"90",X"C2",X"55",X"31",X"C9",X"FF",X"FF",X"1A",X"E6",X"F0",X"F6",
		X"0C",X"12",X"13",X"13",X"2E",X"D8",X"7E",X"12",X"C6",X"10",X"77",X"13",X"2E",X"D4",X"7E",X"12",
		X"23",X"7E",X"02",X"23",X"03",X"7E",X"02",X"13",X"03",X"23",X"35",X"C2",X"63",X"31",X"C9",X"00",
		X"FF",X"FF",X"FF",X"FF",X"21",X"D0",X"4B",X"7E",X"FE",X"02",X"C0",X"34",X"2E",X"D9",X"34",X"C0",
		X"C3",X"DE",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"B9",X"43",X"7E",X"A7",X"C0",X"2E",X"B2",
		X"7E",X"FE",X"1F",X"C0",X"2E",X"C2",X"7E",X"E6",X"07",X"C6",X"66",X"6F",X"26",X"32",X"46",X"3A",
		X"B8",X"43",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"80",X"FE",X"08",X"DA",X"D0",X"31",X"3E",X"00",
		X"47",X"0F",X"0F",X"0F",X"21",X"A5",X"43",X"77",X"2D",X"36",X"07",X"78",X"C6",X"6E",X"6F",X"26",
		X"32",X"7E",X"21",X"9D",X"43",X"77",X"2C",X"36",X"00",X"11",X"79",X"41",X"06",X"04",X"CD",X"C4",
		X"00",X"C3",X"00",X"07",X"C3",X"B4",X"32",X"35",X"CA",X"30",X"32",X"7E",X"E6",X"1F",X"CA",X"80",
		X"03",X"FE",X"1F",X"C2",X"0B",X"32",X"3E",X"10",X"32",X"63",X"43",X"7E",X"0F",X"0F",X"E6",X"07",
		X"4F",X"7E",X"E6",X"E0",X"0F",X"0F",X"0F",X"C6",X"80",X"6F",X"26",X"2B",X"06",X"2B",X"7E",X"81",
		X"4F",X"23",X"56",X"23",X"5E",X"23",X"6E",X"26",X"2B",X"C3",X"40",X"32",X"FF",X"FF",X"FF",X"FF",
		X"2E",X"A4",X"36",X"02",X"2E",X"B8",X"7E",X"E6",X"F0",X"C6",X"10",X"77",X"C3",X"80",X"03",X"FF",
		X"D5",X"3E",X"00",X"12",X"7E",X"FE",X"FF",X"CA",X"50",X"32",X"C5",X"81",X"4F",X"0A",X"12",X"C1",
		X"13",X"23",X"7D",X"E6",X"07",X"C2",X"41",X"32",X"D1",X"CD",X"17",X"02",X"7D",X"E6",X"3F",X"C2",
		X"40",X"32",X"C9",X"FF",X"FF",X"FF",X"01",X"02",X"03",X"03",X"03",X"02",X"01",X"01",X"40",X"05",
		X"10",X"15",X"20",X"25",X"30",X"35",X"21",X"95",X"43",X"7E",X"A7",X"C0",X"2E",X"B9",X"46",X"2D",
		X"7E",X"2F",X"0F",X"E6",X"30",X"4F",X"7E",X"E6",X"10",X"07",X"C6",X"C0",X"6F",X"26",X"2B",X"E5",
		X"CD",X"A0",X"32",X"E1",X"7D",X"C6",X"04",X"6F",X"E6",X"1F",X"C2",X"8F",X"32",X"C9",X"FF",X"FF",
		X"7E",X"B8",X"C0",X"2C",X"3A",X"83",X"43",X"AE",X"A1",X"C0",X"2C",X"56",X"2C",X"5E",X"3E",X"6F",
		X"12",X"C9",X"FF",X"FF",X"21",X"9B",X"43",X"7E",X"0F",X"D8",X"2E",X"A5",X"C3",X"F7",X"31",X"3A",
		X"BB",X"43",X"A7",X"C8",X"07",X"07",X"07",X"4F",X"21",X"70",X"4B",X"06",X"80",X"CD",X"D8",X"05",
		X"16",X"4B",X"26",X"3F",X"3E",X"40",X"91",X"C6",X"70",X"5F",X"C6",X"10",X"6F",X"41",X"3A",X"B8",
		X"43",X"E6",X"10",X"CA",X"E0",X"05",X"7D",X"C6",X"40",X"6F",X"C3",X"E0",X"05",X"CD",X"E0",X"05",
		X"21",X"E2",X"43",X"56",X"2C",X"5E",X"2E",X"B9",X"7E",X"C6",X"04",X"0F",X"0F",X"0F",X"83",X"E6",
		X"1F",X"47",X"7B",X"E6",X"E0",X"B0",X"5F",X"7A",X"C6",X"08",X"57",X"01",X"02",X"02",X"C5",X"D5",
		X"CD",X"2A",X"33",X"D1",X"C1",X"CD",X"9B",X"33",X"05",X"C2",X"0E",X"33",X"CD",X"F0",X"33",X"06",
		X"02",X"0D",X"C2",X"0E",X"33",X"C3",X"90",X"37",X"FF",X"FF",X"1A",X"FE",X"6F",X"D8",X"16",X"A8",
		X"CA",X"70",X"33",X"FE",X"7C",X"D0",X"FE",X"78",X"D2",X"42",X"33",X"E6",X"03",X"07",X"07",X"C6",
		X"AC",X"57",X"CD",X"4C",X"33",X"C8",X"E1",X"E1",X"E1",X"C3",X"C4",X"0C",X"78",X"E6",X"01",X"47",
		X"79",X"E6",X"01",X"07",X"B0",X"47",X"3A",X"B9",X"43",X"E6",X"04",X"B0",X"6F",X"26",X"3E",X"46",
		X"3A",X"C2",X"43",X"0F",X"E6",X"03",X"82",X"6F",X"26",X"33",X"7E",X"A0",X"C9",X"FF",X"FF",X"FF",
		X"CD",X"4C",X"33",X"C8",X"E1",X"E1",X"C1",X"AF",X"77",X"11",X"69",X"43",X"2F",X"12",X"21",X"70",
		X"43",X"36",X"1A",X"2C",X"1E",X"B9",X"1A",X"2F",X"0F",X"E6",X"70",X"C6",X"10",X"77",X"2C",X"1E",
		X"E2",X"1A",X"77",X"2C",X"1C",X"1A",X"3D",X"3D",X"77",X"C9",X"E1",X"2E",X"01",X"7B",X"85",X"E6",
		X"1F",X"6F",X"7B",X"E6",X"E0",X"B5",X"5F",X"C9",X"FB",X"FA",X"EE",X"CC",X"33",X"3B",X"3A",X"EA",
		X"BB",X"BB",X"FE",X"EF",X"1A",X"4A",X"CC",X"CC",X"BB",X"FA",X"EE",X"CC",X"21",X"E2",X"43",X"56",
		X"2C",X"5E",X"13",X"13",X"2E",X"C2",X"7E",X"E6",X"06",X"47",X"2E",X"9B",X"7E",X"07",X"E6",X"08",
		X"80",X"C6",X"70",X"6F",X"26",X"1B",X"CD",X"E6",X"33",X"3A",X"B8",X"43",X"E6",X"0F",X"FE",X"02",
		X"C0",X"2D",X"1C",X"CD",X"10",X"02",X"7E",X"12",X"CD",X"17",X"02",X"2C",X"7E",X"12",X"C9",X"34",
		X"2E",X"FE",X"CD",X"9D",X"33",X"C3",X"17",X"02",X"60",X"32",X"61",X"34",X"62",X"32",X"61",X"34",
		X"CD",X"76",X"08",X"CD",X"00",X"38",X"CD",X"00",X"26",X"CD",X"00",X"38",X"CD",X"80",X"39",X"3A",
		X"BB",X"43",X"A7",X"CA",X"62",X"34",X"FE",X"04",X"D2",X"38",X"34",X"CD",X"74",X"34",X"CD",X"86",
		X"34",X"CD",X"60",X"35",X"CD",X"98",X"34",X"CD",X"AA",X"34",X"3A",X"9B",X"43",X"0F",X"DA",X"78",
		X"0F",X"CD",X"30",X"39",X"C3",X"40",X"0C",X"FF",X"3A",X"9B",X"43",X"0F",X"DA",X"52",X"34",X"CD",
		X"74",X"34",X"CD",X"60",X"35",X"CD",X"98",X"34",X"CD",X"30",X"39",X"C3",X"40",X"0C",X"FF",X"FF",
		X"FF",X"FF",X"CD",X"86",X"34",X"CD",X"60",X"35",X"CD",X"AA",X"34",X"C3",X"78",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"3A",X"9B",X"43",X"0F",X"D8",X"CD",X"40",X"0C",X"CD",X"78",X"0F",X"C3",X"04",X"22",
		X"FF",X"FF",X"FF",X"FF",X"21",X"70",X"4B",X"E5",X"CD",X"C0",X"34",X"E1",X"7D",X"C6",X"08",X"6F",
		X"FE",X"90",X"C2",X"77",X"34",X"C9",X"21",X"90",X"4B",X"E5",X"CD",X"C0",X"34",X"E1",X"7D",X"C6",
		X"08",X"6F",X"FE",X"B0",X"C2",X"89",X"34",X"C9",X"21",X"70",X"4B",X"E5",X"CD",X"B0",X"35",X"E1",
		X"7D",X"C6",X"08",X"6F",X"FE",X"90",X"C2",X"9B",X"34",X"C9",X"21",X"90",X"4B",X"E5",X"CD",X"B0",
		X"35",X"E1",X"7D",X"C6",X"08",X"6F",X"FE",X"B0",X"C2",X"AD",X"34",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"A7",X"C8",X"47",X"C6",X"C0",X"5F",X"16",X"3E",X"1A",X"4F",X"2C",X"56",X"2C",X"5E",X"2C",
		X"78",X"07",X"07",X"07",X"86",X"E6",X"7E",X"6F",X"26",X"3E",X"7E",X"2C",X"6E",X"67",X"7A",X"FE",
		X"4B",X"C2",X"0C",X"35",X"7B",X"FE",X"50",X"DA",X"0C",X"35",X"06",X"08",X"2C",X"2C",X"D6",X"20",
		X"5F",X"FE",X"50",X"DA",X"09",X"35",X"06",X"10",X"2C",X"2C",X"D6",X"20",X"5F",X"FE",X"50",X"DA",
		X"09",X"35",X"06",X"18",X"2C",X"2C",X"D6",X"20",X"5F",X"79",X"80",X"4F",X"06",X"35",X"C5",X"01",
		X"DF",X"FF",X"EB",X"36",X"00",X"23",X"36",X"00",X"09",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",
		X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"36",X"00",X"23",X"36",X"00",X"C9",X"FF",X"FF",
		X"CD",X"58",X"37",X"47",X"07",X"07",X"4F",X"07",X"07",X"B0",X"32",X"6F",X"43",X"3A",X"B8",X"43",
		X"FE",X"40",X"DA",X"77",X"35",X"3E",X"30",X"E6",X"30",X"0F",X"47",X"3A",X"BB",X"43",X"3D",X"FE",
		X"04",X"DA",X"86",X"35",X"3E",X"03",X"07",X"B0",X"47",X"3A",X"9A",X"43",X"07",X"07",X"E6",X"20",
		X"B0",X"C6",X"80",X"6F",X"26",X"3E",X"7E",X"32",X"6E",X"43",X"2C",X"7E",X"81",X"E6",X"F8",X"32",
		X"6D",X"43",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"A7",X"C8",X"47",X"2C",X"2C",X"2C",X"2C",X"7E",X"A7",X"CA",X"BE",X"35",X"35",X"EB",X"D5",
		X"78",X"07",X"07",X"07",X"6F",X"26",X"3F",X"46",X"23",X"4E",X"C5",X"23",X"46",X"23",X"4E",X"C5",
		X"23",X"46",X"23",X"4E",X"C5",X"23",X"46",X"23",X"4E",X"C5",X"EB",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"2C",X"2C",X"7E",X"FE",X"10",X"D2",X"28",X"36",X"47",X"2D",X"86",X"77",X"2D",X"2D",X"78",X"86",
		X"77",X"FE",X"08",X"DA",X"6A",X"36",X"E6",X"07",X"77",X"2D",X"7E",X"D6",X"20",X"77",X"D2",X"04",
		X"36",X"2D",X"35",X"2C",X"2C",X"2C",X"2C",X"4E",X"2C",X"2C",X"7E",X"2D",X"36",X"10",X"91",X"CA",
		X"72",X"36",X"3D",X"0F",X"0F",X"0F",X"E6",X"1F",X"B8",X"3C",X"77",X"D8",X"3A",X"6E",X"43",X"77",
		X"B8",X"C8",X"04",X"70",X"C9",X"FF",X"FF",X"FF",X"E6",X"0F",X"CA",X"44",X"37",X"47",X"2D",X"7E",
		X"90",X"77",X"2D",X"2D",X"7E",X"90",X"77",X"D2",X"95",X"36",X"E6",X"07",X"77",X"2D",X"7E",X"C6",
		X"20",X"77",X"D2",X"48",X"36",X"2D",X"34",X"2C",X"2C",X"2C",X"2C",X"7E",X"2C",X"2C",X"96",X"0F",
		X"0F",X"0F",X"E6",X"1F",X"B8",X"3C",X"2D",X"DA",X"63",X"36",X"3A",X"6E",X"43",X"B8",X"CA",X"63",
		X"36",X"78",X"3C",X"F6",X"10",X"77",X"C9",X"77",X"C9",X"FF",X"78",X"A7",X"C0",X"2C",X"2C",X"2C",
		X"34",X"C9",X"2D",X"46",X"2C",X"2C",X"3A",X"C2",X"43",X"E6",X"F8",X"B8",X"D2",X"80",X"36",X"47",
		X"3A",X"6D",X"43",X"4F",X"C6",X"08",X"32",X"6D",X"43",X"78",X"91",X"36",X"08",X"D8",X"FE",X"08",
		X"D8",X"77",X"C9",X"D8",X"FE",X"2C",X"2C",X"46",X"2C",X"2C",X"7E",X"B8",X"C0",X"2D",X"36",X"00",
		X"2C",X"3A",X"C2",X"43",X"E6",X"F8",X"B8",X"DA",X"AB",X"36",X"47",X"3A",X"6D",X"43",X"C6",X"08",
		X"32",X"6D",X"43",X"80",X"36",X"C8",X"D8",X"FE",X"C8",X"D0",X"77",X"C9",X"77",X"C9",X"FF",X"FF",
		X"7E",X"0F",X"D8",X"2D",X"7E",X"3C",X"E6",X"07",X"77",X"C9",X"FF",X"FF",X"D1",X"C1",X"E1",X"C9",
		X"FF",X"FF",X"D1",X"C1",X"E1",X"7E",X"A7",X"C0",X"70",X"2D",X"2D",X"2D",X"2D",X"72",X"3A",X"68",
		X"43",X"F6",X"01",X"32",X"68",X"43",X"C9",X"FF",X"FF",X"FF",X"D1",X"C1",X"E1",X"7E",X"A7",X"C0",
		X"2C",X"2C",X"7E",X"E6",X"0F",X"C0",X"2D",X"2D",X"70",X"2D",X"2D",X"2D",X"2D",X"72",X"3A",X"68",
		X"43",X"F6",X"02",X"32",X"68",X"43",X"C9",X"FF",X"FF",X"FF",X"D1",X"C1",X"E1",X"7E",X"A7",X"C0",
		X"2C",X"2C",X"7E",X"E6",X"0F",X"C0",X"2D",X"2D",X"70",X"2D",X"2D",X"2D",X"2D",X"72",X"3A",X"68",
		X"43",X"F6",X"04",X"32",X"68",X"43",X"3A",X"6F",X"43",X"A3",X"E6",X"F0",X"C0",X"7B",X"E6",X"0F",
		X"77",X"2C",X"2C",X"2C",X"2C",X"71",X"3A",X"68",X"43",X"F6",X"08",X"32",X"68",X"43",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"36",X"11",X"2D",X"35",X"2D",X"2D",X"36",X"07",X"2D",X"7E",X"C6",X"20",
		X"77",X"D0",X"2D",X"34",X"C9",X"FF",X"FF",X"FF",X"21",X"9B",X"43",X"7E",X"07",X"07",X"07",X"E6",
		X"07",X"2E",X"C2",X"86",X"E6",X"0F",X"C9",X"E6",X"0E",X"07",X"D1",X"C1",X"E1",X"7E",X"A7",X"C0",
		X"2C",X"2C",X"7E",X"E6",X"10",X"C2",X"83",X"37",X"2D",X"2D",X"70",X"2D",X"2D",X"2D",X"2D",X"72",
		X"C9",X"FF",X"FF",X"2D",X"2D",X"71",X"2D",X"2D",X"2D",X"2D",X"7B",X"E6",X"0F",X"77",X"C9",X"FF",
		X"21",X"9B",X"43",X"7E",X"0F",X"D8",X"E6",X"03",X"07",X"07",X"C6",X"C0",X"6F",X"26",X"37",X"56",
		X"23",X"4E",X"23",X"7E",X"23",X"6E",X"67",X"06",X"00",X"7E",X"E6",X"FC",X"FE",X"78",X"C2",X"B6",
		X"37",X"7E",X"3C",X"E6",X"FB",X"77",X"09",X"15",X"C2",X"A9",X"37",X"C3",X"BC",X"33",X"FF",X"FF",
		X"08",X"1F",X"48",X"07",X"08",X"21",X"4A",X"40",X"04",X"1F",X"49",X"1F",X"04",X"21",X"49",X"DC",
		X"3A",X"92",X"43",X"E6",X"0C",X"0F",X"C6",X"F8",X"6F",X"26",X"33",X"7E",X"32",X"E7",X"49",X"32",
		X"67",X"49",X"2C",X"56",X"21",X"6A",X"41",X"01",X"20",X"00",X"1E",X"05",X"3A",X"BC",X"43",X"70",
		X"0F",X"DA",X"F5",X"37",X"72",X"09",X"1D",X"C2",X"EF",X"37",X"C9",X"34",X"62",X"32",X"61",X"34",
		X"3A",X"C4",X"43",X"E6",X"08",X"C8",X"3A",X"E6",X"43",X"C6",X"08",X"57",X"3A",X"D2",X"4B",X"5F",
		X"3A",X"E7",X"43",X"E6",X"E0",X"47",X"3A",X"E7",X"43",X"93",X"00",X"E6",X"1F",X"B0",X"5F",X"1A",
		X"D6",X"90",X"D8",X"47",X"3A",X"C6",X"43",X"E6",X"07",X"C6",X"00",X"6F",X"26",X"3E",X"4E",X"7B",
		X"E6",X"0E",X"07",X"07",X"5F",X"3E",X"A8",X"93",X"5F",X"16",X"4B",X"78",X"FE",X"40",X"DC",X"44",
		X"38",X"C3",X"BA",X"38",X"C6",X"60",X"6F",X"26",X"3B",X"7E",X"A1",X"C8",X"CD",X"A1",X"38",X"EB",
		X"7E",X"36",X"00",X"2C",X"2C",X"2C",X"2C",X"56",X"E1",X"21",X"BB",X"43",X"35",X"FE",X"08",X"DA",
		X"80",X"38",X"5F",X"3E",X"FF",X"32",X"69",X"43",X"01",X"10",X"1F",X"7B",X"FE",X"0D",X"DA",X"FA",
		X"38",X"0E",X"20",X"FE",X"0F",X"C2",X"FA",X"38",X"0E",X"40",X"C3",X"FA",X"38",X"0E",X"CA",X"FB",
		X"01",X"05",X"39",X"3E",X"FF",X"32",X"64",X"43",X"C3",X"FA",X"38",X"C3",X"52",X"05",X"FF",X"FF",
		X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0E",X"0F",
		X"FF",X"D5",X"0E",X"20",X"EB",X"23",X"56",X"23",X"5E",X"3A",X"87",X"19",X"C6",X"E2",X"6F",X"26",
		X"17",X"CD",X"DE",X"34",X"D1",X"C9",X"35",X"D1",X"C9",X"FF",X"78",X"FE",X"10",X"D8",X"C6",X"90",
		X"6F",X"26",X"3B",X"7E",X"A1",X"C8",X"CD",X"A1",X"38",X"1A",X"D6",X"08",X"DA",X"EA",X"38",X"47",
		X"62",X"7B",X"C6",X"05",X"6F",X"3A",X"C6",X"43",X"BE",X"17",X"07",X"07",X"07",X"E6",X"08",X"B0",
		X"C6",X"90",X"6F",X"26",X"38",X"46",X"EB",X"CD",X"E0",X"3C",X"3E",X"FF",X"32",X"66",X"43",X"01",
		X"02",X"53",X"C3",X"FA",X"38",X"53",X"C3",X"FA",X"38",X"FF",X"CD",X"14",X"39",X"70",X"2C",X"71",
		X"2C",X"3A",X"E6",X"43",X"77",X"2C",X"3A",X"E7",X"43",X"77",X"3A",X"C4",X"43",X"E6",X"F7",X"32",
		X"C4",X"43",X"C9",X"FF",X"21",X"70",X"43",X"7E",X"E6",X"1F",X"C8",X"2C",X"2C",X"2C",X"2C",X"7E",
		X"E6",X"1F",X"C8",X"2C",X"2C",X"2C",X"2C",X"7E",X"E6",X"1F",X"C8",X"2C",X"2C",X"2C",X"2C",X"C9",
		X"3A",X"D2",X"4B",X"E6",X"1E",X"C6",X"C0",X"6F",X"26",X"3D",X"5E",X"2C",X"6E",X"26",X"4B",X"CD",
		X"00",X"3A",X"3A",X"9F",X"43",X"82",X"4F",X"3A",X"9E",X"43",X"92",X"47",X"E5",X"CD",X"5C",X"39",
		X"E1",X"7D",X"C6",X"08",X"6F",X"1D",X"C2",X"4C",X"39",X"C9",X"FF",X"FF",X"7E",X"FE",X"05",X"D8",
		X"7D",X"C6",X"05",X"6F",X"7E",X"B8",X"D8",X"B9",X"D0",X"D6",X"04",X"47",X"2D",X"2D",X"2D",X"3A",
		X"D2",X"4B",X"86",X"E6",X"1F",X"07",X"07",X"07",X"C6",X"08",X"4F",X"C3",X"B7",X"25",X"FF",X"FF",
		X"3A",X"D2",X"4B",X"D6",X"0C",X"D8",X"FE",X"10",X"D0",X"21",X"C4",X"43",X"11",X"C0",X"4B",X"06",
		X"04",X"CD",X"E0",X"05",X"2E",X"E6",X"06",X"02",X"CD",X"E0",X"05",X"2E",X"E2",X"11",X"E6",X"43",
		X"06",X"02",X"CD",X"E0",X"05",X"2E",X"C4",X"36",X"08",X"11",X"9E",X"43",X"3A",X"9B",X"43",X"0F",
		X"DA",X"BF",X"39",X"1C",X"2E",X"E7",X"7E",X"D6",X"20",X"77",X"2D",X"7E",X"DE",X"00",X"77",X"1A",
		X"32",X"C6",X"43",X"CD",X"00",X"38",X"21",X"C4",X"43",X"7E",X"E6",X"08",X"CA",X"F0",X"39",X"21",
		X"E7",X"43",X"34",X"7E",X"E6",X"1F",X"FE",X"1D",X"DA",X"C3",X"39",X"21",X"C0",X"4B",X"11",X"C4",
		X"43",X"06",X"04",X"CD",X"E0",X"05",X"1E",X"E6",X"06",X"02",X"C3",X"E0",X"05",X"FF",X"FF",X"FF",
		X"2E",X"A6",X"7E",X"FE",X"C0",X"DA",X"C4",X"0C",X"D6",X"01",X"77",X"C3",X"DB",X"39",X"FF",X"FF",
		X"3A",X"BB",X"43",X"D6",X"0C",X"2F",X"3C",X"57",X"3A",X"9B",X"43",X"0F",X"0F",X"D8",X"E1",X"C9",
		X"21",X"B8",X"11",X"8C",X"43",X"CD",X"2A",X"3A",X"CD",X"48",X"3A",X"21",X"66",X"43",X"7E",X"A7",
		X"C8",X"36",X"00",X"1A",X"F6",X"40",X"12",X"C9",X"FF",X"FF",X"21",X"69",X"43",X"7E",X"A7",X"C8",
		X"E6",X"3F",X"3D",X"77",X"0F",X"0F",X"0F",X"00",X"E6",X"07",X"47",X"7E",X"0F",X"E6",X"03",X"80",
		X"47",X"1A",X"E6",X"F0",X"B0",X"12",X"C9",X"FF",X"21",X"64",X"43",X"7E",X"A7",X"C8",X"E6",X"1F",
		X"3D",X"77",X"0F",X"0F",X"2F",X"E6",X"07",X"47",X"7E",X"07",X"E6",X"06",X"80",X"47",X"1A",X"E6",
		X"F0",X"B0",X"12",X"C9",X"8C",X"77",X"C9",X"FE",X"10",X"DA",X"78",X"3A",X"36",X"10",X"3A",X"B8",
		X"3A",X"A4",X"43",X"FE",X"03",X"C2",X"BD",X"27",X"3A",X"B8",X"43",X"E6",X"07",X"07",X"C6",X"8A",
		X"6F",X"26",X"3A",X"7E",X"2C",X"6E",X"67",X"E9",X"C9",X"FF",X"3A",X"88",X"27",X"E6",X"3A",X"9A",
		X"3A",X"D0",X"3A",X"88",X"27",X"E6",X"3A",X"B4",X"3A",X"E8",X"21",X"8C",X"43",X"36",X"AF",X"3A",
		X"B9",X"43",X"FE",X"FD",X"D0",X"36",X"BF",X"E6",X"07",X"C8",X"36",X"7F",X"E6",X"01",X"C8",X"36",
		X"3F",X"C9",X"21",X"2F",X"3A",X"9A",X"43",X"FE",X"02",X"D0",X"E6",X"0F",X"67",X"3A",X"9B",X"43",
		X"E6",X"FC",X"6F",X"7E",X"E6",X"01",X"C8",X"3E",X"0D",X"32",X"8C",X"43",X"C9",X"FF",X"FF",X"FF",
		X"3A",X"BB",X"43",X"A7",X"C8",X"21",X"8C",X"43",X"36",X"3F",X"3A",X"B9",X"43",X"FE",X"F0",X"D8",
		X"E6",X"07",X"C0",X"36",X"2F",X"C9",X"C9",X"F7",X"CD",X"B4",X"3A",X"3A",X"95",X"43",X"A7",X"CA",
		X"E0",X"3D",X"3A",X"9C",X"43",X"E6",X"7C",X"C8",X"0F",X"0F",X"32",X"8D",X"43",X"C9",X"77",X"C9",
		X"06",X"00",X"21",X"B8",X"43",X"7E",X"E6",X"0E",X"FE",X"00",X"C8",X"06",X"40",X"FE",X"06",X"C8",
		X"06",X"80",X"C9",X"06",X"80",X"C9",X"80",X"B6",X"77",X"C9",X"78",X"21",X"62",X"43",X"7E",X"A7",
		X"C8",X"3D",X"E6",X"3F",X"77",X"07",X"00",X"E6",X"0C",X"47",X"2E",X"8D",X"7E",X"E6",X"F0",X"B0",
		X"77",X"C9",X"C9",X"21",X"6A",X"43",X"7E",X"A7",X"C8",X"35",X"E6",X"08",X"F6",X"07",X"2E",X"8D",
		X"77",X"C9",X"8D",X"CD",X"70",X"3A",X"CD",X"33",X"3B",X"CD",X"1B",X"3B",X"CD",X"12",X"3A",X"CD",
		X"D2",X"27",X"CD",X"00",X"3B",X"2E",X"8D",X"7E",X"E6",X"3F",X"B0",X"77",X"C9",X"3A",X"FF",X"FF",
		X"FE",X"F8",X"0F",X"3F",X"FF",X"FE",X"3F",X"F8",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"E0",X"3F",X"F8",X"0F",X"F8",X"0F",X"FC",X"07",X"FC",X"07",X"FC",X"F8",X"0F",X"F8",X"0F",
		X"F8",X"0F",X"F8",X"0F",X"E0",X"3F",X"E0",X"3F",X"E0",X"3F",X"E0",X"3F",X"FF",X"80",X"FF",X"FF",
		X"80",X"FF",X"FE",X"03",X"FE",X"03",X"FE",X"03",X"FE",X"03",X"07",X"07",X"00",X"00",X"00",X"00",
		X"F0",X"1F",X"C0",X"07",X"F0",X"07",X"F0",X"03",X"F8",X"03",X"F8",X"03",X"07",X"F0",X"07",X"F0",
		X"07",X"F0",X"07",X"F0",X"1F",X"C0",X"1F",X"C0",X"1F",X"C0",X"1F",X"C0",X"00",X"7F",X"00",X"00",
		X"7F",X"00",X"01",X"FC",X"01",X"FC",X"01",X"FC",X"01",X"FC",X"F8",X"F8",X"FF",X"FF",X"00",X"00",
		X"3F",X"FF",X"3F",X"FF",X"FC",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"7F",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F8",X"FF",X"FF",X"7F",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"1F",X"00",X"80",X"E0",X"F8",X"FE",X"03",X"0F",X"3F",X"FF",
		X"00",X"E0",X"F9",X"E1",X"AC",X"AE",X"AD",X"AF",X"00",X"E2",X"00",X"FD",X"00",X"00",X"00",X"E7",
		X"F8",X"FF",X"B4",X"B6",X"B5",X"B7",X"00",X"E8",X"00",X"FE",X"00",X"00",X"FA",X"00",X"FC",X"EC",
		X"FB",X"BD",X"BC",X"BE",X"00",X"ED",X"00",X"EE",X"00",X"00",X"F9",X"00",X"FD",X"F2",X"FA",X"F3",
		X"C2",X"C4",X"C3",X"C5",X"00",X"DF",X"00",X"FC",X"00",X"FB",X"00",X"F5",X"C6",X"C8",X"C7",X"C9",
		X"00",X"FF",X"00",X"F6",X"00",X"00",X"00",X"E3",X"00",X"E4",X"B0",X"B2",X"B1",X"B3",X"FC",X"E5",
		X"00",X"E6",X"00",X"00",X"00",X"F9",X"00",X"E9",X"B8",X"BA",X"B9",X"BB",X"FD",X"EA",X"00",X"EB",
		X"00",X"00",X"00",X"F8",X"00",X"EF",X"F8",X"C0",X"BF",X"C1",X"FE",X"F0",X"F8",X"F1",X"FC",X"00",
		X"00",X"DC",X"00",X"DD",X"A7",X"A9",X"CA",X"AA",X"CC",X"D1",X"D0",X"F4",X"00",X"DC",X"00",X"DD",
		X"A7",X"AB",X"CB",X"AA",X"CD",X"D3",X"D2",X"F4",X"D4",X"DC",X"D5",X"D8",X"A7",X"A9",X"A8",X"AA",
		X"00",X"DE",X"00",X"F4",X"D6",X"DC",X"D7",X"D9",X"A7",X"AB",X"A8",X"AA",X"00",X"DE",X"00",X"F4",
		X"D4",X"DC",X"D5",X"D8",X"A7",X"A9",X"CB",X"AA",X"CD",X"D3",X"D2",X"F4",X"D6",X"DC",X"D7",X"D9",
		X"A7",X"AB",X"CA",X"AA",X"CC",X"D1",X"D0",X"F4",X"00",X"DC",X"00",X"DD",X"A7",X"A9",X"A8",X"AA",
		X"00",X"DE",X"00",X"F4",X"00",X"E3",X"00",X"E4",X"B0",X"B2",X"AD",X"AF",X"00",X"E2",X"00",X"FD",
		X"00",X"E0",X"F9",X"E1",X"AC",X"AE",X"B1",X"B3",X"FC",X"E5",X"00",X"E6",X"B8",X"BB",X"B9",X"BC",
		X"7D",X"C6",X"05",X"6F",X"7E",X"E6",X"F8",X"2C",X"2C",X"BE",X"C8",X"2D",X"7E",X"E6",X"F0",X"77",
		X"2D",X"7E",X"E6",X"F8",X"77",X"2D",X"36",X"80",X"2D",X"36",X"00",X"2D",X"2D",X"2D",X"70",X"C9",
		X"00",X"00",X"00",X"00",X"90",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"91",X"00",X"92",X"00",
		X"00",X"00",X"00",X"00",X"F9",X"00",X"93",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"94",X"00",
		X"00",X"00",X"00",X"00",X"95",X"00",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"00",
		X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"00",X"99",X"00",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"00",X"9A",X"00",X"9B",X"00",X"00",X"00",X"FB",X"00",X"9C",X"00",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"FA",X"00",X"9D",X"00",X"9E",X"00",X"00",X"00",X"00",X"00",X"F9",X"00",
		X"9F",X"00",X"A0",X"00",X"FC",X"00",X"00",X"00",X"F8",X"00",X"A1",X"00",X"A2",X"00",X"FD",X"00",
		X"00",X"00",X"00",X"DA",X"A3",X"A5",X"A4",X"A6",X"00",X"DB",X"00",X"00",X"21",X"D0",X"4B",X"7E",
		X"FE",X"03",X"2E",X"E3",X"C2",X"89",X"3D",X"36",X"10",X"7E",X"A7",X"C8",X"35",X"2F",X"00",X"E6",
		X"0F",X"F6",X"10",X"32",X"8D",X"43",X"E1",X"C9",X"21",X"70",X"4B",X"01",X"00",X"00",X"11",X"08",
		X"08",X"7E",X"2C",X"A2",X"CA",X"AF",X"3D",X"04",X"7E",X"FE",X"30",X"D2",X"AF",X"3D",X"4F",X"2C",
		X"2C",X"2C",X"1D",X"C2",X"A1",X"3D",X"C9",X"00",X"0C",X"0C",X"0E",X"FF",X"0D",X"0E",X"0D",X"FF",
		X"06",X"70",X"07",X"70",X"08",X"70",X"07",X"78",X"06",X"80",X"05",X"88",X"04",X"90",X"03",X"98",
		X"02",X"A0",X"01",X"A8",X"01",X"70",X"01",X"70",X"02",X"70",X"03",X"70",X"04",X"70",X"05",X"70",
		X"21",X"8D",X"43",X"36",X"3F",X"3A",X"B9",X"43",X"FE",X"FC",X"D0",X"36",X"2F",X"E6",X"01",X"C8",
		X"2D",X"7E",X"F6",X"40",X"77",X"C9",X"05",X"04",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"3D",X"00",X"3D",X"08",X"3D",X"10",X"3D",X"18",
		X"3D",X"20",X"3D",X"2A",X"3D",X"34",X"3D",X"3E",X"3D",X"48",X"3D",X"52",X"3D",X"5C",X"3D",X"66",
		X"3D",X"48",X"3D",X"52",X"3D",X"5C",X"3D",X"70",X"3D",X"70",X"3D",X"70",X"3C",X"B8",X"3C",X"B8",
		X"3D",X"70",X"3D",X"5C",X"3D",X"52",X"3D",X"48",X"3C",X"B8",X"3C",X"B8",X"3D",X"70",X"3D",X"70",
		X"3C",X"B8",X"3C",X"C4",X"3C",X"B8",X"3C",X"D0",X"3C",X"46",X"3C",X"B8",X"3C",X"B8",X"3C",X"00",
		X"3C",X"00",X"3C",X"B8",X"3C",X"B8",X"3C",X"46",X"3C",X"00",X"3C",X"0E",X"3C",X"1C",X"3C",X"2A",
		X"3C",X"38",X"3C",X"46",X"3C",X"54",X"3C",X"62",X"3C",X"70",X"3C",X"70",X"3C",X"7C",X"3C",X"7C",
		X"3C",X"88",X"3C",X"88",X"3C",X"94",X"3C",X"94",X"3C",X"A0",X"3C",X"A0",X"3C",X"AC",X"3C",X"AC",
		X"04",X"40",X"03",X"20",X"02",X"30",X"02",X"10",X"05",X"48",X"04",X"28",X"03",X"38",X"02",X"18",
		X"06",X"50",X"05",X"30",X"04",X"40",X"03",X"20",X"07",X"58",X"06",X"38",X"05",X"48",X"04",X"28",
		X"05",X"10",X"04",X"20",X"03",X"30",X"03",X"40",X"06",X"18",X"05",X"28",X"04",X"38",X"03",X"48",
		X"07",X"20",X"06",X"30",X"05",X"40",X"04",X"50",X"08",X"30",X"07",X"40",X"06",X"50",X"05",X"60",
		X"FF",X"38",X"30",X"30",X"30",X"28",X"30",X"28",X"28",X"28",X"28",X"20",X"20",X"28",X"28",X"28",
		X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"01",
		X"14",X"15",X"16",X"10",X"08",X"04",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"04",
		X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"FF",X"02",X"FF",X"36",X"D2",X"35",X"E0",
		X"30",X"FF",X"03",X"FF",X"36",X"D2",X"35",X"E0",X"10",X"FF",X"04",X"FF",X"36",X"EA",X"35",X"E0",
		X"10",X"FF",X"05",X"FF",X"36",X"EA",X"36",X"C0",X"10",X"FF",X"08",X"FF",X"36",X"EA",X"36",X"C0",
		X"30",X"FF",X"03",X"FF",X"36",X"EA",X"36",X"C0",X"10",X"FF",X"06",X"FF",X"36",X"EA",X"36",X"C0",
		X"10",X"10",X"09",X"1A",X"37",X"6A",X"36",X"C0",X"10",X"10",X"0B",X"38",X"37",X"0A",X"36",X"C0",
		X"10",X"10",X"0C",X"38",X"37",X"0A",X"36",X"C0",X"10",X"10",X"0A",X"77",X"37",X"0A",X"35",X"E0",
		X"10",X"10",X"09",X"77",X"37",X"0A",X"35",X"E0",X"10",X"FF",X"08",X"FF",X"36",X"D2",X"36",X"C0",
		X"10",X"FF",X"08",X"FF",X"36",X"D2",X"36",X"C0",X"10",X"FF",X"08",X"FF",X"36",X"D2",X"36",X"C0",
		X"01",X"48",X"6E",X"00",X"10",X"D0",X"10",X"10",X"01",X"4A",X"8C",X"00",X"20",X"48",X"00",X"B8",
		X"01",X"4A",X"2A",X"00",X"30",X"60",X"10",X"28",X"01",X"49",X"68",X"00",X"40",X"90",X"00",X"B0",
		X"01",X"4A",X"E6",X"00",X"50",X"30",X"00",X"60",X"01",X"4A",X"84",X"00",X"60",X"48",X"00",X"A0",
		X"01",X"48",X"C2",X"00",X"70",X"B8",X"10",X"80",X"01",X"49",X"40",X"00",X"80",X"98",X"10",X"40",
		X"01",X"4B",X"2E",X"00",X"10",X"20",X"00",X"40",X"01",X"48",X"6C",X"00",X"20",X"D0",X"10",X"70",
		X"01",X"4A",X"CA",X"00",X"30",X"38",X"00",X"58",X"01",X"48",X"C8",X"00",X"40",X"B8",X"10",X"58",
		X"01",X"4A",X"66",X"00",X"50",X"50",X"00",X"70",X"01",X"49",X"24",X"00",X"60",X"A0",X"10",X"40",
		X"01",X"4A",X"02",X"00",X"70",X"68",X"00",X"88",X"01",X"49",X"80",X"00",X"80",X"88",X"10",X"28");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
