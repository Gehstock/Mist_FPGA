library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_pgm_rom2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_pgm_rom2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"01",X"01",X"01",X"11",X"CB",X"9B",X"17",X"01",X"01",X"01",X"11",X"C1",X"9B",X"07",X"01",
		X"01",X"01",X"11",X"D4",X"9B",X"01",X"01",X"01",X"01",X"11",X"C1",X"9B",X"0D",X"01",X"01",X"01",
		X"11",X"D2",X"9B",X"05",X"01",X"01",X"01",X"11",X"C9",X"9B",X"13",X"01",X"01",X"01",X"11",X"A9",
		X"00",X"AA",X"20",X"5B",X"D8",X"A9",X"5A",X"AA",X"A9",X"2F",X"20",X"E3",X"D7",X"A0",X"60",X"A9",
		X"01",X"20",X"12",X"D8",X"A9",X"00",X"A2",X"00",X"20",X"5B",X"D8",X"A9",X"00",X"38",X"20",X"AF",
		X"D7",X"A0",X"00",X"A9",X"01",X"20",X"12",X"D8",X"20",X"C9",X"D8",X"60",X"A0",X"00",X"B1",X"4C",
		X"91",X"49",X"C8",X"CA",X"D0",X"F8",X"60",X"A4",X"03",X"08",X"A9",X"00",X"A0",X"08",X"46",X"03",
		X"90",X"03",X"18",X"65",X"02",X"6A",X"66",X"01",X"88",X"D0",X"F3",X"28",X"10",X"03",X"38",X"E5",
		X"02",X"60",X"A2",X"0F",X"A0",X"00",X"B1",X"4C",X"91",X"49",X"C8",X"C0",X"10",X"D0",X"F7",X"A5",
		X"49",X"18",X"6D",X"35",X"04",X"85",X"49",X"90",X"02",X"E6",X"4A",X"CA",X"D0",X"E6",X"60",X"A5",
		X"4D",X"30",X"12",X"A5",X"4A",X"30",X"1D",X"A5",X"4C",X"38",X"E5",X"49",X"A5",X"4D",X"E5",X"4A",
		X"10",X"12",X"A9",X"FF",X"60",X"A5",X"4A",X"10",X"F9",X"A5",X"49",X"38",X"E5",X"4C",X"A5",X"4A",
		X"E5",X"4D",X"30",X"EE",X"A9",X"00",X"60",X"A2",X"00",X"A5",X"5E",X"D0",X"01",X"60",X"4A",X"B0",
		X"05",X"E8",X"E8",X"4C",X"CE",X"A0",X"BD",X"E0",X"A0",X"48",X"BD",X"DF",X"A0",X"48",X"60",X"EE",
		X"A0",X"F9",X"A1",X"3C",X"A2",X"72",X"A1",X"64",X"A2",X"65",X"A2",X"66",X"A2",X"67",X"A2",X"A5",
		X"6F",X"29",X"03",X"D0",X"E9",X"A5",X"74",X"85",X"49",X"A5",X"75",X"85",X"4A",X"A9",X"08",X"85",
		X"4C",X"A6",X"4B",X"8A",X"29",X"10",X"D0",X"0D",X"8A",X"29",X"07",X"AA",X"BD",X"6B",X"A1",X"8D",
		X"00",X"25",X"4C",X"3C",X"A1",X"A9",X"A1",X"20",X"5B",X"A1",X"A5",X"49",X"18",X"69",X"4E",X"85",
		X"49",X"A5",X"4A",X"69",X"00",X"85",X"4A",X"E8",X"8A",X"29",X"07",X"AA",X"C6",X"4C",X"D0",X"E5",
		X"A9",X"A1",X"8D",X"00",X"25",X"A5",X"5E",X"29",X"FE",X"85",X"5E",X"60",X"BD",X"6B",X"A1",X"20",
		X"5B",X"A1",X"A5",X"49",X"18",X"69",X"4E",X"85",X"49",X"A5",X"4A",X"69",X"00",X"85",X"4A",X"E8",
		X"8A",X"29",X"07",X"AA",X"C6",X"4C",X"D0",X"E4",X"E6",X"4B",X"60",X"A0",X"04",X"91",X"49",X"48",
		X"98",X"18",X"69",X"06",X"A8",X"68",X"C0",X"4C",X"D0",X"F3",X"60",X"E1",X"E2",X"E3",X"E4",X"E5",
		X"E6",X"E7",X"E4",X"A9",X"0B",X"85",X"19",X"A6",X"19",X"BD",X"29",X"04",X"F0",X"16",X"20",X"CA",
		X"A1",X"BD",X"29",X"04",X"29",X"C0",X"4A",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"B9",X"A2",X"A1",
		X"A0",X"00",X"91",X"49",X"C6",X"19",X"10",X"DF",X"A9",X"00",X"8D",X"01",X"03",X"A9",X"00",X"85",
		X"5E",X"60",X"01",X"02",X"04",X"04",X"04",X"0A",X"10",X"16",X"1C",X"22",X"28",X"2E",X"34",X"3A",
		X"40",X"46",X"00",X"00",X"4E",X"00",X"9C",X"00",X"EA",X"00",X"38",X"01",X"86",X"01",X"D4",X"01",
		X"22",X"02",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"A0",X"00",X"29",X"3F",X"F0",X"06",
		X"C8",X"38",X"E9",X"06",X"D0",X"FA",X"98",X"48",X"0A",X"A8",X"B9",X"B2",X"A1",X"18",X"7D",X"A6",
		X"A1",X"85",X"49",X"A9",X"00",X"79",X"B3",X"A1",X"85",X"4A",X"18",X"A5",X"74",X"65",X"49",X"85",
		X"49",X"A5",X"75",X"65",X"4A",X"85",X"4A",X"68",X"A8",X"60",X"A5",X"6F",X"29",X"02",X"D0",X"F9",
		X"E6",X"A5",X"A5",X"A5",X"29",X"0F",X"D0",X"05",X"A9",X"0D",X"85",X"5E",X"60",X"85",X"1D",X"A9",
		X"00",X"85",X"1B",X"85",X"1E",X"A9",X"00",X"85",X"1C",X"A6",X"1B",X"A4",X"1C",X"20",X"D6",X"A1",
		X"A0",X"00",X"A5",X"1D",X"29",X"07",X"09",X"E0",X"91",X"49",X"E6",X"1C",X"A5",X"1C",X"29",X"07",
		X"D0",X"E7",X"E6",X"1D",X"E6",X"1B",X"A5",X"1B",X"C9",X"0C",X"90",X"D9",X"60",X"AD",X"5D",X"04",
		X"C9",X"0C",X"90",X"06",X"38",X"E9",X"0C",X"4C",X"40",X"A2",X"0A",X"0A",X"85",X"19",X"0A",X"65",
		X"19",X"A8",X"A2",X"00",X"B9",X"17",X"B8",X"9D",X"29",X"04",X"C8",X"E8",X"E0",X"0C",X"D0",X"F4",
		X"A9",X"08",X"85",X"5E",X"60",X"60",X"60",X"60",X"60",X"98",X"10",X"0E",X"49",X"FF",X"18",X"69",
		X"01",X"20",X"7A",X"A2",X"49",X"FF",X"18",X"69",X"01",X"60",X"A8",X"8A",X"10",X"10",X"49",X"FF",
		X"18",X"69",X"01",X"20",X"8E",X"A2",X"49",X"20",X"49",X"FF",X"18",X"69",X"01",X"60",X"85",X"1A",
		X"98",X"C5",X"1A",X"F0",X"2F",X"90",X"11",X"A4",X"1A",X"85",X"1A",X"98",X"20",X"A8",X"A2",X"38",
		X"E9",X"10",X"49",X"FF",X"18",X"69",X"01",X"60",X"A0",X"00",X"84",X"19",X"A0",X"04",X"26",X"19",
		X"2A",X"C5",X"1A",X"90",X"02",X"E5",X"1A",X"88",X"D0",X"F4",X"A5",X"19",X"2A",X"29",X"0F",X"AA",
		X"BD",X"C7",X"A2",X"60",X"A9",X"08",X"60",X"00",X"01",X"02",X"02",X"02",X"03",X"04",X"04",X"05",
		X"05",X"06",X"06",X"06",X"07",X"07",X"07",X"6B",X"00",X"BD",X"01",X"02",X"A8",X"29",X"20",X"F0",
		X"14",X"98",X"38",X"E9",X"40",X"A8",X"29",X"C0",X"F0",X"05",X"98",X"9D",X"01",X"02",X"60",X"98",
		X"29",X"1F",X"4C",X"EB",X"A2",X"98",X"18",X"69",X"40",X"A8",X"29",X"C0",X"C9",X"C0",X"D0",X"EA",
		X"98",X"29",X"1F",X"09",X"60",X"A8",X"29",X"0F",X"C9",X"04",X"D0",X"DE",X"98",X"29",X"1F",X"4C",
		X"EB",X"A2",X"E0",X"00",X"D0",X"05",X"A5",X"71",X"4C",X"1E",X"A3",X"BD",X"06",X"02",X"18",X"69",
		X"02",X"4A",X"4A",X"29",X"0F",X"85",X"19",X"BD",X"01",X"02",X"85",X"1A",X"29",X"0F",X"C9",X"03",
		X"F0",X"0F",X"48",X"A9",X"00",X"9D",X"0A",X"21",X"A9",X"71",X"9D",X"0B",X"21",X"68",X"4C",X"59",
		X"A3",X"BD",X"02",X"02",X"D0",X"09",X"A5",X"1A",X"29",X"F0",X"09",X"02",X"4C",X"55",X"A3",X"A5",
		X"1A",X"29",X"F0",X"09",X"06",X"85",X"1A",X"29",X"0F",X"C9",X"05",X"D0",X"04",X"A9",X"50",X"D0",
		X"21",X"C9",X"0B",X"F0",X"13",X"C9",X"04",X"D0",X"13",X"A5",X"1A",X"29",X"C0",X"4A",X"4A",X"4A",
		X"4A",X"4A",X"4A",X"09",X"40",X"4C",X"82",X"A3",X"A0",X"00",X"84",X"19",X"0A",X"0A",X"0A",X"0A",
		X"05",X"19",X"9D",X"04",X"21",X"A9",X"A4",X"9D",X"05",X"21",X"06",X"19",X"A5",X"1A",X"29",X"C0",
		X"4A",X"05",X"19",X"85",X"19",X"A5",X"1A",X"29",X"0F",X"0A",X"A8",X"B9",X"B3",X"A3",X"30",X"11",
		X"B9",X"B2",X"A3",X"05",X"19",X"9D",X"08",X"21",X"B9",X"B3",X"A3",X"18",X"69",X"A5",X"9D",X"09",
		X"21",X"60",X"00",X"01",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"80",X"01",
		X"80",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"FF",X"FF",X"00",X"01",X"00",X"02",X"80",X"01",
		X"00",X"02",X"A2",X"00",X"A0",X"00",X"BD",X"00",X"02",X"29",X"03",X"C9",X"02",X"90",X"5B",X"C9",
		X"03",X"F0",X"0C",X"E0",X"00",X"F0",X"03",X"4C",X"5C",X"A5",X"A9",X"00",X"4C",X"3A",X"A4",X"A9",
		X"00",X"99",X"00",X"22",X"99",X"01",X"22",X"99",X"02",X"22",X"99",X"03",X"22",X"9D",X"09",X"02",
		X"9D",X"0A",X"02",X"9D",X"0B",X"02",X"9D",X"0C",X"02",X"A9",X"60",X"9D",X"07",X"21",X"A9",X"00",
		X"9D",X"00",X"21",X"9D",X"06",X"21",X"A9",X"A4",X"9D",X"05",X"21",X"A9",X"AF",X"9D",X"09",X"21",
		X"A9",X"00",X"9D",X"08",X"21",X"A9",X"00",X"9D",X"04",X"21",X"A9",X"00",X"9D",X"0A",X"21",X"A9",
		X"71",X"9D",X"0B",X"21",X"9D",X"03",X"21",X"4C",X"6B",X"A5",X"29",X"03",X"F0",X"0C",X"BD",X"01",
		X"02",X"29",X"0F",X"C9",X"0D",X"D0",X"03",X"4C",X"6B",X"A5",X"20",X"12",X"A3",X"8A",X"4A",X"A8",
		X"BD",X"09",X"02",X"85",X"08",X"BD",X"0A",X"02",X"85",X"09",X"30",X"04",X"A9",X"00",X"F0",X"02",
		X"A9",X"FF",X"06",X"08",X"26",X"09",X"2A",X"06",X"08",X"26",X"09",X"2A",X"29",X"1F",X"99",X"03",
		X"22",X"A5",X"09",X"99",X"02",X"22",X"BD",X"0B",X"02",X"85",X"0A",X"BD",X"0C",X"02",X"85",X"0B",
		X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"06",X"0A",X"26",X"0B",X"2A",X"06",X"0A",X"26",
		X"0B",X"2A",X"29",X"1F",X"99",X"01",X"22",X"A5",X"0B",X"99",X"00",X"22",X"BD",X"01",X"02",X"29",
		X"0F",X"C9",X"03",X"D0",X"03",X"4C",X"38",X"A5",X"C9",X"05",X"F0",X"1A",X"C9",X"0E",X"90",X"38",
		X"0A",X"A8",X"BD",X"00",X"02",X"29",X"03",X"C9",X"01",X"D0",X"33",X"A9",X"E6",X"9D",X"00",X"21",
		X"9D",X"06",X"21",X"4C",X"29",X"A5",X"A9",X"70",X"9D",X"03",X"21",X"A9",X"71",X"9D",X"0B",X"21",
		X"A9",X"00",X"9D",X"02",X"21",X"9D",X"0A",X"21",X"A9",X"E2",X"9D",X"00",X"21",X"A9",X"87",X"9D",
		X"06",X"21",X"4C",X"6B",X"A5",X"4C",X"96",X"A5",X"0A",X"A8",X"C9",X"16",X"F0",X"F7",X"C0",X"08",
		X"D0",X"2B",X"AD",X"0A",X"60",X"29",X"07",X"09",X"C0",X"C9",X"C0",X"D0",X"04",X"A9",X"C7",X"D0",
		X"00",X"9D",X"00",X"21",X"B9",X"01",X"01",X"9D",X"06",X"21",X"A5",X"F6",X"C9",X"03",X"D0",X"19",
		X"A9",X"0C",X"9D",X"0F",X"02",X"A9",X"20",X"9D",X"02",X"21",X"4C",X"6B",X"A5",X"B9",X"00",X"01",
		X"9D",X"00",X"21",X"B9",X"01",X"01",X"9D",X"06",X"21",X"B9",X"D6",X"A5",X"9D",X"0F",X"02",X"B9",
		X"D5",X"A5",X"9D",X"02",X"21",X"4C",X"6B",X"A5",X"AD",X"62",X"56",X"9D",X"0A",X"21",X"AD",X"63",
		X"56",X"9D",X"0B",X"21",X"A0",X"04",X"BD",X"02",X"02",X"F0",X"02",X"A0",X"0C",X"B9",X"00",X"01",
		X"9D",X"00",X"21",X"B9",X"01",X"01",X"9D",X"06",X"21",X"4C",X"6B",X"A5",X"C9",X"01",X"F0",X"0B",
		X"BD",X"01",X"02",X"29",X"0F",X"A8",X"B9",X"13",X"B0",X"10",X"0C",X"8A",X"18",X"69",X"10",X"AA",
		X"4A",X"A8",X"F0",X"18",X"4C",X"D6",X"A3",X"A5",X"6F",X"29",X"03",X"D0",X"EE",X"AD",X"0A",X"60",
		X"29",X"07",X"A8",X"B9",X"8D",X"A5",X"9D",X"00",X"21",X"4C",X"6B",X"A5",X"60",X"E7",X"E1",X"E1",
		X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"BD",X"0D",X"02",X"29",X"18",X"4A",X"4A",X"4A",X"84",X"19",
		X"A8",X"B9",X"B1",X"A5",X"9D",X"00",X"21",X"A9",X"00",X"9D",X"06",X"21",X"A4",X"19",X"4C",X"29",
		X"A5",X"E1",X"E2",X"E3",X"E7",X"C5",X"C2",X"E4",X"E4",X"A4",X"A6",X"E5",X"00",X"C7",X"00",X"E2",
		X"87",X"E5",X"A4",X"E1",X"84",X"C7",X"E4",X"E6",X"E4",X"E4",X"E1",X"E2",X"00",X"00",X"00",X"E4",
		X"E2",X"C5",X"A2",X"C7",X"E4",X"7F",X"02",X"20",X"03",X"60",X"03",X"00",X"04",X"60",X"02",X"00",
		X"04",X"00",X"04",X"00",X"04",X"60",X"03",X"3F",X"04",X"3F",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"A2",X"00",X"8E",X"3A",X"04",X"86",X"82",X"8E",X"04",X"03",X"86",
		X"40",X"BD",X"00",X"02",X"29",X"03",X"C9",X"02",X"90",X"05",X"F0",X"1F",X"4C",X"5C",X"A6",X"BD",
		X"01",X"02",X"29",X"0F",X"A8",X"B9",X"13",X"B0",X"29",X"20",X"D0",X"03",X"EE",X"3A",X"04",X"98",
		X"0A",X"A8",X"B9",X"2A",X"A7",X"48",X"B9",X"29",X"A7",X"48",X"60",X"8A",X"F0",X"DE",X"BD",X"01",
		X"02",X"29",X"0F",X"A8",X"B9",X"13",X"B0",X"30",X"20",X"BD",X"02",X"21",X"18",X"69",X"10",X"9D",
		X"02",X"21",X"10",X"18",X"A9",X"00",X"9D",X"02",X"21",X"FE",X"03",X"21",X"BD",X"03",X"21",X"C9",
		X"74",X"90",X"09",X"20",X"FE",X"A6",X"4C",X"5C",X"A6",X"20",X"C2",X"A6",X"A5",X"40",X"18",X"69",
		X"10",X"AA",X"B0",X"03",X"4C",X"FF",X"A5",X"AD",X"01",X"03",X"D0",X"15",X"AD",X"04",X"03",X"F0",
		X"1B",X"AD",X"3A",X"04",X"0D",X"36",X"04",X"D0",X"13",X"A9",X"FF",X"8D",X"01",X"03",X"4C",X"8C",
		X"A6",X"AD",X"04",X"03",X"0D",X"3A",X"04",X"D0",X"03",X"8D",X"01",X"03",X"AD",X"00",X"02",X"C9",
		X"02",X"D0",X"2E",X"A9",X"01",X"8D",X"01",X"03",X"AD",X"0A",X"60",X"09",X"E0",X"8D",X"00",X"21",
		X"AD",X"06",X"02",X"18",X"69",X"03",X"29",X"3F",X"8D",X"06",X"02",X"A2",X"00",X"20",X"1B",X"A3",
		X"AD",X"3A",X"04",X"0D",X"04",X"03",X"D0",X"09",X"A5",X"BA",X"D0",X"05",X"A9",X"03",X"8D",X"00",
		X"02",X"60",X"BD",X"03",X"02",X"0A",X"0A",X"A8",X"B9",X"88",X"B1",X"9D",X"00",X"21",X"B9",X"89",
		X"B1",X"9D",X"01",X"21",X"B9",X"8A",X"B1",X"9D",X"02",X"21",X"B9",X"8B",X"B1",X"9D",X"03",X"21",
		X"BD",X"03",X"02",X"18",X"7D",X"02",X"02",X"29",X"07",X"9D",X"03",X"02",X"D0",X"0F",X"BD",X"02",
		X"02",X"30",X"0B",X"A9",X"FF",X"9D",X"02",X"02",X"A9",X"08",X"9D",X"03",X"02",X"60",X"78",X"A4",
		X"40",X"A9",X"00",X"99",X"00",X"21",X"99",X"06",X"21",X"A9",X"60",X"99",X"05",X"21",X"A9",X"00",
		X"99",X"04",X"21",X"A9",X"A4",X"99",X"05",X"21",X"A9",X"60",X"99",X"07",X"21",X"A9",X"71",X"99",
		X"03",X"21",X"A9",X"03",X"9D",X"00",X"02",X"58",X"60",X"64",X"A8",X"48",X"A7",X"E3",X"A8",X"0F",
		X"A9",X"02",X"AA",X"E5",X"A9",X"9B",X"A9",X"20",X"AA",X"44",X"AA",X"89",X"AB",X"ED",X"AC",X"7F",
		X"A9",X"78",X"AF",X"4C",X"AD",X"6E",X"AE",X"17",X"AE",X"A5",X"73",X"F0",X"13",X"A9",X"0A",X"8D",
		X"05",X"02",X"A0",X"50",X"20",X"87",X"B0",X"AD",X"0E",X"02",X"8D",X"06",X"02",X"4C",X"83",X"A7",
		X"A9",X"03",X"8D",X"05",X"02",X"24",X"EF",X"10",X"33",X"A9",X"05",X"8D",X"05",X"02",X"A0",X"50",
		X"20",X"87",X"B0",X"A5",X"47",X"30",X"22",X"AD",X"0E",X"02",X"8D",X"06",X"02",X"A5",X"F7",X"C9",
		X"06",X"B0",X"13",X"A2",X"00",X"20",X"B4",X"C9",X"A5",X"73",X"D0",X"07",X"AD",X"0A",X"60",X"29",
		X"03",X"F0",X"03",X"20",X"DE",X"C3",X"20",X"DE",X"A7",X"4C",X"5C",X"A6",X"AD",X"5C",X"04",X"8D",
		X"05",X"02",X"AD",X"00",X"80",X"29",X"0F",X"49",X"0F",X"F0",X"0F",X"A8",X"B9",X"C0",X"A7",X"30",
		X"09",X"8D",X"06",X"02",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"20",X"DE",X"A7",X"4C",X"5C",X"A6",
		X"80",X"10",X"30",X"80",X"20",X"18",X"28",X"80",X"00",X"08",X"38",X"80",X"80",X"80",X"80",X"80",
		X"8A",X"18",X"69",X"10",X"AA",X"C9",X"50",X"D0",X"44",X"A9",X"00",X"85",X"4F",X"60",X"A5",X"73",
		X"D0",X"1A",X"24",X"EF",X"10",X"17",X"AD",X"0E",X"02",X"85",X"71",X"A5",X"F7",X"C9",X"07",X"F0",
		X"2A",X"C9",X"02",X"90",X"07",X"C9",X"04",X"B0",X"03",X"4C",X"1B",X"A8",X"60",X"AD",X"00",X"88",
		X"29",X"0F",X"49",X"0F",X"D0",X"05",X"A9",X"00",X"85",X"4F",X"60",X"A8",X"B9",X"C0",X"A7",X"30",
		X"EB",X"85",X"71",X"C6",X"4F",X"10",X"E5",X"A9",X"02",X"85",X"4F",X"A2",X"10",X"BD",X"00",X"02",
		X"29",X"03",X"F0",X"AC",X"86",X"40",X"A5",X"71",X"8D",X"04",X"02",X"9D",X"06",X"02",X"24",X"EF",
		X"10",X"06",X"AD",X"06",X"02",X"9D",X"06",X"02",X"20",X"22",X"BD",X"A9",X"01",X"9D",X"0D",X"02",
		X"AD",X"09",X"02",X"9D",X"09",X"02",X"AD",X"0A",X"02",X"9D",X"0A",X"02",X"AD",X"0B",X"02",X"9D",
		X"0B",X"02",X"AD",X"0C",X"02",X"9D",X"0C",X"02",X"A9",X"00",X"9D",X"00",X"02",X"20",X"B4",X"C9",
		X"A9",X"00",X"85",X"40",X"60",X"20",X"7C",X"AF",X"A5",X"82",X"F0",X"33",X"A8",X"DE",X"0D",X"02",
		X"10",X"2A",X"AD",X"3F",X"04",X"09",X"01",X"9D",X"0D",X"02",X"A9",X"FF",X"85",X"47",X"4A",X"85",
		X"46",X"20",X"03",X"CE",X"A6",X"40",X"9D",X"0E",X"02",X"A5",X"83",X"9D",X"01",X"02",X"A5",X"84",
		X"18",X"69",X"01",X"29",X"0F",X"D0",X"02",X"A9",X"0F",X"9D",X"05",X"02",X"4C",X"D8",X"A8",X"86",
		X"82",X"DE",X"0D",X"02",X"10",X"28",X"AD",X"0A",X"60",X"10",X"11",X"A9",X"FF",X"85",X"47",X"4A",
		X"85",X"46",X"A0",X"00",X"20",X"03",X"CE",X"A6",X"40",X"4C",X"C1",X"A8",X"AD",X"0A",X"60",X"29",
		X"3F",X"9D",X"0E",X"02",X"AD",X"3F",X"04",X"0A",X"0A",X"09",X"01",X"9D",X"0D",X"02",X"BD",X"01",
		X"02",X"85",X"83",X"BD",X"05",X"02",X"85",X"84",X"20",X"31",X"B1",X"20",X"B4",X"C9",X"20",X"DE",
		X"C3",X"4C",X"5C",X"A6",X"20",X"7C",X"AF",X"DE",X"0D",X"02",X"D0",X"18",X"BD",X"00",X"02",X"29",
		X"F7",X"9D",X"00",X"02",X"AD",X"3F",X"04",X"09",X"01",X"9D",X"0D",X"02",X"20",X"23",X"B0",X"A6",
		X"40",X"9D",X"0E",X"02",X"20",X"31",X"B1",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"4C",X"5C",X"A6",
		X"24",X"EF",X"30",X"27",X"A5",X"6C",X"F0",X"08",X"A9",X"20",X"9D",X"0D",X"02",X"4C",X"30",X"A9",
		X"AD",X"01",X"03",X"D0",X"58",X"A5",X"6F",X"29",X"0E",X"D0",X"52",X"DE",X"0D",X"02",X"30",X"2A",
		X"BD",X"02",X"02",X"F0",X"06",X"BD",X"0D",X"02",X"4C",X"41",X"A9",X"BD",X"0D",X"02",X"18",X"69",
		X"0C",X"A8",X"29",X"30",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"71",X"9D",X"03",X"21",X"98",X"29",
		X"0F",X"0A",X"0A",X"0A",X"9D",X"02",X"21",X"4C",X"CA",X"AF",X"A9",X"02",X"9D",X"01",X"02",X"BD",
		X"02",X"02",X"F0",X"05",X"A9",X"06",X"9D",X"01",X"02",X"A9",X"01",X"9D",X"0D",X"02",X"A9",X"00",
		X"9D",X"00",X"02",X"A9",X"71",X"9D",X"0B",X"21",X"A9",X"00",X"9D",X"0A",X"21",X"4C",X"5C",X"A6",
		X"24",X"EF",X"30",X"F9",X"A9",X"00",X"9D",X"05",X"02",X"A5",X"6F",X"29",X"07",X"D0",X"0A",X"DE",
		X"0D",X"02",X"10",X"05",X"A9",X"03",X"9D",X"00",X"02",X"4C",X"5C",X"A6",X"20",X"7C",X"AF",X"AD",
		X"04",X"03",X"0D",X"56",X"04",X"0D",X"57",X"04",X"D0",X"09",X"AD",X"05",X"02",X"9D",X"05",X"02",
		X"4C",X"DA",X"A9",X"DE",X"0D",X"02",X"30",X"03",X"4C",X"DA",X"A9",X"AD",X"05",X"02",X"38",X"E9",
		X"01",X"9D",X"05",X"02",X"AD",X"3F",X"04",X"09",X"01",X"9D",X"0D",X"02",X"A9",X"FF",X"85",X"46",
		X"A0",X"00",X"20",X"03",X"CE",X"A6",X"40",X"9D",X"0E",X"02",X"20",X"31",X"B1",X"20",X"B4",X"C9",
		X"20",X"DE",X"C3",X"4C",X"5C",X"A6",X"20",X"7C",X"AF",X"DE",X"0D",X"02",X"10",X"09",X"AD",X"3F",
		X"04",X"9D",X"0D",X"02",X"20",X"C5",X"B0",X"20",X"31",X"B1",X"20",X"B4",X"C9",X"20",X"DE",X"C3",
		X"4C",X"5C",X"A6",X"FE",X"0D",X"02",X"BD",X"0D",X"02",X"C9",X"18",X"90",X"08",X"A9",X"03",X"9D",
		X"00",X"02",X"4C",X"5C",X"A6",X"BD",X"06",X"02",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"4C",X"5C",
		X"A6",X"20",X"7C",X"AF",X"DE",X"0D",X"02",X"D0",X"10",X"AD",X"3F",X"04",X"09",X"01",X"9D",X"0D",
		X"02",X"20",X"56",X"B0",X"A6",X"40",X"9D",X"0E",X"02",X"20",X"31",X"B1",X"20",X"B4",X"C9",X"20",
		X"DE",X"C3",X"4C",X"5C",X"A6",X"20",X"7C",X"AF",X"FE",X"05",X"02",X"BD",X"05",X"02",X"C9",X"10",
		X"90",X"03",X"DE",X"05",X"02",X"AD",X"5D",X"04",X"C9",X"1C",X"B0",X"1E",X"BD",X"02",X"02",X"10",
		X"10",X"A9",X"02",X"9D",X"02",X"02",X"A9",X"00",X"9D",X"03",X"02",X"20",X"3B",X"AB",X"9D",X"06",
		X"02",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"4C",X"5C",X"A6",X"BD",X"04",X"02",X"10",X"40",X"A9",
		X"00",X"9D",X"04",X"02",X"9D",X"03",X"02",X"20",X"3B",X"AB",X"9D",X"0E",X"02",X"AD",X"5D",X"04",
		X"C9",X"2D",X"90",X"0C",X"AD",X"0A",X"60",X"29",X"8F",X"10",X"13",X"29",X"0F",X"4C",X"A9",X"AA",
		X"AD",X"0A",X"60",X"29",X"87",X"10",X"07",X"29",X"07",X"49",X"FF",X"18",X"69",X"01",X"18",X"7D",
		X"0E",X"02",X"29",X"3F",X"9D",X"06",X"02",X"A9",X"08",X"9D",X"0D",X"02",X"4C",X"71",X"AA",X"BD",
		X"02",X"02",X"10",X"20",X"DE",X"0D",X"02",X"10",X"A8",X"A9",X"01",X"9D",X"02",X"02",X"A9",X"00",
		X"9D",X"03",X"02",X"AD",X"5D",X"04",X"38",X"E9",X"25",X"30",X"4A",X"C9",X"20",X"90",X"02",X"A9",
		X"1F",X"9D",X"03",X"02",X"DE",X"0D",X"02",X"10",X"3C",X"FE",X"04",X"02",X"BD",X"04",X"02",X"C9",
		X"05",X"90",X"19",X"A9",X"00",X"9D",X"04",X"02",X"BD",X"03",X"02",X"18",X"69",X"20",X"90",X"09",
		X"18",X"69",X"01",X"29",X"1F",X"D0",X"02",X"A9",X"1F",X"9D",X"03",X"02",X"BD",X"03",X"02",X"29",
		X"1F",X"0A",X"A8",X"B9",X"4A",X"AB",X"9D",X"0D",X"02",X"B9",X"4B",X"AB",X"9D",X"02",X"02",X"20",
		X"3B",X"AB",X"9D",X"0E",X"02",X"BD",X"02",X"02",X"85",X"1B",X"20",X"38",X"B1",X"A9",X"00",X"9D",
		X"02",X"02",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"4C",X"5C",X"A6",X"A9",X"FF",X"85",X"47",X"4A",
		X"85",X"46",X"A0",X"00",X"20",X"03",X"CE",X"A6",X"40",X"60",X"07",X"01",X"07",X"01",X"06",X"01",
		X"06",X"01",X"05",X"01",X"05",X"01",X"04",X"01",X"04",X"01",X"04",X"02",X"04",X"02",X"04",X"03",
		X"04",X"03",X"04",X"04",X"04",X"04",X"04",X"05",X"04",X"05",X"04",X"06",X"03",X"06",X"03",X"07",
		X"03",X"08",X"03",X"09",X"03",X"0A",X"02",X"08",X"02",X"09",X"01",X"07",X"01",X"08",X"01",X"09",
		X"01",X"0A",X"01",X"0B",X"01",X"0C",X"01",X"0D",X"01",X"0E",X"A5",X"6C",X"D0",X"04",X"A5",X"73",
		X"F0",X"0D",X"A9",X"0F",X"9D",X"05",X"02",X"A9",X"01",X"1D",X"00",X"02",X"9D",X"00",X"02",X"DE",
		X"0D",X"02",X"F0",X"20",X"BD",X"00",X"02",X"10",X"06",X"20",X"31",X"B1",X"4C",X"BB",X"AB",X"BD",
		X"06",X"02",X"18",X"7D",X"04",X"02",X"29",X"3F",X"9D",X"06",X"02",X"20",X"B4",X"C9",X"20",X"DE",
		X"C3",X"4C",X"5C",X"A6",X"BD",X"02",X"02",X"85",X"4C",X"BD",X"03",X"02",X"85",X"4D",X"20",X"CF",
		X"AC",X"BD",X"00",X"02",X"10",X"5E",X"8A",X"A8",X"84",X"19",X"98",X"18",X"69",X"10",X"D0",X"0C",
		X"E4",X"19",X"D0",X"37",X"A9",X"00",X"8D",X"34",X"01",X"4C",X"1B",X"AC",X"A8",X"B9",X"01",X"02",
		X"29",X"0F",X"C9",X"09",X"D0",X"E4",X"B9",X"00",X"02",X"29",X"03",X"F0",X"DB",X"4C",X"DA",X"AB",
		X"9D",X"0D",X"02",X"C8",X"B1",X"4C",X"9D",X"04",X"02",X"A9",X"02",X"18",X"65",X"4C",X"9D",X"02",
		X"02",X"A9",X"00",X"65",X"4D",X"9D",X"03",X"02",X"4C",X"AF",X"AB",X"BD",X"00",X"02",X"29",X"7F",
		X"9D",X"00",X"02",X"AD",X"27",X"04",X"C5",X"40",X"F0",X"3B",X"AD",X"25",X"04",X"85",X"4C",X"AD",
		X"26",X"04",X"85",X"4D",X"A0",X"00",X"B1",X"4C",X"10",X"C6",X"A9",X"80",X"1D",X"00",X"02",X"9D",
		X"00",X"02",X"FE",X"05",X"02",X"BD",X"05",X"02",X"C9",X"10",X"D0",X"0B",X"DE",X"05",X"02",X"A9",
		X"01",X"1D",X"00",X"02",X"9D",X"00",X"02",X"EC",X"27",X"04",X"F0",X"44",X"AD",X"35",X"01",X"9D",
		X"0E",X"02",X"4C",X"B6",X"AC",X"A0",X"00",X"B1",X"4C",X"D0",X"11",X"A9",X"C6",X"85",X"4C",X"8D",
		X"25",X"04",X"A9",X"B1",X"85",X"4D",X"8D",X"26",X"04",X"4C",X"65",X"AC",X"30",X"0D",X"A5",X"4C",
		X"8D",X"25",X"04",X"A5",X"4D",X"8D",X"26",X"04",X"4C",X"34",X"AC",X"AD",X"34",X"01",X"F0",X"EE",
		X"A9",X"02",X"18",X"65",X"4C",X"85",X"4C",X"A9",X"00",X"65",X"4D",X"85",X"4D",X"4C",X"65",X"AC",
		X"A9",X"7F",X"8D",X"34",X"01",X"85",X"46",X"A0",X"00",X"20",X"03",X"CE",X"29",X"3F",X"A6",X"40",
		X"9D",X"0E",X"02",X"8D",X"35",X"01",X"A0",X"01",X"B1",X"4C",X"9D",X"0D",X"02",X"A9",X"02",X"18",
		X"65",X"4C",X"9D",X"02",X"02",X"A9",X"00",X"65",X"4D",X"9D",X"03",X"02",X"4C",X"A9",X"AB",X"A0",
		X"50",X"E0",X"50",X"F0",X"15",X"B9",X"00",X"02",X"19",X"01",X"02",X"29",X"0F",X"C9",X"09",X"F0",
		X"09",X"98",X"18",X"69",X"10",X"A8",X"C4",X"40",X"90",X"EB",X"8C",X"27",X"04",X"60",X"20",X"7C",
		X"AF",X"A0",X"50",X"B9",X"01",X"02",X"19",X"00",X"02",X"29",X"0F",X"C9",X"09",X"F0",X"0A",X"98",
		X"18",X"69",X"10",X"A8",X"D0",X"ED",X"4C",X"DE",X"AF",X"DE",X"0D",X"02",X"10",X"18",X"AD",X"3F",
		X"04",X"09",X"01",X"9D",X"0D",X"02",X"A9",X"7F",X"85",X"46",X"A0",X"00",X"20",X"03",X"CE",X"29",
		X"3F",X"A6",X"40",X"9D",X"0E",X"02",X"20",X"31",X"B1",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"4C",
		X"5C",X"A6",X"BD",X"03",X"02",X"C5",X"19",X"B0",X"5E",X"0A",X"7D",X"03",X"02",X"A8",X"B9",X"AD",
		X"B1",X"9D",X"02",X"21",X"B9",X"AE",X"B1",X"9D",X"03",X"21",X"4C",X"5C",X"A6",X"A5",X"F6",X"C9",
		X"03",X"D0",X"02",X"A9",X"01",X"18",X"69",X"06",X"85",X"19",X"A5",X"6C",X"F0",X"0C",X"BD",X"00",
		X"02",X"29",X"03",X"C9",X"01",X"F0",X"11",X"4C",X"DE",X"AF",X"A5",X"73",X"D0",X"F0",X"BD",X"00",
		X"02",X"29",X"03",X"D0",X"03",X"4C",X"FE",X"AD",X"DE",X"0D",X"02",X"10",X"B5",X"A5",X"F6",X"C9",
		X"03",X"D0",X"05",X"A9",X"04",X"4C",X"8D",X"AD",X"38",X"A9",X"05",X"E5",X"F6",X"9D",X"0D",X"02",
		X"BD",X"03",X"02",X"C5",X"19",X"90",X"06",X"20",X"FE",X"A6",X"4C",X"5C",X"A6",X"0A",X"7D",X"03",
		X"02",X"A8",X"B9",X"AC",X"B1",X"85",X"46",X"A9",X"60",X"9D",X"01",X"21",X"AD",X"0A",X"60",X"29",
		X"07",X"A8",X"B9",X"8D",X"A5",X"9D",X"00",X"21",X"FE",X"03",X"02",X"A9",X"80",X"8D",X"00",X"03",
		X"A9",X"00",X"A8",X"48",X"C4",X"40",X"F0",X"24",X"B9",X"01",X"02",X"29",X"0F",X"C9",X"04",X"F0",
		X"1B",X"B9",X"00",X"02",X"29",X"03",X"C9",X"02",X"B0",X"12",X"C9",X"01",X"D0",X"09",X"B9",X"01",
		X"02",X"29",X"0F",X"C9",X"0D",X"F0",X"05",X"A6",X"40",X"20",X"03",X"CE",X"68",X"18",X"69",X"10",
		X"A8",X"D0",X"CF",X"A9",X"00",X"8D",X"00",X"03",X"20",X"46",X"BD",X"4C",X"5C",X"A6",X"DE",X"0D",
		X"02",X"10",X"09",X"AD",X"3F",X"04",X"9D",X"0D",X"02",X"20",X"C5",X"B0",X"20",X"31",X"B1",X"20",
		X"B4",X"C9",X"20",X"DE",X"C3",X"4C",X"5C",X"A6",X"EE",X"04",X"03",X"AC",X"04",X"03",X"8A",X"99",
		X"04",X"03",X"AD",X"01",X"03",X"F0",X"0A",X"10",X"05",X"A9",X"01",X"9D",X"00",X"02",X"4C",X"DE",
		X"AF",X"DE",X"0D",X"02",X"10",X"13",X"AD",X"3F",X"04",X"4A",X"09",X"01",X"9D",X"0D",X"02",X"A9",
		X"FF",X"85",X"47",X"4A",X"85",X"46",X"20",X"D5",X"B0",X"A5",X"6F",X"D0",X"0D",X"BD",X"05",X"02",
		X"18",X"69",X"01",X"C9",X"10",X"B0",X"03",X"9D",X"05",X"02",X"BD",X"05",X"02",X"85",X"19",X"20",
		X"31",X"B1",X"C6",X"19",X"10",X"F9",X"20",X"B4",X"C9",X"20",X"DE",X"C3",X"4C",X"5C",X"A6",X"EE",
		X"04",X"03",X"AC",X"04",X"03",X"8A",X"99",X"04",X"03",X"AD",X"01",X"03",X"F0",X"0A",X"10",X"05",
		X"A9",X"01",X"9D",X"00",X"02",X"4C",X"DE",X"AF",X"BD",X"02",X"02",X"D0",X"58",X"A9",X"00",X"9D",
		X"05",X"02",X"DE",X"0D",X"02",X"30",X"12",X"AD",X"0A",X"60",X"29",X"3F",X"D0",X"08",X"AD",X"0A",
		X"60",X"29",X"3F",X"9D",X"0E",X"02",X"4C",X"2C",X"AF",X"A9",X"30",X"9D",X"0D",X"02",X"A9",X"50",
		X"9D",X"02",X"02",X"A8",X"20",X"49",X"AF",X"B0",X"18",X"98",X"18",X"69",X"10",X"90",X"F1",X"A9",
		X"00",X"9D",X"02",X"02",X"9D",X"05",X"02",X"AD",X"3F",X"04",X"0A",X"9D",X"0D",X"02",X"4C",X"5C",
		X"A6",X"A9",X"FF",X"85",X"47",X"4A",X"85",X"46",X"20",X"03",X"CE",X"A6",X"40",X"A5",X"47",X"9D",
		X"06",X"02",X"4C",X"35",X"AF",X"A8",X"20",X"49",X"AF",X"90",X"D4",X"DE",X"0D",X"02",X"30",X"0E",
		X"BD",X"06",X"02",X"18",X"69",X"01",X"29",X"3F",X"9D",X"06",X"02",X"4C",X"2F",X"AF",X"A9",X"FF",
		X"9D",X"0D",X"02",X"A5",X"6F",X"29",X"01",X"D0",X"23",X"BD",X"05",X"02",X"18",X"69",X"01",X"C9",
		X"10",X"B0",X"03",X"9D",X"05",X"02",X"A9",X"FF",X"85",X"47",X"4A",X"85",X"46",X"20",X"03",X"CE",
		X"A6",X"40",X"A5",X"47",X"29",X"3F",X"9D",X"06",X"02",X"9D",X"0E",X"02",X"20",X"31",X"B1",X"20",
		X"B4",X"C9",X"20",X"DE",X"C3",X"BD",X"02",X"02",X"F0",X"0C",X"A8",X"A5",X"6F",X"29",X"02",X"D0",
		X"05",X"A9",X"E7",X"99",X"00",X"21",X"4C",X"5C",X"A6",X"C4",X"40",X"F0",X"28",X"B9",X"00",X"02",
		X"29",X"03",X"C9",X"02",X"B0",X"1F",X"B9",X"01",X"02",X"29",X"0F",X"C9",X"03",X"F0",X"16",X"C9",
		X"05",X"F0",X"0C",X"C9",X"08",X"F0",X"0E",X"C9",X"0F",X"F0",X"0A",X"C9",X"0D",X"D0",X"08",X"A5",
		X"79",X"C9",X"1E",X"B0",X"02",X"18",X"60",X"38",X"60",X"4C",X"5C",X"A6",X"A5",X"6C",X"05",X"73",
		X"0D",X"00",X"02",X"D0",X"52",X"BD",X"00",X"02",X"29",X"03",X"C9",X"01",X"D0",X"39",X"BD",X"01",
		X"02",X"29",X"0F",X"A8",X"B9",X"13",X"B0",X"29",X"08",X"D0",X"3C",X"A5",X"6F",X"29",X"07",X"D0",
		X"27",X"B9",X"13",X"B0",X"29",X"02",X"D0",X"03",X"DE",X"0D",X"02",X"98",X"0A",X"A8",X"B9",X"00",
		X"01",X"9D",X"06",X"21",X"B9",X"01",X"01",X"9D",X"00",X"21",X"BD",X"0D",X"02",X"10",X"09",X"A9",
		X"00",X"9D",X"00",X"02",X"9D",X"0D",X"02",X"60",X"68",X"68",X"BD",X"0D",X"02",X"C9",X"08",X"B0",
		X"03",X"20",X"D9",X"A2",X"4C",X"5C",X"A6",X"68",X"68",X"A9",X"00",X"9D",X"00",X"02",X"A5",X"6F",
		X"29",X"03",X"D0",X"23",X"A0",X"00",X"A9",X"FF",X"85",X"47",X"4A",X"85",X"46",X"20",X"03",X"CE",
		X"A6",X"40",X"18",X"69",X"20",X"29",X"3F",X"9D",X"0E",X"02",X"BD",X"05",X"02",X"18",X"69",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
