library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",
		X"00",X"44",X"6C",X"38",X"38",X"6C",X"44",X"00",X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",
		X"00",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",
		X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",
		X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",
		X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",
		X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",
		X"00",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",
		X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",
		X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",
		X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",
		X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"16",X"0E",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",
		X"00",X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",
		X"00",X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",
		X"00",X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",
		X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",
		X"00",X"00",X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"3E",X"FE",X"70",X"38",X"70",X"FE",X"3E",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"06",X"1E",X"F0",X"F0",X"1E",X"06",
		X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",
		X"00",X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",
		X"00",X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",
		X"00",X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",
		X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",
		X"00",X"00",X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"3E",X"FE",X"70",X"38",X"70",X"FE",X"3E",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"06",X"1E",X"F0",X"F0",X"1E",X"06",
		X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"60",X"60",X"08",X"1C",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"50",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"7E",X"81",X"BD",X"BD",X"A5",X"A5",X"81",X"7E",
		X"00",X"FF",X"FF",X"C3",X"C3",X"E7",X"7E",X"7E",X"FF",X"DB",X"DB",X"DB",X"7E",X"FF",X"C3",X"C3",
		X"F7",X"76",X"7E",X"FF",X"C3",X"C3",X"FF",X"7E",X"FF",X"89",X"7E",X"7E",X"7E",X"7E",X"7E",X"89",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"8F",X"76",X"76",X"76",X"76",X"76",X"F9",
		X"FF",X"FF",X"7E",X"76",X"76",X"76",X"76",X"89",X"FF",X"F9",X"F7",X"F7",X"F7",X"F7",X"08",X"FF",
		X"FF",X"F9",X"76",X"76",X"76",X"76",X"76",X"8F",X"FF",X"89",X"76",X"76",X"76",X"76",X"76",X"8F",
		X"FF",X"F9",X"FE",X"FE",X"FE",X"FE",X"FE",X"89",X"FF",X"89",X"76",X"76",X"76",X"76",X"76",X"89",
		X"FF",X"F9",X"76",X"76",X"76",X"76",X"76",X"89",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"50",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"76",X"76",X"00",X"00",X"EE",
		X"00",X"6C",X"82",X"6C",X"00",X"6C",X"82",X"6C",X"00",X"00",X"00",X"EE",X"00",X"6C",X"82",X"6C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"E2",X"92",X"8C",
		X"00",X"00",X"00",X"00",X"82",X"92",X"92",X"6C",X"00",X"00",X"00",X"00",X"0E",X"10",X"10",X"EC",
		X"00",X"00",X"00",X"00",X"8E",X"92",X"92",X"E2",X"00",X"00",X"00",X"00",X"7C",X"92",X"92",X"60",
		X"00",X"00",X"00",X"00",X"82",X"42",X"22",X"1E",X"00",X"00",X"00",X"00",X"6C",X"92",X"92",X"6C",
		X"00",X"00",X"00",X"00",X"4C",X"92",X"92",X"7C",X"00",X"6C",X"82",X"6C",X"00",X"00",X"00",X"00",
		X"C2",X"94",X"6A",X"FC",X"FE",X"FF",X"FF",X"FE",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"D8",X"00",
		X"00",X"46",X"7F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"3F",X"7E",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"84",X"28",X"D4",X"F8",X"FC",X"FE",X"FE",X"FC",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"B0",X"00",
		X"01",X"8D",X"FE",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"7F",X"FD",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"50",X"A8",X"F0",X"F8",X"FC",X"FC",X"F8",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"60",X"00",
		X"03",X"1A",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FB",X"90",
		X"00",X"01",X"01",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"01",X"00",
		X"10",X"A0",X"50",X"E0",X"F0",X"F8",X"F8",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"06",X"34",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"20",
		X"00",X"02",X"03",X"01",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"00",X"01",X"03",X"01",
		X"20",X"40",X"A0",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",
		X"0C",X"69",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"40",
		X"00",X"04",X"07",X"03",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"01",X"03",X"07",X"02",
		X"40",X"80",X"40",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"18",X"D2",X"ED",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",X"80",
		X"00",X"08",X"0F",X"07",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"03",X"07",X"0F",X"04",
		X"80",X"00",X"80",X"00",X"80",X"C0",X"C0",X"80",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"30",X"A5",X"DA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B6",X"00",
		X"00",X"11",X"1F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"07",X"0F",X"1F",X"09",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"61",X"4A",X"B5",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"6C",X"00",
		X"00",X"23",X"3F",X"1F",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"0F",X"1F",X"3F",X"12",
		X"78",X"FC",X"FC",X"70",X"02",X"00",X"7D",X"7D",X"7D",X"7D",X"00",X"02",X"FC",X"FC",X"78",X"00",
		X"00",X"7C",X"FE",X"FE",X"40",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"40",X"38",X"FE",X"FE",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"80",X"A0",X"A0",
		X"00",X"00",X"00",X"00",X"0E",X"1F",X"1F",X"1F",X"1F",X"1E",X"40",X"80",X"3F",X"7F",X"7F",X"7F",
		X"A0",X"A0",X"80",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"3F",X"80",X"40",X"1E",X"1F",X"1F",X"1F",X"1F",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"78",X"7F",X"78",X"00",X"7E",X"5E",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"25",X"00",X"04",X"10",X"00",X"68",X"1F",X"76",X"3C",
		X"5E",X"7E",X"00",X"78",X"7F",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"46",X"0F",X"28",X"00",X"00",X"04",X"00",X"24",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"FE",X"03",X"01",X"F8",X"F8",X"F8",X"F9",X"F9",X"F9",
		X"00",X"03",X"07",X"07",X"07",X"07",X"03",X"3F",X"C0",X"00",X"00",X"0F",X"7F",X"7F",X"7F",X"7F",
		X"F9",X"F9",X"F9",X"F8",X"F8",X"F8",X"01",X"02",X"FC",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"7F",X"7F",X"7F",X"7F",X"0F",X"00",X"00",X"C0",X"3F",X"03",X"07",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"FF",X"FE",X"0C",X"FE",X"FE",X"FE",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"01",X"12",X"00",X"60",X"00",X"9C",
		X"BE",X"FE",X"FE",X"FE",X"0C",X"FE",X"FF",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"9C",X"00",X"60",X"00",X"12",X"01",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"02",X"01",X"F9",X"F9",X"F9",X"F9",X"F8",X"F8",X"F8",
		X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"F0",X"00",X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"F8",X"F8",X"F8",X"F9",X"F9",X"F9",X"F9",X"01",X"02",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"E0",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"1F",X"00",X"F0",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"FF",X"D8",X"B0",X"00",X"FF",X"FF",X"FF",X"FD",X"DD",X"DC",
		X"00",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"7F",X"7F",X"3C",X"2F",X"27",X"27",X"27",X"25",X"25",
		X"DC",X"DD",X"FD",X"FF",X"FF",X"FF",X"00",X"B0",X"D8",X"FF",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"25",X"25",X"27",X"27",X"27",X"2F",X"3C",X"7F",X"7F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"70",X"00",X"E0",X"E0",X"E0",X"E8",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"1E",X"E0",X"07",X"3F",X"FF",X"FF",X"FF",
		X"E8",X"E8",X"E0",X"E0",X"E0",X"00",X"70",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"3F",X"07",X"E0",X"1E",X"3F",X"3F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"BE",X"3B",X"F8",X"FE",X"FE",X"FA",X"9A",X"B8",
		X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"10",X"21",X"23",X"27",X"27",X"27",X"26",
		X"B8",X"9A",X"FA",X"FE",X"FE",X"F8",X"3B",X"BE",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",
		X"26",X"27",X"27",X"27",X"23",X"21",X"10",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"B8",X"7C",X"7C",X"7C",X"78",X"02",X"FD",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FD",X"02",X"78",X"7C",X"7C",X"7C",X"B8",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"08",X"FA",X"FC",X"F9",X"F8",X"F0",X"03",X"78",X"FE",X"FE",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"02",
		X"BE",X"FE",X"FE",X"78",X"03",X"F0",X"F8",X"F9",X"FC",X"F8",X"08",X"00",X"40",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"1C",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"1C",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"3C",X"3C",X"3C",X"1C",X"00",X"3E",X"3E",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"80",X"04",X"00",X"00",X"12",X"00",X"80",
		X"3E",X"3E",X"3E",X"00",X"1C",X"3C",X"3C",X"3C",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"02",X"88",X"01",X"04",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"7C",X"F8",X"02",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"F8",X"02",X"F8",X"7C",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"18",X"3C",X"3C",X"3D",X"40",X"BE",X"BE",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"04",X"02",X"00",
		X"BE",X"BE",X"BE",X"40",X"3D",X"3C",X"3C",X"18",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"04",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"3E",X"18",X"FF",X"FC",X"84",X"84",X"84",X"84",X"FC",X"FF",X"18",X"3E",X"3E",X"3E",
		X"FE",X"FE",X"FE",X"18",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"18",X"FE",X"FE",X"FE",
		X"18",X"7E",X"7E",X"7E",X"1C",X"00",X"FC",X"03",X"03",X"FC",X"1C",X"7E",X"7E",X"7E",X"18",X"00",
		X"00",X"30",X"FC",X"FC",X"FC",X"78",X"FF",X"80",X"80",X"FF",X"00",X"58",X"FC",X"FC",X"FC",X"30",
		X"1C",X"3E",X"3E",X"20",X"FE",X"F1",X"E3",X"FF",X"FF",X"E3",X"F1",X"FE",X"3E",X"3E",X"1C",X"00",
		X"00",X"78",X"FC",X"FC",X"7D",X"3F",X"67",X"5F",X"5F",X"67",X"3F",X"41",X"FC",X"FC",X"FC",X"78",
		X"FE",X"FE",X"FE",X"38",X"FC",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FC",X"38",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"FE",X"FE",
		X"18",X"BC",X"BC",X"FE",X"FE",X"FF",X"FA",X"F2",X"02",X"37",X"FF",X"FE",X"FE",X"BC",X"BC",X"18",
		X"63",X"F7",X"F7",X"FF",X"FF",X"5F",X"7F",X"73",X"72",X"6D",X"7F",X"FF",X"FF",X"F7",X"F7",X"63",
		X"FC",X"FE",X"FE",X"FE",X"00",X"08",X"08",X"00",X"00",X"20",X"20",X"00",X"FE",X"FE",X"FE",X"FC",
		X"7F",X"FF",X"FF",X"FF",X"20",X"80",X"87",X"8F",X"8F",X"87",X"80",X"20",X"FF",X"FF",X"FF",X"7F",
		X"EF",X"EF",X"FF",X"1F",X"DF",X"1F",X"7F",X"5F",X"7F",X"5F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",
		X"F3",X"F3",X"F3",X"42",X"40",X"4C",X"5E",X"7F",X"7F",X"5E",X"4C",X"40",X"42",X"F3",X"F3",X"F3",
		X"E0",X"00",X"00",X"8E",X"CE",X"C0",X"E2",X"C2",X"E2",X"E2",X"C0",X"8E",X"8E",X"00",X"00",X"E0",
		X"79",X"00",X"02",X"07",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"15",X"00",X"00",X"79",
		X"E0",X"E0",X"00",X"EE",X"0E",X"E0",X"F2",X"12",X"12",X"F2",X"E0",X"0E",X"EE",X"00",X"E0",X"E0",
		X"79",X"00",X"00",X"FC",X"FE",X"BE",X"FC",X"FE",X"FE",X"FC",X"FE",X"FE",X"3C",X"08",X"00",X"79",
		X"E0",X"E0",X"00",X"EE",X"0E",X"E0",X"F2",X"12",X"12",X"F2",X"E0",X"0E",X"EE",X"00",X"E0",X"E0",
		X"79",X"01",X"30",X"F1",X"F0",X"87",X"F7",X"F1",X"F1",X"F7",X"C7",X"F0",X"31",X"30",X"01",X"79",
		X"E0",X"E0",X"00",X"EE",X"0E",X"E0",X"F2",X"12",X"12",X"F2",X"E0",X"0E",X"EE",X"00",X"E0",X"E0",
		X"79",X"09",X"60",X"69",X"68",X"0F",X"6F",X"61",X"61",X"6F",X"0F",X"68",X"69",X"60",X"09",X"79",
		X"00",X"78",X"FC",X"EC",X"EC",X"60",X"80",X"30",X"30",X"80",X"70",X"F4",X"F4",X"FC",X"78",X"00",
		X"00",X"78",X"FC",X"EC",X"EC",X"42",X"84",X"29",X"29",X"84",X"42",X"F4",X"F4",X"FC",X"78",X"00",
		X"3C",X"3C",X"38",X"40",X"80",X"00",X"E0",X"E1",X"E1",X"E0",X"00",X"80",X"40",X"38",X"3C",X"3C",
		X"10",X"7C",X"7C",X"7C",X"18",X"40",X"5F",X"5F",X"5F",X"5F",X"40",X"18",X"7C",X"7C",X"7C",X"10",
		X"80",X"60",X"04",X"9A",X"E8",X"FC",X"F8",X"70",X"F8",X"F4",X"E0",X"52",X"B0",X"00",X"50",X"20",
		X"00",X"80",X"05",X"E7",X"0D",X"BF",X"3F",X"2F",X"96",X"BF",X"BF",X"9F",X"06",X"20",X"12",X"00",
		X"00",X"A8",X"40",X"E8",X"1C",X"90",X"40",X"88",X"D0",X"E0",X"F0",X"F8",X"70",X"28",X"C0",X"00",
		X"21",X"44",X"32",X"C4",X"2A",X"6D",X"97",X"53",X"37",X"57",X"17",X"9F",X"2F",X"B2",X"24",X"41",
		X"42",X"04",X"40",X"E4",X"F2",X"F0",X"C8",X"12",X"99",X"A2",X"F4",X"F8",X"F4",X"7A",X"74",X"80",
		X"0A",X"8B",X"45",X"0B",X"9F",X"7F",X"BF",X"DF",X"5F",X"3F",X"8F",X"23",X"49",X"13",X"04",X"02",
		X"20",X"20",X"10",X"F8",X"FC",X"FC",X"FE",X"FF",X"FC",X"FE",X"FC",X"F8",X"F0",X"F0",X"C0",X"00",
		X"33",X"14",X"8D",X"8F",X"3B",X"DF",X"BF",X"7F",X"3F",X"5F",X"BF",X"FF",X"5F",X"3F",X"15",X"08",
		X"00",X"00",X"00",X"00",X"30",X"78",X"3C",X"38",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"7C",X"EC",X"DE",X"9C",X"CA",X"E7",X"72",X"AE",
		X"00",X"40",X"80",X"00",X"00",X"00",X"B0",X"60",X"70",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"F2",X"8E",X"3A",X"2C",X"F6",X"7B",X"7E",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"02",X"B6",X"95",X"16",X"A0",X"77",X"77",X"CF",X"E7",
		X"00",X"00",X"02",X"06",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2B",X"43",X"D3",X"6C",X"8C",X"16",X"3E",X"3F",X"08",X"20",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"02",X"01",X"06",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"A6",X"C2",X"FA",X"E8",X"F8",X"F0",X"C8",X"80",X"00",X"20",X"60",X"00",X"00",X"00",
		X"02",X"0C",X"1B",X"41",X"13",X"3D",X"F8",X"9F",X"CF",X"9F",X"0E",X"DE",X"C8",X"EA",X"F4",X"FE",
		X"00",X"C0",X"70",X"80",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"3E",X"DF",X"EE",X"DA",X"C4",X"A9",X"F0",X"32",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"38",X"36",X"46",X"8F",X"9E",X"7F",X"7C",X"60",X"FE",X"F3",X"3F",X"9F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"03",X"50",X"A2",X"4D",X"02",X"01",
		X"C3",X"7B",X"FD",X"FF",X"3A",X"B3",X"3A",X"AC",X"1D",X"51",X"82",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"02",X"04",X"0A",X"00",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"C4",X"F0",X"FA",X"F8",X"F8",X"F4",X"60",X"84",X"88",X"80",X"20",X"20",X"40",X"00",
		X"01",X"08",X"01",X"27",X"1F",X"3F",X"F1",X"FA",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FE",X"FF",
		X"00",X"00",X"60",X"F0",X"F8",X"F4",X"E0",X"F0",X"F0",X"FA",X"F0",X"C8",X"58",X"80",X"00",X"00",
		X"FC",X"FE",X"FE",X"FD",X"DB",X"F7",X"FB",X"FF",X"7F",X"BF",X"FF",X"AF",X"F6",X"61",X"01",X"00",
		X"80",X"28",X"2B",X"00",X"FE",X"FE",X"FF",X"FE",X"77",X"FE",X"F5",X"FB",X"FF",X"5F",X"3F",X"3F",
		X"01",X"02",X"05",X"08",X"00",X"09",X"0B",X"0F",X"95",X"6E",X"4F",X"FF",X"2F",X"20",X"46",X"59",
		X"FF",X"FF",X"F5",X"FB",X"FF",X"FF",X"EE",X"FB",X"FF",X"FF",X"7F",X"EE",X"4D",X"C8",X"04",X"00",
		X"27",X"8B",X"A7",X"2F",X"2F",X"2B",X"4F",X"0F",X"9B",X"0D",X"A7",X"40",X"A4",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"D0",X"B8",X"18",X"14",X"0C",X"22",X"70",X"0A",X"F0",X"80",X"58",X"00",
		X"05",X"10",X"BC",X"EC",X"00",X"40",X"8B",X"26",X"68",X"48",X"20",X"00",X"01",X"01",X"06",X"00",
		X"00",X"00",X"40",X"A0",X"42",X"08",X"08",X"00",X"20",X"40",X"80",X"00",X"80",X"40",X"00",X"40",
		X"00",X"04",X"01",X"01",X"06",X"00",X"00",X"10",X"88",X"75",X"7A",X"60",X"4A",X"0C",X"14",X"1E",
		X"00",X"40",X"14",X"30",X"35",X"02",X"80",X"08",X"9C",X"2B",X"01",X"00",X"80",X"00",X"20",X"F0",
		X"00",X"0A",X"00",X"00",X"04",X"00",X"11",X"01",X"00",X"04",X"0A",X"00",X"00",X"0A",X"0A",X"03",
		X"00",X"80",X"80",X"20",X"00",X"C4",X"84",X"20",X"24",X"28",X"80",X"C4",X"E0",X"60",X"58",X"60",
		X"00",X"00",X"4C",X"00",X"00",X"14",X"4E",X"08",X"00",X"18",X"38",X"82",X"C6",X"40",X"14",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"78",X"38",X"FC",X"FA",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F4",X"F0",X"74",X"30",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"08",X"16",X"1C",X"1F",X"1F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"21",X"1D",X"0F",X"0C",X"08",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"20",X"20",X"80",X"00",X"40",
		X"00",X"00",X"00",X"04",X"20",X"04",X"00",X"93",X"40",X"29",X"68",X"7A",X"F5",X"FA",X"F4",X"F8",
		X"00",X"20",X"20",X"00",X"80",X"00",X"20",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F4",X"FC",X"75",X"28",X"78",X"30",X"10",X"00",X"22",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"5E",X"2E",X"56",X"1C",X"0F",X"BB",X"37",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"06",X"02",X"01",X"05",X"08",X"02",
		X"07",X"25",X"8F",X"0F",X"2C",X"8A",X"49",X"04",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"20",X"40",X"20",X"10",X"00",X"00",X"C0",X"80",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"01",X"00",X"00",X"A0",X"12",X"14",X"02",X"01",X"20",X"40",X"01",X"80",X"40",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"22",X"01",X"81",X"40",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",X"00",X"08",X"10",X"00",X"80",X"48",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",
		X"80",X"80",X"C0",X"40",X"20",X"40",X"C0",X"A0",X"05",X"0A",X"04",X"04",X"14",X"08",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"80",X"CE",X"CE",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"CE",X"CE",X"80",X"00",X"E0",
		X"79",X"00",X"3F",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"3F",X"00",X"79",
		X"CF",X"03",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"03",X"CF",
		X"03",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"00",X"03",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",
		X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"C0",X"48",X"7C",X"FC",X"7D",X"E6",X"75",X"D2",X"BC",X"6C",X"FA",X"EC",X"AA",X"B0",X"76",X"10",
		X"00",X"82",X"15",X"0C",X"4E",X"07",X"ED",X"FF",X"FE",X"FF",X"8F",X"07",X"21",X"04",X"01",X"00",
		X"00",X"F0",X"08",X"F4",X"14",X"14",X"F4",X"08",X"F0",X"60",X"60",X"60",X"E0",X"E0",X"00",X"00",
		X"FC",X"FF",X"C0",X"C9",X"C1",X"C1",X"C9",X"C0",X"FF",X"FC",X"04",X"04",X"3F",X"3F",X"40",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"90",X"48",X"64",X"98",X"80",X"00",X"00",
		X"20",X"90",X"C8",X"E4",X"F2",X"69",X"34",X"62",X"EB",X"F7",X"22",X"22",X"F7",X"EB",X"63",X"36",
		X"00",X"F0",X"0C",X"00",X"E4",X"E0",X"E0",X"0C",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"C3",X"C0",X"C8",X"C7",X"C1",X"C8",X"C6",X"C3",X"FA",X"FA",X"0A",X"3E",X"3A",X"44",X"20",
		X"00",X"04",X"D4",X"54",X"34",X"79",X"F9",X"E0",X"80",X"C4",X"64",X"34",X"90",X"E0",X"60",X"00",
		X"00",X"80",X"80",X"0E",X"86",X"07",X"07",X"FF",X"FF",X"FF",X"06",X"03",X"C1",X"90",X"00",X"00",
		X"80",X"80",X"80",X"80",X"BC",X"44",X"44",X"FC",X"90",X"B0",X"60",X"C0",X"80",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"E3",X"F7",X"88",X"FF",X"88",X"00",X"00",X"39",X"3F",X"06",X"28",
		X"02",X"15",X"6C",X"E2",X"F2",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"70",X"00",X"80",X"80",X"00",
		X"03",X"9E",X"BE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",X"9F",X"81",X"00",X"00",
		X"E0",X"60",X"70",X"60",X"60",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"83",X"21",X"01",X"09",X"09",X"07",X"9F",X"03",X"06",X"06",X"06",X"1E",X"1E",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"78",X"3E",X"06",X"00",X"00",X"00",X"81",X"C3",X"7E",X"3C",
		X"80",X"80",X"80",X"B0",X"BE",X"8F",X"81",X"80",X"80",X"80",X"C0",X"71",X"3F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"00",
		X"C0",X"80",X"90",X"AE",X"83",X"80",X"80",X"80",X"80",X"C0",X"70",X"0E",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"78",X"3E",X"06",X"00",X"00",X"00",X"81",X"C3",X"7E",X"3C",
		X"80",X"80",X"80",X"F0",X"7E",X"0F",X"01",X"00",X"00",X"80",X"80",X"81",X"8E",X"80",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"00",X"01",X"FE",X"00",X"00",X"00",X"C0",X"38",X"07",
		X"00",X"80",X"80",X"70",X"0E",X"01",X"00",X"02",X"10",X"80",X"80",X"70",X"0E",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"F0",X"7E",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"78",X"3C",X"06",X"82",X"02",X"02",X"02",X"02",X"03",X"00",
		X"80",X"80",X"80",X"B0",X"BE",X"8F",X"83",X"81",X"81",X"81",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"24",X"20",X"3C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"00",X"04",X"04",X"04",X"04",X"C0",X"F8",X"3C",X"07",X"03",X"00",
		X"10",X"20",X"4E",X"9F",X"91",X"80",X"C0",X"C0",X"70",X"3E",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"78",X"3E",X"06",X"00",X"00",X"00",X"81",X"C3",X"7E",X"3C",
		X"80",X"80",X"80",X"F0",X"3E",X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"07",X"1F",X"18",X"C0",X"C0",X"00",X"00",X"C0",X"F8",X"3F",
		X"80",X"80",X"F0",X"FE",X"0F",X"00",X"03",X"06",X"03",X"80",X"80",X"F0",X"FE",X"0F",X"01",X"00",
		X"00",X"00",X"08",X"08",X"F8",X"08",X"08",X"00",X"F8",X"10",X"20",X"10",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"81",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",
		X"00",X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
