library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_3H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_3H is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"5F",X"16",X"00",X"19",X"C9",X"FF",X"FF",
		X"DF",X"EB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"5E",X"23",X"56",X"23",X"C9",X"FF",X"FF",X"FF",
		X"E1",X"CF",X"D7",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"7E",X"23",
		X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"D9",X"21",X"90",X"43",X"CB",X"C6",X"3A",X"00",X"60",
		X"32",X"91",X"43",X"D9",X"08",X"ED",X"45",X"31",X"00",X"44",X"3A",X"00",X"60",X"21",X"00",X"40",
		X"01",X"00",X"04",X"36",X"00",X"23",X"0B",X"78",X"B1",X"20",X"F8",X"CD",X"9F",X"00",X"CD",X"37",
		X"01",X"CD",X"9B",X"04",X"21",X"90",X"43",X"CB",X"46",X"28",X"FC",X"CB",X"86",X"18",X"EC",X"3A",
		X"91",X"43",X"B7",X"C8",X"FE",X"10",X"30",X"09",X"3D",X"21",X"AF",X"00",X"CF",X"D7",X"E9",X"77",
		X"00",X"0E",X"00",X"D6",X"10",X"CB",X"7F",X"28",X"03",X"0C",X"E6",X"7F",X"21",X"B2",X"06",X"CF",
		X"D7",X"7E",X"23",X"FD",X"21",X"00",X"40",X"B7",X"28",X"04",X"FD",X"21",X"B0",X"41",X"0D",X"28",
		X"44",X"7E",X"FE",X"FF",X"C8",X"23",X"DF",X"E5",X"6F",X"26",X"00",X"29",X"29",X"29",X"29",X"4D",
		X"44",X"29",X"09",X"4D",X"44",X"FD",X"E5",X"DD",X"E1",X"DD",X"09",X"DD",X"36",X"00",X"80",X"DD",
		X"73",X"0C",X"DD",X"72",X"0D",X"21",X"02",X"06",X"DF",X"DD",X"73",X"10",X"DD",X"72",X"11",X"DD",
		X"36",X"01",X"03",X"DD",X"36",X"2C",X"40",X"DD",X"36",X"2D",X"00",X"DD",X"36",X"0A",X"00",X"CD",
		X"CF",X"01",X"E1",X"18",X"BC",X"7E",X"FE",X"FF",X"C8",X"23",X"23",X"23",X"E5",X"6F",X"26",X"00",
		X"29",X"29",X"29",X"29",X"5D",X"54",X"29",X"19",X"EB",X"FD",X"E5",X"E1",X"19",X"06",X"30",X"36",
		X"00",X"23",X"10",X"FB",X"E1",X"18",X"DE",X"06",X"12",X"DD",X"21",X"00",X"40",X"C5",X"3E",X"12",
		X"90",X"32",X"92",X"43",X"DD",X"CB",X"00",X"7E",X"C4",X"54",X"01",X"11",X"30",X"00",X"DD",X"19",
		X"C1",X"10",X"EA",X"C9",X"DD",X"6E",X"14",X"DD",X"66",X"15",X"2B",X"DD",X"75",X"14",X"DD",X"74",
		X"15",X"7C",X"B5",X"CC",X"CF",X"01",X"DD",X"CB",X"00",X"5E",X"28",X"09",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"03",X"00",X"C9",X"DD",X"CB",X"00",X"56",X"28",X"15",X"DD",X"6E",X"28",X"DD",X"66",
		X"29",X"2B",X"DD",X"75",X"28",X"DD",X"74",X"29",X"7C",X"B5",X"20",X"04",X"DD",X"CB",X"00",X"96",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"19",X"DD",X"75",X"02",
		X"DD",X"74",X"03",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"08",X"DD",X"56",X"09",X"19",
		X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"CB",X"00",X"76",X"C0",X"DD",X"6E",X"0E",X"DD",X"66",
		X"0F",X"2B",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"7D",X"B4",X"C0",X"CD",X"D1",X"03",X"C9",X"DD",
		X"CB",X"00",X"76",X"C2",X"35",X"04",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"DD",X"7E",
		X"00",X"E6",X"E6",X"DD",X"77",X"00",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"DD",X"75",X"16",X"DD",
		X"74",X"17",X"DD",X"6E",X"2E",X"DD",X"66",X"2F",X"DD",X"75",X"14",X"DD",X"74",X"15",X"FF",X"FE",
		X"80",X"30",X"59",X"DD",X"CB",X"00",X"46",X"28",X"10",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"2B",
		X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C3",X"AE",X"02",X"DD",X"CB",X"00",X"C6",X"47",X"E6",X"0F",
		X"FE",X"0C",X"20",X"06",X"DD",X"CB",X"00",X"DE",X"18",X"D4",X"21",X"B0",X"05",X"CF",X"DF",X"CB",
		X"38",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"DD",X"7E",X"01",X"CB",X"2F",X"CB",X"2F",X"80",X"28",
		X"13",X"47",X"FE",X"08",X"38",X"08",X"DD",X"CB",X"01",X"46",X"20",X"08",X"06",X"07",X"CB",X"3A",
		X"CB",X"1B",X"10",X"FA",X"DD",X"73",X"06",X"DD",X"72",X"07",X"18",X"A2",X"FE",X"F0",X"38",X"27",
		X"E6",X"0F",X"21",X"FE",X"01",X"E5",X"E7",X"08",X"03",X"0D",X"03",X"1A",X"03",X"28",X"03",X"38",
		X"03",X"46",X"03",X"56",X"03",X"6D",X"03",X"72",X"03",X"77",X"03",X"7C",X"03",X"87",X"03",X"9B",
		X"03",X"A4",X"03",X"AD",X"03",X"B5",X"03",X"E6",X"7F",X"21",X"E0",X"05",X"CF",X"DF",X"DD",X"6E",
		X"2C",X"DD",X"66",X"2D",X"CD",X"17",X"04",X"06",X"06",X"CB",X"3C",X"CB",X"1D",X"10",X"FA",X"DD",
		X"75",X"14",X"DD",X"74",X"15",X"DD",X"75",X"2E",X"DD",X"74",X"2F",X"C3",X"FE",X"01",X"DD",X"6E",
		X"10",X"DD",X"66",X"11",X"DF",X"DD",X"73",X"02",X"DD",X"72",X"03",X"DD",X"75",X"12",X"DD",X"74",
		X"13",X"CD",X"D1",X"03",X"DD",X"CB",X"00",X"66",X"20",X"05",X"DD",X"CB",X"00",X"6E",X"C8",X"DD",
		X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"17",X"DD",X"56",X"18",X"DD",X"4E",X"14",X"DD",X"46",
		X"15",X"CD",X"EB",X"02",X"DD",X"75",X"08",X"DD",X"74",X"09",X"C9",X"B7",X"ED",X"52",X"30",X"08",
		X"EB",X"21",X"00",X"00",X"B7",X"ED",X"52",X"37",X"F5",X"59",X"50",X"CD",X"F8",X"03",X"F1",X"D0",
		X"EB",X"21",X"00",X"00",X"B7",X"ED",X"52",X"C9",X"FF",X"DD",X"77",X"01",X"C9",X"FF",X"21",X"02",
		X"06",X"CF",X"D7",X"DD",X"75",X"10",X"DD",X"74",X"11",X"C9",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",
		X"DF",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"C9",X"CD",X"C1",X"03",X"E5",X"CD",X"1A",X"03",X"EB",
		X"E1",X"73",X"23",X"72",X"DD",X"34",X"0A",X"C9",X"DD",X"35",X"0A",X"CD",X"C1",X"03",X"DF",X"DD",
		X"73",X"0C",X"DD",X"72",X"0D",X"C9",X"FF",X"DD",X"77",X"0B",X"E5",X"CD",X"C1",X"03",X"D1",X"73",
		X"23",X"72",X"DD",X"34",X"0A",X"C9",X"DD",X"35",X"0A",X"DD",X"35",X"0B",X"20",X"01",X"C9",X"CD",
		X"C1",X"03",X"DD",X"34",X"0A",X"DF",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"C9",X"DD",X"CB",X"00",
		X"E6",X"C9",X"DD",X"CB",X"00",X"EE",X"C9",X"DD",X"CB",X"00",X"AE",X"C9",X"FF",X"87",X"47",X"DD",
		X"7E",X"01",X"B0",X"DD",X"77",X"01",X"C9",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"DF",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"73",X"2C",X"DD",X"72",X"2D",X"C9",X"DD",X"7E",X"01",X"E6",X"03",
		X"DD",X"77",X"01",X"C9",X"DD",X"36",X"2C",X"40",X"DD",X"36",X"2D",X"00",X"C9",X"DD",X"CB",X"00",
		X"F6",X"E1",X"C3",X"35",X"04",X"E1",X"DD",X"E5",X"E1",X"06",X"20",X"36",X"00",X"23",X"10",X"FB",
		X"C9",X"DD",X"E5",X"E1",X"11",X"18",X"00",X"19",X"DD",X"7E",X"0A",X"87",X"5F",X"16",X"00",X"19",
		X"C9",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"DF",X"4B",X"42",X"DD",X"73",X"0E",X"DD",X"72",X"0F",
		X"DF",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"EB",X"CD",X"EB",
		X"02",X"DD",X"75",X"04",X"DD",X"74",X"05",X"C9",X"F5",X"C5",X"EB",X"4D",X"44",X"21",X"00",X"00",
		X"3E",X"10",X"EB",X"29",X"EB",X"ED",X"6A",X"B7",X"ED",X"42",X"30",X"03",X"09",X"18",X"01",X"13",
		X"3D",X"20",X"EF",X"EB",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"4D",X"44",X"21",X"00",X"00",X"7A",
		X"B3",X"28",X"0E",X"CB",X"38",X"CB",X"19",X"30",X"01",X"19",X"EB",X"29",X"EB",X"79",X"B0",X"20",
		X"F2",X"D1",X"C1",X"F1",X"C9",X"FF",X"CB",X"7F",X"28",X"07",X"DD",X"CB",X"00",X"B6",X"C3",X"CF",
		X"01",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"DF",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"73",
		X"14",X"DD",X"72",X"15",X"CB",X"47",X"28",X"07",X"DF",X"DD",X"73",X"06",X"DD",X"72",X"07",X"CB",
		X"4F",X"28",X"07",X"DF",X"DD",X"73",X"08",X"DD",X"72",X"09",X"CB",X"57",X"28",X"07",X"DF",X"DD",
		X"73",X"02",X"DD",X"72",X"03",X"CB",X"5F",X"28",X"07",X"DF",X"DD",X"73",X"04",X"DD",X"72",X"05",
		X"CB",X"67",X"28",X"10",X"7E",X"DD",X"77",X"2A",X"23",X"DF",X"DD",X"73",X"28",X"DD",X"72",X"29",
		X"DD",X"CB",X"00",X"D6",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",X"DD",X"21",X"B0",X"41",X"FD",
		X"21",X"60",X"43",X"06",X"03",X"C5",X"DD",X"E5",X"CD",X"F6",X"04",X"FD",X"71",X"07",X"11",X"50",
		X"FE",X"DD",X"19",X"CD",X"F6",X"04",X"FD",X"7E",X"07",X"B1",X"2F",X"FD",X"77",X"07",X"DD",X"E1",
		X"C1",X"11",X"90",X"00",X"DD",X"19",X"11",X"10",X"00",X"FD",X"19",X"10",X"D8",X"21",X"60",X"43",
		X"0E",X"00",X"CD",X"E6",X"04",X"21",X"70",X"43",X"0E",X"10",X"CD",X"E6",X"04",X"21",X"80",X"43",
		X"0E",X"80",X"CD",X"E6",X"04",X"C9",X"06",X"10",X"3E",X"10",X"90",X"ED",X"79",X"0C",X"7E",X"23",
		X"ED",X"79",X"0D",X"10",X"F3",X"C9",X"0E",X"00",X"DD",X"CB",X"00",X"7E",X"28",X"25",X"CB",X"C1",
		X"11",X"00",X"00",X"CD",X"8F",X"05",X"FD",X"75",X"00",X"FD",X"74",X"01",X"FD",X"77",X"08",X"DD",
		X"7E",X"01",X"E6",X"03",X"47",X"DD",X"CB",X"00",X"56",X"28",X"08",X"CB",X"D9",X"DD",X"7E",X"2A",
		X"FD",X"77",X"06",X"DD",X"CB",X"30",X"7E",X"28",X"28",X"CB",X"C9",X"11",X"30",X"00",X"CD",X"8F",
		X"05",X"FD",X"75",X"02",X"FD",X"74",X"03",X"FD",X"77",X"09",X"DD",X"7E",X"31",X"87",X"87",X"E6",
		X"0C",X"B0",X"47",X"DD",X"CB",X"30",X"56",X"28",X"08",X"CB",X"E1",X"DD",X"7E",X"58",X"FD",X"77",
		X"06",X"DD",X"CB",X"60",X"7E",X"28",X"34",X"CB",X"D1",X"11",X"60",X"00",X"CD",X"8F",X"05",X"FD",
		X"75",X"04",X"FD",X"74",X"05",X"FD",X"77",X"0A",X"DD",X"7E",X"61",X"87",X"87",X"87",X"87",X"E6",
		X"30",X"B0",X"47",X"DD",X"CB",X"60",X"56",X"28",X"12",X"CB",X"E9",X"11",X"88",X"00",X"DD",X"19",
		X"DD",X"7E",X"00",X"11",X"78",X"FF",X"DD",X"19",X"FD",X"77",X"06",X"FD",X"70",X"0E",X"C9",X"C5",
		X"DD",X"19",X"21",X"00",X"00",X"B7",X"ED",X"52",X"EB",X"DD",X"7E",X"03",X"DD",X"6E",X"06",X"DD",
		X"66",X"07",X"DD",X"19",X"06",X"04",X"CB",X"3F",X"CB",X"3C",X"CB",X"1D",X"10",X"F8",X"C1",X"C9",
		X"2B",X"B3",X"1D",X"A9",X"9F",X"9F",X"A9",X"96",X"35",X"8E",X"39",X"86",X"B1",X"7E",X"95",X"77",
		X"DE",X"70",X"89",X"6A",X"8E",X"64",X"E9",X"5E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"02",X"00",X"04",X"00",X"06",X"00",X"08",X"00",X"0C",X"00",X"10",X"00",X"18",X"00",
		X"20",X"00",X"30",X"00",X"40",X"00",X"60",X"00",X"80",X"00",X"C0",X"00",X"00",X"01",X"80",X"01",
		X"00",X"02",X"18",X"06",X"26",X"06",X"34",X"06",X"42",X"06",X"50",X"06",X"5E",X"06",X"6C",X"06",
		X"7A",X"06",X"88",X"06",X"96",X"06",X"A4",X"06",X"FF",X"FF",X"02",X"00",X"FF",X"FF",X"08",X"00",
		X"00",X"80",X"0A",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"FF",X"FF",X"08",X"00",X"00",X"80",
		X"14",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"FF",X"FF",X"3C",X"00",X"FF",X"FF",X"80",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"F0",X"00",X"00",X"80",X"F0",X"00",X"01",X"00",
		X"01",X"00",X"0A",X"00",X"00",X"F0",X"0A",X"00",X"00",X"80",X"14",X"00",X"01",X"00",X"FF",X"FF",
		X"02",X"00",X"FF",X"FF",X"14",X"00",X"00",X"60",X"32",X"00",X"00",X"00",X"00",X"80",X"02",X"00",
		X"FF",X"FF",X"08",X"00",X"00",X"80",X"1E",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"FF",X"FF",
		X"3C",X"00",X"00",X"80",X"B0",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"FF",X"FF",X"1E",X"00",
		X"00",X"80",X"60",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"FF",X"FF",X"60",X"00",X"00",X"80",
		X"3C",X"00",X"00",X"00",X"00",X"50",X"04",X"00",X"FF",X"FF",X"B0",X"00",X"00",X"80",X"A0",X"00",
		X"00",X"50",X"F2",X"06",X"3A",X"07",X"F0",X"06",X"8A",X"07",X"BE",X"07",X"D1",X"07",X"F8",X"07",
		X"50",X"08",X"8C",X"08",X"B6",X"08",X"87",X"17",X"00",X"09",X"F0",X"06",X"A2",X"09",X"FA",X"09",
		X"1E",X"0A",X"02",X"0B",X"F0",X"06",X"82",X"0C",X"38",X"0D",X"D7",X"13",X"0E",X"16",X"D7",X"16",
		X"44",X"0A",X"4F",X"18",X"E7",X"1A",X"A9",X"19",X"4F",X"1D",X"92",X"0A",X"CA",X"0A",X"1E",X"1E",
		X"00",X"FF",X"00",X"07",X"FA",X"06",X"08",X"1A",X"07",X"FF",X"F0",X"03",X"F1",X"03",X"FA",X"01",
		X"FB",X"40",X"00",X"20",X"80",X"24",X"27",X"30",X"34",X"37",X"40",X"44",X"47",X"50",X"54",X"57",
		X"60",X"64",X"80",X"F1",X"08",X"69",X"80",X"70",X"88",X"FF",X"F0",X"03",X"F1",X"00",X"FA",X"01",
		X"FB",X"40",X"00",X"21",X"80",X"25",X"28",X"31",X"35",X"38",X"41",X"45",X"48",X"51",X"55",X"58",
		X"61",X"65",X"80",X"F1",X"08",X"6A",X"80",X"71",X"86",X"FF",X"00",X"05",X"42",X"07",X"06",X"66",
		X"07",X"FF",X"FE",X"0F",X"05",X"00",X"00",X"10",X"00",X"FE",X"FF",X"FF",X"00",X"FF",X"0F",X"05",
		X"00",X"00",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"0F",X"20",X"00",X"00",X"05",X"F0",X"FF",
		X"FF",X"FF",X"00",X"F9",X"80",X"FF",X"FE",X"0F",X"05",X"00",X"00",X"12",X"00",X"FF",X"FF",X"FF",
		X"00",X"F9",X"0F",X"05",X"00",X"00",X"0B",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"0F",X"20",X"00",
		X"00",X"07",X"F0",X"FF",X"FF",X"FF",X"DD",X"F9",X"80",X"FF",X"01",X"05",X"92",X"07",X"06",X"A8",
		X"07",X"FF",X"F0",X"03",X"F1",X"05",X"FA",X"01",X"FB",X"10",X"00",X"F8",X"60",X"86",X"0C",X"84",
		X"50",X"86",X"0C",X"84",X"F2",X"92",X"07",X"FF",X"F0",X"03",X"F1",X"05",X"FA",X"01",X"FB",X"10",
		X"00",X"F8",X"61",X"86",X"0C",X"84",X"51",X"86",X"0C",X"84",X"F2",X"B1",X"07",X"FF",X"00",X"05",
		X"C3",X"07",X"FF",X"F8",X"50",X"82",X"54",X"57",X"60",X"64",X"67",X"82",X"F1",X"03",X"69",X"90",
		X"FF",X"01",X"07",X"D9",X"07",X"08",X"EA",X"07",X"FF",X"FB",X"1F",X"10",X"00",X"00",X"10",X"00",
		X"00",X"FF",X"FF",X"00",X"10",X"15",X"10",X"00",X"80",X"FF",X"FE",X"0F",X"10",X"00",X"00",X"05",
		X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"00",X"07",X"00",X"08",X"08",X"28",X"08",X"FF",
		X"F0",X"03",X"F1",X"0C",X"FA",X"01",X"FB",X"30",X"00",X"70",X"84",X"6B",X"60",X"5B",X"82",X"5A",
		X"59",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4B",X"4A",X"49",X"48",X"47",X"46",
		X"45",X"44",X"43",X"42",X"41",X"40",X"82",X"FF",X"F0",X"03",X"F1",X"0C",X"FA",X"01",X"FB",X"30",
		X"00",X"6B",X"84",X"6A",X"6B",X"5A",X"82",X"59",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",
		X"50",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"40",X"3B",X"82",X"FF",
		X"01",X"07",X"58",X"08",X"08",X"7C",X"08",X"FF",X"FE",X"0F",X"03",X"00",X"00",X"25",X"FF",X"FF",
		X"FF",X"FF",X"00",X"F2",X"0F",X"03",X"00",X"00",X"20",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"0F",
		X"20",X"00",X"00",X"20",X"FC",X"FF",X"FF",X"FF",X"00",X"FB",X"80",X"FF",X"FE",X"0F",X"0A",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"FF",X"FF",X"FF",X"F9",X"80",X"FF",X"00",X"05",X"94",X"08",
		X"06",X"A5",X"08",X"FF",X"F5",X"03",X"FE",X"0F",X"06",X"00",X"00",X"03",X"C0",X"FF",X"DD",X"DD",
		X"00",X"FF",X"80",X"F6",X"FF",X"F5",X"03",X"FE",X"0F",X"06",X"00",X"00",X"03",X"D0",X"FF",X"DD",
		X"DD",X"00",X"FF",X"80",X"F6",X"FF",X"00",X"05",X"BE",X"08",X"06",X"D1",X"08",X"FF",X"FE",X"0F",
		X"10",X"00",X"00",X"02",X"E0",X"FF",X"DD",X"DD",X"00",X"EF",X"F0",X"03",X"F1",X"00",X"71",X"85",
		X"FF",X"FE",X"0F",X"03",X"00",X"00",X"04",X"00",X"00",X"DD",X"DD",X"FF",X"E0",X"0F",X"03",X"00",
		X"00",X"03",X"00",X"00",X"FF",X"FF",X"FF",X"E0",X"0F",X"03",X"00",X"00",X"02",X"00",X"00",X"FF",
		X"FF",X"FF",X"E0",X"0F",X"05",X"00",X"00",X"03",X"00",X"00",X"FF",X"FF",X"FF",X"E0",X"80",X"FF",
		X"00",X"00",X"0E",X"09",X"01",X"4A",X"09",X"02",X"82",X"09",X"03",X"92",X"09",X"FF",X"F0",X"00",
		X"F1",X"02",X"FA",X"01",X"FB",X"20",X"00",X"40",X"82",X"41",X"42",X"43",X"44",X"45",X"46",X"47",
		X"48",X"49",X"4A",X"4B",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"59",
		X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",
		X"44",X"43",X"42",X"41",X"40",X"82",X"F2",X"0E",X"09",X"FF",X"F0",X"00",X"F1",X"03",X"FA",X"01",
		X"FB",X"20",X"00",X"60",X"82",X"61",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"70",
		X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"79",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",
		X"72",X"71",X"70",X"6B",X"6A",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"82",X"F2",X"4A",
		X"09",X"FF",X"FE",X"0F",X"09",X"00",X"00",X"03",X"E0",X"FF",X"DD",X"DD",X"FF",X"FF",X"80",X"F2",
		X"82",X"09",X"FE",X"0F",X"09",X"00",X"00",X"05",X"E0",X"FF",X"DD",X"DD",X"FF",X"FF",X"80",X"F2",
		X"92",X"09",X"00",X"07",X"B0",X"09",X"08",X"C1",X"09",X"04",X"D4",X"09",X"05",X"E7",X"09",X"FF",
		X"F1",X"08",X"FB",X"10",X"00",X"65",X"83",X"63",X"61",X"63",X"82",X"65",X"80",X"67",X"69",X"86",
		X"FF",X"F1",X"08",X"FB",X"10",X"00",X"61",X"83",X"5B",X"82",X"59",X"83",X"5B",X"82",X"61",X"81",
		X"63",X"65",X"86",X"FF",X"F1",X"08",X"FB",X"10",X"00",X"0C",X"88",X"65",X"83",X"63",X"61",X"63",
		X"82",X"65",X"81",X"67",X"69",X"86",X"FF",X"F1",X"08",X"FB",X"10",X"00",X"0C",X"88",X"61",X"83",
		X"5B",X"59",X"5B",X"82",X"61",X"81",X"63",X"65",X"86",X"FF",X"00",X"05",X"02",X"0A",X"06",X"10",
		X"0A",X"FF",X"FE",X"0F",X"10",X"00",X"00",X"05",X"C0",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"FF",
		X"FE",X"0F",X"09",X"00",X"00",X"04",X"C0",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"FF",X"00",X"04",
		X"26",X"0A",X"08",X"35",X"0A",X"FF",X"F1",X"01",X"FB",X"30",X"00",X"F8",X"60",X"86",X"70",X"88",
		X"69",X"85",X"67",X"83",X"FF",X"F1",X"02",X"FB",X"30",X"00",X"F8",X"50",X"86",X"60",X"88",X"70",
		X"85",X"71",X"83",X"FF",X"00",X"00",X"4C",X"0A",X"01",X"73",X"0A",X"FF",X"F5",X"02",X"F1",X"08",
		X"FB",X"15",X"00",X"57",X"84",X"54",X"56",X"82",X"58",X"59",X"5B",X"61",X"63",X"65",X"67",X"83",
		X"69",X"82",X"F6",X"FE",X"1F",X"80",X"00",X"00",X"03",X"FC",X"FF",X"FF",X"FF",X"FE",X"FF",X"10",
		X"80",X"00",X"FF",X"FE",X"1F",X"0B",X"00",X"00",X"04",X"C0",X"FF",X"FF",X"FF",X"F0",X"FF",X"08",
		X"10",X"00",X"1F",X"20",X"00",X"00",X"02",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"05",X"09",X"00",
		X"80",X"FF",X"00",X"07",X"9A",X"0A",X"08",X"B9",X"0A",X"FF",X"FE",X"1F",X"0B",X"00",X"00",X"04",
		X"C0",X"FF",X"FF",X"FF",X"F0",X"FF",X"08",X"10",X"00",X"1F",X"40",X"00",X"00",X"02",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"05",X"40",X"00",X"80",X"FF",X"FE",X"1F",X"20",X"00",X"00",X"05",X"00",
		X"00",X"FF",X"FF",X"00",X"F8",X"10",X"20",X"00",X"80",X"FF",X"00",X"07",X"D2",X"0A",X"08",X"EC",
		X"0A",X"FF",X"F1",X"0C",X"FA",X"03",X"FB",X"40",X"00",X"20",X"80",X"24",X"27",X"30",X"34",X"37",
		X"40",X"44",X"47",X"50",X"54",X"57",X"60",X"64",X"67",X"70",X"82",X"FF",X"F1",X"0C",X"FA",X"03",
		X"FB",X"40",X"00",X"70",X"80",X"67",X"64",X"60",X"57",X"54",X"57",X"60",X"30",X"27",X"24",X"20",
		X"80",X"FF",X"00",X"00",X"13",X"0B",X"01",X"5C",X"0B",X"02",X"A5",X"0B",X"03",X"EE",X"0B",X"04",
		X"37",X"0C",X"FF",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"20",X"00",X"54",X"86",X"57",X"0C",
		X"50",X"54",X"0C",X"49",X"50",X"0C",X"49",X"50",X"0C",X"49",X"0C",X"47",X"0C",X"52",X"55",X"0C",
		X"4B",X"52",X"0C",X"47",X"4B",X"0C",X"47",X"4B",X"0C",X"50",X"0C",X"52",X"0C",X"49",X"48",X"49",
		X"4B",X"50",X"4B",X"50",X"52",X"54",X"0C",X"57",X"59",X"0C",X"57",X"54",X"50",X"57",X"52",X"0C",
		X"55",X"54",X"52",X"50",X"4B",X"54",X"88",X"0C",X"50",X"0C",X"88",X"FF",X"F0",X"03",X"F1",X"00",
		X"FA",X"00",X"FB",X"20",X"00",X"44",X"86",X"47",X"0C",X"40",X"44",X"0C",X"39",X"40",X"0C",X"39",
		X"40",X"0C",X"39",X"0C",X"37",X"0C",X"42",X"45",X"0C",X"3B",X"42",X"0C",X"37",X"3B",X"0C",X"37",
		X"3B",X"0C",X"40",X"0C",X"42",X"0C",X"39",X"38",X"39",X"3B",X"40",X"3B",X"40",X"42",X"44",X"0C",
		X"47",X"49",X"0C",X"47",X"44",X"40",X"47",X"42",X"0C",X"45",X"44",X"42",X"40",X"3B",X"44",X"88",
		X"0C",X"40",X"0C",X"88",X"FF",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"20",X"00",X"50",X"86",
		X"54",X"0C",X"49",X"50",X"0C",X"45",X"49",X"0C",X"45",X"49",X"0C",X"45",X"0C",X"44",X"0C",X"4B",
		X"52",X"0C",X"47",X"4B",X"0C",X"42",X"45",X"0C",X"42",X"47",X"0C",X"49",X"0C",X"4B",X"0C",X"45",
		X"44",X"45",X"47",X"49",X"48",X"49",X"4B",X"50",X"0C",X"54",X"55",X"0C",X"54",X"50",X"49",X"54",
		X"4B",X"0C",X"52",X"50",X"4B",X"49",X"47",X"50",X"88",X"0C",X"47",X"0C",X"88",X"FF",X"F0",X"03",
		X"F1",X"00",X"FA",X"00",X"FB",X"20",X"00",X"40",X"86",X"44",X"0C",X"39",X"40",X"0C",X"35",X"39",
		X"0C",X"39",X"35",X"0C",X"35",X"0C",X"34",X"0C",X"3B",X"42",X"0C",X"37",X"3B",X"0C",X"32",X"35",
		X"0C",X"32",X"37",X"0C",X"39",X"0C",X"3B",X"0C",X"35",X"34",X"35",X"37",X"39",X"38",X"39",X"3B",
		X"45",X"0C",X"44",X"45",X"0C",X"44",X"40",X"39",X"44",X"3B",X"0C",X"42",X"40",X"3B",X"39",X"37",
		X"40",X"88",X"0C",X"37",X"0C",X"88",X"FF",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"20",X"00",
		X"24",X"86",X"0C",X"27",X"0C",X"24",X"24",X"27",X"0C",X"20",X"0C",X"24",X"0C",X"20",X"20",X"24",
		X"0C",X"22",X"0C",X"25",X"0C",X"22",X"22",X"25",X"0C",X"1B",X"0C",X"22",X"0C",X"1B",X"1B",X"22",
		X"0C",X"19",X"0C",X"17",X"0C",X"15",X"0C",X"14",X"0C",X"15",X"0C",X"17",X"0C",X"19",X"0C",X"1B",
		X"0C",X"20",X"0C",X"24",X"0C",X"1B",X"1B",X"22",X"0C",X"20",X"20",X"24",X"0C",X"20",X"88",X"0C",
		X"88",X"FF",X"01",X"00",X"90",X"0C",X"01",X"BD",X"0C",X"02",X"EA",X"0C",X"03",X"17",X"0D",X"FF",
		X"F0",X"01",X"F1",X"05",X"FA",X"00",X"FB",X"28",X"00",X"54",X"87",X"47",X"84",X"54",X"87",X"47",
		X"84",X"52",X"87",X"45",X"84",X"52",X"87",X"45",X"84",X"50",X"87",X"44",X"84",X"50",X"87",X"44",
		X"84",X"50",X"86",X"0C",X"84",X"4B",X"50",X"87",X"52",X"84",X"F2",X"AE",X"0D",X"F0",X"01",X"F1",
		X"05",X"FA",X"00",X"FB",X"28",X"00",X"50",X"87",X"44",X"84",X"50",X"87",X"44",X"84",X"4B",X"87",
		X"42",X"84",X"4B",X"87",X"42",X"84",X"47",X"87",X"40",X"84",X"47",X"87",X"40",X"84",X"47",X"86",
		X"0C",X"84",X"47",X"49",X"87",X"4B",X"84",X"F2",X"BA",X"0E",X"F0",X"01",X"F1",X"05",X"FA",X"00",
		X"FB",X"28",X"00",X"40",X"87",X"47",X"84",X"45",X"87",X"44",X"84",X"39",X"87",X"3B",X"84",X"40",
		X"87",X"42",X"84",X"37",X"87",X"39",X"84",X"3B",X"87",X"40",X"84",X"42",X"86",X"0C",X"84",X"42",
		X"44",X"87",X"45",X"84",X"F2",X"C7",X"0F",X"F0",X"01",X"F1",X"01",X"FA",X"00",X"FB",X"28",X"00",
		X"24",X"88",X"17",X"88",X"22",X"88",X"15",X"88",X"20",X"88",X"17",X"88",X"20",X"86",X"0C",X"84",
		X"1B",X"20",X"87",X"22",X"84",X"F2",X"D3",X"10",X"01",X"00",X"46",X"0D",X"01",X"5B",X"0D",X"02",
		X"73",X"0D",X"03",X"8B",X"0D",X"FF",X"F0",X"02",X"F1",X"08",X"FA",X"00",X"FB",X"30",X"00",X"55",
		X"88",X"54",X"52",X"50",X"49",X"8A",X"50",X"86",X"F2",X"87",X"11",X"F0",X"02",X"F1",X"08",X"FA",
		X"00",X"FB",X"30",X"00",X"0C",X"84",X"59",X"88",X"57",X"55",X"54",X"87",X"52",X"8A",X"57",X"86",
		X"F2",X"41",X"12",X"F0",X"02",X"F1",X"08",X"FA",X"00",X"FB",X"30",X"00",X"0C",X"86",X"60",X"88",
		X"5B",X"59",X"57",X"86",X"55",X"8A",X"57",X"86",X"F2",X"AF",X"12",X"F0",X"02",X"F1",X"07",X"FA",
		X"00",X"FB",X"30",X"00",X"17",X"88",X"15",X"14",X"12",X"10",X"8A",X"10",X"86",X"F2",X"21",X"13",
		X"01",X"00",X"AE",X"0D",X"01",X"BA",X"0E",X"02",X"C7",X"0F",X"03",X"D3",X"10",X"FF",X"F0",X"01",
		X"F1",X"05",X"FB",X"28",X"00",X"F3",X"DC",X"0D",X"F3",X"29",X"0E",X"F3",X"DC",X"0D",X"F3",X"37",
		X"0E",X"F3",X"3E",X"0E",X"F3",X"57",X"0E",X"F3",X"7C",X"0E",X"F3",X"95",X"0E",X"F3",X"3E",X"0E",
		X"F3",X"6A",X"0E",X"F3",X"7C",X"0E",X"F3",X"A7",X"0E",X"F2",X"AE",X"0D",X"54",X"87",X"53",X"84",
		X"54",X"87",X"53",X"84",X"54",X"86",X"50",X"0C",X"50",X"54",X"87",X"53",X"84",X"54",X"86",X"50",
		X"0C",X"50",X"0C",X"50",X"52",X"87",X"51",X"84",X"52",X"87",X"51",X"84",X"52",X"86",X"4B",X"0C",
		X"4B",X"52",X"87",X"51",X"84",X"52",X"86",X"4B",X"0C",X"4B",X"0C",X"4B",X"0C",X"88",X"50",X"4B",
		X"49",X"47",X"50",X"86",X"54",X"8A",X"0C",X"84",X"54",X"54",X"86",X"47",X"88",X"0C",X"84",X"54",
		X"52",X"86",X"45",X"88",X"0C",X"84",X"52",X"84",X"F4",X"50",X"88",X"4B",X"86",X"50",X"88",X"0C",
		X"84",X"4B",X"50",X"87",X"52",X"84",X"F4",X"50",X"88",X"50",X"4B",X"49",X"88",X"F4",X"54",X"87",
		X"53",X"84",X"54",X"87",X"53",X"84",X"54",X"86",X"4B",X"0C",X"4B",X"54",X"87",X"53",X"84",X"54",
		X"86",X"55",X"88",X"54",X"0C",X"86",X"F4",X"49",X"88",X"54",X"52",X"50",X"4B",X"86",X"50",X"88",
		X"49",X"88",X"0C",X"84",X"49",X"4B",X"87",X"50",X"84",X"F4",X"59",X"88",X"5B",X"60",X"86",X"5B",
		X"88",X"0C",X"84",X"59",X"89",X"0C",X"87",X"59",X"88",X"54",X"88",X"F4",X"52",X"87",X"51",X"84",
		X"52",X"87",X"51",X"84",X"52",X"86",X"49",X"0C",X"49",X"52",X"87",X"51",X"84",X"52",X"86",X"54",
		X"88",X"52",X"0C",X"86",X"F4",X"57",X"88",X"57",X"55",X"86",X"54",X"88",X"0C",X"84",X"52",X"89",
		X"0C",X"87",X"53",X"89",X"0C",X"86",X"F4",X"57",X"88",X"57",X"58",X"86",X"59",X"88",X"0C",X"86",
		X"5B",X"89",X"0C",X"84",X"4B",X"50",X"88",X"52",X"88",X"F4",X"F0",X"01",X"F1",X"05",X"FB",X"28",
		X"00",X"F3",X"E8",X"0E",X"F3",X"35",X"0F",X"F3",X"E8",X"0E",X"F3",X"43",X"0F",X"F3",X"4A",X"0F",
		X"F3",X"63",X"0F",X"F3",X"88",X"0F",X"F3",X"A1",X"0F",X"F3",X"4A",X"0F",X"F3",X"76",X"0F",X"F3",
		X"88",X"0F",X"F3",X"B3",X"0F",X"F2",X"BA",X"0E",X"50",X"87",X"4B",X"84",X"50",X"87",X"4B",X"84",
		X"50",X"86",X"49",X"0C",X"49",X"50",X"87",X"4B",X"84",X"50",X"86",X"47",X"0C",X"47",X"0C",X"47",
		X"4B",X"87",X"4A",X"84",X"4B",X"87",X"4A",X"84",X"4B",X"86",X"45",X"0C",X"45",X"4B",X"87",X"4A",
		X"84",X"4B",X"86",X"45",X"0C",X"45",X"0C",X"45",X"0C",X"88",X"49",X"47",X"45",X"44",X"47",X"86",
		X"50",X"8A",X"0C",X"84",X"50",X"50",X"86",X"44",X"88",X"0C",X"84",X"50",X"4B",X"86",X"42",X"88",
		X"0C",X"84",X"4B",X"84",X"F4",X"49",X"88",X"47",X"86",X"47",X"88",X"0C",X"84",X"47",X"49",X"87",
		X"4B",X"84",X"F4",X"47",X"88",X"47",X"47",X"45",X"88",X"F4",X"4B",X"87",X"4A",X"84",X"4B",X"87",
		X"4A",X"84",X"4B",X"86",X"48",X"0C",X"48",X"4B",X"87",X"4A",X"84",X"4B",X"86",X"50",X"88",X"4B",
		X"0C",X"86",X"F4",X"44",X"88",X"50",X"4B",X"49",X"47",X"86",X"49",X"88",X"44",X"0C",X"84",X"44",
		X"84",X"47",X"87",X"49",X"84",X"F4",X"54",X"88",X"57",X"59",X"86",X"57",X"88",X"0C",X"84",X"54",
		X"89",X"0C",X"87",X"54",X"88",X"49",X"88",X"F4",X"49",X"87",X"48",X"84",X"49",X"87",X"48",X"84",
		X"49",X"86",X"45",X"0C",X"45",X"49",X"87",X"48",X"84",X"49",X"86",X"50",X"88",X"49",X"0C",X"86",
		X"F4",X"54",X"88",X"54",X"52",X"86",X"50",X"88",X"0C",X"84",X"4B",X"89",X"0C",X"87",X"4A",X"89",
		X"0C",X"86",X"F4",X"52",X"88",X"52",X"54",X"86",X"55",X"88",X"0C",X"86",X"55",X"89",X"0C",X"84",
		X"47",X"84",X"49",X"88",X"4B",X"88",X"F4",X"F0",X"01",X"F1",X"00",X"FB",X"28",X"00",X"F3",X"F5",
		X"0F",X"F3",X"42",X"10",X"F3",X"F5",X"0F",X"F3",X"50",X"10",X"F3",X"57",X"10",X"F3",X"70",X"10",
		X"F3",X"94",X"10",X"F3",X"AD",X"10",X"F3",X"57",X"10",X"F3",X"82",X"10",X"F3",X"94",X"10",X"F3",
		X"BF",X"10",X"F2",X"C7",X"0F",X"44",X"87",X"43",X"84",X"44",X"87",X"43",X"84",X"44",X"86",X"40",
		X"0C",X"40",X"44",X"87",X"43",X"84",X"44",X"86",X"40",X"0C",X"40",X"0C",X"40",X"42",X"87",X"41",
		X"84",X"42",X"87",X"41",X"84",X"42",X"86",X"3B",X"0C",X"3B",X"42",X"87",X"41",X"84",X"42",X"86",
		X"3B",X"0C",X"3B",X"0C",X"3B",X"0C",X"88",X"40",X"3B",X"39",X"37",X"40",X"86",X"44",X"8A",X"0C",
		X"84",X"44",X"44",X"86",X"37",X"88",X"0C",X"84",X"44",X"42",X"86",X"45",X"88",X"0C",X"84",X"42",
		X"84",X"F4",X"40",X"88",X"3B",X"86",X"40",X"88",X"0C",X"84",X"3B",X"40",X"87",X"42",X"84",X"F4",
		X"40",X"88",X"40",X"3B",X"39",X"88",X"F4",X"44",X"87",X"43",X"84",X"44",X"87",X"43",X"84",X"44",
		X"86",X"3B",X"0C",X"3B",X"44",X"87",X"43",X"84",X"44",X"86",X"45",X"88",X"44",X"0C",X"86",X"F4",
		X"39",X"88",X"44",X"42",X"44",X"4B",X"86",X"40",X"88",X"39",X"0C",X"84",X"39",X"3B",X"87",X"40",
		X"84",X"F4",X"49",X"88",X"4B",X"50",X"86",X"4B",X"88",X"0C",X"84",X"49",X"89",X"0C",X"87",X"49",
		X"88",X"44",X"88",X"F4",X"42",X"87",X"41",X"84",X"42",X"87",X"41",X"84",X"42",X"86",X"49",X"0C",
		X"49",X"42",X"87",X"41",X"84",X"42",X"86",X"44",X"88",X"42",X"0C",X"86",X"F4",X"47",X"88",X"47",
		X"45",X"86",X"44",X"88",X"0C",X"84",X"42",X"89",X"0C",X"87",X"43",X"89",X"0C",X"86",X"F4",X"47",
		X"88",X"47",X"48",X"86",X"49",X"88",X"0C",X"86",X"4B",X"89",X"0C",X"84",X"3B",X"84",X"40",X"88",
		X"42",X"88",X"F4",X"F0",X"00",X"F1",X"01",X"FB",X"28",X"00",X"F3",X"01",X"11",X"F3",X"20",X"11",
		X"F3",X"01",X"11",X"F3",X"2D",X"11",X"F3",X"34",X"11",X"F3",X"3F",X"11",X"F3",X"55",X"11",X"F3",
		X"60",X"11",X"F3",X"34",X"11",X"F3",X"4A",X"11",X"F3",X"55",X"11",X"F3",X"6B",X"11",X"F2",X"D3",
		X"10",X"20",X"88",X"0C",X"17",X"0C",X"20",X"17",X"19",X"1B",X"19",X"0C",X"14",X"0C",X"19",X"14",
		X"15",X"17",X"20",X"0C",X"1B",X"0C",X"19",X"17",X"15",X"14",X"12",X"17",X"19",X"1B",X"88",X"F4",
		X"20",X"88",X"0C",X"89",X"0C",X"84",X"22",X"84",X"24",X"87",X"25",X"84",X"F4",X"20",X"88",X"20",
		X"1B",X"19",X"88",X"F4",X"24",X"88",X"0C",X"1B",X"0C",X"24",X"22",X"20",X"1B",X"88",X"F4",X"19",
		X"88",X"1B",X"20",X"1B",X"19",X"17",X"19",X"1B",X"88",X"F4",X"19",X"88",X"18",X"19",X"1B",X"20",
		X"0C",X"21",X"0C",X"88",X"F4",X"22",X"88",X"0C",X"19",X"0C",X"22",X"20",X"1B",X"19",X"88",X"F4",
		X"17",X"88",X"0C",X"1B",X"20",X"22",X"0C",X"23",X"0C",X"88",X"F4",X"17",X"89",X"17",X"86",X"1B",
		X"88",X"24",X"27",X"88",X"25",X"24",X"22",X"88",X"F4",X"01",X"00",X"87",X"11",X"01",X"41",X"12",
		X"02",X"AF",X"12",X"03",X"21",X"13",X"FF",X"F0",X"01",X"F1",X"00",X"FB",X"30",X"00",X"F3",X"A0",
		X"11",X"F3",X"B4",X"11",X"F3",X"A0",X"11",X"F3",X"C7",X"11",X"F3",X"E2",X"11",X"F2",X"87",X"11",
		X"40",X"86",X"42",X"44",X"47",X"45",X"44",X"45",X"47",X"45",X"44",X"45",X"4A",X"88",X"49",X"86",
		X"49",X"0C",X"86",X"F4",X"49",X"86",X"49",X"49",X"49",X"45",X"45",X"42",X"42",X"3A",X"3A",X"37",
		X"37",X"3A",X"42",X"40",X"0C",X"86",X"F4",X"52",X"86",X"52",X"52",X"52",X"49",X"49",X"45",X"45",
		X"42",X"45",X"49",X"50",X"88",X"49",X"86",X"45",X"0C",X"84",X"45",X"45",X"0C",X"45",X"86",X"0C",
		X"86",X"F4",X"39",X"88",X"40",X"47",X"89",X"45",X"86",X"44",X"45",X"40",X"39",X"40",X"84",X"0C",
		X"39",X"86",X"3A",X"40",X"3A",X"39",X"39",X"37",X"37",X"36",X"37",X"3A",X"47",X"8A",X"0C",X"3A",
		X"88",X"42",X"49",X"89",X"47",X"86",X"46",X"47",X"42",X"3A",X"42",X"84",X"0C",X"3A",X"86",X"40",
		X"42",X"44",X"42",X"42",X"40",X"40",X"42",X"44",X"40",X"49",X"8A",X"0C",X"88",X"40",X"50",X"0C",
		X"86",X"49",X"4A",X"49",X"88",X"4A",X"86",X"49",X"47",X"46",X"47",X"4A",X"88",X"0C",X"42",X"86",
		X"44",X"0C",X"42",X"44",X"0C",X"42",X"42",X"45",X"47",X"0C",X"45",X"47",X"8A",X"0C",X"0C",X"86",
		X"F4",X"F0",X"01",X"F1",X"00",X"FB",X"30",X"00",X"F3",X"5A",X"12",X"F3",X"6C",X"12",X"F3",X"5A",
		X"12",X"F3",X"74",X"12",X"F3",X"83",X"12",X"F2",X"41",X"12",X"0C",X"8A",X"35",X"86",X"0C",X"35",
		X"0C",X"35",X"0C",X"35",X"F5",X"08",X"0C",X"86",X"32",X"86",X"F6",X"F4",X"0C",X"86",X"34",X"0C",
		X"34",X"0C",X"86",X"F4",X"0C",X"86",X"34",X"0C",X"34",X"0C",X"84",X"40",X"40",X"0C",X"40",X"86",
		X"0C",X"86",X"F4",X"F5",X"08",X"0C",X"86",X"35",X"F6",X"F5",X"10",X"0C",X"32",X"F6",X"F5",X"04",
		X"0C",X"34",X"F6",X"F5",X"08",X"0C",X"35",X"F6",X"F5",X"04",X"0C",X"32",X"F6",X"3A",X"40",X"0C",
		X"3A",X"40",X"0C",X"3A",X"40",X"42",X"44",X"0C",X"42",X"44",X"8A",X"0C",X"0C",X"86",X"F4",X"F0",
		X"01",X"F1",X"00",X"FB",X"30",X"00",X"F3",X"C8",X"12",X"F3",X"D9",X"12",X"F3",X"C8",X"12",X"F3",
		X"E1",X"12",X"F3",X"F0",X"12",X"F2",X"AF",X"12",X"0C",X"8A",X"29",X"86",X"0C",X"29",X"F5",X"06",
		X"0C",X"29",X"F6",X"F5",X"04",X"0C",X"2A",X"F6",X"F4",X"0C",X"86",X"27",X"0C",X"27",X"0C",X"86",
		X"F4",X"0C",X"86",X"27",X"0C",X"27",X"0C",X"84",X"39",X"39",X"0C",X"39",X"86",X"0C",X"86",X"F4",
		X"F5",X"08",X"0C",X"86",X"29",X"F6",X"F5",X"08",X"0C",X"27",X"F6",X"F5",X"08",X"0C",X"2A",X"F6",
		X"F5",X"04",X"0C",X"27",X"F6",X"F5",X"08",X"0C",X"29",X"F6",X"F5",X"04",X"0C",X"27",X"F6",X"37",
		X"39",X"0C",X"37",X"39",X"0C",X"37",X"39",X"3A",X"40",X"0C",X"3A",X"40",X"8A",X"0C",X"0C",X"86",
		X"F4",X"F0",X"00",X"F1",X"00",X"FA",X"01",X"FB",X"30",X"00",X"F3",X"3C",X"13",X"F3",X"4F",X"13",
		X"F3",X"3C",X"13",X"F3",X"5E",X"13",X"F3",X"74",X"13",X"F2",X"21",X"13",X"10",X"86",X"12",X"14",
		X"15",X"88",X"10",X"10",X"09",X"12",X"09",X"12",X"86",X"12",X"15",X"19",X"1A",X"88",X"F4",X"15",
		X"88",X"1A",X"87",X"19",X"84",X"17",X"86",X"15",X"14",X"88",X"10",X"10",X"86",X"F4",X"12",X"88",
		X"1A",X"86",X"12",X"15",X"19",X"10",X"88",X"10",X"86",X"15",X"0C",X"84",X"15",X"15",X"0C",X"15",
		X"86",X"0C",X"86",X"F4",X"15",X"88",X"10",X"15",X"17",X"86",X"19",X"15",X"88",X"15",X"16",X"17",
		X"86",X"19",X"17",X"88",X"12",X"17",X"21",X"86",X"22",X"17",X"88",X"12",X"87",X"12",X"84",X"17",
		X"86",X"15",X"14",X"12",X"17",X"88",X"12",X"17",X"19",X"86",X"1A",X"17",X"88",X"12",X"0A",X"10",
		X"86",X"12",X"14",X"88",X"10",X"09",X"10",X"86",X"0A",X"09",X"88",X"05",X"09",X"07",X"86",X"09",
		X"07",X"09",X"0A",X"10",X"15",X"88",X"14",X"86",X"15",X"12",X"88",X"17",X"1A",X"86",X"17",X"14",
		X"12",X"0A",X"10",X"0C",X"0A",X"10",X"0C",X"0A",X"10",X"0A",X"10",X"0C",X"0A",X"10",X"8A",X"20",
		X"86",X"1A",X"17",X"14",X"10",X"86",X"F4",X"01",X"00",X"E5",X"13",X"01",X"1A",X"15",X"02",X"92",
		X"15",X"03",X"87",X"14",X"FF",X"F0",X"01",X"F1",X"05",X"FB",X"30",X"00",X"F3",X"0F",X"14",X"F3",
		X"2F",X"14",X"F3",X"2F",X"14",X"F0",X"02",X"F3",X"54",X"14",X"F3",X"6A",X"14",X"F3",X"54",X"14",
		X"F0",X"01",X"F1",X"08",X"F3",X"7D",X"14",X"F1",X"00",X"F3",X"2F",X"14",X"F2",X"E5",X"13",X"45",
		X"86",X"45",X"88",X"45",X"86",X"45",X"89",X"0C",X"86",X"45",X"45",X"45",X"45",X"43",X"89",X"0C",
		X"86",X"45",X"45",X"45",X"45",X"43",X"88",X"43",X"42",X"42",X"42",X"89",X"0C",X"86",X"F4",X"52",
		X"86",X"52",X"88",X"50",X"86",X"4A",X"88",X"0C",X"52",X"86",X"52",X"88",X"47",X"86",X"4A",X"88",
		X"0C",X"52",X"86",X"52",X"55",X"52",X"57",X"55",X"52",X"50",X"4A",X"4A",X"88",X"51",X"86",X"4A",
		X"88",X"0C",X"88",X"F4",X"53",X"86",X"53",X"84",X"53",X"87",X"51",X"86",X"53",X"53",X"84",X"53",
		X"87",X"51",X"86",X"53",X"88",X"48",X"8A",X"0C",X"88",X"F4",X"51",X"86",X"51",X"84",X"51",X"87",
		X"51",X"86",X"51",X"51",X"53",X"55",X"51",X"88",X"4A",X"8A",X"0C",X"88",X"F4",X"55",X"8A",X"57",
		X"88",X"57",X"55",X"8B",X"0C",X"88",X"F4",X"F0",X"00",X"F1",X"05",X"FA",X"01",X"FB",X"30",X"00",
		X"F3",X"AF",X"14",X"F3",X"CD",X"14",X"F3",X"CD",X"14",X"F3",X"ED",X"14",X"F3",X"00",X"15",X"F3",
		X"ED",X"14",X"F1",X"08",X"F3",X"13",X"15",X"F1",X"00",X"F3",X"CD",X"14",X"F2",X"87",X"14",X"F5",
		X"02",X"1A",X"86",X"2A",X"21",X"22",X"23",X"33",X"19",X"2A",X"F6",X"1A",X"2A",X"21",X"22",X"23",
		X"33",X"25",X"35",X"26",X"36",X"28",X"38",X"1A",X"1A",X"1A",X"1A",X"86",X"F4",X"F1",X"00",X"F5",
		X"02",X"0A",X"86",X"0A",X"11",X"12",X"13",X"13",X"19",X"1A",X"F6",X"0A",X"0A",X"11",X"12",X"13",
		X"13",X"15",X"15",X"16",X"16",X"18",X"18",X"1A",X"1A",X"1A",X"1A",X"86",X"F4",X"23",X"86",X"23",
		X"21",X"21",X"20",X"20",X"1A",X"1A",X"18",X"18",X"16",X"16",X"15",X"15",X"13",X"13",X"86",X"F4",
		X"11",X"86",X"11",X"10",X"10",X"0A",X"0A",X"08",X"08",X"0A",X"0A",X"10",X"10",X"11",X"11",X"12",
		X"12",X"86",X"F4",X"15",X"8A",X"10",X"15",X"15",X"8A",X"F4",X"F0",X"01",X"F1",X"05",X"FB",X"30",
		X"00",X"F3",X"40",X"15",X"F3",X"40",X"15",X"F3",X"40",X"15",X"F3",X"61",X"15",X"F3",X"72",X"15",
		X"F3",X"61",X"15",X"F1",X"08",X"F3",X"88",X"15",X"F1",X"05",X"F3",X"40",X"15",X"F2",X"1A",X"15",
		X"4A",X"86",X"4A",X"88",X"49",X"86",X"4A",X"89",X"0C",X"86",X"4A",X"4A",X"4A",X"49",X"86",X"45",
		X"89",X"0C",X"86",X"4A",X"4A",X"4A",X"49",X"45",X"88",X"45",X"45",X"45",X"45",X"89",X"0C",X"86",
		X"F4",X"4A",X"86",X"4A",X"4A",X"4A",X"88",X"0C",X"86",X"46",X"48",X"4A",X"4A",X"4A",X"8A",X"0C",
		X"88",X"F4",X"48",X"86",X"48",X"48",X"48",X"88",X"0C",X"86",X"48",X"48",X"51",X"88",X"50",X"86",
		X"48",X"88",X"0C",X"86",X"4A",X"45",X"86",X"F4",X"50",X"8A",X"53",X"88",X"53",X"50",X"8B",X"0C",
		X"88",X"F4",X"F0",X"01",X"F1",X"05",X"FA",X"00",X"FB",X"30",X"00",X"F3",X"BA",X"15",X"F3",X"BA",
		X"15",X"F3",X"BA",X"15",X"F3",X"DD",X"15",X"F3",X"EE",X"15",X"F3",X"DD",X"15",X"F1",X"08",X"F3",
		X"04",X"16",X"F1",X"05",X"F3",X"BA",X"15",X"F2",X"92",X"15",X"52",X"86",X"52",X"88",X"50",X"86",
		X"4A",X"47",X"4A",X"84",X"50",X"87",X"52",X"86",X"52",X"51",X"50",X"4A",X"89",X"0C",X"86",X"52",
		X"52",X"51",X"50",X"4A",X"88",X"4A",X"4A",X"4A",X"4A",X"89",X"0C",X"86",X"F4",X"46",X"86",X"46",
		X"46",X"46",X"88",X"0C",X"86",X"43",X"45",X"46",X"46",X"46",X"8A",X"0C",X"88",X"F4",X"45",X"86",
		X"45",X"45",X"45",X"88",X"0C",X"86",X"45",X"45",X"4A",X"88",X"48",X"86",X"45",X"88",X"0C",X"86",
		X"46",X"41",X"86",X"F4",X"49",X"8A",X"4A",X"88",X"4A",X"49",X"8B",X"0C",X"88",X"F4",X"00",X"00",
		X"22",X"16",X"01",X"42",X"16",X"02",X"62",X"16",X"03",X"82",X"16",X"04",X"9D",X"16",X"05",X"B9",
		X"16",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"1A",X"00",X"0C",X"89",X"47",X"8A",X"49",X"4B",X"50",
		X"86",X"F1",X"05",X"FB",X"34",X"00",X"49",X"86",X"4B",X"50",X"52",X"54",X"0C",X"84",X"50",X"0C",
		X"82",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"1A",X"00",X"0C",X"88",X"44",X"8A",X"45",X"47",X"49",
		X"88",X"F1",X"05",X"FB",X"34",X"00",X"39",X"86",X"3B",X"40",X"42",X"40",X"0C",X"84",X"40",X"0C",
		X"82",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"1A",X"00",X"0C",X"86",X"40",X"8A",X"42",X"44",X"45",
		X"89",X"F1",X"05",X"FB",X"34",X"00",X"35",X"86",X"37",X"39",X"3B",X"37",X"0C",X"84",X"37",X"0C",
		X"82",X"FF",X"F0",X"07",X"F1",X"00",X"FB",X"1A",X"00",X"0C",X"8C",X"0C",X"F1",X"01",X"FB",X"34",
		X"00",X"17",X"86",X"15",X"14",X"12",X"10",X"0C",X"84",X"10",X"0C",X"82",X"FF",X"F0",X"07",X"F1",
		X"00",X"FB",X"1A",X"00",X"0C",X"8C",X"0C",X"8C",X"F1",X"01",X"FB",X"34",X"00",X"27",X"86",X"25",
		X"24",X"22",X"20",X"0C",X"84",X"20",X"0C",X"82",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"1A",X"00",
		X"39",X"8A",X"3B",X"40",X"42",X"F1",X"05",X"FB",X"34",X"00",X"32",X"86",X"34",X"35",X"37",X"37",
		X"86",X"0C",X"84",X"34",X"0C",X"82",X"FF",X"00",X"00",X"EE",X"16",X"01",X"02",X"17",X"02",X"1B",
		X"17",X"03",X"32",X"17",X"04",X"46",X"17",X"05",X"5F",X"17",X"06",X"73",X"17",X"FF",X"F0",X"03",
		X"F1",X"07",X"FB",X"30",X"00",X"0C",X"88",X"54",X"54",X"52",X"52",X"49",X"4B",X"50",X"8A",X"0C",
		X"8F",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"30",X"00",X"0C",X"88",X"0C",X"86",X"50",X"88",X"50",
		X"4B",X"4B",X"86",X"45",X"88",X"47",X"47",X"8A",X"0C",X"8F",X"FF",X"F0",X"03",X"F1",X"07",X"FB",
		X"30",X"00",X"0C",X"88",X"F5",X"04",X"47",X"88",X"F6",X"42",X"88",X"44",X"88",X"44",X"8A",X"0C",
		X"8F",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"30",X"00",X"0C",X"88",X"44",X"44",X"42",X"42",X"40",
		X"3B",X"40",X"8A",X"0C",X"8F",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"30",X"00",X"0C",X"88",X"0C",
		X"86",X"40",X"88",X"40",X"3B",X"3B",X"86",X"39",X"88",X"37",X"37",X"8A",X"0C",X"8F",X"FF",X"F0",
		X"03",X"F1",X"07",X"FB",X"30",X"00",X"0C",X"88",X"20",X"20",X"1B",X"1B",X"19",X"1B",X"20",X"8A",
		X"0C",X"8F",X"FF",X"F0",X"03",X"F1",X"07",X"FB",X"30",X"00",X"0C",X"88",X"15",X"15",X"14",X"14",
		X"12",X"14",X"17",X"8A",X"0C",X"8F",X"FF",X"00",X"00",X"95",X"17",X"01",X"E3",X"17",X"02",X"04",
		X"18",X"03",X"25",X"18",X"FF",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"28",X"00",X"50",X"84",
		X"0C",X"50",X"54",X"57",X"0C",X"59",X"0C",X"60",X"0C",X"59",X"0C",X"57",X"0C",X"54",X"0C",X"49",
		X"0C",X"49",X"50",X"54",X"0C",X"57",X"0C",X"59",X"0C",X"57",X"0C",X"54",X"0C",X"50",X"0C",X"45",
		X"0C",X"45",X"49",X"50",X"0C",X"55",X"0C",X"57",X"0C",X"55",X"0C",X"50",X"0C",X"49",X"0C",X"47",
		X"0C",X"47",X"4B",X"52",X"0C",X"55",X"0C",X"57",X"0C",X"55",X"0C",X"52",X"0C",X"4B",X"0C",X"47",
		X"0C",X"8A",X"FF",X"F0",X"03",X"F1",X"09",X"FA",X"00",X"FB",X"28",X"00",X"47",X"8B",X"0C",X"86",
		X"47",X"49",X"8B",X"0C",X"86",X"44",X"40",X"8B",X"0C",X"86",X"3B",X"84",X"40",X"42",X"8B",X"0C",
		X"84",X"0C",X"8A",X"FF",X"F0",X"03",X"F1",X"09",X"FA",X"00",X"FB",X"28",X"00",X"40",X"8B",X"0C",
		X"86",X"40",X"39",X"8B",X"0C",X"86",X"39",X"35",X"8B",X"0C",X"86",X"34",X"84",X"35",X"37",X"8B",
		X"0C",X"84",X"0C",X"8A",X"FF",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"28",X"00",X"20",X"88",
		X"24",X"27",X"29",X"86",X"27",X"19",X"88",X"20",X"24",X"27",X"86",X"24",X"15",X"88",X"19",X"20",
		X"15",X"86",X"20",X"17",X"88",X"1B",X"22",X"25",X"86",X"22",X"17",X"84",X"0C",X"8A",X"FF",X"00",
		X"00",X"5D",X"18",X"01",X"BB",X"18",X"02",X"12",X"19",X"03",X"70",X"19",X"FF",X"F0",X"03",X"F1",
		X"09",X"FB",X"30",X"00",X"47",X"89",X"40",X"84",X"44",X"47",X"89",X"40",X"84",X"44",X"47",X"0C",
		X"47",X"0C",X"47",X"46",X"47",X"49",X"47",X"88",X"44",X"F1",X"00",X"59",X"84",X"58",X"59",X"86",
		X"5B",X"87",X"59",X"84",X"57",X"56",X"57",X"86",X"59",X"87",X"57",X"84",X"55",X"54",X"55",X"86",
		X"57",X"87",X"55",X"84",X"54",X"86",X"55",X"57",X"0C",X"59",X"84",X"58",X"59",X"86",X"5B",X"87",
		X"59",X"84",X"57",X"56",X"57",X"86",X"59",X"87",X"57",X"84",X"55",X"54",X"52",X"0C",X"5B",X"60",
		X"62",X"0C",X"60",X"86",X"0C",X"84",X"60",X"86",X"0C",X"86",X"FF",X"F0",X"03",X"F1",X"09",X"FB",
		X"30",X"00",X"44",X"89",X"37",X"84",X"40",X"44",X"89",X"37",X"84",X"40",X"44",X"0C",X"44",X"0C",
		X"44",X"43",X"44",X"45",X"44",X"88",X"40",X"F1",X"00",X"40",X"86",X"39",X"40",X"84",X"3B",X"39",
		X"86",X"3B",X"37",X"3B",X"84",X"39",X"37",X"86",X"39",X"35",X"39",X"84",X"37",X"35",X"86",X"0C",
		X"84",X"34",X"86",X"35",X"37",X"39",X"84",X"40",X"86",X"39",X"40",X"84",X"3B",X"39",X"86",X"3B",
		X"37",X"3B",X"84",X"39",X"37",X"86",X"39",X"35",X"3B",X"37",X"37",X"0C",X"84",X"37",X"86",X"0C",
		X"86",X"FF",X"F0",X"03",X"F1",X"09",X"FB",X"30",X"00",X"40",X"89",X"34",X"84",X"37",X"40",X"89",
		X"34",X"84",X"37",X"40",X"0C",X"40",X"0C",X"40",X"3B",X"40",X"42",X"40",X"88",X"37",X"F1",X"00",
		X"55",X"84",X"54",X"55",X"86",X"57",X"87",X"55",X"84",X"54",X"53",X"54",X"86",X"55",X"87",X"54",
		X"84",X"52",X"51",X"52",X"86",X"54",X"87",X"52",X"84",X"50",X"86",X"52",X"54",X"0C",X"55",X"84",
		X"54",X"55",X"86",X"57",X"87",X"55",X"84",X"54",X"53",X"54",X"86",X"55",X"87",X"54",X"84",X"52",
		X"50",X"4B",X"0C",X"57",X"59",X"5B",X"0C",X"57",X"86",X"0C",X"84",X"57",X"86",X"0C",X"86",X"FF",
		X"F0",X"03",X"F1",X"09",X"FB",X"30",X"00",X"37",X"89",X"30",X"84",X"34",X"37",X"89",X"30",X"84",
		X"34",X"37",X"0C",X"37",X"0C",X"37",X"36",X"37",X"39",X"37",X"88",X"34",X"F1",X"00",X"25",X"25",
		X"24",X"24",X"22",X"22",X"20",X"86",X"22",X"24",X"25",X"25",X"88",X"25",X"24",X"24",X"22",X"22",
		X"20",X"86",X"0C",X"84",X"20",X"86",X"0C",X"86",X"FF",X"00",X"00",X"BD",X"19",X"01",X"0A",X"1A",
		X"02",X"54",X"1A",X"03",X"99",X"1A",X"04",X"B3",X"1A",X"05",X"CD",X"1A",X"FF",X"F0",X"03",X"F1",
		X"08",X"FA",X"00",X"FB",X"30",X"00",X"40",X"86",X"40",X"88",X"47",X"45",X"86",X"44",X"42",X"40",
		X"47",X"88",X"45",X"44",X"42",X"86",X"42",X"42",X"88",X"49",X"47",X"86",X"45",X"44",X"42",X"49",
		X"47",X"88",X"45",X"44",X"44",X"86",X"47",X"88",X"4B",X"44",X"86",X"47",X"4B",X"45",X"49",X"88",
		X"50",X"45",X"86",X"49",X"50",X"52",X"52",X"0C",X"55",X"88",X"54",X"86",X"52",X"50",X"52",X"52",
		X"0C",X"89",X"52",X"86",X"50",X"4B",X"86",X"F2",X"BD",X"19",X"F0",X"03",X"F1",X"08",X"FA",X"00",
		X"FB",X"30",X"00",X"37",X"86",X"37",X"88",X"44",X"42",X"86",X"40",X"3B",X"37",X"44",X"88",X"42",
		X"40",X"3B",X"86",X"39",X"39",X"88",X"45",X"44",X"86",X"42",X"40",X"39",X"45",X"44",X"88",X"42",
		X"40",X"3B",X"86",X"44",X"88",X"47",X"3B",X"86",X"44",X"47",X"40",X"45",X"88",X"49",X"40",X"86",
		X"45",X"49",X"49",X"49",X"89",X"0C",X"8A",X"49",X"86",X"49",X"0C",X"89",X"4B",X"86",X"50",X"52",
		X"86",X"F2",X"0A",X"1A",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"30",X"00",X"F5",X"0D",X"20",
		X"86",X"F6",X"19",X"86",X"1B",X"20",X"86",X"F5",X"0D",X"22",X"86",X"F6",X"1B",X"86",X"20",X"22",
		X"86",X"F5",X"05",X"24",X"86",X"F6",X"20",X"86",X"22",X"24",X"86",X"F5",X"05",X"25",X"86",X"F6",
		X"22",X"86",X"24",X"25",X"22",X"22",X"0C",X"17",X"88",X"19",X"86",X"1B",X"20",X"22",X"22",X"0C",
		X"89",X"17",X"86",X"19",X"1B",X"86",X"F2",X"54",X"1A",X"F0",X"02",X"F1",X"0A",X"FB",X"30",X"00",
		X"30",X"8E",X"32",X"34",X"8C",X"35",X"37",X"86",X"37",X"0C",X"8B",X"37",X"86",X"37",X"0C",X"8B",
		X"F2",X"99",X"1A",X"F0",X"02",X"F1",X"0A",X"FB",X"30",X"00",X"34",X"8E",X"35",X"37",X"8C",X"39",
		X"3B",X"86",X"3B",X"0C",X"8B",X"3B",X"86",X"3B",X"0C",X"8B",X"F2",X"B3",X"1A",X"F0",X"02",X"F1",
		X"0A",X"FB",X"30",X"00",X"37",X"8E",X"39",X"3B",X"8C",X"40",X"42",X"86",X"42",X"0C",X"8B",X"42",
		X"86",X"42",X"0C",X"8B",X"F2",X"CD",X"1A",X"00",X"00",X"FE",X"1A",X"01",X"65",X"1B",X"02",X"24",
		X"1C",X"03",X"89",X"1C",X"04",X"DB",X"1C",X"05",X"F4",X"1C",X"06",X"0D",X"1D",X"FF",X"F0",X"03",
		X"F1",X"01",X"FA",X"00",X"FB",X"30",X"00",X"F5",X"04",X"50",X"88",X"F6",X"F5",X"04",X"4B",X"88",
		X"F6",X"F5",X"04",X"49",X"88",X"F6",X"0C",X"86",X"47",X"88",X"49",X"4B",X"50",X"86",X"F5",X"04",
		X"50",X"88",X"F6",X"F5",X"04",X"4B",X"88",X"F6",X"49",X"88",X"45",X"4B",X"47",X"50",X"49",X"52",
		X"52",X"55",X"55",X"88",X"F5",X"04",X"54",X"88",X"F6",X"F5",X"04",X"52",X"88",X"F6",X"F5",X"04",
		X"50",X"88",X"F6",X"4B",X"88",X"4B",X"4B",X"86",X"4B",X"50",X"52",X"86",X"F5",X"04",X"54",X"88",
		X"F6",X"F5",X"04",X"52",X"88",X"F6",X"50",X"88",X"49",X"52",X"4B",X"54",X"50",X"55",X"55",X"57",
		X"57",X"88",X"F2",X"FE",X"1A",X"F0",X"03",X"F1",X"00",X"FA",X"00",X"FB",X"30",X"00",X"F3",X"89",
		X"1B",X"F3",X"A2",X"1B",X"F3",X"89",X"1B",X"F3",X"B7",X"1B",X"F3",X"D7",X"1B",X"F3",X"F0",X"1B",
		X"F3",X"D7",X"1B",X"F3",X"06",X"1C",X"F2",X"65",X"1B",X"F5",X"03",X"0C",X"86",X"49",X"86",X"F6",
		X"50",X"84",X"4B",X"49",X"86",X"F5",X"03",X"0C",X"86",X"47",X"86",X"F6",X"4B",X"84",X"49",X"47",
		X"86",X"F4",X"F5",X"03",X"0C",X"86",X"45",X"86",X"F6",X"49",X"84",X"47",X"45",X"86",X"44",X"44",
		X"45",X"45",X"47",X"47",X"49",X"49",X"F4",X"0C",X"86",X"45",X"45",X"84",X"47",X"49",X"86",X"0C",
		X"47",X"47",X"84",X"49",X"4B",X"86",X"0C",X"49",X"49",X"84",X"4B",X"50",X"86",X"0C",X"4B",X"0C",
		X"4B",X"0C",X"52",X"0C",X"52",X"86",X"F4",X"F5",X"03",X"0C",X"86",X"50",X"86",X"F6",X"54",X"84",
		X"52",X"50",X"86",X"F5",X"03",X"0C",X"86",X"4B",X"86",X"F6",X"52",X"84",X"50",X"4B",X"86",X"F4",
		X"F5",X"03",X"0C",X"86",X"49",X"86",X"F6",X"50",X"84",X"4B",X"49",X"86",X"0C",X"47",X"0C",X"47",
		X"47",X"47",X"49",X"4B",X"86",X"F4",X"0C",X"86",X"49",X"49",X"84",X"4B",X"50",X"86",X"0C",X"4B",
		X"4B",X"84",X"50",X"52",X"86",X"0C",X"50",X"50",X"84",X"52",X"54",X"86",X"F5",X"04",X"0C",X"86",
		X"52",X"86",X"F6",X"F4",X"F0",X"03",X"F1",X"01",X"FA",X"00",X"FB",X"30",X"00",X"F5",X"04",X"45",
		X"88",X"F6",X"F5",X"04",X"44",X"88",X"F6",X"F5",X"04",X"42",X"88",X"F6",X"40",X"88",X"42",X"44",
		X"45",X"88",X"F5",X"04",X"45",X"88",X"F6",X"F5",X"04",X"44",X"88",X"F6",X"42",X"88",X"42",X"44",
		X"44",X"45",X"45",X"47",X"47",X"4B",X"4B",X"F5",X"04",X"49",X"88",X"F6",X"F5",X"04",X"47",X"88",
		X"F6",X"F5",X"04",X"45",X"88",X"F6",X"44",X"88",X"44",X"44",X"86",X"44",X"45",X"47",X"86",X"F5",
		X"04",X"49",X"88",X"F6",X"F5",X"04",X"47",X"88",X"F6",X"45",X"88",X"45",X"47",X"47",X"49",X"49",
		X"88",X"F5",X"04",X"4B",X"88",X"F6",X"F2",X"24",X"1C",X"F0",X"03",X"F1",X"01",X"FA",X"00",X"FB",
		X"30",X"00",X"F5",X"06",X"25",X"86",X"F6",X"27",X"86",X"25",X"86",X"F5",X"06",X"24",X"86",X"F6",
		X"25",X"86",X"24",X"86",X"F5",X"06",X"22",X"86",X"F6",X"24",X"86",X"22",X"20",X"20",X"22",X"22",
		X"24",X"24",X"25",X"25",X"F5",X"06",X"25",X"86",X"F6",X"27",X"86",X"25",X"86",X"F5",X"06",X"24",
		X"86",X"00",X"F6",X"25",X"86",X"24",X"22",X"22",X"20",X"22",X"24",X"24",X"22",X"24",X"25",X"25",
		X"24",X"25",X"86",X"F5",X"08",X"27",X"86",X"F6",X"F2",X"89",X"1C",X"F0",X"03",X"F1",X"09",X"FA",
		X"FF",X"FB",X"30",X"00",X"35",X"8C",X"34",X"32",X"30",X"35",X"34",X"32",X"8A",X"34",X"35",X"37",
		X"8C",X"F2",X"DB",X"1C",X"F0",X"03",X"F1",X"09",X"FA",X"00",X"FB",X"30",X"00",X"30",X"8C",X"2B",
		X"29",X"27",X"30",X"2B",X"29",X"8A",X"2B",X"30",X"32",X"8C",X"F2",X"F4",X"1C",X"F0",X"03",X"F1",
		X"00",X"FA",X"00",X"FB",X"30",X"00",X"F5",X"08",X"20",X"86",X"F6",X"F5",X"08",X"1B",X"86",X"F6",
		X"F5",X"08",X"19",X"86",X"F6",X"17",X"88",X"19",X"1B",X"86",X"17",X"19",X"86",X"1B",X"F5",X"08",
		X"20",X"86",X"F6",X"F5",X"08",X"1B",X"86",X"F6",X"F5",X"04",X"19",X"86",X"F6",X"F5",X"04",X"1B",
		X"86",X"F6",X"F5",X"04",X"20",X"86",X"F6",X"F5",X"08",X"22",X"86",X"F6",X"F2",X"0D",X"1D",X"00",
		X"00",X"66",X"1D",X"01",X"7C",X"1D",X"02",X"A2",X"1D",X"03",X"C7",X"1D",X"04",X"E3",X"1D",X"05",
		X"F1",X"1D",X"06",X"FF",X"1D",X"FF",X"F0",X"03",X"F1",X"08",X"FA",X"00",X"FB",X"28",X"00",X"F5",
		X"04",X"50",X"8B",X"F6",X"F5",X"04",X"52",X"8B",X"F6",X"F2",X"66",X"1D",X"F0",X"03",X"F1",X"08",
		X"FA",X"00",X"FB",X"28",X"00",X"0C",X"86",X"F5",X"03",X"54",X"8A",X"54",X"88",X"F6",X"54",X"8A",
		X"54",X"86",X"0C",X"86",X"F5",X"03",X"55",X"8A",X"55",X"88",X"F6",X"55",X"8A",X"55",X"86",X"F2",
		X"7C",X"1D",X"F0",X"03",X"F1",X"08",X"FA",X"00",X"FB",X"28",X"00",X"0C",X"88",X"F5",X"03",X"57",
		X"88",X"57",X"8A",X"F6",X"57",X"88",X"57",X"0C",X"88",X"F5",X"03",X"59",X"88",X"59",X"8A",X"F6",
		X"59",X"88",X"59",X"88",X"F2",X"A2",X"1D",X"F0",X"03",X"F1",X"08",X"FA",X"00",X"FB",X"28",X"00",
		X"0C",X"89",X"59",X"8B",X"59",X"59",X"59",X"89",X"0C",X"5B",X"8B",X"5B",X"5B",X"8B",X"5B",X"89",
		X"F2",X"C7",X"1D",X"F0",X"02",X"F1",X"03",X"FB",X"28",X"00",X"20",X"8F",X"22",X"8F",X"F2",X"E3",
		X"1D",X"F0",X"01",X"F1",X"03",X"FB",X"28",X"00",X"30",X"8F",X"32",X"8F",X"F2",X"F1",X"1D",X"F0",
		X"02",X"F1",X"08",X"FB",X"28",X"00",X"F5",X"04",X"40",X"86",X"44",X"47",X"49",X"47",X"44",X"F6",
		X"F5",X"04",X"42",X"86",X"45",X"49",X"4B",X"49",X"45",X"86",X"F6",X"F2",X"FF",X"1D",X"00",X"00",
		X"44",X"1E",X"01",X"64",X"1E",X"02",X"2C",X"1E",X"03",X"8C",X"1E",X"FF",X"F0",X"01",X"F1",X"07",
		X"FB",X"38",X"00",X"45",X"8A",X"F5",X"06",X"45",X"88",X"F6",X"47",X"8A",X"F5",X"06",X"47",X"88",
		X"F6",X"F2",X"2C",X"1E",X"F0",X"01",X"F1",X"07",X"FB",X"38",X"00",X"50",X"89",X"49",X"86",X"F5",
		X"06",X"50",X"86",X"49",X"86",X"F6",X"52",X"89",X"4B",X"86",X"F5",X"06",X"52",X"86",X"4B",X"86",
		X"F6",X"F2",X"44",X"1E",X"F0",X"01",X"F1",X"07",X"FB",X"38",X"00",X"0C",X"88",X"0C",X"84",X"F5",
		X"06",X"4B",X"86",X"47",X"86",X"F6",X"4B",X"86",X"47",X"84",X"0C",X"88",X"0C",X"84",X"F5",X"06",
		X"50",X"86",X"49",X"86",X"F6",X"50",X"86",X"49",X"84",X"F2",X"64",X"1E",X"F0",X"01",X"F1",X"01",
		X"FB",X"38",X"00",X"F5",X"02",X"15",X"86",X"15",X"19",X"19",X"20",X"20",X"19",X"19",X"86",X"F6",
		X"F5",X"02",X"17",X"86",X"17",X"1B",X"1B",X"22",X"22",X"1B",X"1B",X"86",X"F6",X"F2",X"8C",X"1E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
