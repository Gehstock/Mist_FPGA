library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"04",X"37",X"C5",X"E5",X"86",X"03",X"14",X"6A",X"A5",X"B5",X"85",X"8A",X"80",X"B9",X"10",
		X"BB",X"40",X"BA",X"06",X"54",X"62",X"FB",X"47",X"E7",X"53",X"1F",X"6B",X"AB",X"EA",X"14",X"BA",
		X"06",X"54",X"62",X"FB",X"47",X"E7",X"53",X"1F",X"37",X"17",X"6B",X"AB",X"EA",X"21",X"F9",X"03",
		X"FB",X"F6",X"35",X"9A",X"7F",X"E9",X"12",X"05",X"85",X"A5",X"B8",X"20",X"B0",X"00",X"D5",X"27",
		X"AE",X"AF",X"C5",X"8A",X"80",X"A5",X"26",X"A3",X"46",X"C9",X"0A",X"37",X"92",X"79",X"B2",X"77",
		X"D2",X"7B",X"80",X"53",X"0F",X"03",X"FD",X"96",X"5B",X"24",X"64",X"03",X"FD",X"96",X"61",X"24",
		X"8F",X"27",X"AE",X"AF",X"B4",X"24",X"14",X"6A",X"04",X"43",X"93",X"83",X"26",X"A3",X"46",X"C9",
		X"0A",X"37",X"D2",X"7B",X"92",X"79",X"83",X"24",X"00",X"44",X"00",X"B8",X"07",X"A5",X"B5",X"D4",
		X"1A",X"D4",X"3A",X"8A",X"80",X"96",X"89",X"04",X"43",X"B9",X"04",X"B4",X"24",X"26",X"A3",X"E9",
		X"8B",X"FA",X"03",X"FC",X"A9",X"C6",X"81",X"9A",X"7F",X"B4",X"24",X"26",X"A1",X"E9",X"99",X"04",
		X"81",X"8A",X"80",X"BA",X"E0",X"FA",X"AB",X"54",X"48",X"FA",X"77",X"77",X"53",X"3F",X"37",X"17",
		X"6A",X"AB",X"54",X"48",X"FA",X"AB",X"54",X"48",X"46",X"C9",X"FA",X"47",X"E7",X"53",X"1F",X"37",
		X"17",X"6A",X"AA",X"03",X"C0",X"F6",X"A5",X"04",X"43",X"BA",X"06",X"FA",X"AB",X"54",X"55",X"54",
		X"55",X"FA",X"97",X"67",X"6A",X"AB",X"54",X"55",X"54",X"55",X"FA",X"AB",X"54",X"55",X"54",X"55",
		X"FA",X"77",X"77",X"53",X"3F",X"6A",X"AA",X"03",X"C0",X"E6",X"CB",X"04",X"43",X"AB",X"54",X"3C",
		X"54",X"3C",X"FA",X"77",X"77",X"53",X"3F",X"6A",X"AA",X"03",X"C0",X"E6",X"DD",X"04",X"59",X"FF",
		X"BB",X"02",X"B9",X"88",X"BA",X"88",X"27",X"A8",X"AC",X"AD",X"D5",X"AC",X"AD",X"C5",X"97",X"A5",
		X"B5",X"34",X"DA",X"F9",X"53",X"3F",X"AF",X"FA",X"AE",X"D5",X"53",X"1F",X"AF",X"C5",X"F9",X"D5",
		X"AE",X"23",X"FF",X"62",X"D4",X"B7",X"34",X"5B",X"E8",X"11",X"9A",X"7F",X"EB",X"11",X"BB",X"08",
		X"8A",X"80",X"FC",X"D5",X"AC",X"C5",X"FD",X"D5",X"AD",X"C5",X"34",X"DA",X"F9",X"53",X"7F",X"AF",
		X"D5",X"AF",X"C5",X"FA",X"AE",X"D5",X"AE",X"23",X"FF",X"62",X"D4",X"B7",X"34",X"5B",X"E8",X"3A",
		X"9A",X"7F",X"EB",X"3A",X"D5",X"27",X"AE",X"AF",X"C5",X"04",X"43",X"0A",X"B2",X"62",X"76",X"63",
		X"24",X"00",X"A5",X"83",X"F9",X"96",X"6C",X"FC",X"AA",X"96",X"6C",X"19",X"34",X"DA",X"37",X"AB",
		X"FA",X"37",X"5B",X"AB",X"54",X"19",X"54",X"22",X"FA",X"AB",X"54",X"19",X"54",X"22",X"34",X"DA",
		X"F9",X"AB",X"54",X"19",X"54",X"22",X"80",X"53",X"0F",X"03",X"FD",X"C6",X"6C",X"04",X"43",X"BB",
		X"90",X"D5",X"B9",X"01",X"BA",X"04",X"BB",X"30",X"C5",X"54",X"7C",X"F2",X"AC",X"96",X"A1",X"04",
		X"37",X"AA",X"54",X"7C",X"37",X"96",X"AB",X"FA",X"A9",X"24",X"C0",X"37",X"D4",X"65",X"B9",X"03",
		X"D4",X"83",X"34",X"C9",X"E9",X"B0",X"FA",X"03",X"FA",X"A9",X"34",X"C9",X"E9",X"BA",X"B9",X"03",
		X"27",X"AE",X"AF",X"34",X"C9",X"E9",X"C3",X"24",X"99",X"D5",X"E9",X"D2",X"B9",X"08",X"FA",X"37",
		X"17",X"AA",X"FB",X"6A",X"AB",X"54",X"70",X"F5",X"C4",X"40",X"F9",X"F7",X"A9",X"FA",X"F7",X"AA",
		X"F9",X"F6",X"EA",X"32",X"EC",X"F9",X"53",X"FE",X"A9",X"83",X"32",X"E5",X"F9",X"43",X"01",X"A9",
		X"83",X"32",X"EC",X"F9",X"43",X"01",X"A9",X"83",X"54",X"41",X"14",X"6B",X"54",X"41",X"14",X"6B",
		X"B9",X"20",X"BA",X"40",X"FA",X"AB",X"54",X"62",X"FA",X"97",X"67",X"AB",X"54",X"62",X"FA",X"47",
		X"E7",X"53",X"1F",X"6A",X"AA",X"E6",X"04",X"04",X"43",X"54",X"48",X"14",X"6C",X"54",X"48",X"14",
		X"6C",X"83",X"54",X"33",X"14",X"6C",X"54",X"33",X"14",X"6C",X"54",X"33",X"14",X"6C",X"54",X"33",
		X"14",X"6C",X"83",X"27",X"AE",X"AF",X"D5",X"AE",X"AF",X"A4",X"24",X"FB",X"47",X"E7",X"AE",X"53",
		X"1F",X"AF",X"FE",X"53",X"E0",X"AE",X"A4",X"24",X"FB",X"77",X"77",X"AE",X"53",X"3F",X"AF",X"FE",
		X"53",X"C0",X"AE",X"A4",X"24",X"FB",X"77",X"AE",X"53",X"7F",X"AF",X"FE",X"53",X"80",X"AE",X"D5",
		X"A4",X"24",X"FB",X"77",X"77",X"AE",X"53",X"3F",X"AF",X"FE",X"53",X"C0",X"AE",X"D5",X"A4",X"6E",
		X"FB",X"77",X"77",X"AE",X"53",X"3F",X"AF",X"FE",X"53",X"C0",X"AE",X"83",X"FB",X"1B",X"A3",X"A8",
		X"83",X"98",X"30",X"A0",X"0C",X"A2",X"A6",X"A4",X"A2",X"18",X"A8",X"A8",X"0C",X"A8",X"AA",X"A4",
		X"18",X"A0",X"30",X"A6",X"0C",X"A8",X"AB",X"AA",X"A8",X"18",X"B0",X"B0",X"0C",X"B0",X"B2",X"AA",
		X"AB",X"18",X"A8",X"A8",X"0C",X"A8",X"AB",X"AA",X"A8",X"A6",X"B6",X"B4",X"B2",X"B0",X"AB",X"AA",
		X"A8",X"30",X"A6",X"0C",X"A8",X"AB",X"AA",X"A8",X"18",X"B0",X"B0",X"0C",X"B0",X"B2",X"AA",X"AB",
		X"18",X"A8",X"A8",X"0C",X"A8",X"AB",X"AA",X"A8",X"A6",X"B0",X"A8",X"AA",X"18",X"A6",X"18",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"86",X"82",X"80",X"0C",X"82",X"18",X"86",X"86",X"0C",X"82",X"18",X"80",X"82",X"18",X"88",
		X"84",X"82",X"0C",X"84",X"18",X"88",X"88",X"0C",X"84",X"18",X"82",X"84",X"00",X"10",X"86",X"20",
		X"86",X"10",X"80",X"86",X"20",X"86",X"10",X"80",X"86",X"20",X"86",X"10",X"80",X"86",X"84",X"86",
		X"87",X"88",X"20",X"88",X"10",X"82",X"88",X"20",X"88",X"10",X"82",X"88",X"20",X"88",X"10",X"82",
		X"88",X"87",X"88",X"89",X"00",X"00",X"00",X"00",X"0C",X"90",X"90",X"90",X"90",X"92",X"94",X"96",
		X"96",X"96",X"96",X"94",X"92",X"00",X"04",X"A4",X"10",X"A6",X"04",X"AC",X"10",X"B0",X"04",X"B4",
		X"10",X"B6",X"00",X"09",X"EA",X"8A",X"E8",X"88",X"6C",X"EA",X"8A",X"09",X"E8",X"88",X"E6",X"86",
		X"E4",X"84",X"E2",X"82",X"24",X"E1",X"81",X"48",X"E2",X"82",X"24",X"FF",X"09",X"DA",X"8A",X"D8",
		X"88",X"6C",X"DA",X"8A",X"0C",X"D4",X"84",X"D6",X"86",X"D1",X"81",X"6C",X"D2",X"82",X"24",X"FF",
		X"12",X"82",X"C6",X"82",X"C9",X"86",X"CC",X"89",X"D2",X"8C",X"D6",X"92",X"D9",X"96",X"DC",X"99",
		X"09",X"E2",X"9C",X"E1",X"9C",X"E2",X"9C",X"E1",X"9C",X"09",X"E2",X"9C",X"E1",X"9C",X"E2",X"9C",
		X"E1",X"9C",X"24",X"E2",X"9C",X"00",X"0F",X"E8",X"90",X"B0",X"94",X"A8",X"1E",X"F0",X"98",X"E8",
		X"94",X"0F",X"E7",X"90",X"B0",X"93",X"A7",X"1E",X"F0",X"97",X"E7",X"93",X"0F",X"E6",X"92",X"B0",
		X"96",X"A6",X"1E",X"F0",X"9A",X"F4",X"A0",X"B8",X"06",X"97",X"18",X"98",X"3C",X"88",X"00",X"1E",
		X"E0",X"98",X"0F",X"E2",X"9A",X"E4",X"9C",X"1E",X"E6",X"A0",X"E4",X"A0",X"1E",X"E2",X"A0",X"0F",
		X"E0",X"9A",X"1E",X"DC",X"98",X"0F",X"DA",X"96",X"1E",X"D8",X"94",X"1E",X"E0",X"98",X"0F",X"E2",
		X"9A",X"E4",X"9C",X"1E",X"E6",X"A0",X"E4",X"A0",X"1E",X"E2",X"A0",X"0F",X"E0",X"9A",X"38",X"DC",
		X"98",X"00",X"12",X"E4",X"94",X"A9",X"EC",X"8C",X"B2",X"E7",X"87",X"AA",X"F0",X"83",X"B3",X"09",
		X"F6",X"92",X"B2",X"B4",X"B0",X"F2",X"8C",X"AC",X"B0",X"AA",X"EC",X"88",X"A8",X"AA",X"A6",X"E8",
		X"84",X"A4",X"A6",X"A2",X"12",X"E0",X"80",X"82",X"84",X"24",X"88",X"12",X"8A",X"90",X"92",X"48",
		X"90",X"00",X"1E",X"E0",X"90",X"E8",X"88",X"0F",X"E4",X"80",X"A0",X"1E",X"88",X"DC",X"94",X"E8",
		X"8C",X"0F",X"E4",X"94",X"9C",X"1E",X"8C",X"DA",X"86",X"E0",X"80",X"0F",X"E6",X"86",X"A8",X"80",
		X"A6",X"1E",X"E4",X"90",X"88",X"E2",X"98",X"92",X"E0",X"90",X"E8",X"88",X"0F",X"E4",X"80",X"A0",
		X"1E",X"88",X"DC",X"94",X"E8",X"8C",X"0F",X"E4",X"94",X"9C",X"1E",X"8C",X"DA",X"86",X"E0",X"80",
		X"0F",X"E4",X"94",X"A8",X"8C",X"A4",X"1E",X"E2",X"88",X"82",X"3C",X"E0",X"90",X"00",X"20",X"80",
		X"10",X"E4",X"A0",X"E4",X"A0",X"E6",X"A2",X"E6",X"A2",X"E8",X"A4",X"E8",X"A4",X"10",X"EA",X"86",
		X"80",X"EA",X"86",X"80",X"E8",X"86",X"E6",X"80",X"E6",X"82",X"84",X"90",X"E8",X"88",X"E8",X"90",
		X"E8",X"88",X"E6",X"90",X"E8",X"98",X"96",X"94",X"E6",X"92",X"8A",X"E6",X"92",X"E6",X"8A",X"E6",
		X"92",X"E4",X"8A",X"92",X"E2",X"8A",X"E0",X"86",X"8A",X"8B",X"90",X"E6",X"86",X"8B",X"EA",X"90",
		X"92",X"E8",X"98",X"96",X"94",X"92",X"90",X"8B",X"8A",X"E4",X"88",X"E6",X"86",X"20",X"86",X"10",
		X"86",X"90",X"8B",X"8A",X"88",X"40",X"86",X"00",X"86",X"90",X"8B",X"8A",X"88",X"40",X"86",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A3",X"83",
		X"00",X"01",X"80",X"00",X"02",X"06",X"00",X"40",X"20",X"12",X"14",X"16",X"18",X"1A",X"1C",X"00",
		X"08",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",X"FF",X"00",X"0E",X"00",
		X"08",X"00",X"A3",X"83",X"D5",X"B6",X"90",X"B8",X"20",X"80",X"53",X"0F",X"20",X"37",X"17",X"60",
		X"96",X"4D",X"F0",X"A3",X"C6",X"4B",X"F2",X"73",X"D4",X"83",X"E9",X"4B",X"FF",X"96",X"42",X"FE",
		X"C6",X"5E",X"FA",X"03",X"F8",X"C6",X"5E",X"A9",X"27",X"AE",X"AF",X"C4",X"90",X"F0",X"A3",X"C6",
		X"6E",X"92",X"66",X"B2",X"6A",X"D2",X"89",X"F2",X"75",X"8A",X"80",X"A8",X"D4",X"1A",X"D4",X"3A",
		X"C6",X"4D",X"B9",X"08",X"C4",X"90",X"F4",X"04",X"04",X"37",X"F4",X"3B",X"04",X"37",X"27",X"AE",
		X"AF",X"C4",X"90",X"E9",X"79",X"B9",X"10",X"BB",X"73",X"FB",X"47",X"E7",X"53",X"1F",X"6B",X"AB",
		X"77",X"77",X"AE",X"53",X"3F",X"AF",X"F5",X"C4",X"40",X"B9",X"48",X"95",X"BA",X"06",X"BB",X"C0",
		X"E9",X"9B",X"B8",X"20",X"27",X"A0",X"AE",X"AF",X"85",X"A4",X"24",X"EA",X"AC",X"BA",X"06",X"FB",
		X"47",X"E7",X"53",X"1F",X"A8",X"97",X"67",X"68",X"37",X"17",X"6B",X"AB",X"FB",X"77",X"77",X"53",
		X"3F",X"AF",X"80",X"53",X"0F",X"03",X"F6",X"C6",X"98",X"F5",X"C4",X"40",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"28",X"00",X"2A",X"61",X"2C",X"E6",X"2F",X"91",X"32",X"66",X"FF",X"FF",X"35",X"65",X"38",X"92",
		X"3B",X"EF",X"3F",X"75",X"43",X"46",X"47",X"46",X"4B",X"83",X"BB",X"00",X"B9",X"30",X"B1",X"FF",
		X"C4",X"26",X"D4",X"29",X"96",X"22",X"E8",X"22",X"83",X"B9",X"30",X"FB",X"96",X"2F",X"11",X"F1",
		X"96",X"36",X"FB",X"1B",X"E3",X"83",X"FB",X"1B",X"84",X"FE",X"D4",X"29",X"C6",X"64",X"F2",X"43",
		X"AA",X"D4",X"29",X"A8",X"37",X"96",X"4F",X"AE",X"AF",X"D5",X"AE",X"AF",X"C5",X"17",X"83",X"D4",
		X"65",X"F8",X"83",X"D2",X"5C",X"D5",X"BE",X"00",X"BF",X"00",X"C5",X"83",X"D4",X"29",X"D5",X"A8",
		X"D4",X"65",X"C5",X"F8",X"83",X"F8",X"53",X"0F",X"E7",X"AC",X"A3",X"AF",X"FC",X"17",X"A3",X"AE",
		X"F8",X"53",X"30",X"47",X"AC",X"FF",X"97",X"67",X"AF",X"FE",X"67",X"AE",X"1C",X"FC",X"03",X"FC",
		X"96",X"75",X"83",X"FE",X"6F",X"E6",X"88",X"1F",X"6F",X"E6",X"8C",X"1F",X"AE",X"83",X"FF",X"FF",
		X"42",X"03",X"78",X"62",X"76",X"B7",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",
		X"A3",X"A8",X"C5",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",X"A3",X"D5",X"68",
		X"39",X"16",X"B5",X"C4",X"96",X"C5",X"83",X"F5",X"E4",X"40",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"06",X"09",X"0C",X"0F",X"12",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",
		X"30",X"33",X"36",X"39",X"3C",X"3F",X"42",X"45",X"48",X"4B",X"4E",X"51",X"54",X"57",X"5A",X"5D",
		X"60",X"5D",X"5A",X"57",X"54",X"51",X"4E",X"4B",X"48",X"45",X"42",X"3F",X"3C",X"39",X"36",X"33",
		X"30",X"2D",X"2A",X"27",X"24",X"21",X"1E",X"1B",X"18",X"15",X"12",X"0F",X"0C",X"09",X"06",X"03",
		X"E2",X"FC",X"04",X"1E",X"AB",X"D5",X"FB",X"1B",X"C5",X"B4",X"22",X"C6",X"5E",X"A8",X"92",X"5A",
		X"D4",X"1A",X"D4",X"3A",X"D4",X"53",X"C6",X"05",X"B9",X"03",X"8A",X"80",X"D4",X"83",X"D5",X"D4",
		X"83",X"D4",X"90",X"E9",X"1C",X"B9",X"03",X"D5",X"D4",X"90",X"E9",X"27",X"FA",X"03",X"FA",X"A9",
		X"C6",X"12",X"9A",X"7F",X"D5",X"D4",X"90",X"E9",X"34",X"E4",X"12",X"AB",X"D5",X"FB",X"1B",X"C5",
		X"B4",X"22",X"C6",X"5E",X"A8",X"D4",X"1A",X"D4",X"3A",X"D4",X"53",X"C6",X"3C",X"FA",X"A9",X"D4",
		X"83",X"D4",X"83",X"D5",X"D4",X"90",X"E9",X"53",X"E4",X"47",X"F4",X"5F",X"E4",X"05",X"83",X"BF",
		X"80",X"B9",X"F0",X"B8",X"02",X"F4",X"76",X"E5",X"00",X"F4",X"82",X"18",X"F8",X"96",X"65",X"19",
		X"F9",X"03",X"0D",X"96",X"63",X"83",X"F9",X"B3",X"BE",X"08",X"EE",X"7A",X"FB",X"77",X"77",X"AB",
		X"E4",X"85",X"BA",X"04",X"AB",X"53",X"03",X"A3",X"F2",X"94",X"6F",X"E6",X"8F",X"23",X"FF",X"AF",
		X"39",X"EA",X"78",X"83",X"6F",X"F6",X"8F",X"27",X"E4",X"8F",X"9E",X"BA",X"04",X"AB",X"53",X"03",
		X"A3",X"F2",X"AD",X"6F",X"E6",X"A8",X"23",X"FF",X"AF",X"39",X"EA",X"91",X"83",X"6F",X"F6",X"A8",
		X"27",X"E4",X"A8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F5",X"04",X"00",X"F8",X"F5",X"24",X"00",X"F8",X"F5",X"44",X"00",X"F8",X"F5",X"64",X"00",
		X"F8",X"F5",X"84",X"00",X"F8",X"F5",X"A4",X"00",X"F8",X"F5",X"C4",X"00",X"F8",X"F5",X"E4",X"00",
		X"D0",X"D4",X"D8",X"DC",X"E0",X"E4",X"E8",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A3",X"83",X"70",X"7C",X"0F",X"E0",X"E3",X"80",X"5F",X"0F",X"FC",X"F0",X"C0",X"8F",X"02",X"7F",
		X"04",X"FF",X"03",X"FC",X"3C",X"C0",X"4B",X"0F",X"BD",X"08",X"F8",X"C3",X"0B",X"3F",X"90",X"FE",
		X"41",X"4B",X"0F",X"F8",X"11",X"F8",X"0B",X"0E",X"EF",X"81",X"3F",X"B0",X"F0",X"0B",X"F0",X"1B",
		X"48",X"7F",X"90",X"FE",X"40",X"8F",X"0F",X"FC",X"E0",X"C0",X"4F",X"C1",X"2F",X"7C",X"F0",X"0F",
		X"F0",X"83",X"07",X"3F",X"09",X"FF",X"D0",X"D0",X"1F",X"C0",X"8B",X"09",X"3F",X"0F",X"FC",X"C1",
		X"F0",X"57",X"C0",X"2F",X"24",X"FF",X"40",X"F7",X"02",X"3F",X"3C",X"F0",X"07",X"A9",X"6E",X"D0",
		X"67",X"C0",X"1F",X"29",X"9F",X"03",X"7E",X"1C",X"BC",X"0B",X"F8",X"3C",X"F0",X"83",X"C0",X"7F",
		X"D0",X"2F",X"80",X"BF",X"01",X"FE",X"00",X"FF",X"02",X"FC",X"07",X"FC",X"0B",X"B8",X"1E",X"F0",
		X"1F",X"D0",X"3B",X"D0",X"1F",X"C0",X"BF",X"80",X"FF",X"00",X"FE",X"00",X"FF",X"01",X"BE",X"03",
		X"FC",X"07",X"F8",X"06",X"F4",X"0B",X"F0",X"1F",X"F0",X"2F",X"C0",X"3F",X"00",X"FF",X"C0",X"CF",
		X"00",X"FF",X"00",X"FF",X"03",X"FC",X"00",X"FD",X"06",X"F4",X"0F",X"F0",X"2B",X"B0",X"0F",X"BC",
		X"3D",X"F0",X"2D",X"C0",X"3F",X"C0",X"7F",X"E0",X"F1",X"80",X"7F",X"40",X"FF",X"00",X"FF",X"02",
		X"FC",X"00",X"FE",X"03",X"D3",X"07",X"FC",X"03",X"F4",X"07",X"8E",X"1F",X"E8",X"07",X"DE",X"07",
		X"3C",X"0F",X"E4",X"0F",X"F8",X"0F",X"A0",X"3F",X"20",X"2F",X"B8",X"35",X"F8",X"34",X"F4",X"0E",
		X"F8",X"52",X"F0",X"47",X"F0",X"2F",X"F0",X"53",X"C0",X"3F",X"D0",X"BF",X"C0",X"7B",X"C0",X"0F",
		X"41",X"BF",X"C0",X"AF",X"C0",X"3E",X"80",X"BF",X"80",X"FF",X"40",X"FF",X"00",X"BF",X"40",X"BF",
		X"A3",X"83",X"00",X"7F",X"01",X"FF",X"03",X"AF",X"01",X"EF",X"03",X"FC",X"02",X"FC",X"03",X"FC",
		X"0F",X"74",X"0E",X"E8",X"03",X"5F",X"0F",X"7C",X"06",X"7D",X"0A",X"6E",X"0F",X"7C",X"1C",X"BC",
		X"08",X"FD",X"09",X"FC",X"64",X"F8",X"50",X"5F",X"74",X"F8",X"80",X"FF",X"00",X"FF",X"00",X"BF",
		X"01",X"FE",X"01",X"AF",X"03",X"FC",X"01",X"FF",X"00",X"FF",X"01",X"CF",X"0F",X"FC",X"01",X"FC",
		X"03",X"FC",X"81",X"EB",X"81",X"D7",X"03",X"FD",X"00",X"FC",X"82",X"FF",X"03",X"FC",X"00",X"AE",
		X"0B",X"5F",X"E1",X"D2",X"91",X"1F",X"84",X"FF",X"00",X"FF",X"40",X"2F",X"05",X"FE",X"01",X"FE",
		X"01",X"FF",X"40",X"7F",X"00",X"FF",X"40",X"FF",X"40",X"3F",X"C0",X"F7",X"40",X"5F",X"E1",X"D2",
		X"46",X"1F",X"F8",X"81",X"0F",X"9E",X"07",X"BF",X"50",X"7D",X"D0",X"3E",X"30",X"FC",X"01",X"BE",
		X"78",X"F0",X"C1",X"C7",X"83",X"F4",X"03",X"FE",X"41",X"F1",X"43",X"5E",X"3F",X"F0",X"92",X"C0",
		X"1F",X"F0",X"1F",X"F0",X"1F",X"F0",X"0F",X"F0",X"0F",X"F0",X"0B",X"F0",X"0F",X"F4",X"0F",X"F0",
		X"03",X"F4",X"0F",X"F0",X"0F",X"F8",X"0B",X"28",X"FD",X"80",X"3F",X"F0",X"2F",X"C0",X"3F",X"40",
		X"FF",X"00",X"3F",X"00",X"FE",X"42",X"FF",X"00",X"FD",X"01",X"BF",X"E0",X"C3",X"0B",X"F9",X"D1",
		X"74",X"E5",X"06",X"8F",X"03",X"3F",X"3D",X"F0",X"0F",X"D0",X"0F",X"F0",X"1F",X"E0",X"3F",X"D0",
		X"0F",X"C0",X"1F",X"F4",X"7D",X"C0",X"0F",X"0D",X"2F",X"F0",X"07",X"E6",X"1F",X"E0",X"1F",X"C0",
		X"6F",X"80",X"3F",X"F0",X"2F",X"C0",X"7F",X"80",X"AF",X"C0",X"BF",X"00",X"FF",X"00",X"3F",X"40",
		X"FF",X"C0",X"FA",X"80",X"77",X"B4",X"F0",X"E1",X"C1",X"E3",X"82",X"CF",X"06",X"BC",X"0F",X"F4",
		X"A3",X"83",X"03",X"BC",X"0F",X"F0",X"3A",X"E0",X"0F",X"F0",X"0F",X"F0",X"1F",X"C0",X"BF",X"80",
		X"3F",X"40",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FD",X"03",X"FB",X"02",X"FC",X"03",
		X"E9",X"0B",X"FC",X"03",X"B9",X"43",X"A7",X"A4",X"0B",X"BC",X"0F",X"F0",X"0F",X"F0",X"0B",X"F0",
		X"0F",X"F0",X"0F",X"F0",X"0B",X"F8",X"4B",X"D0",X"0F",X"6A",X"CB",X"42",X"0F",X"7F",X"70",X"6E",
		X"70",X"2F",X"B0",X"EE",X"80",X"7F",X"00",X"BF",X"00",X"FF",X"00",X"FF",X"01",X"BF",X"90",X"5D",
		X"E1",X"0A",X"E5",X"0B",X"FD",X"03",X"FC",X"0B",X"F0",X"0B",X"E0",X"2F",X"C0",X"7F",X"40",X"7F",
		X"04",X"FC",X"03",X"FD",X"07",X"F4",X"07",X"CB",X"0F",X"1D",X"3D",X"3C",X"E4",X"B7",X"40",X"7F",
		X"00",X"7F",X"40",X"7F",X"3D",X"F0",X"C3",X"81",X"FF",X"00",X"FD",X"03",X"F8",X"0B",X"F0",X"0F",
		X"D0",X"2F",X"08",X"FF",X"06",X"F8",X"3E",X"C0",X"1F",X"C0",X"3F",X"38",X"F8",X"F0",X"D0",X"D7",
		X"03",X"FC",X"42",X"F8",X"43",X"0B",X"FD",X"30",X"E8",X"0F",X"B0",X"6F",X"40",X"FF",X"10",X"FC",
		X"BA",X"C0",X"2F",X"00",X"FF",X"02",X"FC",X"52",X"A9",X"92",X"2F",X"E0",X"5F",X"E0",X"9E",X"01",
		X"FD",X"C2",X"61",X"FD",X"01",X"FC",X"16",X"F0",X"1F",X"D0",X"1F",X"B5",X"15",X"F5",X"03",X"FC",
		X"07",X"E8",X"6B",X"90",X"6B",X"85",X"4F",X"B2",X"A5",X"96",X"55",X"3E",X"90",X"BE",X"0A",X"F8",
		X"17",X"D0",X"8F",X"03",X"FD",X"62",X"94",X"6F",X"41",X"7E",X"09",X"7E",X"55",X"A5",X"6A",X"F4",
		X"C1",X"57",X"81",X"AF",X"91",X"E9",X"03",X"FD",X"01",X"FF",X"00",X"FE",X"81",X"3A",X"89",X"1F",
		X"B4",X"3D",X"A0",X"7E",X"D0",X"07",X"F9",X"15",X"F8",X"B6",X"90",X"1B",X"AA",X"D1",X"D3",X"42",
		X"A3",X"83",X"7E",X"15",X"8E",X"0B",X"FD",X"02",X"E9",X"2F",X"90",X"2F",X"A4",X"7D",X"E0",X"6A",
		X"D0",X"7E",X"81",X"4B",X"57",X"E5",X"51",X"9B",X"0A",X"7E",X"28",X"F9",X"41",X"2F",X"94",X"7F",
		X"80",X"6F",X"A0",X"5F",X"A1",X"59",X"6E",X"54",X"FE",X"01",X"E7",X"03",X"F9",X"0A",X"F8",X"46",
		X"B9",X"95",X"16",X"7D",X"A4",X"B5",X"82",X"BA",X"38",X"B8",X"29",X"B9",X"55",X"69",X"95",X"47",
		X"1E",X"2E",X"A5",X"2B",X"B8",X"2A",X"B4",X"17",X"6D",X"1A",X"B9",X"55",X"96",X"A6",X"95",X"69",
		X"59",X"E6",X"82",X"9B",X"16",X"2E",X"6D",X"F4",X"81",X"9B",X"25",X"BD",X"51",X"A9",X"57",X"E4",
		X"A9",X"A0",X"5F",X"91",X"7A",X"C1",X"6B",X"51",X"7E",X"A0",X"FA",X"80",X"AF",X"10",X"FD",X"03",
		X"F9",X"07",X"B8",X"2A",X"A4",X"5F",X"51",X"6E",X"55",X"6D",X"59",X"1A",X"AA",X"5A",X"A5",X"1E",
		X"B8",X"65",X"B5",X"52",X"B9",X"46",X"A5",X"0F",X"E5",X"59",X"65",X"5E",X"E1",X"46",X"9E",X"92",
		X"6A",X"5A",X"4A",X"7E",X"64",X"A5",X"4E",X"56",X"2E",X"96",X"66",X"A5",X"76",X"54",X"AE",X"45",
		X"EA",X"25",X"F8",X"D1",X"E1",X"07",X"B9",X"55",X"9A",X"A5",X"E5",X"91",X"4B",X"A9",X"57",X"D4",
		X"0B",X"6D",X"69",X"A5",X"53",X"B9",X"05",X"BE",X"05",X"FD",X"54",X"EA",X"42",X"BA",X"55",X"69",
		X"1A",X"AA",X"56",X"5A",X"AA",X"A1",X"5B",X"E1",X"A5",X"55",X"5E",X"69",X"55",X"AA",X"56",X"A5",
		X"5A",X"95",X"1B",X"A9",X"6A",X"A4",X"5B",X"F4",X"91",X"96",X"47",X"96",X"5B",X"55",X"1E",X"B5",
		X"95",X"96",X"56",X"6A",X"2A",X"A9",X"2A",X"A9",X"AA",X"D0",X"6B",X"E0",X"6A",X"45",X"2F",X"A5",
		X"69",X"E5",X"52",X"A9",X"0B",X"AA",X"5A",X"95",X"1E",X"A9",X"79",X"D4",X"B2",X"D4",X"96",X"91",
		X"A3",X"83",X"70",X"7C",X"0F",X"E0",X"E3",X"80",X"5F",X"0F",X"FC",X"F0",X"C0",X"8F",X"02",X"7F",
		X"04",X"FF",X"03",X"FC",X"3C",X"C0",X"4B",X"0F",X"BD",X"08",X"F8",X"C3",X"0B",X"3F",X"90",X"FE",
		X"41",X"4B",X"0F",X"F8",X"11",X"F8",X"0B",X"0E",X"EF",X"81",X"3F",X"B0",X"F0",X"0B",X"F0",X"1B",
		X"48",X"7F",X"90",X"FE",X"40",X"8F",X"0F",X"FC",X"E0",X"C0",X"4F",X"C1",X"2F",X"7C",X"F0",X"0F",
		X"F0",X"83",X"07",X"3F",X"09",X"FF",X"D0",X"D0",X"1F",X"C0",X"8B",X"09",X"3F",X"0F",X"FC",X"C1",
		X"F0",X"57",X"C0",X"2F",X"24",X"FF",X"40",X"F7",X"02",X"3F",X"3C",X"F0",X"07",X"A9",X"6E",X"D0",
		X"67",X"C0",X"1F",X"29",X"9F",X"03",X"7E",X"1C",X"BC",X"0B",X"F8",X"3C",X"F0",X"83",X"C0",X"7F",
		X"D0",X"2F",X"80",X"BF",X"01",X"FE",X"00",X"FF",X"02",X"FC",X"07",X"FC",X"0B",X"B8",X"1E",X"F0",
		X"1F",X"D0",X"3B",X"D0",X"1F",X"C0",X"BF",X"80",X"FF",X"00",X"FE",X"00",X"FF",X"01",X"BE",X"03",
		X"FC",X"07",X"F8",X"06",X"F4",X"0B",X"F0",X"1F",X"F0",X"2F",X"C0",X"3F",X"00",X"FF",X"C0",X"CF",
		X"00",X"FF",X"00",X"FF",X"03",X"FC",X"00",X"FD",X"06",X"F4",X"0F",X"F0",X"2B",X"B0",X"0F",X"BC",
		X"3D",X"F0",X"2D",X"C0",X"3F",X"C0",X"7F",X"E0",X"F1",X"80",X"7F",X"40",X"FF",X"00",X"FF",X"02",
		X"FC",X"00",X"FE",X"03",X"D3",X"07",X"FC",X"03",X"F4",X"07",X"8E",X"1F",X"E8",X"07",X"DE",X"07",
		X"3C",X"0F",X"E4",X"0F",X"F8",X"0F",X"A0",X"3F",X"20",X"2F",X"B8",X"35",X"F8",X"34",X"F4",X"0E",
		X"F8",X"52",X"F0",X"47",X"F0",X"2F",X"F0",X"53",X"C0",X"3F",X"D0",X"BF",X"C0",X"7B",X"C0",X"0F",
		X"41",X"BF",X"C0",X"AF",X"C0",X"3E",X"80",X"BF",X"80",X"FF",X"40",X"FF",X"00",X"BF",X"40",X"BF",
		X"A3",X"83",X"00",X"7F",X"01",X"FF",X"03",X"AF",X"01",X"EF",X"03",X"FC",X"02",X"FC",X"03",X"FC",
		X"0F",X"74",X"0E",X"E8",X"03",X"5F",X"0F",X"7C",X"06",X"7D",X"0A",X"6E",X"0F",X"7C",X"1C",X"BC",
		X"08",X"FD",X"09",X"FC",X"64",X"F8",X"50",X"5F",X"74",X"F8",X"80",X"FF",X"00",X"FF",X"00",X"BF",
		X"01",X"FE",X"01",X"AF",X"03",X"FC",X"01",X"FF",X"00",X"FF",X"01",X"CF",X"0F",X"FC",X"01",X"FC",
		X"03",X"FC",X"81",X"EB",X"81",X"D7",X"03",X"FD",X"00",X"FC",X"82",X"FF",X"03",X"FC",X"00",X"AE",
		X"0B",X"5F",X"E1",X"D2",X"91",X"1F",X"84",X"FF",X"00",X"FF",X"40",X"2F",X"05",X"FE",X"01",X"FE",
		X"01",X"FF",X"40",X"7F",X"00",X"FF",X"40",X"FF",X"40",X"3F",X"C0",X"F7",X"40",X"5F",X"E1",X"D2",
		X"46",X"1F",X"F8",X"81",X"0F",X"9E",X"07",X"BF",X"50",X"7D",X"D0",X"3E",X"30",X"FC",X"01",X"BE",
		X"78",X"F0",X"C1",X"C7",X"83",X"F4",X"03",X"FE",X"41",X"F1",X"43",X"5E",X"3F",X"F0",X"92",X"C0",
		X"1F",X"F0",X"1F",X"F0",X"1F",X"F0",X"0F",X"F0",X"0F",X"F0",X"0B",X"F0",X"0F",X"F4",X"0F",X"F0",
		X"03",X"F4",X"0F",X"F0",X"0F",X"F8",X"0B",X"28",X"FD",X"80",X"3F",X"F0",X"2F",X"C0",X"3F",X"40",
		X"FF",X"00",X"3F",X"00",X"FE",X"42",X"FF",X"00",X"FD",X"01",X"BF",X"E0",X"C3",X"0B",X"F9",X"D1",
		X"74",X"E5",X"06",X"8F",X"03",X"3F",X"3D",X"F0",X"0F",X"D0",X"0F",X"F0",X"1F",X"E0",X"3F",X"D0",
		X"0F",X"C0",X"1F",X"F4",X"7D",X"C0",X"0F",X"0D",X"2F",X"F0",X"07",X"E6",X"1F",X"E0",X"1F",X"C0",
		X"6F",X"80",X"3F",X"F0",X"2F",X"C0",X"7F",X"80",X"AF",X"C0",X"BF",X"00",X"FF",X"00",X"3F",X"40",
		X"FF",X"C0",X"FA",X"80",X"77",X"B4",X"F0",X"E1",X"C1",X"E3",X"82",X"CF",X"06",X"BC",X"0F",X"F4",
		X"00",X"03",X"06",X"09",X"0C",X"0F",X"12",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",
		X"30",X"33",X"36",X"39",X"3C",X"3F",X"42",X"45",X"48",X"4B",X"4E",X"51",X"54",X"57",X"5A",X"5D",
		X"60",X"5D",X"5A",X"57",X"54",X"51",X"4E",X"4B",X"48",X"45",X"42",X"3F",X"3C",X"39",X"36",X"33",
		X"30",X"2D",X"2A",X"27",X"24",X"21",X"1E",X"1B",X"18",X"15",X"12",X"0F",X"0C",X"09",X"06",X"03",
		X"42",X"03",X"78",X"62",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",X"A3",X"A8",
		X"C5",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"53",X"3F",X"A3",X"D5",X"68",X"39",X"16",
		X"63",X"C4",X"44",X"C5",X"E5",X"83",X"07",X"CB",X"0F",X"1D",X"3D",X"3C",X"E4",X"B7",X"40",X"7F",
		X"00",X"7F",X"40",X"7F",X"3D",X"F0",X"C3",X"81",X"FF",X"00",X"FD",X"03",X"F8",X"0B",X"F0",X"0F",
		X"D0",X"2F",X"08",X"FF",X"06",X"F8",X"3E",X"C0",X"1F",X"C0",X"3F",X"38",X"F8",X"F0",X"D0",X"D7",
		X"03",X"FC",X"42",X"F8",X"43",X"0B",X"FD",X"30",X"E8",X"0F",X"B0",X"6F",X"40",X"FF",X"10",X"FC",
		X"BA",X"C0",X"2F",X"00",X"FF",X"02",X"FC",X"52",X"A9",X"92",X"2F",X"E0",X"5F",X"E0",X"9E",X"01",
		X"FD",X"C2",X"61",X"FD",X"01",X"FC",X"16",X"F0",X"1F",X"D0",X"1F",X"B5",X"15",X"F5",X"03",X"FC",
		X"00",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0E",X"10",X"12",X"14",X"16",X"18",X"1A",X"1C",X"1E",
		X"20",X"22",X"24",X"26",X"28",X"2A",X"2C",X"2E",X"30",X"32",X"34",X"36",X"38",X"3A",X"3C",X"3E",
		X"40",X"3E",X"3C",X"3A",X"38",X"36",X"34",X"32",X"30",X"2E",X"2C",X"2A",X"28",X"26",X"24",X"22",
		X"20",X"1E",X"1C",X"1A",X"18",X"16",X"14",X"12",X"10",X"0E",X"0C",X"0A",X"08",X"06",X"04",X"02",
		X"00",X"03",X"06",X"09",X"0C",X"0F",X"12",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",
		X"30",X"33",X"36",X"39",X"3C",X"3F",X"42",X"45",X"48",X"4B",X"4E",X"51",X"54",X"57",X"5A",X"5D",
		X"60",X"5D",X"5A",X"57",X"54",X"51",X"4E",X"4B",X"48",X"45",X"42",X"3F",X"3C",X"39",X"36",X"33",
		X"30",X"2D",X"2A",X"27",X"24",X"21",X"1E",X"1B",X"18",X"15",X"12",X"0F",X"0C",X"09",X"06",X"03",
		X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"53",X"3F",X"A3",X"A8",X"C5",X"FC",X"6E",X"AC",
		X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",X"A3",X"D5",X"68",X"39",X"16",X"5F",X"E4",X"40",X"C5",
		X"E5",X"83",X"5F",X"91",X"7A",X"C1",X"6B",X"51",X"7E",X"A0",X"FA",X"80",X"AF",X"10",X"FD",X"03",
		X"F9",X"07",X"B8",X"2A",X"A4",X"5F",X"51",X"6E",X"55",X"6D",X"59",X"1A",X"AA",X"5A",X"A5",X"1E",
		X"B8",X"65",X"B5",X"52",X"B9",X"46",X"A5",X"0F",X"E5",X"59",X"65",X"5E",X"E1",X"46",X"9E",X"92",
		X"6A",X"5A",X"4A",X"7E",X"64",X"A5",X"4E",X"56",X"2E",X"96",X"66",X"A5",X"76",X"54",X"AE",X"45",
		X"EA",X"25",X"F8",X"D1",X"E1",X"07",X"B9",X"55",X"9A",X"A5",X"E5",X"91",X"4B",X"A9",X"57",X"D4",
		X"0B",X"6D",X"69",X"A5",X"53",X"B9",X"05",X"BE",X"05",X"FD",X"54",X"EA",X"42",X"BA",X"55",X"69",
		X"00",X"05",X"0A",X"0F",X"14",X"19",X"1E",X"23",X"28",X"2D",X"32",X"37",X"3C",X"41",X"46",X"4B",
		X"50",X"55",X"5A",X"5F",X"64",X"69",X"6E",X"73",X"78",X"7D",X"82",X"87",X"8C",X"91",X"96",X"9B",
		X"9F",X"9B",X"96",X"91",X"8C",X"87",X"82",X"7D",X"78",X"73",X"6E",X"69",X"64",X"5F",X"5A",X"55",
		X"50",X"4B",X"46",X"41",X"3C",X"37",X"32",X"2D",X"28",X"23",X"1E",X"19",X"14",X"0F",X"0A",X"05");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
