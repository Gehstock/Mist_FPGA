library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bagman_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bagman_tile_bit0 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"18",X"0C",X"1C",X"5C",X"F8",
		X"60",X"74",X"7D",X"79",X"3E",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"EC",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"1C",X"1F",X"1F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"60",X"F8",X"F8",X"F8",X"F0",
		X"7F",X"7F",X"7F",X"1B",X"03",X"01",X"00",X"00",X"F0",X"FC",X"FC",X"FC",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"74",X"00",X"00",X"00",X"18",X"0C",X"5C",X"DC",X"F8",
		X"7D",X"79",X"3E",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"EC",X"C0",X"80",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"3F",X"3F",X"3F",X"07",X"0F",X"1F",X"07",X"0F",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"03",X"0F",
		X"04",X"04",X"00",X"20",X"70",X"21",X"00",X"80",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"0F",X"8F",
		X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"EF",X"FF",X"0F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"00",X"00",X"18",X"3C",X"3C",X"3C",X"3F",
		X"07",X"07",X"06",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"7E",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"7C",X"FC",
		X"3F",X"3F",X"79",X"3E",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"60",X"75",X"7D",X"79",X"3E",X"00",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"07",X"07",X"07",X"0F",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"3F",X"07",X"47",X"C3",X"EB",X"FB",X"F2",X"7C",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1D",X"00",X"00",X"00",X"70",X"70",X"E0",X"E0",X"EC",
		X"0F",X"07",X"43",X"C1",X"E9",X"FB",X"F6",X"7C",X"F8",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C1",X"00",X"00",X"00",X"00",X"38",X"78",X"F8",X"F0",
		X"E9",X"FB",X"F3",X"7D",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"F8",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"3A",X"00",X"00",X"00",X"00",X"08",X"1C",X"3C",X"7C",
		X"3E",X"3C",X"1F",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"78",X"7C",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"0C",X"1C",X"DC",X"F8",
		X"74",X"7D",X"79",X"3E",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"4C",X"5C",
		X"74",X"7D",X"79",X"3E",X"00",X"00",X"00",X"00",X"D8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"3F",X"3F",X"3F",X"07",X"0F",X"1F",X"07",X"07",
		X"02",X"20",X"70",X"20",X"00",X"04",X"0E",X"04",X"07",X"03",X"00",X"06",X"02",X"07",X"7F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"3F",X"3F",X"3F",X"07",X"07",X"0F",X"03",X"0F",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"03",X"00",X"06",X"02",X"07",X"7F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"07",X"0F",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"06",X"02",X"07",X"7F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"3F",X"3F",X"07",X"0F",X"8F",X"8F",X"8F",
		X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"CF",X"FF",X"3F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"0C",X"00",X"00",X"00",X"18",X"1C",X"3C",X"3C",X"3F",
		X"07",X"07",X"0F",X"07",X"01",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"FF",X"FE",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"7C",X"FC",
		X"3F",X"3F",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"1F",X"1F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"F0",
		X"7F",X"7F",X"7F",X"1B",X"03",X"01",X"00",X"00",X"F0",X"FC",X"FC",X"FC",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"00",X"00",X"10",X"18",X"1C",X"0C",X"5C",X"D8",
		X"60",X"74",X"70",X"71",X"3E",X"08",X"00",X"00",X"FC",X"FC",X"FC",X"EC",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"74",X"00",X"00",X"10",X"18",X"1C",X"4C",X"DC",X"D8",
		X"7D",X"71",X"3E",X"08",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"E0",X"C0",X"80",X"00",X"00",
		X"08",X"04",X"02",X"01",X"20",X"20",X"20",X"60",X"00",X"00",X"00",X"00",X"08",X"3C",X"FC",X"FC",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"80",X"80",X"5C",X"FC",X"FC",
		X"60",X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"F8",X"F8",X"FC",X"FC",X"F8",X"68",X"00",X"00",
		X"08",X"04",X"02",X"01",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"08",X"1C",X"7C",X"FC",
		X"60",X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"F8",X"F8",X"FC",X"FC",X"F8",X"68",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"20",X"20",X"20",X"00",X"28",X"1C",X"FC",X"FC",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"3A",X"10",X"10",X"10",X"00",X"18",X"1C",X"3C",X"7C",
		X"3E",X"38",X"1F",X"07",X"01",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"7C",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"80",X"80",X"80",X"00",X"9C",X"3C",X"7C",X"F8",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"F8",X"FC",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"40",X"40",X"40",X"00",X"4C",X"1C",X"DC",X"F8",
		X"74",X"7D",X"71",X"3E",X"0E",X"02",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"00",X"00",X"00",X"10",X"18",X"3C",X"4C",X"DC",
		X"74",X"70",X"71",X"3E",X"0E",X"02",X"00",X"00",X"D8",X"FC",X"FC",X"FC",X"6C",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"00",X"09",X"25",X"D4",X"B5",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"02",X"03",X"01",X"07",X"0F",X"0D",X"08",X"00",X"1C",X"7E",X"A3",X"FF",X"AB",X"FF",X"AB",X"8B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"08",X"08",X"0E",X"0F",X"0E",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0E",X"0F",X"0E",X"08",X"08",X"1C",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1C",X"1E",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"9F",X"8F",X"8F",X"87",X"83",X"81",X"80",
		X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"BF",
		X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"87",X"87",X"87",X"87",X"83",X"83",X"83",X"83",
		X"9F",X"9F",X"8F",X"8F",X"8F",X"8F",X"8F",X"87",X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",
		X"9F",X"9F",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"8F",X"8F",X"8F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"81",X"83",X"83",X"87",X"87",X"87",X"8F",X"8F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"9F",X"8F",X"87",X"87",X"83",X"81",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"87",X"83",X"83",X"81",X"81",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"8F",X"8F",X"8F",X"8F",X"87",X"87",X"87",X"87",X"8F",X"8F",X"8F",X"8F",X"9F",X"9F",X"9F",
		X"80",X"80",X"81",X"81",X"83",X"83",X"87",X"87",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"B8",X"B0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"BF",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"0C",X"10",X"30",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"26",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"64",X"74",X"7C",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"3A",X"18",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"64",X"74",X"7C",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"3A",X"09",X"08",X"08",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"01",X"01",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"A0",X"B8",X"B4",X"EA",X"AE",X"9A",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"10",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"10",X"30",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"30",X"30",X"30",X"70",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"70",X"70",X"70",X"70",X"70",X"70",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"03",X"06",X"0C",X"18",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F8",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"3C",X"7E",X"FF",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"FF",X"7E",X"3C",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"01",X"03",X"07",X"1F",X"1F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"0E",X"1E",X"1E",
		X"1E",X"1E",X"1E",X"10",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",
		X"00",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"00",X"10",X"18",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"47",X"57",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"18",X"00",X"00",X"00",
		X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"18",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"04",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"18",X"00",X"00",X"00",X"00",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"18",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"18",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"04",X"00",X"00",X"10",X"18",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"02",X"00",X"00",X"00",X"00",X"08",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"06",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"02",X"00",X"00",X"00",X"00",X"08",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"06",X"06",X"06",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"71",X"89",X"89",X"89",X"89",X"89",X"67",X"00",X"6E",X"91",X"91",X"91",X"91",X"91",X"6E",X"00",
		X"7E",X"91",X"91",X"91",X"91",X"91",X"61",X"00",X"FF",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"C3",X"A5",X"A5",X"A5",X"BD",X"C3",X"7E",X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",
		X"00",X"7F",X"02",X"04",X"08",X"10",X"20",X"7F",X"00",X"06",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",
		X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"8F",X"2F",X"EF",X"EF",X"EF",X"EF",X"8F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E3",
		X"8F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"37",X"77",X"77",X"37",X"87",X"E7",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"F8",X"F3",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F3",X"F8",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"2F",X"0F",X"7F",X"7F",
		X"3F",X"8F",X"E7",X"F7",X"F7",X"F7",X"F7",X"F7",X"0F",X"EF",X"EF",X"EF",X"CF",X"DF",X"DF",X"9F",
		X"87",X"BF",X"BF",X"BF",X"9F",X"DF",X"DF",X"CF",X"BF",X"BF",X"3F",X"7F",X"7F",X"7F",X"0F",X"EF",
		X"EF",X"EF",X"E7",X"F7",X"F7",X"F7",X"87",X"BF",X"EF",X"0F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"1F",X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"8F",X"1F",X"7F",X"FF",
		X"BF",X"87",X"F7",X"77",X"17",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"C7",X"F1",X"FC",X"FE",X"FE",
		X"FC",X"F1",X"C7",X"1F",X"7F",X"FF",X"FC",X"F9",X"C7",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F1",X"F4",X"F7",X"F7",X"F7",X"F7",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",X"F7",X"F7",X"F7",X"F7",X"F4",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"80",X"41",X"AA",X"00",X"00",X"00",X"02",X"15",X"2A",X"55",X"AA",
		X"00",X"00",X"00",X"80",X"40",X"A8",X"55",X"AA",X"01",X"02",X"15",X"AA",X"55",X"AA",X"55",X"AA",
		X"40",X"80",X"50",X"A8",X"55",X"AA",X"55",X"AA",X"15",X"2A",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"50",X"A8",X"54",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"07",
		X"F0",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"03",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"FC",X"FC",X"FC",X"FC",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"00",X"01",X"01",X"01",X"00",X"00",X"10",X"10",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"78",X"38",X"00",X"00",X"10",X"10",X"1F",X"3F",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"1C",X"1E",X"1F",X"1F",X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"01",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7E",X"7C",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"7F",X"7F",X"7F",X"7F",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"01",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",
		X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"10",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"C0",X"FF",X"FF",X"FE",X"FE",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"00",X"00",X"10",X"10",
		X"80",X"80",X"80",X"80",X"00",X"00",X"10",X"10",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"0F",X"0F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",
		X"01",X"03",X"03",X"07",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"FE",X"FE",X"FF",X"FF",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"FE",X"FE",X"FF",X"FF",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"7F",X"3F",X"1F",X"0F",X"07",X"07",X"03",X"01",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"FF",X"7F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"00",X"01",X"03",X"03",X"07",X"0F",X"0F",X"1F",
		X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1E",X"1C",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"3F",X"3F",X"3F",X"7F",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",
		X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"60",X"20",X"00",X"00",X"10",X"10",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"0E",X"0C",X"00",X"00",X"10",X"10",
		X"00",X"00",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",
		X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FC",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",
		X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FE",X"FE",X"FE",X"00",X"00",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"F0",X"F8",X"F8",X"FC",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
