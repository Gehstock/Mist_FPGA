library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_pgm_rom4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_pgm_rom4 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"2A",X"03",X"3C",X"00",X"84",X"03",X"42",X"00",X"DE",X"03",X"48",X"00",X"38",X"04",X"4E",X"00",
		X"92",X"04",X"54",X"00",X"EC",X"04",X"5A",X"00",X"46",X"05",X"60",X"00",X"A0",X"05",X"12",X"00",
		X"5A",X"00",X"24",X"00",X"B4",X"00",X"36",X"00",X"0E",X"01",X"48",X"00",X"68",X"01",X"5A",X"00",
		X"C2",X"01",X"6C",X"00",X"1C",X"02",X"7E",X"00",X"76",X"02",X"90",X"00",X"D0",X"02",X"A2",X"00",
		X"2A",X"03",X"B4",X"00",X"84",X"03",X"C6",X"00",X"DE",X"03",X"D8",X"00",X"38",X"04",X"EA",X"00",
		X"92",X"04",X"FC",X"00",X"EC",X"04",X"0E",X"01",X"46",X"05",X"20",X"01",X"A0",X"05",X"18",X"00",
		X"54",X"00",X"30",X"00",X"A8",X"00",X"48",X"00",X"FC",X"00",X"60",X"00",X"50",X"01",X"78",X"00",
		X"A4",X"01",X"90",X"00",X"F8",X"01",X"A8",X"00",X"4C",X"02",X"C0",X"00",X"A0",X"02",X"D8",X"00",
		X"F4",X"02",X"F0",X"00",X"48",X"03",X"08",X"01",X"9C",X"03",X"20",X"01",X"F0",X"03",X"38",X"01",
		X"44",X"04",X"50",X"01",X"98",X"04",X"68",X"01",X"EC",X"04",X"80",X"01",X"40",X"05",X"24",X"00",
		X"54",X"00",X"48",X"00",X"A8",X"00",X"6C",X"00",X"FC",X"00",X"90",X"00",X"50",X"01",X"B4",X"00",
		X"A4",X"01",X"D8",X"00",X"F8",X"01",X"FC",X"00",X"4C",X"02",X"20",X"01",X"A0",X"02",X"44",X"01",
		X"F4",X"02",X"68",X"01",X"48",X"03",X"8C",X"01",X"9C",X"03",X"B0",X"01",X"F0",X"03",X"D4",X"01",
		X"44",X"04",X"F8",X"01",X"98",X"04",X"1C",X"02",X"EC",X"04",X"40",X"02",X"40",X"05",X"2A",X"00",
		X"4E",X"00",X"54",X"00",X"9C",X"00",X"7E",X"00",X"EA",X"00",X"A8",X"00",X"38",X"01",X"D2",X"00",
		X"86",X"01",X"FC",X"00",X"D4",X"01",X"26",X"01",X"22",X"02",X"50",X"01",X"70",X"02",X"7A",X"01",
		X"BE",X"02",X"A4",X"01",X"0C",X"03",X"CE",X"01",X"5A",X"03",X"F8",X"01",X"A8",X"03",X"22",X"02",
		X"F6",X"03",X"4C",X"02",X"44",X"04",X"76",X"02",X"92",X"04",X"A0",X"02",X"E0",X"04",X"30",X"00",
		X"48",X"00",X"60",X"00",X"90",X"00",X"90",X"00",X"D8",X"00",X"C0",X"00",X"20",X"01",X"F0",X"00",
		X"68",X"01",X"20",X"01",X"B0",X"01",X"50",X"01",X"F8",X"01",X"80",X"01",X"40",X"02",X"B0",X"01",
		X"88",X"02",X"E0",X"01",X"D0",X"02",X"10",X"02",X"18",X"03",X"40",X"02",X"60",X"03",X"70",X"02",
		X"A8",X"03",X"A0",X"02",X"F0",X"03",X"D0",X"02",X"38",X"04",X"00",X"03",X"80",X"04",X"3C",X"00",
		X"48",X"00",X"78",X"00",X"90",X"00",X"B4",X"00",X"D8",X"00",X"F0",X"00",X"20",X"01",X"2C",X"01",
		X"68",X"01",X"68",X"01",X"B0",X"01",X"A4",X"01",X"F8",X"01",X"E0",X"01",X"40",X"02",X"1C",X"02",
		X"88",X"02",X"58",X"02",X"D0",X"02",X"94",X"02",X"18",X"03",X"D0",X"02",X"60",X"03",X"0C",X"03",
		X"A8",X"03",X"48",X"03",X"F0",X"03",X"84",X"03",X"38",X"04",X"C0",X"03",X"80",X"04",X"42",X"00",
		X"42",X"00",X"84",X"00",X"84",X"00",X"C6",X"00",X"C6",X"00",X"08",X"01",X"08",X"01",X"4A",X"01",
		X"4A",X"01",X"8C",X"01",X"8C",X"01",X"CE",X"01",X"CE",X"01",X"10",X"02",X"10",X"02",X"52",X"02",
		X"52",X"02",X"94",X"02",X"94",X"02",X"D6",X"02",X"D6",X"02",X"18",X"03",X"18",X"03",X"5A",X"03",
		X"5A",X"03",X"9C",X"03",X"9C",X"03",X"DE",X"03",X"DE",X"03",X"20",X"04",X"20",X"04",X"48",X"00",
		X"3C",X"00",X"90",X"00",X"78",X"00",X"D8",X"00",X"B4",X"00",X"20",X"01",X"F0",X"00",X"68",X"01",
		X"2C",X"01",X"B0",X"01",X"68",X"01",X"F8",X"01",X"A4",X"01",X"40",X"02",X"E0",X"01",X"88",X"02",
		X"1C",X"02",X"D0",X"02",X"58",X"02",X"18",X"03",X"94",X"02",X"60",X"03",X"D0",X"02",X"A8",X"03",
		X"0C",X"03",X"F0",X"03",X"48",X"03",X"38",X"04",X"84",X"03",X"80",X"04",X"C0",X"03",X"48",X"00",
		X"30",X"00",X"90",X"00",X"60",X"00",X"D8",X"00",X"90",X"00",X"20",X"01",X"C0",X"00",X"68",X"01",
		X"F0",X"00",X"B0",X"01",X"20",X"01",X"F8",X"01",X"50",X"01",X"40",X"02",X"80",X"01",X"88",X"02",
		X"B0",X"01",X"D0",X"02",X"E0",X"01",X"18",X"03",X"10",X"02",X"60",X"03",X"40",X"02",X"A8",X"03",
		X"70",X"02",X"F0",X"03",X"A0",X"02",X"38",X"04",X"D0",X"02",X"80",X"04",X"00",X"03",X"4E",X"00",
		X"2A",X"00",X"9C",X"00",X"54",X"00",X"EA",X"00",X"7E",X"00",X"38",X"01",X"A8",X"00",X"86",X"01",
		X"D2",X"00",X"D4",X"01",X"FC",X"00",X"22",X"02",X"26",X"01",X"70",X"02",X"50",X"01",X"BE",X"02",
		X"7A",X"01",X"0C",X"03",X"A4",X"01",X"5A",X"03",X"CE",X"01",X"A8",X"03",X"F8",X"01",X"F6",X"03",
		X"22",X"02",X"44",X"04",X"4C",X"02",X"92",X"04",X"76",X"02",X"E0",X"04",X"A0",X"02",X"54",X"00",
		X"24",X"00",X"A8",X"00",X"48",X"00",X"FC",X"00",X"6C",X"00",X"50",X"01",X"90",X"00",X"A4",X"01",
		X"B4",X"00",X"F8",X"01",X"D8",X"00",X"4C",X"02",X"FC",X"00",X"A0",X"02",X"20",X"01",X"F4",X"02",
		X"44",X"01",X"48",X"03",X"68",X"01",X"9C",X"03",X"8C",X"01",X"F0",X"03",X"B0",X"01",X"44",X"04",
		X"D4",X"01",X"98",X"04",X"F8",X"01",X"EC",X"04",X"1C",X"02",X"40",X"05",X"40",X"02",X"54",X"00",
		X"18",X"00",X"A8",X"00",X"30",X"00",X"FC",X"00",X"48",X"00",X"50",X"01",X"60",X"00",X"A4",X"01",
		X"78",X"00",X"F8",X"01",X"90",X"00",X"4C",X"02",X"A8",X"00",X"A0",X"02",X"C0",X"00",X"F4",X"02",
		X"D8",X"00",X"48",X"03",X"F0",X"00",X"9C",X"03",X"08",X"01",X"F0",X"03",X"20",X"01",X"44",X"04",
		X"38",X"01",X"98",X"04",X"50",X"01",X"EC",X"04",X"68",X"01",X"40",X"05",X"80",X"01",X"5A",X"00",
		X"12",X"00",X"B4",X"00",X"24",X"00",X"0E",X"01",X"36",X"00",X"68",X"01",X"48",X"00",X"C2",X"01",
		X"5A",X"00",X"1C",X"02",X"6C",X"00",X"76",X"02",X"7E",X"00",X"D0",X"02",X"90",X"00",X"2A",X"03",
		X"A2",X"00",X"84",X"03",X"B4",X"00",X"DE",X"03",X"C6",X"00",X"38",X"04",X"D8",X"00",X"92",X"04",
		X"EA",X"00",X"EC",X"04",X"FC",X"00",X"46",X"05",X"0E",X"01",X"A0",X"05",X"20",X"01",X"5A",X"00",
		X"06",X"00",X"B4",X"00",X"0C",X"00",X"0E",X"01",X"12",X"00",X"68",X"01",X"18",X"00",X"C2",X"01",
		X"1E",X"00",X"1C",X"02",X"24",X"00",X"76",X"02",X"2A",X"00",X"D0",X"02",X"30",X"00",X"2A",X"03",
		X"36",X"00",X"84",X"03",X"3C",X"00",X"DE",X"03",X"42",X"00",X"38",X"04",X"48",X"00",X"92",X"04",
		X"4E",X"00",X"EC",X"04",X"54",X"00",X"46",X"05",X"5A",X"00",X"A0",X"05",X"60",X"00",X"5A",X"00",
		X"00",X"00",X"B4",X"00",X"00",X"00",X"0E",X"01",X"00",X"00",X"68",X"01",X"00",X"00",X"C2",X"01",
		X"00",X"00",X"1C",X"02",X"00",X"00",X"76",X"02",X"00",X"00",X"D0",X"02",X"00",X"00",X"2A",X"03",
		X"00",X"00",X"84",X"03",X"00",X"00",X"DE",X"03",X"00",X"00",X"38",X"04",X"00",X"00",X"92",X"04",
		X"00",X"00",X"EC",X"04",X"00",X"00",X"46",X"05",X"00",X"00",X"A0",X"05",X"00",X"00",X"A6",X"40",
		X"D0",X"06",X"AD",X"04",X"02",X"4C",X"EB",X"C3",X"BD",X"06",X"02",X"20",X"D9",X"A2",X"A6",X"40",
		X"BD",X"01",X"02",X"29",X"0F",X"A8",X"B9",X"13",X"B0",X"29",X"40",X"F0",X"03",X"4C",X"12",X"C6",
		X"BD",X"00",X"02",X"29",X"03",X"D0",X"0A",X"A5",X"6C",X"D0",X"06",X"A6",X"40",X"A5",X"73",X"F0",
		X"03",X"4C",X"5B",X"C6",X"20",X"7A",X"C5",X"20",X"8C",X"C4",X"A6",X"40",X"D0",X"06",X"AD",X"22",
		X"01",X"8D",X"D1",X"03",X"AC",X"22",X"01",X"B9",X"29",X"04",X"F0",X"2F",X"A8",X"29",X"C0",X"C9",
		X"40",X"F0",X"03",X"4C",X"3D",X"C4",X"E0",X"00",X"D0",X"03",X"4C",X"12",X"C6",X"98",X"29",X"3F",
		X"18",X"65",X"59",X"AA",X"A5",X"5B",X"DD",X"6E",X"BF",X"A5",X"5C",X"FD",X"6F",X"BF",X"F0",X"10",
		X"10",X"05",X"49",X"FF",X"18",X"69",X"01",X"C9",X"04",X"90",X"05",X"A6",X"40",X"4C",X"12",X"C6",
		X"A6",X"40",X"BD",X"01",X"02",X"29",X"0F",X"C9",X"06",X"D0",X"03",X"4C",X"C5",X"C5",X"98",X"29",
		X"C0",X"C9",X"C0",X"D0",X"03",X"4C",X"B7",X"C5",X"20",X"42",X"BD",X"AC",X"22",X"01",X"B9",X"56",
		X"D5",X"A6",X"40",X"9D",X"06",X"02",X"20",X"B4",X"C9",X"4C",X"5B",X"C6",X"A5",X"59",X"0A",X"85",
		X"19",X"A5",X"5A",X"2A",X"85",X"1B",X"A5",X"5B",X"C5",X"19",X"A5",X"5C",X"E5",X"1B",X"90",X"10",
		X"A0",X"05",X"A5",X"44",X"30",X"02",X"A0",X"0B",X"8C",X"22",X"01",X"A9",X"02",X"85",X"59",X"60",
		X"A5",X"59",X"18",X"65",X"19",X"85",X"19",X"A5",X"1B",X"65",X"5A",X"6A",X"66",X"19",X"4A",X"66",
		X"19",X"85",X"1B",X"A5",X"19",X"C5",X"5B",X"A5",X"1B",X"E5",X"5C",X"B0",X"30",X"A0",X"00",X"A5",
		X"42",X"10",X"0B",X"A0",X"0A",X"A5",X"44",X"10",X"0B",X"A0",X"06",X"4C",X"E4",X"C4",X"A5",X"44",
		X"10",X"02",X"A0",X"04",X"8C",X"22",X"01",X"46",X"5A",X"66",X"59",X"18",X"A5",X"59",X"65",X"5B",
		X"85",X"5B",X"A5",X"5A",X"65",X"5C",X"85",X"5C",X"A9",X"00",X"85",X"59",X"60",X"A5",X"5B",X"85",
		X"19",X"A5",X"5C",X"85",X"1B",X"06",X"19",X"26",X"1B",X"06",X"19",X"26",X"1B",X"B0",X"30",X"A5",
		X"19",X"65",X"5B",X"85",X"19",X"A5",X"1B",X"65",X"5C",X"85",X"1B",X"B0",X"22",X"A5",X"59",X"C5",
		X"19",X"A5",X"5A",X"E5",X"1B",X"90",X"18",X"A0",X"02",X"A5",X"42",X"10",X"02",X"A0",X"08",X"8C",
		X"22",X"01",X"A5",X"59",X"85",X"5B",X"A5",X"5A",X"85",X"5C",X"A9",X"00",X"85",X"59",X"60",X"A0",
		X"01",X"A5",X"42",X"10",X"0B",X"A0",X"07",X"A5",X"44",X"30",X"0B",X"A0",X"09",X"4C",X"56",X"C5",
		X"A5",X"44",X"10",X"02",X"A0",X"03",X"8C",X"22",X"01",X"06",X"59",X"26",X"5A",X"18",X"A5",X"59",
		X"65",X"5B",X"85",X"5B",X"A5",X"5A",X"65",X"5C",X"85",X"5C",X"B0",X"05",X"A9",X"04",X"85",X"59",
		X"60",X"A9",X"FF",X"85",X"5B",X"85",X"5C",X"4C",X"6C",X"C5",X"BD",X"09",X"02",X"85",X"59",X"BD",
		X"0A",X"02",X"85",X"5A",X"85",X"42",X"10",X"10",X"49",X"FF",X"85",X"5A",X"A5",X"59",X"49",X"FF",
		X"85",X"59",X"E6",X"59",X"D0",X"02",X"E6",X"5A",X"BD",X"0B",X"02",X"85",X"5B",X"BD",X"0C",X"02",
		X"85",X"5C",X"85",X"44",X"10",X"10",X"49",X"FF",X"85",X"5C",X"A5",X"5B",X"49",X"FF",X"85",X"5B",
		X"E6",X"5B",X"D0",X"02",X"E6",X"5C",X"60",X"AC",X"22",X"01",X"A6",X"40",X"BD",X"01",X"02",X"29",
		X"0F",X"C9",X"06",X"D0",X"1F",X"20",X"36",X"BD",X"AE",X"22",X"01",X"BD",X"29",X"04",X"20",X"CA",
		X"A1",X"A9",X"A1",X"A0",X"00",X"91",X"49",X"AC",X"22",X"01",X"A9",X"00",X"99",X"29",X"04",X"A6",
		X"40",X"4C",X"5B",X"C6",X"B9",X"62",X"BF",X"38",X"FD",X"06",X"02",X"38",X"E9",X"01",X"10",X"07",
		X"85",X"19",X"A9",X"40",X"18",X"65",X"19",X"29",X"3F",X"9D",X"06",X"02",X"BD",X"01",X"02",X"29",
		X"0F",X"D0",X"07",X"BD",X"06",X"02",X"09",X"80",X"85",X"82",X"20",X"B4",X"C9",X"20",X"42",X"BD",
		X"A6",X"40",X"BD",X"00",X"02",X"29",X"08",X"F0",X"01",X"60",X"E0",X"00",X"F0",X"09",X"BD",X"01",
		X"02",X"29",X"0F",X"C9",X"07",X"D0",X"34",X"BD",X"0A",X"02",X"85",X"59",X"BD",X"0C",X"02",X"85",
		X"5B",X"A9",X"07",X"85",X"5D",X"20",X"03",X"D5",X"A6",X"40",X"90",X"1F",X"BD",X"06",X"02",X"48",
		X"AC",X"22",X"01",X"B9",X"56",X"D5",X"A6",X"40",X"9D",X"06",X"02",X"20",X"B4",X"C9",X"20",X"70",
		X"C7",X"A6",X"40",X"68",X"9D",X"06",X"02",X"20",X"42",X"BD",X"60",X"20",X"70",X"C7",X"BD",X"00",
		X"02",X"29",X"02",X"F0",X"01",X"60",X"8A",X"D0",X"03",X"4C",X"CE",X"C6",X"BD",X"01",X"02",X"29",
		X"0F",X"C9",X"03",X"D0",X"20",X"A9",X"07",X"85",X"5D",X"BD",X"0A",X"02",X"85",X"59",X"BD",X"0C",
		X"02",X"85",X"5B",X"20",X"03",X"D5",X"90",X"03",X"4C",X"ED",X"C7",X"A9",X"00",X"85",X"5D",X"20",
		X"1F",X"D5",X"90",X"F4",X"60",X"BD",X"0A",X"02",X"10",X"05",X"49",X"FF",X"18",X"69",X"01",X"C9",
		X"70",X"90",X"17",X"A0",X"6E",X"BD",X"0A",X"02",X"10",X"02",X"A0",X"92",X"98",X"9D",X"0A",X"02",
		X"A9",X"00",X"9D",X"09",X"02",X"85",X"19",X"4C",X"E5",X"C6",X"BD",X"0C",X"02",X"10",X"05",X"49",
		X"FF",X"18",X"69",X"01",X"C9",X"60",X"B0",X"07",X"60",X"A9",X"03",X"9D",X"00",X"02",X"60",X"A0",
		X"5E",X"BD",X"0C",X"02",X"10",X"02",X"A0",X"A2",X"98",X"9D",X"0C",X"02",X"A9",X"00",X"9D",X"0B",
		X"02",X"A9",X"20",X"85",X"19",X"A5",X"6C",X"F0",X"29",X"8A",X"A8",X"BD",X"01",X"02",X"29",X"0F",
		X"AA",X"C9",X"04",X"F0",X"15",X"C9",X"08",X"F0",X"11",X"C9",X"09",X"F0",X"0D",X"C9",X"0A",X"F0",
		X"09",X"C9",X"06",X"D0",X"02",X"A2",X"02",X"FE",X"48",X"04",X"98",X"AA",X"A9",X"03",X"9D",X"00",
		X"02",X"60",X"E0",X"50",X"B0",X"03",X"4C",X"C9",X"C6",X"BD",X"01",X"02",X"29",X"0F",X"A8",X"B9",
		X"13",X"B0",X"A8",X"29",X"01",X"D0",X"A2",X"98",X"29",X"08",X"F0",X"2A",X"BD",X"00",X"02",X"29",
		X"03",X"F0",X"23",X"BD",X"01",X"02",X"29",X"0F",X"C9",X"09",X"D0",X"8D",X"CE",X"03",X"03",X"AD",
		X"03",X"03",X"C9",X"F5",X"D0",X"83",X"86",X"19",X"A9",X"01",X"85",X"59",X"A9",X"00",X"85",X"5A",
		X"85",X"5B",X"20",X"80",X"D1",X"60",X"A5",X"19",X"38",X"FD",X"06",X"02",X"38",X"E9",X"01",X"10",
		X"03",X"18",X"69",X"40",X"29",X"3F",X"9D",X"06",X"02",X"20",X"B4",X"C9",X"20",X"5B",X"C6",X"60",
		X"86",X"19",X"BD",X"07",X"02",X"85",X"4C",X"BD",X"08",X"02",X"85",X"4D",X"A2",X"03",X"A0",X"03",
		X"B1",X"4C",X"95",X"1B",X"88",X"CA",X"10",X"F8",X"A6",X"19",X"BD",X"06",X"02",X"C9",X"11",X"B0",
		X"15",X"20",X"AD",X"C7",X"18",X"BD",X"0B",X"02",X"65",X"1D",X"9D",X"0B",X"02",X"BD",X"0C",X"02",
		X"65",X"1E",X"9D",X"0C",X"02",X"60",X"C9",X"21",X"B0",X"15",X"20",X"C6",X"C7",X"18",X"BD",X"09",
		X"02",X"65",X"1B",X"9D",X"09",X"02",X"BD",X"0A",X"02",X"65",X"1C",X"9D",X"0A",X"02",X"60",X"C9",
		X"31",X"B0",X"15",X"20",X"DB",X"C7",X"38",X"BD",X"0B",X"02",X"E5",X"1D",X"9D",X"0B",X"02",X"BD",
		X"0C",X"02",X"E5",X"1E",X"9D",X"0C",X"02",X"60",X"20",X"94",X"C7",X"38",X"BD",X"09",X"02",X"E5",
		X"1B",X"9D",X"09",X"02",X"BD",X"0A",X"02",X"E5",X"1C",X"9D",X"0A",X"02",X"60",X"A9",X"00",X"85",
		X"59",X"9D",X"01",X"02",X"86",X"19",X"A9",X"13",X"0A",X"AA",X"BD",X"72",X"C9",X"85",X"5A",X"BD",
		X"73",X"C9",X"85",X"5B",X"8A",X"48",X"20",X"4E",X"BD",X"68",X"AA",X"AC",X"03",X"03",X"C0",X"04",
		X"B0",X"03",X"EE",X"03",X"03",X"F8",X"88",X"30",X"0B",X"BD",X"72",X"C9",X"18",X"65",X"5A",X"85",
		X"5A",X"4C",X"16",X"C8",X"D8",X"A5",X"5A",X"A8",X"A6",X"19",X"A9",X"60",X"9D",X"01",X"21",X"A9",
		X"00",X"9D",X"00",X"21",X"9D",X"06",X"21",X"A9",X"71",X"9D",X"0B",X"21",X"A9",X"00",X"9D",X"0A",
		X"21",X"A5",X"5B",X"4C",X"9D",X"C8",X"86",X"19",X"48",X"A5",X"79",X"8D",X"3E",X"04",X"A9",X"60",
		X"9D",X"01",X"21",X"A9",X"00",X"9D",X"00",X"21",X"9D",X"06",X"21",X"68",X"C9",X"22",X"D0",X"2C",
		X"24",X"EF",X"30",X"25",X"AD",X"39",X"04",X"F8",X"18",X"6D",X"43",X"04",X"8D",X"43",X"04",X"AD",
		X"38",X"04",X"6D",X"42",X"04",X"8D",X"42",X"04",X"AD",X"37",X"04",X"6D",X"41",X"04",X"8D",X"41",
		X"04",X"D8",X"A9",X"00",X"A0",X"00",X"20",X"1B",X"CA",X"4C",X"FD",X"C8",X"0A",X"AA",X"A9",X"00",
		X"85",X"59",X"BD",X"72",X"C9",X"A8",X"85",X"5A",X"BD",X"73",X"C9",X"85",X"5B",X"20",X"1B",X"CA",
		X"A6",X"19",X"BD",X"01",X"02",X"29",X"0F",X"A8",X"B9",X"13",X"B0",X"30",X"40",X"20",X"2E",X"BD",
		X"A9",X"00",X"85",X"1C",X"A5",X"19",X"18",X"69",X"04",X"85",X"11",X"A9",X"20",X"18",X"69",X"03",
		X"85",X"12",X"20",X"1D",X"C9",X"A6",X"19",X"8A",X"4A",X"4A",X"4A",X"38",X"E9",X"0A",X"A8",X"78",
		X"B9",X"B3",X"D8",X"9D",X"04",X"21",X"B9",X"B4",X"D8",X"9D",X"05",X"21",X"A9",X"00",X"9D",X"02",
		X"21",X"A9",X"70",X"9D",X"03",X"21",X"A9",X"02",X"9D",X"00",X"02",X"58",X"60",X"78",X"C0",X"0D",
		X"D0",X"0B",X"A0",X"05",X"A9",X"00",X"20",X"1B",X"CA",X"A9",X"01",X"D0",X"02",X"A9",X"02",X"9D",
		X"00",X"02",X"A9",X"00",X"9D",X"03",X"02",X"A9",X"01",X"9D",X"02",X"02",X"AD",X"64",X"56",X"9D",
		X"04",X"21",X"AD",X"65",X"56",X"9D",X"05",X"21",X"58",X"20",X"4A",X"BD",X"60",X"A5",X"59",X"29",
		X"0F",X"38",X"F0",X"03",X"18",X"C6",X"1C",X"20",X"AF",X"D7",X"A5",X"5A",X"4A",X"4A",X"4A",X"4A",
		X"20",X"4B",X"C9",X"A5",X"5A",X"29",X"0F",X"20",X"4B",X"C9",X"A5",X"5B",X"4A",X"4A",X"4A",X"4A",
		X"18",X"20",X"AF",X"D7",X"A5",X"5B",X"18",X"20",X"AF",X"D7",X"60",X"18",X"F0",X"05",X"C6",X"1C",
		X"4C",X"AF",X"D7",X"24",X"1C",X"30",X"01",X"38",X"4C",X"AF",X"D7",X"A6",X"40",X"A5",X"08",X"9D",
		X"09",X"02",X"A5",X"09",X"9D",X"0A",X"02",X"A5",X"0A",X"9D",X"0B",X"02",X"A5",X"0B",X"9D",X"0C",
		X"02",X"60",X"00",X"25",X"00",X"50",X"00",X"75",X"01",X"00",X"01",X"25",X"01",X"50",X"01",X"75",
		X"02",X"00",X"02",X"25",X"02",X"50",X"02",X"75",X"03",X"00",X"03",X"25",X"03",X"50",X"03",X"75",
		X"04",X"00",X"04",X"25",X"04",X"50",X"04",X"75",X"05",X"00",X"05",X"25",X"05",X"50",X"05",X"75",
		X"06",X"00",X"06",X"25",X"06",X"50",X"06",X"75",X"07",X"00",X"07",X"25",X"07",X"50",X"07",X"75",
		X"08",X"00",X"10",X"00",X"E0",X"50",X"B0",X"13",X"24",X"EF",X"30",X"0F",X"A5",X"73",X"D0",X"0B",
		X"BD",X"06",X"02",X"18",X"69",X"04",X"29",X"38",X"9D",X"06",X"02",X"BD",X"06",X"02",X"85",X"1D",
		X"C9",X"11",X"90",X"20",X"C9",X"21",X"B0",X"0A",X"A9",X"20",X"38",X"E5",X"1D",X"85",X"1D",X"4C",
		X"F4",X"C9",X"C9",X"31",X"B0",X"08",X"38",X"E9",X"20",X"85",X"1D",X"4C",X"F4",X"C9",X"A9",X"40",
		X"E5",X"1D",X"85",X"1D",X"BD",X"05",X"02",X"0A",X"0A",X"0A",X"0A",X"85",X"1C",X"A5",X"1D",X"29",
		X"1F",X"4A",X"66",X"1C",X"4A",X"66",X"1C",X"85",X"1B",X"A9",X"9E",X"18",X"65",X"1C",X"9D",X"07",
		X"02",X"A9",X"BF",X"65",X"1B",X"9D",X"08",X"02",X"60",X"D4",X"00",X"24",X"EF",X"30",X"67",X"18",
		X"F8",X"6D",X"43",X"04",X"8D",X"43",X"04",X"98",X"6D",X"42",X"04",X"8D",X"42",X"04",X"90",X"08",
		X"AD",X"41",X"04",X"69",X"00",X"8D",X"41",X"04",X"D8",X"AC",X"45",X"04",X"F0",X"48",X"F8",X"A0",
		X"00",X"AD",X"41",X"04",X"C8",X"38",X"ED",X"45",X"04",X"10",X"F9",X"D8",X"88",X"CC",X"47",X"04",
		X"F0",X"34",X"8C",X"47",X"04",X"8A",X"48",X"98",X"48",X"AD",X"40",X"04",X"C9",X"06",X"B0",X"1F",
		X"EE",X"40",X"04",X"AD",X"C8",X"04",X"F0",X"0E",X"AD",X"C9",X"04",X"F0",X"09",X"AD",X"40",X"04",
		X"8D",X"AA",X"04",X"4C",X"7C",X"CA",X"AD",X"40",X"04",X"8D",X"75",X"04",X"20",X"3B",X"9C",X"20",
		X"3A",X"BD",X"68",X"A8",X"68",X"AA",X"60",X"AD",X"C9",X"04",X"F0",X"15",X"AD",X"41",X"04",X"8D",
		X"AB",X"04",X"AD",X"42",X"04",X"8D",X"AC",X"04",X"AD",X"43",X"04",X"8D",X"AD",X"04",X"4C",X"B3",
		X"CA",X"AD",X"41",X"04",X"8D",X"76",X"04",X"AD",X"42",X"04",X"8D",X"77",X"04",X"AD",X"43",X"04",
		X"8D",X"78",X"04",X"AD",X"76",X"04",X"8D",X"41",X"04",X"AD",X"77",X"04",X"8D",X"42",X"04",X"AD",
		X"78",X"04",X"8D",X"43",X"04",X"A5",X"54",X"85",X"12",X"A5",X"53",X"85",X"11",X"A0",X"00",X"A2",
		X"C4",X"24",X"EF",X"30",X"0C",X"AD",X"C9",X"04",X"D0",X"07",X"2C",X"D0",X"03",X"10",X"02",X"A2",
		X"C7",X"8A",X"91",X"11",X"20",X"33",X"CB",X"AD",X"AB",X"04",X"8D",X"41",X"04",X"AD",X"AC",X"04",
		X"8D",X"42",X"04",X"AD",X"AD",X"04",X"8D",X"43",X"04",X"A5",X"55",X"85",X"11",X"A5",X"56",X"85",
		X"12",X"A0",X"00",X"A2",X"C4",X"24",X"EF",X"30",X"0C",X"AD",X"C9",X"04",X"F0",X"07",X"2C",X"D0",
		X"03",X"10",X"02",X"A2",X"C7",X"8A",X"91",X"11",X"20",X"33",X"CB",X"AD",X"C9",X"04",X"D0",X"12",
		X"AD",X"76",X"04",X"8D",X"41",X"04",X"AD",X"77",X"04",X"8D",X"42",X"04",X"AD",X"78",X"04",X"8D",
		X"43",X"04",X"60",X"A9",X"06",X"18",X"65",X"11",X"85",X"11",X"A2",X"00",X"A0",X"00",X"84",X"19",
		X"BD",X"41",X"04",X"4A",X"4A",X"4A",X"4A",X"F0",X"02",X"C6",X"19",X"24",X"19",X"18",X"30",X"01",
		X"38",X"86",X"1B",X"20",X"AF",X"D7",X"A6",X"1B",X"BD",X"41",X"04",X"29",X"0F",X"F0",X"02",X"C6",
		X"19",X"24",X"19",X"18",X"30",X"01",X"38",X"20",X"AF",X"D7",X"A6",X"1B",X"E8",X"E0",X"03",X"D0",
		X"CF",X"60",X"CE",X"50",X"0B",X"E4",X"00",X"01",X"90",X"E0",X"10",X"0B",X"E1",X"00",X"01",X"AD",
		X"20",X"04",X"C9",X"03",X"F0",X"16",X"AD",X"C8",X"04",X"F0",X"11",X"A2",X"02",X"20",X"B7",X"DC",
		X"AD",X"C9",X"04",X"18",X"69",X"01",X"20",X"AF",X"D7",X"4C",X"A1",X"CB",X"A2",X"10",X"20",X"B7",
		X"DC",X"AD",X"72",X"CB",X"85",X"59",X"AD",X"73",X"CB",X"85",X"5B",X"AD",X"74",X"CB",X"85",X"65",
		X"AD",X"75",X"CB",X"85",X"63",X"AD",X"76",X"CB",X"85",X"5A",X"AD",X"77",X"CB",X"85",X"5C",X"A9",
		X"00",X"85",X"19",X"85",X"1D",X"85",X"0C",X"A9",X"01",X"85",X"1C",X"20",X"3B",X"CD",X"A9",X"00",
		X"20",X"2C",X"CC",X"A6",X"19",X"BD",X"16",X"03",X"20",X"3F",X"CC",X"88",X"20",X"05",X"D8",X"A5",
		X"5B",X"38",X"E5",X"65",X"85",X"5B",X"A5",X"19",X"18",X"69",X"07",X"85",X"19",X"E6",X"1D",X"A5",
		X"1C",X"C9",X"11",X"D0",X"21",X"AD",X"78",X"CB",X"85",X"59",X"AD",X"79",X"CB",X"85",X"5B",X"AD",
		X"7B",X"CB",X"85",X"65",X"AD",X"7C",X"CB",X"85",X"63",X"AD",X"7D",X"CB",X"85",X"5A",X"AD",X"7E",
		X"CB",X"85",X"5C",X"4C",X"CB",X"CB",X"C9",X"21",X"90",X"01",X"60",X"C9",X"16",X"D0",X"F4",X"AD",
		X"7A",X"CB",X"85",X"59",X"AD",X"79",X"CB",X"85",X"5B",X"4C",X"13",X"CC",X"AA",X"F0",X"04",X"0A",
		X"69",X"14",X"AA",X"BD",X"C4",X"5D",X"20",X"6F",X"CC",X"BD",X"C5",X"5D",X"4C",X"6F",X"CC",X"A2",
		X"00",X"86",X"64",X"48",X"29",X"F0",X"4A",X"4A",X"4A",X"20",X"50",X"CC",X"68",X"29",X"0F",X"0A",
		X"F0",X"07",X"A2",X"FF",X"86",X"64",X"4C",X"62",X"CC",X"24",X"64",X"30",X"05",X"A2",X"00",X"4C",
		X"66",X"CC",X"18",X"69",X"02",X"AA",X"BD",X"C4",X"5D",X"20",X"6F",X"CC",X"BD",X"C5",X"5D",X"91",
		X"11",X"C8",X"D0",X"02",X"E6",X"12",X"60",X"E6",X"A3",X"A5",X"19",X"18",X"69",X"07",X"C9",X"8C",
		X"90",X"14",X"A9",X"01",X"8D",X"21",X"04",X"A9",X"FF",X"85",X"A3",X"A9",X"00",X"85",X"A4",X"60",
		X"A9",X"00",X"85",X"A3",X"85",X"A4",X"85",X"19",X"38",X"A6",X"19",X"BD",X"15",X"03",X"ED",X"43",
		X"04",X"BD",X"14",X"03",X"ED",X"42",X"04",X"BD",X"13",X"03",X"ED",X"41",X"04",X"B0",X"C8",X"E0",
		X"85",X"F0",X"51",X"A0",X"85",X"B9",X"16",X"03",X"D0",X"0C",X"98",X"38",X"E9",X"07",X"A8",X"10",
		X"F4",X"A2",X"00",X"4C",X"04",X"CD",X"98",X"18",X"69",X"07",X"AA",X"C5",X"19",X"F0",X"35",X"A8",
		X"38",X"E9",X"07",X"AA",X"BD",X"10",X"03",X"99",X"10",X"03",X"BD",X"11",X"03",X"99",X"11",X"03",
		X"BD",X"12",X"03",X"99",X"12",X"03",X"BD",X"13",X"03",X"99",X"13",X"03",X"BD",X"14",X"03",X"99",
		X"14",X"03",X"BD",X"15",X"03",X"99",X"15",X"03",X"BD",X"16",X"03",X"99",X"16",X"03",X"8A",X"A8",
		X"E4",X"19",X"D0",X"CC",X"86",X"A9",X"AD",X"41",X"04",X"9D",X"13",X"03",X"AD",X"42",X"04",X"9D",
		X"14",X"03",X"AD",X"43",X"04",X"9D",X"15",X"03",X"A9",X"00",X"9D",X"10",X"03",X"9D",X"11",X"03",
		X"9D",X"12",X"03",X"AD",X"5D",X"04",X"18",X"69",X"01",X"20",X"A1",X"DC",X"9D",X"16",X"03",X"20",
		X"0E",X"BE",X"20",X"5A",X"BD",X"A9",X"04",X"8D",X"21",X"04",X"60",X"20",X"C9",X"D8",X"A0",X"00",
		X"A9",X"01",X"20",X"12",X"D8",X"A5",X"59",X"A6",X"5B",X"20",X"1D",X"D8",X"A4",X"5A",X"A5",X"5C",
		X"20",X"12",X"D8",X"A5",X"1D",X"C5",X"A3",X"D0",X"08",X"A5",X"11",X"85",X"A3",X"A5",X"12",X"85",
		X"A4",X"A4",X"63",X"A9",X"00",X"20",X"EF",X"D7",X"A0",X"00",X"AD",X"20",X"04",X"F0",X"17",X"C9",
		X"01",X"F0",X"13",X"A5",X"1C",X"20",X"3F",X"CC",X"A9",X"00",X"20",X"2C",X"CC",X"F8",X"18",X"A9",
		X"01",X"65",X"1C",X"85",X"1C",X"D8",X"A6",X"19",X"BD",X"10",X"03",X"20",X"DD",X"CD",X"BD",X"10",
		X"03",X"29",X"1F",X"20",X"2C",X"CC",X"A6",X"19",X"BD",X"11",X"03",X"20",X"DD",X"CD",X"BD",X"11",
		X"03",X"29",X"1F",X"20",X"2C",X"CC",X"A6",X"19",X"BD",X"12",X"03",X"20",X"DD",X"CD",X"BD",X"12",
		X"03",X"29",X"1F",X"20",X"2C",X"CC",X"A5",X"63",X"20",X"6F",X"CC",X"A9",X"60",X"20",X"6F",X"CC",
		X"A9",X"00",X"20",X"2C",X"CC",X"A6",X"19",X"BD",X"13",X"03",X"20",X"3F",X"CC",X"A6",X"19",X"BD",
		X"14",X"03",X"20",X"43",X"CC",X"A6",X"19",X"BD",X"15",X"03",X"4C",X"43",X"CC",X"4A",X"4A",X"4A",
		X"4A",X"4A",X"4A",X"AA",X"BD",X"F2",X"CD",X"A6",X"19",X"20",X"6F",X"CC",X"A9",X"60",X"20",X"6F",
		X"CC",X"60",X"C4",X"C2",X"C1",X"C7",X"A2",X"00",X"A9",X"00",X"9D",X"10",X"03",X"E8",X"E0",X"8C",
		X"D0",X"F6",X"60",X"BD",X"0A",X"02",X"C9",X"80",X"6A",X"85",X"67",X"B9",X"0A",X"02",X"C9",X"80",
		X"6A",X"38",X"E5",X"67",X"85",X"42",X"10",X"05",X"49",X"FF",X"18",X"69",X"01",X"85",X"43",X"4A",
		X"85",X"67",X"BD",X"0C",X"02",X"C9",X"80",X"6A",X"85",X"69",X"B9",X"0C",X"02",X"C9",X"80",X"6A",
		X"38",X"E5",X"69",X"85",X"44",X"10",X"05",X"49",X"FF",X"18",X"69",X"01",X"85",X"45",X"4A",X"85",
		X"69",X"C5",X"67",X"90",X"0E",X"A5",X"67",X"18",X"65",X"43",X"4A",X"4A",X"4A",X"18",X"65",X"69",
		X"4C",X"5E",X"CE",X"A5",X"69",X"18",X"65",X"45",X"4A",X"4A",X"4A",X"18",X"65",X"67",X"C5",X"46",
		X"B0",X"50",X"2C",X"00",X"03",X"10",X"3C",X"98",X"AA",X"D0",X"11",X"A5",X"F6",X"C9",X"03",X"F0",
		X"0A",X"A5",X"1B",X"85",X"6C",X"20",X"0E",X"BE",X"20",X"52",X"BD",X"60",X"BD",X"01",X"02",X"29",
		X"0F",X"C9",X"0E",X"90",X"06",X"A8",X"A9",X"01",X"99",X"48",X"04",X"BD",X"01",X"02",X"29",X"0F",
		X"C9",X"05",X"D0",X"0A",X"A9",X"01",X"9D",X"0D",X"02",X"A9",X"22",X"4C",X"46",X"C8",X"A9",X"13",
		X"4C",X"46",X"C8",X"84",X"48",X"85",X"46",X"A6",X"44",X"A4",X"42",X"20",X"69",X"A2",X"29",X"3F",
		X"85",X"47",X"60",X"A6",X"40",X"A9",X"00",X"85",X"21",X"BD",X"00",X"02",X"29",X"02",X"F0",X"04",
		X"60",X"4C",X"25",X"CF",X"B9",X"00",X"02",X"29",X"02",X"D0",X"F6",X"C4",X"40",X"F0",X"F2",X"A6",
		X"40",X"38",X"BD",X"0A",X"02",X"F9",X"0A",X"02",X"85",X"42",X"10",X"06",X"49",X"FF",X"85",X"42",
		X"E6",X"42",X"38",X"BD",X"0C",X"02",X"F9",X"0C",X"02",X"85",X"44",X"10",X"06",X"49",X"FF",X"85",
		X"44",X"E6",X"44",X"18",X"B9",X"0F",X"02",X"7D",X"0F",X"02",X"C5",X"42",X"90",X"27",X"C5",X"44",
		X"90",X"23",X"85",X"46",X"0A",X"65",X"46",X"4A",X"85",X"46",X"A5",X"42",X"18",X"65",X"44",X"B0",
		X"14",X"C5",X"46",X"B0",X"10",X"A6",X"21",X"E8",X"98",X"95",X"21",X"E8",X"B9",X"01",X"02",X"29",
		X"0F",X"95",X"21",X"86",X"21",X"98",X"18",X"69",X"10",X"A8",X"B0",X"03",X"4C",X"C4",X"CE",X"60",
		X"A5",X"40",X"85",X"6E",X"4C",X"3F",X"CF",X"C6",X"21",X"C6",X"21",X"A5",X"6E",X"85",X"40",X"A8",
		X"A6",X"21",X"F0",X"65",X"B5",X"21",X"85",X"19",X"B9",X"00",X"02",X"29",X"02",X"D0",X"E8",X"B9",
		X"01",X"02",X"29",X"0F",X"85",X"1B",X"C5",X"19",X"D0",X"18",X"84",X"40",X"A8",X"CA",X"B5",X"21",
		X"85",X"41",X"98",X"0A",X"AA",X"BD",X"AB",X"CF",X"48",X"BD",X"AA",X"CF",X"48",X"A4",X"41",X"A6",
		X"40",X"60",X"B0",X"0E",X"85",X"19",X"B5",X"21",X"85",X"1B",X"CA",X"B5",X"21",X"85",X"41",X"4C",
		X"89",X"CF",X"84",X"41",X"CA",X"B5",X"21",X"85",X"40",X"C6",X"1B",X"A5",X"1B",X"38",X"E5",X"19",
		X"85",X"1B",X"A5",X"19",X"AA",X"BD",X"CA",X"CF",X"06",X"1B",X"65",X"1B",X"AA",X"BD",X"DA",X"CF",
		X"48",X"BD",X"D9",X"CF",X"48",X"A4",X"41",X"A6",X"40",X"60",X"CF",X"D3",X"36",X"CF",X"CF",X"D3",
		X"E0",X"D3",X"36",X"CF",X"36",X"CF",X"CF",X"D3",X"CF",X"D3",X"36",X"CF",X"36",X"CF",X"CF",X"D3",
		X"36",X"CF",X"36",X"CF",X"36",X"CF",X"90",X"D4",X"36",X"CF",X"00",X"1E",X"3A",X"54",X"6C",X"82",
		X"96",X"A8",X"B8",X"C6",X"D2",X"DC",X"E4",X"EA",X"EE",X"C8",X"D0",X"CD",X"D0",X"36",X"CF",X"D0",
		X"D0",X"36",X"CF",X"36",X"CF",X"2B",X"D1",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"90",X"D4",X"BC",X"D4",X"12",X"D2",X"15",X"D3",X"41",X"D3",X"36",X"CF",X"12");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
