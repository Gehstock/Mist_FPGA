library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"0B",X"0E",X"0B",X"0F",X"01",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"CC",X"FF",X"FF",X"F3",X"F0",X"F0",X"F3",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"F0",
		X"F0",X"F0",X"F3",X"FF",X"FF",X"CC",X"88",X"88",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F3",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"0C",X"00",X"0E",X"0F",X"0F",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"11",X"11",X"33",X"FF",X"FF",X"FC",X"F0",X"F0",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"F0",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"F0",X"F0",X"FC",X"FF",X"FF",X"33",X"11",X"11",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"87",X"C3",X"C3",X"C3",X"C0",X"00",X"00",X"E1",X"F0",X"F0",X"30",X"10",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"0F",X"0F",X"00",X"00",X"00",X"F8",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"FF",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"FF",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"0F",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",
		X"00",X"00",X"C0",X"C3",X"C3",X"C3",X"87",X"0F",X"00",X"00",X"00",X"10",X"30",X"F0",X"F0",X"E1",
		X"00",X"00",X"00",X"0F",X"0F",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"F8",
		X"FF",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"FF",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"0F",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"33",X"00",X"00",X"00",
		X"F0",X"F0",X"70",X"70",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"30",X"10",X"10",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"10",X"10",X"30",X"30",X"70",X"70",X"F0",X"F0",
		X"10",X"10",X"30",X"30",X"70",X"70",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"F0",
		X"EE",X"FF",X"11",X"99",X"55",X"FF",X"EE",X"00",X"33",X"77",X"55",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",
		X"33",X"99",X"99",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"11",X"33",X"22",X"00",X"33",X"77",X"44",X"44",X"44",X"66",X"22",X"00",
		X"55",X"FF",X"FF",X"55",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"BB",X"AA",X"00",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"44",X"66",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"EE",X"FF",X"99",X"99",X"99",X"BB",X"22",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"0F",X"08",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"0F",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",
		X"88",X"88",X"88",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"77",X"33",X"11",X"00",X"00",
		X"99",X"AA",X"CC",X"FF",X"CC",X"AA",X"99",X"00",X"44",X"22",X"11",X"77",X"11",X"22",X"44",X"00",
		X"88",X"CC",X"EE",X"FF",X"88",X"88",X"88",X"00",X"00",X"11",X"33",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"15",X"15",X"19",X"22",X"CC",X"33",X"44",X"88",X"8A",X"8A",X"89",X"44",X"33",
		X"00",X"FF",X"FF",X"44",X"44",X"FF",X"FF",X"00",X"00",X"11",X"33",X"66",X"66",X"33",X"11",X"00",
		X"66",X"FF",X"99",X"99",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"EE",X"FF",X"11",X"11",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"33",X"11",X"DD",X"99",X"FF",X"FF",X"11",X"00",X"66",X"44",X"55",X"44",X"77",X"77",X"44",X"00",
		X"00",X"00",X"CC",X"99",X"FF",X"FF",X"11",X"00",X"66",X"44",X"55",X"44",X"77",X"77",X"44",X"00",
		X"FF",X"FF",X"99",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"44",X"77",X"77",X"44",X"00",X"00",
		X"00",X"00",X"EE",X"FF",X"11",X"77",X"66",X"00",X"44",X"44",X"77",X"77",X"44",X"44",X"00",X"00",
		X"11",X"33",X"EE",X"CC",X"FF",X"FF",X"11",X"00",X"66",X"77",X"11",X"00",X"77",X"77",X"44",X"00",
		X"33",X"11",X"11",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"44",X"77",X"77",X"44",X"00",
		X"FF",X"FF",X"88",X"CC",X"88",X"FF",X"FF",X"00",X"77",X"77",X"33",X"11",X"33",X"77",X"77",X"00",
		X"FF",X"FF",X"CC",X"88",X"00",X"FF",X"FF",X"00",X"77",X"77",X"00",X"11",X"33",X"77",X"77",X"00",
		X"CC",X"EE",X"33",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"66",X"33",X"11",X"00",
		X"00",X"88",X"88",X"99",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"DD",X"EE",X"55",X"11",X"11",X"FF",X"EE",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"11",X"BB",X"EE",X"CC",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"BB",X"22",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"66",X"44",X"77",X"77",X"44",X"66",X"00",
		X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"88",X"CC",X"66",X"33",X"66",X"CC",X"88",X"00",X"77",X"77",X"00",X"00",X"00",X"77",X"77",X"00",
		X"CC",X"FF",X"33",X"EE",X"33",X"FF",X"CC",X"00",X"77",X"77",X"00",X"11",X"00",X"77",X"77",X"00",
		X"11",X"33",X"66",X"CC",X"66",X"33",X"11",X"00",X"44",X"66",X"33",X"11",X"33",X"66",X"44",X"00",
		X"00",X"00",X"99",X"FF",X"FF",X"99",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"33",X"11",X"99",X"99",X"DD",X"77",X"33",X"00",X"66",X"77",X"55",X"44",X"44",X"44",X"66",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"FF",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"FF",X"77",X"03",X"03",X"03",X"03",X"03",X"03",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"22",X"11",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FB",X"66",X"44",X"88",X"99",X"00",X"00",X"00",X"00",X"11",X"22",X"CC",X"00",X"11",X"00",X"00",
		X"00",X"88",X"44",X"22",X"22",X"66",X"FB",X"FF",X"00",X"00",X"00",X"00",X"CC",X"33",X"00",X"0F",
		X"00",X"88",X"77",X"00",X"CC",X"00",X"00",X"00",X"FB",X"66",X"AA",X"99",X"44",X"44",X"00",X"00",
		X"00",X"00",X"44",X"88",X"00",X"FF",X"00",X"00",X"00",X"44",X"88",X"99",X"AA",X"66",X"FB",X"FF",
		X"FB",X"66",X"22",X"22",X"11",X"11",X"00",X"00",X"00",X"11",X"22",X"22",X"11",X"00",X"00",X"00",
		X"00",X"99",X"11",X"22",X"AA",X"66",X"FB",X"FF",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"0F",
		X"22",X"AA",X"44",X"00",X"00",X"CC",X"00",X"00",X"FB",X"66",X"AA",X"22",X"99",X"44",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"44",X"AA",X"11",X"00",X"00",X"00",X"00",X"99",X"22",X"66",X"FB",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",
		X"66",X"6E",X"E6",X"E6",X"6E",X"66",X"EE",X"EE",X"A5",X"D2",X"3C",X"03",X"92",X"69",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"44",X"88",X"00",X"00",
		X"22",X"33",X"44",X"88",X"11",X"66",X"88",X"0F",X"1D",X"2E",X"2E",X"0C",X"1D",X"2E",X"1D",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"0C",X"2E",X"2E",X"2E",X"1D",X"1D",X"0C",X"1D",
		X"00",X"00",X"04",X"22",X"FB",X"F0",X"9F",X"AA",X"00",X"00",X"46",X"11",X"30",X"17",X"10",X"04",
		X"00",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"26",X"9B",X"F0",X"F5",X"D5",X"04",X"00",X"00",X"76",X"33",X"97",X"70",X"11",X"02",X"00",X"00",
		X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"0C",X"1D",X"1D",X"2E",X"2E",X"2E",X"0C",
		X"0F",X"CC",X"33",X"00",X"CC",X"22",X"11",X"22",X"0F",X"1D",X"2E",X"1D",X"2E",X"2E",X"2E",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"88",X"77",X"0F",X"00",X"00",X"88",X"44",X"AA",X"11",X"66",X"0F",
		X"00",X"88",X"04",X"02",X"B3",X"E1",X"0F",X"4C",X"00",X"00",X"8C",X"31",X"00",X"11",X"71",X"18",
		X"00",X"00",X"00",X"00",X"00",X"48",X"F0",X"F0",X"00",X"00",X"00",X"C0",X"E1",X"D3",X"A7",X"5E",
		X"00",X"88",X"66",X"99",X"03",X"0F",X"0F",X"0F",X"2E",X"1D",X"0C",X"0C",X"1D",X"2E",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"03",X"44",X"88",X"00",X"00",X"0F",X"0F",X"0C",X"2E",X"1D",X"0C",X"3F",X"0C",
		X"F0",X"F8",X"C4",X"00",X"00",X"00",X"00",X"00",X"F9",X"F4",X"F2",X"F1",X"C0",X"00",X"00",X"00",
		X"C6",X"8F",X"D3",X"16",X"64",X"88",X"00",X"00",X"44",X"1F",X"30",X"61",X"88",X"00",X"11",X"00",
		X"0F",X"33",X"CC",X"00",X"00",X"00",X"00",X"00",X"0F",X"11",X"00",X"FF",X"44",X"88",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"B8",X"30",X"30",X"10",X"31",X"31",X"73",X"73",X"F7",X"C0",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"E7",X"F7",X"F7",X"73",X"73",X"31",X"31",X"31",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"31",X"31",X"31",X"73",X"73",X"F7",X"F7",X"E7",
		X"10",X"30",X"30",X"B8",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"C0",X"F7",X"73",X"73",X"31",X"31",
		X"08",X"08",X"08",X"08",X"F0",X"00",X"00",X"00",X"EF",X"EF",X"EF",X"EF",X"F0",X"00",X"80",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"EF",X"EF",X"EF",X"EF",X"0F",X"EF",X"EF",X"EF",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"EF",X"EF",X"EF",X"0F",X"EF",X"EF",X"EF",X"EF",
		X"00",X"00",X"00",X"F0",X"08",X"08",X"08",X"08",X"00",X"80",X"00",X"F0",X"EF",X"EF",X"EF",X"EF",
		X"10",X"10",X"10",X"10",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"FC",X"FE",X"76",X"10",X"10",X"00",X"E0",X"76",X"77",X"11",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"3C",X"00",X"00",X"3F",X"3F",X"3F",X"B7",X"87",X"87",X"80",X"00",
		X"00",X"00",X"00",X"30",X"C0",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"80",X"F0",X"0F",X"0F",X"3F",
		X"00",X"FF",X"00",X"00",X"11",X"EE",X"00",X"00",X"88",X"FF",X"44",X"44",X"22",X"11",X"00",X"00",
		X"00",X"00",X"EE",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"22",X"44",X"44",X"FF",X"88",
		X"44",X"44",X"44",X"CC",X"77",X"00",X"00",X"00",X"60",X"E8",X"60",X"71",X"E8",X"60",X"00",X"00",
		X"00",X"00",X"00",X"77",X"CC",X"44",X"44",X"44",X"00",X"00",X"60",X"E8",X"71",X"60",X"E8",X"60",
		X"00",X"1E",X"10",X"10",X"1E",X"10",X"08",X"07",X"08",X"0F",X"04",X"04",X"07",X"02",X"01",X"00",
		X"07",X"08",X"10",X"1E",X"10",X"10",X"1E",X"00",X"00",X"01",X"02",X"07",X"04",X"04",X"0F",X"08",
		X"78",X"3C",X"B4",X"96",X"D2",X"C3",X"E1",X"69",X"F0",X"B4",X"B4",X"1E",X"5A",X"4B",X"E1",X"E9",
		X"78",X"3C",X"B4",X"96",X"D2",X"C3",X"E1",X"69",X"F8",X"B4",X"B4",X"1E",X"5A",X"4B",X"E1",X"E1",
		X"FE",X"FC",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"F1",X"70",X"70",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FC",X"FE",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"F1",
		X"00",X"00",X"88",X"EE",X"33",X"00",X"00",X"00",X"E2",X"E2",X"73",X"E2",X"E2",X"22",X"22",X"00",
		X"00",X"00",X"00",X"33",X"EE",X"88",X"00",X"00",X"00",X"22",X"22",X"E2",X"E2",X"73",X"E2",X"E2",
		X"00",X"0F",X"00",X"0F",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",
		X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",X"00",X"30",X"3C",X"30",X"3C",X"30",X"3C",X"30",X"00",
		X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"30",X"3C",X"30",X"3C",X"30",X"3C",X"30",X"3C",
		X"E1",X"E1",X"E1",X"F0",X"F0",X"FF",X"F0",X"00",X"5E",X"5E",X"5E",X"DE",X"FE",X"FF",X"FE",X"00",
		X"F0",X"FF",X"F0",X"F0",X"E1",X"E1",X"E1",X"E1",X"FE",X"FF",X"FE",X"DE",X"5E",X"5E",X"5E",X"5E",
		X"FF",X"FF",X"F3",X"30",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"F3",X"FF",X"FF",X"EF",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"BF",X"BF",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"F0",X"FF",X"FF",X"BF",X"BF",X"0F",
		X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"FE",X"FE",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",
		X"93",X"93",X"93",X"93",X"93",X"93",X"F0",X"00",X"DD",X"88",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"F0",X"91",X"F7",X"F7",X"83",X"B3",X"80",X"00",X"30",X"00",X"00",X"00",X"88",X"DD",X"FF",
		X"00",X"0F",X"07",X"FF",X"BF",X"FF",X"F0",X"00",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"F0",X"00",
		X"00",X"F0",X"0F",X"B3",X"C0",X"60",X"30",X"07",X"00",X"F0",X"2C",X"3C",X"2C",X"2C",X"2C",X"EC",
		X"EC",X"EC",X"2C",X"2C",X"EC",X"2C",X"F0",X"00",X"B3",X"B3",X"80",X"80",X"91",X"83",X"F0",X"00",
		X"00",X"F0",X"EC",X"2C",X"EC",X"E0",X"2C",X"EC",X"00",X"F0",X"91",X"81",X"B3",X"90",X"83",X"91",
		X"FC",X"76",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"64",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"22",X"22",X"55",X"88",X"00",X"00",X"00",X"E6",X"EE",X"CC",X"88",X"77",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"44",X"00",X"00",X"00",X"00",X"20",X"71",X"71",X"F3",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"33",X"11",X"88",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"07",X"8F",X"07",X"00",X"00",X"00",X"00",X"00",X"88",X"33",X"CC",
		X"32",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"76",X"76",X"76",X"76",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"44",X"AA",X"33",X"11",X"00",X"00",X"00",X"CC",X"88",X"88",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"99",X"00",X"00",X"00",X"C4",X"E6",X"E6",X"E6",X"C4",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"0C",X"0C",X"0C",X"0C",X"F0",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"1F",X"0C",X"F0",X"8C",X"44",X"F0",X"00",X"00",X"04",X"00",X"F0",X"01",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"0C",X"F0",X"0E",X"00",X"00",X"00",X"F0",X"02",X"03",X"F0",X"07",
		X"80",X"70",X"00",X"80",X"70",X"00",X"00",X"00",X"70",X"20",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"80",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",
		X"1F",X"0E",X"F0",X"0C",X"00",X"F0",X"00",X"00",X"00",X"01",X"F0",X"13",X"11",X"F0",X"00",X"00",
		X"00",X"00",X"0C",X"F0",X"0C",X"0C",X"F0",X"0E",X"00",X"00",X"00",X"F0",X"01",X"03",X"F0",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"3C",X"2C",X"2C",X"0C",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"2C",X"2C",X"3C",
		X"78",X"70",X"70",X"30",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",
		X"13",X"0B",X"09",X"18",X"F0",X"00",X"00",X"00",X"6B",X"6B",X"73",X"71",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"36",X"17",X"13",X"00",X"00",X"00",X"00",X"70",X"60",X"43",X"6B",
		X"C8",X"C8",X"C8",X"C0",X"F0",X"00",X"00",X"00",X"F7",X"F7",X"F7",X"F3",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"F0",X"A0",X"F0",X"F3",
		X"1D",X"15",X"04",X"16",X"F0",X"00",X"00",X"00",X"6A",X"6A",X"73",X"71",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"3A",X"3B",X"19",X"00",X"00",X"00",X"00",X"70",X"61",X"40",X"6A",
		X"00",X"00",X"CC",X"3C",X"88",X"00",X"00",X"00",X"11",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"3C",X"CC",X"00",X"88",X"78",X"00",X"00",X"00",X"11",X"00",X"00",X"13",X"67",
		X"02",X"01",X"88",X"CF",X"88",X"00",X"00",X"00",X"11",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CF",X"88",X"01",X"02",X"8F",X"00",X"00",X"00",X"F0",X"00",X"00",X"11",X"F1",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"3C",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"7C",X"88",X"00",X"00",X"00",X"47",X"00",X"33",X"47",X"11",X"00",X"00",X"00",
		X"00",X"00",X"08",X"7C",X"88",X"00",X"00",X"78",X"00",X"00",X"01",X"13",X"11",X"00",X"11",X"EF",
		X"01",X"23",X"01",X"89",X"01",X"01",X"00",X"00",X"11",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"81",X"41",X"21",X"89",X"01",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"22",
		X"F0",X"5A",X"1E",X"8F",X"CE",X"3F",X"DD",X"00",X"CF",X"8F",X"FF",X"EF",X"DF",X"77",X"23",X"00",
		X"00",X"DF",X"6F",X"8E",X"FC",X"1E",X"B4",X"78",X"00",X"33",X"47",X"FF",X"FF",X"8F",X"EF",X"0F",
		X"23",X"01",X"45",X"01",X"89",X"01",X"00",X"00",X"44",X"11",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"81",X"41",X"21",X"01",X"01",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"E1",X"87",X"DE",X"9E",X"68",X"1F",X"00",X"CF",X"78",X"DF",X"FF",X"FF",X"47",X"33",X"00",
		X"00",X"C0",X"79",X"BC",X"1E",X"C3",X"68",X"1E",X"00",X"12",X"77",X"FF",X"FE",X"F8",X"DE",X"EF",
		X"F1",X"F0",X"F0",X"78",X"3C",X"3C",X"78",X"0F",X"78",X"78",X"78",X"69",X"4B",X"4B",X"69",X"0F",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"78",X"78",X"78",X"78",X"78",X"78",X"78",
		X"6F",X"EF",X"EF",X"6F",X"EF",X"E1",X"E1",X"0F",X"BF",X"FF",X"F1",X"F3",X"F3",X"F0",X"F0",X"0F",
		X"0F",X"E1",X"E1",X"EF",X"EF",X"6F",X"EF",X"EF",X"0F",X"F0",X"F0",X"F0",X"F7",X"F7",X"F1",X"FF",
		X"B5",X"5A",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"69",X"1E",X"3C",X"3C",X"78",X"78",X"78",X"0F",
		X"0F",X"E1",X"D2",X"D2",X"B4",X"87",X"78",X"F0",X"0F",X"78",X"78",X"78",X"78",X"5A",X"5A",X"69",
		X"67",X"EF",X"EF",X"67",X"EF",X"E1",X"E1",X"0F",X"BB",X"FF",X"F1",X"F3",X"F3",X"F0",X"F0",X"0F",
		X"0F",X"E1",X"E1",X"EF",X"EF",X"67",X"EF",X"EF",X"0F",X"78",X"F0",X"F0",X"F7",X"F7",X"F1",X"FF",
		X"00",X"01",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0D",X"06",X"00",X"10",X"10",X"00",X"0C",X"02",X"01",X"02",X"0C",X"00",X"00",X"00",
		X"04",X"03",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"08",X"04",X"02",X"01",X"01",X"01",X"02",X"20",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"00",X"79",X"71",X"79",X"51",X"91",X"11",X"00",X"80",
		X"EE",X"CF",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"11",X"11",X"11",X"11",X"FF",X"FF",X"FB",X"71",
		X"00",X"11",X"77",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"11",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"EE",X"EE",X"EE",X"CC",X"CC",X"C8",X"70",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",
		X"6E",X"6E",X"E6",X"6E",X"6E",X"66",X"EE",X"EE",X"69",X"1E",X"0B",X"01",X"2D",X"07",X"FF",X"FF",
		X"10",X"70",X"C8",X"CC",X"CC",X"EE",X"EE",X"66",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",
		X"00",X"0D",X"07",X"08",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"00",X"03",X"00",X"00",X"00",
		X"03",X"0C",X"00",X"09",X"06",X"10",X"10",X"00",X"00",X"0D",X"03",X"0C",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"04",X"02",X"01",X"01",X"01",X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C1",X"E3",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"C8",X"F8",X"F8",X"98",X"88",X"88",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"1D",X"1F",X"1F",X"1F",X"1D",X"11",X"11",X"11",
		X"88",X"88",X"98",X"F8",X"F8",X"C8",X"88",X"88",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"C0",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"10",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"10",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"A0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",
		X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"76",X"FE",X"FC",X"FC",X"EF",X"44",X"00",X"00",X"01",X"01",X"03",X"0F",X"03",X"01",X"01",X"00",
		X"30",X"28",X"2C",X"0F",X"0F",X"06",X"00",X"00",X"87",X"C3",X"C3",X"0D",X"1D",X"17",X"03",X"11",
		X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"80",X"80",X"33",X"33",X"33",X"91",X"91",X"81",
		X"F8",X"F8",X"F8",X"8F",X"0F",X"0F",X"00",X"00",X"F8",X"8F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",
		X"20",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"0F",X"0F",X"2C",X"28",X"00",X"00",X"01",X"01",X"03",X"0F",X"03",X"01",
		X"00",X"00",X"00",X"44",X"EF",X"E9",X"F8",X"FC",X"11",X"11",X"03",X"17",X"1D",X"C1",X"87",X"87",
		X"30",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"01",X"00",X"00",X"00",X"10",X"10",X"30",X"20",
		X"30",X"70",X"F0",X"F0",X"F0",X"D0",X"40",X"60",X"07",X"03",X"91",X"91",X"F3",X"F3",X"F3",X"40",
		X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"2C",X"00",X"00",X"01",X"01",X"03",X"0F",X"03",X"01",
		X"00",X"00",X"00",X"44",X"EF",X"E9",X"F8",X"FC",X"11",X"03",X"17",X"1D",X"59",X"C1",X"87",X"87",
		X"28",X"30",X"00",X"00",X"88",X"88",X"88",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"90",X"07",X"83",X"91",X"D1",X"F3",X"F3",X"71",X"20",
		X"00",X"80",X"C0",X"C0",X"1C",X"3C",X"08",X"08",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",
		X"76",X"47",X"03",X"01",X"30",X"ED",X"77",X"DD",X"E0",X"F0",X"78",X"78",X"80",X"C3",X"4B",X"0F",
		X"08",X"3C",X"1C",X"E0",X"C0",X"80",X"00",X"00",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"77",X"ED",X"30",X"01",X"03",X"47",X"76",X"00",X"4B",X"C3",X"80",X"38",X"78",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"00",X"33",X"77",X"66",X"7F",X"FF",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"66",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"33",X"66",X"77",X"66",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"66",X"77",X"66",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0D",X"05",X"07",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0F",X"05",X"05",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0F",X"04",X"0C",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"07",X"05",X"0D",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"07",X"05",X"0F",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0F",X"05",X"0F",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"CD",
		X"0F",X"00",X"0F",X"04",X"0C",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"0F",X"01",X"0F",X"00",X"0F",X"01",X"0F",X"00",X"00",X"11",X"00",X"00",X"22",X"11",X"11",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"7F",X"FF",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"CD",
		X"00",X"0F",X"01",X"0F",X"00",X"0F",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"00",X"00",X"00",
		X"7F",X"66",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"00",X"00",X"22",X"11",X"11",X"77",X"FF",X"77",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"09",X"0F",X"06",X"0E",X"0C",X"08",X"0E",X"07",X"0B",X"07",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"11",X"11",X"22",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"0B",X"07",X"0E",X"08",X"0C",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"22",X"11",X"11",X"77",X"FF",X"77",X"FF",X"77",
		X"00",X"01",X"07",X"0F",X"09",X"0F",X"09",X"0F",X"06",X"0E",X"08",X"0E",X"0B",X"0B",X"07",X"0F",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"22",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"0C",X"06",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"22",X"11",X"11",X"77",X"FF",X"77",X"FF",X"77",
		X"00",X"00",X"01",X"0F",X"09",X"0F",X"09",X"0F",X"00",X"06",X"0E",X"08",X"0E",X"07",X"07",X"0F",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"22",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"0E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"0E",X"00",X"00",X"22",X"11",X"11",X"77",X"FF",X"77",
		X"01",X"01",X"00",X"01",X"07",X"0F",X"09",X"0F",X"0C",X"0C",X"08",X"08",X"0E",X"0F",X"0F",X"03",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"11",X"11",X"22",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"00",X"01",X"01",X"00",X"0F",X"0F",X"0E",X"08",X"08",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"02",X"01",X"03",X"0F",X"0E",X"00",X"00",X"22",X"11",X"11",X"77",X"FF",X"77",
		X"0E",X"0F",X"07",X"01",X"07",X"0F",X"09",X"0F",X"00",X"00",X"08",X"08",X"0C",X"0F",X"0B",X"01",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"11",X"11",X"22",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"07",X"0F",X"0E",X"00",X"0B",X"0F",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"FF",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"32",X"76",X"77",X"00",X"00",X"00",X"00",X"FF",X"E6",X"44",X"EC",
		X"77",X"FF",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"76",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"E6",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"EE",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"32",X"76",X"77",X"32",X"10",X"00",X"00",X"FF",X"D5",X"64",X"CC",X"55",X"F7",
		X"FF",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"32",X"77",X"76",X"32",X"00",X"00",X"00",X"F7",X"55",X"CC",X"64",X"D5",X"FF",
		X"FF",X"77",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"FF",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"32",X"77",X"76",X"32",X"11",X"00",X"00",X"F7",X"55",X"EC",X"44",X"D5",X"FF",
		X"FF",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"EE",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"74",X"EC",X"FF",X"00",X"00",X"00",X"00",X"FF",X"DD",X"88",X"C8",
		X"EE",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EC",X"74",X"11",X"00",X"00",X"00",X"00",X"00",X"88",X"DD",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"FF",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"74",X"EC",X"FF",X"00",X"44",X"EE",X"44",X"FF",X"DD",X"88",X"98",
		X"EE",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EC",X"74",X"11",X"00",X"00",X"00",X"00",X"00",X"88",X"DD",X"FF",X"22",X"77",X"22",X"00",X"00",
		X"00",X"00",X"88",X"00",X"99",X"FF",X"77",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"32",X"76",X"77",X"00",X"11",X"33",X"11",X"FF",X"E6",X"44",X"CC",
		X"66",X"EE",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"76",X"32",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"E6",X"FF",X"88",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"AA",X"11",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"00",X"00",X"00",X"00",X"33",X"F9",X"D9",X"FF",
		X"11",X"AA",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D9",X"F9",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"74",X"DC",X"FF",X"00",X"00",X"00",X"00",X"CC",X"FF",X"99",X"B8",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DC",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"99",X"FF",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"E2",X"B3",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"77",X"77",X"00",X"44",X"EE",X"44",X"FF",X"BB",X"11",X"91",
		X"B3",X"E2",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"BB",X"FF",X"22",X"77",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"00",X"00",X"00",X"00",X"11",X"71",X"F1",X"F1",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"09",X"0F",X"06",X"0E",X"0C",X"08",X"0E",X"07",X"0B",X"07",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"73",X"55",X"88",X"88",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"0B",X"07",X"0E",X"08",X"0C",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"00",X"00",X"11",X"71",X"F1",X"F1",X"F1",X"73",
		X"00",X"01",X"07",X"0F",X"09",X"0F",X"09",X"0F",X"06",X"0E",X"08",X"0E",X"0B",X"0B",X"07",X"0F",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"0C",X"06",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"00",X"00",X"11",X"71",X"F1",X"F1",X"F1",X"73",
		X"00",X"00",X"01",X"0F",X"09",X"0F",X"09",X"0F",X"00",X"06",X"0E",X"08",X"0E",X"07",X"07",X"0F",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"55",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"0E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"0E",X"00",X"00",X"88",X"88",X"55",X"73",X"F1",X"F1",
		X"01",X"01",X"00",X"01",X"07",X"0F",X"09",X"0F",X"0C",X"0C",X"08",X"08",X"0E",X"0F",X"0F",X"03",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"71",X"11",X"00",X"00",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"00",X"01",X"01",X"00",X"0F",X"0F",X"0E",X"08",X"08",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"02",X"01",X"03",X"0F",X"0E",X"00",X"00",X"88",X"88",X"55",X"73",X"F1",X"F1",
		X"0E",X"0F",X"07",X"01",X"07",X"0F",X"09",X"0F",X"00",X"00",X"08",X"08",X"0C",X"0F",X"0B",X"01",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"71",X"11",X"00",X"00",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"07",X"0F",X"0E",X"00",X"0B",X"0F",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"70",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"CC",X"22",X"10",X"FC",X"30",X"00",X"00",X"00",X"00",X"2C",X"38",X"E0",X"E0",
		X"F0",X"30",X"60",X"60",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"10",X"66",X"88",X"00",X"00",X"00",X"00",X"00",X"38",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"33",X"44",X"00",X"33",X"44",
		X"00",X"00",X"00",X"00",X"8B",X"42",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"F0",X"90",X"90",
		X"C0",X"C0",X"60",X"60",X"30",X"10",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"00",X"00",X"00",
		X"42",X"8B",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"33",X"00",X"77",X"00",X"00",
		X"00",X"00",X"00",X"8B",X"42",X"F0",X"F0",X"42",X"00",X"00",X"00",X"80",X"F0",X"90",X"90",X"F0",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"30",X"30",X"20",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"60",X"70",X"F0",X"70",X"11",X"00",X"00",X"22",X"11",X"00",X"11",X"00",
		X"88",X"44",X"22",X"10",X"FC",X"30",X"10",X"EE",X"00",X"00",X"2C",X"38",X"E0",X"E0",X"38",X"2C",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"10",X"00",X"00",X"00",X"60",X"30",X"10",X"2C",X"38",
		X"60",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"11",X"00",X"00",X"00",X"00",
		X"30",X"FC",X"10",X"EE",X"00",X"00",X"00",X"00",X"E0",X"E0",X"38",X"2C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"44",X"22",X"11",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"16",X"94",X"F0",X"00",X"00",X"40",X"E0",X"40",X"60",X"F0",X"30",
		X"F0",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"33",X"44",X"00",X"00",X"00",X"00",
		X"F0",X"94",X"16",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"60",X"20",X"70",X"20",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"10",
		X"00",X"00",X"00",X"00",X"00",X"16",X"94",X"F0",X"00",X"00",X"10",X"30",X"10",X"30",X"F0",X"30",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"94",X"16",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"60",X"40",X"E0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"48",X"60",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"11",X"10",X"F3",X"00",X"00",X"00",X"00",X"00",X"ED",X"E1",X"F0",
		X"F0",X"60",X"48",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"10",X"00",X"77",X"00",X"00",X"00",X"00",X"F8",X"E1",X"ED",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"8B",X"42",X"F0",X"00",X"00",X"00",X"70",X"40",X"E0",X"F0",X"90",
		X"C0",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"42",X"8B",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"E0",X"40",X"70",X"00",X"00",X"00",
		X"00",X"00",X"88",X"44",X"22",X"2A",X"48",X"E0",X"00",X"00",X"00",X"20",X"30",X"30",X"10",X"10",
		X"00",X"00",X"10",X"00",X"00",X"80",X"F0",X"E0",X"00",X"80",X"C0",X"80",X"C0",X"E1",X"E0",X"70",
		X"F1",X"D1",X"D5",X"55",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"30",X"20",X"70",X"20",X"00",X"00",X"70",X"C1",X"43",X"00",X"00",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"00",X"00",X"00",X"10",X"10",X"F0",X"F0",X"F2",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"09",X"0F",X"06",X"0E",X"0C",X"08",X"0E",X"07",X"0B",X"07",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"10",X"10",X"00",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"0B",X"07",X"0E",X"08",X"0C",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"00",X"10",X"10",X"F0",X"F0",X"F2",X"F0",X"F0",
		X"00",X"01",X"07",X"0F",X"09",X"0F",X"09",X"0F",X"06",X"0E",X"08",X"0E",X"0B",X"0B",X"07",X"0F",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"0C",X"06",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"00",X"10",X"10",X"F0",X"F0",X"F2",X"F0",X"F0",
		X"00",X"00",X"01",X"0F",X"09",X"0F",X"09",X"0F",X"00",X"06",X"0E",X"08",X"0E",X"07",X"07",X"0F",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"0E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"0E",X"00",X"00",X"00",X"10",X"10",X"F0",X"F0",X"F2",
		X"01",X"01",X"00",X"01",X"07",X"0F",X"09",X"0F",X"0C",X"0C",X"08",X"08",X"0E",X"0F",X"0F",X"03",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"10",X"10",X"00",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"00",X"01",X"01",X"00",X"0F",X"0F",X"0E",X"08",X"08",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"02",X"01",X"03",X"0F",X"0E",X"00",X"00",X"00",X"10",X"10",X"F0",X"F0",X"F2",
		X"0E",X"0F",X"07",X"01",X"07",X"0F",X"09",X"0F",X"00",X"00",X"08",X"08",X"0C",X"0F",X"0B",X"01",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"10",X"10",X"00",X"00",X"00",X"00",
		X"09",X"0F",X"07",X"01",X"07",X"0F",X"0E",X"00",X"0B",X"0F",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"08",X"0C",X"15",X"B7",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"30",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F7",X"80",X"00",X"33",X"33",X"22",X"03",X"07",X"0C",X"18",
		X"04",X"37",X"15",X"0C",X"08",X"00",X"CC",X"88",X"00",X"30",X"20",X"30",X"00",X"00",X"00",X"00",
		X"00",X"80",X"F7",X"80",X"00",X"00",X"00",X"00",X"08",X"68",X"0C",X"07",X"03",X"22",X"33",X"11",
		X"00",X"66",X"CC",X"00",X"08",X"0C",X"04",X"95",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"62",X"D1",X"00",X"00",X"00",X"11",X"33",X"03",X"07",X"0E",X"1C",
		X"37",X"04",X"37",X"1D",X"08",X"00",X"88",X"00",X"30",X"20",X"30",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C4",X"B3",X"00",X"00",X"00",X"00",X"00",X"0C",X"3C",X"0E",X"07",X"03",X"22",X"77",X"66",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"2E",X"2E",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"30",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F7",X"80",X"33",X"66",X"66",X"22",X"03",X"07",X"0C",X"1C",
		X"0C",X"2E",X"2E",X"0C",X"08",X"00",X"00",X"00",X"00",X"30",X"20",X"30",X"00",X"00",X"00",X"00",
		X"00",X"80",X"F7",X"80",X"00",X"00",X"00",X"00",X"0C",X"2C",X"0C",X"07",X"03",X"22",X"77",X"66",
		X"00",X"88",X"CC",X"00",X"08",X"1D",X"3F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B3",X"C4",X"00",X"11",X"33",X"22",X"03",X"07",X"0C",X"18",
		X"3F",X"1D",X"0C",X"0C",X"08",X"00",X"00",X"00",X"30",X"00",X"10",X"10",X"10",X"00",X"00",X"00",
		X"80",X"00",X"D1",X"62",X"C0",X"00",X"00",X"11",X"08",X"68",X"0C",X"07",X"03",X"22",X"EE",X"CC",
		X"00",X"88",X"CC",X"00",X"08",X"1D",X"3F",X"84",X"00",X"00",X"00",X"00",X"00",X"70",X"50",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"33",X"22",X"22",X"03",X"07",X"0F",X"18",
		X"04",X"04",X"3F",X"1D",X"08",X"00",X"44",X"CC",X"00",X"70",X"50",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"68",X"0F",X"07",X"03",X"22",X"33",X"11",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"15",X"B7",X"00",X"00",X"00",X"00",X"70",X"50",X"70",X"00",
		X"00",X"22",X"33",X"00",X"00",X"CC",X"33",X"00",X"44",X"66",X"FF",X"22",X"03",X"07",X"0C",X"18",
		X"04",X"37",X"15",X"0C",X"08",X"00",X"00",X"CC",X"00",X"00",X"30",X"20",X"30",X"00",X"00",X"00",
		X"00",X"00",X"B3",X"C4",X"80",X"00",X"00",X"00",X"08",X"68",X"0C",X"07",X"03",X"EE",X"33",X"FF",
		X"88",X"00",X"00",X"00",X"08",X"0C",X"15",X"B7",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",
		X"11",X"11",X"00",X"00",X"00",X"00",X"B3",X"C4",X"11",X"FF",X"22",X"22",X"03",X"06",X"0C",X"18",
		X"04",X"37",X"15",X"0C",X"08",X"00",X"00",X"00",X"30",X"20",X"30",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C4",X"B3",X"00",X"00",X"33",X"11",X"77",X"08",X"68",X"0C",X"06",X"03",X"22",X"22",X"EE",
		X"00",X"00",X"00",X"00",X"08",X"2E",X"2E",X"0C",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"33",X"00",X"11",X"00",X"00",X"C0",X"73",X"C0",X"CC",X"44",X"EE",X"22",X"03",X"07",X"0D",X"68",
		X"04",X"0C",X"2E",X"2E",X"08",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"73",X"C0",X"00",X"00",X"33",X"77",X"08",X"38",X"0D",X"07",X"03",X"22",X"EE",X"88",
		X"00",X"00",X"CC",X"00",X"00",X"08",X"19",X"6E",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"30",
		X"00",X"00",X"00",X"00",X"00",X"80",X"E7",X"81",X"00",X"33",X"33",X"66",X"07",X"0F",X"08",X"C0",
		X"08",X"6E",X"19",X"08",X"00",X"00",X"CC",X"00",X"00",X"30",X"20",X"30",X"00",X"00",X"00",X"00",
		X"01",X"81",X"E7",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"08",X"0F",X"07",X"66",X"33",X"11",
		X"00",X"00",X"E0",X"A0",X"E0",X"44",X"88",X"00",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"00",
		X"CC",X"77",X"33",X"22",X"03",X"02",X"8E",X"14",X"88",X"88",X"00",X"00",X"0C",X"06",X"06",X"97",
		X"00",X"00",X"CC",X"44",X"44",X"70",X"50",X"70",X"00",X"33",X"22",X"00",X"00",X"00",X"00",X"00",
		X"04",X"9C",X"16",X"03",X"00",X"00",X"11",X"33",X"06",X"06",X"17",X"0C",X"88",X"88",X"FF",X"88",
		X"70",X"50",X"50",X"D0",X"00",X"F0",X"10",X"F0",X"08",X"0F",X"0F",X"08",X"08",X"00",X"00",X"0F",
		X"00",X"0E",X"0E",X"02",X"02",X"0E",X"00",X"0C",X"54",X"54",X"54",X"54",X"CC",X"DC",X"DC",X"DC",
		X"00",X"C0",X"40",X"F0",X"00",X"50",X"50",X"F0",X"09",X"09",X"0D",X"03",X"08",X"0F",X"0F",X"08",
		X"19",X"19",X"19",X"1D",X"33",X"3B",X"3B",X"33",X"CC",X"DC",X"DC",X"DC",X"CC",X"DC",X"DC",X"DC",
		X"EF",X"13",X"15",X"19",X"99",X"99",X"99",X"99",X"F7",X"C8",X"A8",X"98",X"99",X"99",X"99",X"99",
		X"FF",X"00",X"00",X"FF",X"80",X"40",X"31",X"32",X"FF",X"00",X"00",X"FF",X"01",X"02",X"8C",X"4C",
		X"99",X"99",X"99",X"99",X"91",X"51",X"31",X"FE",X"99",X"99",X"99",X"99",X"89",X"8A",X"8C",X"7F",
		X"23",X"13",X"04",X"08",X"FF",X"00",X"00",X"FF",X"C4",X"C8",X"20",X"10",X"FF",X"00",X"00",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
