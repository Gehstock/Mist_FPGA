library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dderby_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dderby_sp_bits_3 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"79",X"99",X"99",X"00",X"97",X"99",X"22",X"00",X"33",X"26",X"76",
		X"00",X"E9",X"22",X"69",X"00",X"E9",X"99",X"62",X"00",X"E9",X"27",X"66",X"00",X"99",X"29",X"66",
		X"00",X"99",X"29",X"66",X"00",X"99",X"29",X"66",X"00",X"77",X"29",X"66",X"00",X"77",X"99",X"66",
		X"00",X"77",X"99",X"66",X"00",X"77",X"29",X"66",X"00",X"99",X"29",X"66",X"00",X"99",X"29",X"66",
		X"00",X"39",X"29",X"66",X"00",X"E9",X"27",X"66",X"00",X"E9",X"99",X"62",X"00",X"E9",X"22",X"69",
		X"00",X"33",X"26",X"76",X"00",X"97",X"99",X"22",X"00",X"79",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"97",X"99",X"99",X"00",X"22",X"77",X"99",X"00",X"92",X"66",X"69",X"00",
		X"26",X"99",X"99",X"00",X"69",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",
		X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"62",X"99",X"00",
		X"29",X"26",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",
		X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"69",X"22",X"99",X"00",X"26",X"99",X"99",X"00",
		X"92",X"66",X"69",X"00",X"22",X"77",X"99",X"00",X"97",X"99",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"26",X"00",
		X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"79",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"72",X"99",X"00",X"00",X"77",X"27",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"09",X"69",X"97",X"00",X"09",X"29",X"96",X"00",X"E3",X"29",X"76",X"00",X"E3",X"22",X"66",
		X"00",X"33",X"79",X"66",X"00",X"96",X"29",X"66",X"00",X"92",X"29",X"66",X"00",X"07",X"99",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"96",X"00",X"00",X"00",X"99",X"79",X"00",X"00",X"99",X"99",X"00",X"00",X"62",X"29",X"00",X"00",
		X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"62",X"99",X"00",X"00",X"62",X"92",X"70",X"00",
		X"00",X"00",X"79",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"72",X"66",X"00",X"00",X"97",X"22",
		X"00",X"00",X"99",X"97",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"67",X"92",X"66",X"00",X"29",X"92",X"09",X"00",X"29",X"22",X"09",X"00",X"79",X"22",X"09",X"00",
		X"99",X"62",X"90",X"00",X"99",X"66",X"90",X"00",X"99",X"27",X"90",X"00",X"99",X"62",X"00",X"00",
		X"99",X"22",X"00",X"00",X"79",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"72",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"62",X"00",X"00",
		X"00",X"76",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",
		X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"29",X"00",X"00",X"77",X"29",X"00",X"00",X"22",X"62",
		X"00",X"00",X"62",X"26",X"00",X"00",X"26",X"92",X"00",X"00",X"26",X"99",X"00",X"0E",X"22",X"92",
		X"00",X"0E",X"22",X"22",X"00",X"07",X"72",X"92",X"00",X"00",X"72",X"29",X"00",X"09",X"27",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"79",X"96",X"00",X"00",X"79",X"66",
		X"00",X"00",X"29",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"72",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"79",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"92",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"07",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"70",X"00",X"00",X"62",X"79",X"00",X"00",X"29",X"77",X"00",X"00",X"99",X"77",X"00",X"00",
		X"99",X"27",X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"92",X"97",X"00",X"00",X"92",X"97",X"00",X"00",
		X"29",X"70",X"00",X"00",X"62",X"00",X"00",X"00",X"22",X"09",X"00",X"00",X"76",X"99",X"00",X"00",
		X"77",X"90",X"00",X"00",X"77",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"70",X"00",X"00",X"09",X"27",X"00",X"00",X"E9",X"27",
		X"00",X"00",X"E0",X"27",X"00",X"00",X"30",X"22",X"00",X"00",X"37",X"62",X"00",X"00",X"62",X"22",
		X"00",X"00",X"62",X"92",X"00",X"00",X"26",X"92",X"00",X"00",X"26",X"99",X"00",X"00",X"22",X"97",
		X"00",X"00",X"22",X"72",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"62",X"00",X"00",X"92",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"09",X"66",
		X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"72",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",
		X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"72",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"29",X"79",X"00",X"00",X"92",X"29",X"00",X"00",X"66",X"69",X"00",X"00",X"26",X"67",X"00",X"00",
		X"26",X"62",X"00",X"00",X"26",X"26",X"00",X"00",X"22",X"06",X"00",X"00",X"22",X"99",X"00",X"00",
		X"77",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"90",X"EE",X"00",
		X"00",X"99",X"99",X"00",X"00",X"07",X"09",X"00",X"00",X"97",X"92",X"00",X"00",X"22",X"92",X"00",
		X"00",X"27",X"92",X"00",X"00",X"27",X"92",X"00",X"00",X"27",X"92",X"00",X"00",X"27",X"92",X"00",
		X"00",X"27",X"92",X"00",X"00",X"22",X"92",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"99",X"00",
		X"00",X"77",X"22",X"00",X"00",X"62",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",X"00",
		X"00",X"99",X"99",X"00",X"00",X"77",X"79",X"00",X"00",X"66",X"27",X"00",X"00",X"66",X"22",X"00",
		X"00",X"66",X"27",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",
		X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",
		X"00",X"66",X"29",X"00",X"00",X"22",X"62",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"77",X"72",X"00",
		X"00",X"22",X"22",X"00",X"00",X"92",X"99",X"00",X"00",X"27",X"29",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"77",X"77",X"00",X"00",X"90",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",
		X"00",X"00",X"AB",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"AD",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"99",X"90",X"00",X"00",X"91",X"90",X"00",X"00",X"11",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"41",X"00",X"00",X"09",X"11",X"00",X"00",
		X"91",X"10",X"00",X"00",X"11",X"09",X"00",X"00",X"14",X"99",X"00",X"00",X"11",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"90",X"90",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"9A",X"90",X"00",X"00",X"AD",X"90",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"AD",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"99",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"AA",X"90",X"00",
		X"09",X"AD",X"00",X"00",X"09",X"DA",X"00",X"00",X"9D",X"AD",X"00",X"00",X"9D",X"DA",X"00",X"00",
		X"9D",X"DD",X"00",X"00",X"9D",X"DD",X"00",X"00",X"9D",X"DD",X"00",X"00",X"09",X"DD",X"00",X"00",
		X"F9",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"97",X"99",X"99",X"00",X"22",X"77",X"99",X"00",X"92",X"99",X"69",X"00",
		X"26",X"22",X"99",X"00",X"69",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",
		X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"62",X"99",X"00",
		X"29",X"26",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"29",X"99",X"00",
		X"29",X"29",X"99",X"00",X"29",X"99",X"99",X"00",X"69",X"99",X"99",X"00",X"26",X"99",X"99",X"00",
		X"92",X"69",X"99",X"00",X"22",X"76",X"99",X"00",X"97",X"99",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"96",X"00",X"00",X"00",X"99",X"79",X"00",X"00",X"99",X"99",X"00",X"00",X"62",X"29",X"00",X"00",
		X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"62",X"99",X"00",X"00",X"62",X"92",X"70",X"00",
		X"67",X"92",X"66",X"00",X"29",X"92",X"09",X"00",X"29",X"22",X"09",X"00",X"79",X"22",X"09",X"00",
		X"99",X"62",X"90",X"00",X"99",X"66",X"90",X"00",X"99",X"29",X"00",X"00",X"99",X"69",X"00",X"00",
		X"99",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"72",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"69",X"00",X"00",
		X"00",X"76",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"70",X"00",X"00",X"62",X"79",X"00",X"00",X"29",X"77",X"00",X"00",X"99",X"77",X"00",X"00",
		X"99",X"27",X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"97",X"00",X"00",
		X"29",X"70",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"09",X"00",X"00",X"69",X"99",X"00",X"00",
		X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"29",X"79",X"00",X"00",X"92",X"29",X"00",X"00",X"66",X"69",X"00",X"00",X"99",X"62",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"06",X"00",X"00",X"99",X"99",X"00",X"00",
		X"77",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",
		X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",
		X"00",X"66",X"29",X"00",X"00",X"22",X"62",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"77",X"72",X"00",
		X"00",X"22",X"22",X"00",X"00",X"92",X"99",X"00",X"00",X"27",X"29",X"00",X"00",X"22",X"22",X"00",
		X"00",X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",
		X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"77",X"77",X"00",X"00",X"90",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"79",X"99",X"99",X"00",X"9E",X"99",X"22",X"00",X"9E",X"99",X"76",
		X"00",X"9E",X"22",X"69",X"00",X"99",X"29",X"62",X"00",X"09",X"92",X"66",X"00",X"09",X"92",X"66",
		X"00",X"99",X"92",X"66",X"00",X"99",X"D2",X"66",X"00",X"99",X"D2",X"66",X"00",X"99",X"92",X"66",
		X"00",X"09",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"D2",X"66",X"00",X"09",X"D2",X"66",
		X"00",X"99",X"92",X"66",X"00",X"99",X"99",X"66",X"00",X"E9",X"29",X"62",X"00",X"E9",X"22",X"69",
		X"00",X"E3",X"26",X"76",X"00",X"97",X"99",X"22",X"00",X"79",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E2",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"62",X"00",X"00",X"00",X"26",X"79",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"27",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"99",
		X"00",X"00",X"9D",X"97",X"00",X"09",X"DD",X"96",X"00",X"EE",X"D9",X"76",X"00",X"EE",X"DD",X"66",
		X"00",X"EE",X"99",X"66",X"00",X"93",X"99",X"66",X"00",X"92",X"99",X"66",X"00",X"07",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"9D",X"29",
		X"00",X"00",X"9D",X"26",X"00",X"00",X"DD",X"22",X"00",X"00",X"D9",X"29",X"00",X"0E",X"DD",X"92",
		X"00",X"0E",X"DD",X"22",X"00",X"0E",X"DD",X"92",X"00",X"00",X"9D",X"29",X"00",X"09",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"96",X"00",X"00",X"79",X"66",
		X"00",X"00",X"29",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"72",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"72",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"70",X"00",X"00",X"09",X"97",X"00",X"00",X"99",X"DD",
		X"00",X"00",X"E0",X"DD",X"00",X"00",X"E0",X"9D",X"00",X"00",X"33",X"DD",X"00",X"00",X"32",X"99",
		X"00",X"00",X"62",X"DD",X"00",X"00",X"26",X"22",X"00",X"00",X"26",X"29",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"62",X"00",X"00",X"92",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"07",X"09",X"00",X"00",X"97",X"99",X"00",X"00",X"DD",X"99",X"00",
		X"00",X"9D",X"92",X"00",X"00",X"9D",X"26",X"00",X"00",X"9D",X"22",X"00",X"00",X"9D",X"62",X"00",
		X"00",X"9D",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"22",X"00",
		X"00",X"77",X"22",X"00",X"00",X"62",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",X"00",
		X"00",X"99",X"99",X"00",X"00",X"77",X"79",X"00",X"00",X"66",X"27",X"00",X"00",X"66",X"22",X"00",
		X"00",X"66",X"27",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"79",X"00",X"99",X"00",X"9E",X"99",X"22",X"00",X"9E",X"99",X"76",
		X"00",X"99",X"22",X"69",X"00",X"99",X"29",X"62",X"00",X"09",X"92",X"66",X"00",X"09",X"92",X"66",
		X"00",X"99",X"92",X"66",X"00",X"99",X"D2",X"66",X"00",X"99",X"D2",X"66",X"00",X"99",X"92",X"66",
		X"00",X"09",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"D2",X"66",X"00",X"09",X"D2",X"66",
		X"00",X"99",X"92",X"66",X"00",X"9E",X"99",X"66",X"00",X"EE",X"29",X"62",X"00",X"EE",X"22",X"69",
		X"00",X"E3",X"26",X"76",X"00",X"93",X"99",X"22",X"00",X"79",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"96",X"00",X"00",X"00",X"99",X"70",X"00",X"00",X"99",X"99",X"00",X"00",X"62",X"29",X"00",X"00",
		X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"62",X"99",X"00",X"00",X"62",X"92",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E3",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"62",X"00",X"00",X"00",X"26",X"79",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"27",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"99",
		X"00",X"00",X"9D",X"97",X"00",X"0E",X"DD",X"96",X"00",X"EE",X"D9",X"76",X"00",X"EE",X"DD",X"66",
		X"00",X"EE",X"99",X"66",X"00",X"E3",X"99",X"66",X"00",X"93",X"99",X"66",X"00",X"07",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"79",X"99",X"00",X"00",X"9D",X"29",
		X"00",X"00",X"9D",X"26",X"00",X"00",X"DD",X"22",X"00",X"00",X"D9",X"29",X"00",X"00",X"DD",X"92",
		X"00",X"07",X"DD",X"22",X"00",X"02",X"DD",X"92",X"00",X"00",X"9D",X"29",X"00",X"09",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"96",X"00",X"00",X"79",X"66",
		X"00",X"00",X"29",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"72",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"72",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"70",X"00",X"00",X"09",X"97",X"00",X"00",X"99",X"DD",
		X"00",X"00",X"90",X"DD",X"00",X"00",X"30",X"9D",X"00",X"00",X"77",X"DD",X"00",X"00",X"62",X"99",
		X"00",X"00",X"62",X"DD",X"00",X"00",X"26",X"22",X"00",X"00",X"26",X"29",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"62",X"00",X"00",X"92",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"66",
		X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"07",X"09",X"00",X"00",X"97",X"99",X"00",X"00",X"DD",X"99",X"00",
		X"00",X"9D",X"92",X"00",X"00",X"9D",X"26",X"00",X"00",X"9D",X"22",X"00",X"09",X"9D",X"62",X"00",
		X"09",X"9D",X"22",X"00",X"09",X"92",X"22",X"00",X"09",X"22",X"99",X"00",X"09",X"99",X"22",X"00",
		X"09",X"77",X"22",X"00",X"09",X"62",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",X"00",
		X"00",X"99",X"99",X"00",X"00",X"77",X"79",X"00",X"00",X"66",X"27",X"00",X"00",X"66",X"22",X"00",
		X"00",X"66",X"27",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"97",X"99",X"99",X"00",X"22",X"77",X"99",X"00",X"92",X"07",X"99",X"00",
		X"26",X"99",X"99",X"00",X"69",X"92",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",
		X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"26",X"99",X"00",X"29",X"62",X"99",X"00",
		X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",X"29",X"22",X"99",X"00",
		X"29",X"29",X"99",X"00",X"29",X"29",X"99",X"00",X"69",X"99",X"99",X"00",X"26",X"99",X"99",X"00",
		X"92",X"69",X"99",X"00",X"22",X"76",X"99",X"00",X"97",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"67",X"92",X"66",X"00",X"29",X"92",X"09",X"00",X"29",X"22",X"09",X"00",X"79",X"22",X"09",X"00",
		X"99",X"62",X"90",X"00",X"99",X"62",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"79",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"72",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",
		X"00",X"76",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"72",X"66",X"00",X"00",X"97",X"22",
		X"00",X"00",X"99",X"97",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"70",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"26",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"97",X"00",X"00",X"29",X"70",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"09",X"00",X"00",X"69",X"99",X"00",X"00",X"76",X"00",X"00",X"00",
		X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"29",X"79",X"00",X"00",X"92",X"29",X"00",X"00",X"66",X"69",X"00",X"00",X"22",X"60",X"00",X"00",
		X"29",X"22",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",
		X"77",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",
		X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",
		X"00",X"66",X"29",X"00",X"00",X"22",X"62",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"77",X"72",X"00",
		X"00",X"22",X"22",X"00",X"00",X"92",X"99",X"00",X"00",X"27",X"29",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"77",X"77",X"00",X"00",X"90",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"11",X"09",X"00",
		X"00",X"91",X"09",X"00",X"00",X"91",X"91",X"00",X"01",X"01",X"11",X"00",X"00",X"01",X"02",X"00",
		X"00",X"01",X"12",X"00",X"00",X"10",X"11",X"00",X"00",X"11",X"22",X"00",X"09",X"10",X"00",X"00",
		X"09",X"00",X"00",X"11",X"00",X"90",X"00",X"11",X"00",X"90",X"09",X"10",X"00",X"90",X"00",X"00",
		X"00",X"91",X"20",X"09",X"00",X"10",X"00",X"19",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",
		X"00",X"10",X"11",X"00",X"00",X"10",X"11",X"00",X"10",X"11",X"10",X"00",X"01",X"11",X"11",X"00",
		X"01",X"11",X"22",X"11",X"99",X"99",X"21",X"11",X"00",X"00",X"11",X"10",X"09",X"00",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"99",X"11",X"00",X"20",X"90",
		X"11",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"99",X"10",X"22",X"00",X"99",X"12",X"22",X"00",
		X"01",X"12",X"11",X"00",X"11",X"10",X"11",X"00",X"01",X"21",X"10",X"00",X"01",X"00",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"90",X"00",X"99",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"21",X"10",X"11",X"00",X"01",X"01",X"11",X"00",X"11",X"09",X"11",X"00",X"01",X"11",X"11",
		X"00",X"19",X"10",X"20",X"00",X"10",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"01",X"91",X"00",
		X"00",X"00",X"09",X"00",X"09",X"01",X"99",X"99",X"19",X"01",X"99",X"99",X"11",X"01",X"00",X"99",
		X"11",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"11",X"00",X"99",X"00",
		X"11",X"10",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"11",X"00",X"00",X"91",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"21",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"01",X"00",X"19",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"11",X"00",X"01",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"09",X"00",X"11",X"00",X"99",X"00",X"90",X"09",X"10",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"10",X"00",X"99",X"09",X"10",X"01",X"99",X"09",X"00",X"10",
		X"09",X"99",X"11",X"10",X"99",X"99",X"00",X"11",X"90",X"90",X"00",X"90",X"99",X"99",X"11",X"90",
		X"90",X"90",X"99",X"99",X"00",X"90",X"19",X"99",X"00",X"90",X"10",X"90",X"00",X"91",X"90",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"90",X"11",X"00",X"00",X"90",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"00",X"09",X"00",
		X"01",X"10",X"91",X"00",X"00",X"01",X"91",X"00",X"01",X"11",X"00",X"00",X"00",X"11",X"20",X"00",
		X"99",X"11",X"00",X"00",X"99",X"01",X"00",X"00",X"90",X"11",X"92",X"10",X"99",X"11",X"99",X"10",
		X"00",X"11",X"91",X"11",X"00",X"10",X"99",X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",
		X"00",X"12",X"09",X"00",X"01",X"01",X"09",X"10",X"00",X"00",X"09",X"10",X"00",X"11",X"99",X"00",
		X"11",X"00",X"99",X"09",X"10",X"99",X"99",X"19",X"00",X"99",X"99",X"01",X"09",X"99",X"00",X"90",
		X"00",X"99",X"99",X"99",X"00",X"99",X"00",X"90",X"00",X"90",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"01",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"10",X"00",X"00",
		X"00",X"01",X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"10",X"11",X"00",X"00",X"02",X"10",X"00",
		X"00",X"10",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"10",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"10",X"19",X"09",X"00",X"11",X"11",X"00",X"09",X"99",
		X"11",X"00",X"09",X"99",X"01",X"11",X"09",X"00",X"90",X"01",X"10",X"00",X"91",X"00",X"10",X"00",
		X"91",X"00",X"10",X"00",X"91",X"99",X"01",X"00",X"19",X"99",X"10",X"00",X"01",X"09",X"11",X"00",
		X"00",X"99",X"01",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"90",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"19",X"00",X"00",
		X"11",X"90",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"01",X"04",X"90",
		X"00",X"14",X"11",X"90",X"00",X"41",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"10",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"11",X"11",X"99",
		X"00",X"11",X"11",X"00",X"01",X"11",X"00",X"00",X"19",X"11",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"12",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"12",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"12",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"12",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"12",X"10",X"00",X"00",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"F9",X"9F",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"F9",X"00",X"00",X"F0",X"F9",X"00",X"00",X"F0",X"99",X"F0",X"00",X"9F",X"9F",X"90",
		X"00",X"90",X"9F",X"F0",X"00",X"F0",X"09",X"FF",X"00",X"00",X"90",X"09",X"00",X"F0",X"90",X"0F",
		X"00",X"FF",X"F9",X"F0",X"00",X"9F",X"F0",X"90",X"00",X"9F",X"FF",X"09",X"00",X"90",X"99",X"99",
		X"0F",X"9F",X"09",X"90",X"09",X"FF",X"FF",X"90",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"9F",X"00",X"00",X"9F",X"0F",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"0F",X"9F",X"00",X"00",
		X"9F",X"F0",X"00",X"00",X"F0",X"FF",X"00",X"00",X"FF",X"F9",X"F0",X"00",X"9F",X"99",X"90",X"00",
		X"09",X"99",X"FF",X"00",X"09",X"0F",X"09",X"00",X"09",X"F0",X"F0",X"00",X"00",X"99",X"09",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"90",X"00",X"90",X"09",X"90",X"00",X"F9",X"9F",X"00",X"00",
		X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"FF",X"00",X"00",X"F9",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"9F",X"00",X"0F",X"00",X"9F",X"00",X"09",X"F0",X"0F",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"CA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",
		X"00",X"9A",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"AA",X"D9",X"00",X"00",X"AA",X"99",X"00",X"00",X"A9",X"90",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"93",X"99",X"99",X"00",X"EE",X"99",X"22",X"00",X"EE",X"22",X"99",
		X"00",X"EE",X"66",X"99",X"00",X"EE",X"22",X"29",X"00",X"EE",X"22",X"92",X"00",X"99",X"22",X"96",
		X"00",X"99",X"22",X"96",X"00",X"92",X"77",X"96",X"00",X"92",X"66",X"96",X"00",X"22",X"22",X"96",
		X"00",X"22",X"22",X"96",X"00",X"92",X"66",X"96",X"00",X"92",X"77",X"96",X"00",X"99",X"22",X"96",
		X"00",X"99",X"22",X"96",X"00",X"EE",X"22",X"92",X"00",X"EE",X"22",X"29",X"00",X"EE",X"66",X"99",
		X"00",X"EE",X"22",X"99",X"00",X"EE",X"99",X"22",X"00",X"37",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"22",X"99",X"90",X"00",X"99",X"77",X"90",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"92",X"77",X"99",X"00",X"29",X"72",X"99",X"00",
		X"69",X"72",X"99",X"00",X"69",X"72",X"99",X"00",X"69",X"72",X"99",X"00",X"69",X"72",X"99",X"00",
		X"69",X"72",X"99",X"00",X"69",X"72",X"99",X"00",X"69",X"72",X"99",X"00",X"69",X"72",X"99",X"00",
		X"29",X"72",X"99",X"00",X"92",X"77",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"77",X"90",X"00",X"22",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",
		X"00",X"09",X"62",X"90",X"00",X"99",X"26",X"90",X"00",X"99",X"26",X"99",X"00",X"99",X"22",X"29",
		X"00",X"99",X"72",X"22",X"00",X"99",X"77",X"99",X"00",X"99",X"62",X"29",X"00",X"99",X"22",X"92",
		X"00",X"99",X"22",X"92",X"00",X"99",X"22",X"99",X"00",X"E3",X"22",X"99",X"00",X"E3",X"22",X"92",
		X"00",X"E9",X"97",X"96",X"00",X"E9",X"27",X"96",X"00",X"92",X"22",X"26",X"00",X"92",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",
		X"67",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"00",
		X"00",X"99",X"62",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"96",
		X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"29",X"00",X"00",X"69",X"29",X"00",X"00",X"69",X"29",X"09",X"00",X"69",X"92",X"09",X"00",
		X"99",X"92",X"99",X"00",X"99",X"92",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"29",X"22",X"99",X"00",X"29",X"22",X"90",X"00",X"22",X"22",X"90",X"00",X"22",X"29",X"00",X"00",
		X"77",X"29",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"90",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",
		X"00",X"09",X"22",X"22",X"00",X"99",X"22",X"66",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"22",
		X"00",X"99",X"22",X"99",X"00",X"9E",X"76",X"92",X"00",X"9E",X"77",X"29",X"00",X"EE",X"27",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"99",
		X"00",X"00",X"62",X"96",X"00",X"00",X"22",X"96",X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"29",X"00",X"00",X"69",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"26",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"90",X"00",
		X"22",X"29",X"90",X"00",X"29",X"96",X"90",X"00",X"90",X"96",X"00",X"00",X"29",X"69",X"00",X"00",
		X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"09",X"00",X"00",X"97",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"EE",
		X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",
		X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"72",X"00",X"00",X"27",X"72",
		X"00",X"00",X"27",X"72",X"00",X"00",X"22",X"27",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"62",X"97",X"00",X"00",X"26",X"62",X"00",X"00",X"26",X"69",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"09",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"97",X"90",X"00",X"00",
		X"22",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"79",X"00",X"00",X"22",X"70",X"00",X"00",
		X"22",X"70",X"00",X"00",X"22",X"90",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"09",X"00",X"00",
		X"99",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"77",X"99",X"00",X"00",X"90",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"93",X"00",
		X"00",X"97",X"EE",X"00",X"00",X"22",X"3E",X"00",X"00",X"76",X"33",X"00",X"00",X"76",X"22",X"00",
		X"00",X"76",X"22",X"00",X"00",X"26",X"22",X"00",X"00",X"27",X"22",X"00",X"00",X"27",X"22",X"00",
		X"00",X"27",X"22",X"00",X"00",X"27",X"22",X"00",X"00",X"27",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"92",X"00",X"00",X"29",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"66",X"99",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"26",X"69",X"00",X"00",X"26",X"69",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"72",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"27",X"00",
		X"00",X"29",X"72",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"69",X"00",
		X"00",X"22",X"69",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"69",X"00",
		X"00",X"99",X"99",X"00",X"00",X"66",X"96",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"79",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"D9",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"39",X"00",
		X"00",X"99",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"39",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"05",X"00",X"00",X"05",X"50",X"00",
		X"00",X"05",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"09",X"00",X"00",X"00",X"99",X"BB",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9D",X"B0",X"00",X"B0",X"99",X"BB",X"00",X"0B",X"D9",X"0B",X"00",X"00",X"99",X"0B",X"00",
		X"00",X"99",X"0B",X"00",X"B0",X"95",X"0B",X"00",X"BB",X"55",X"BB",X"00",X"BB",X"99",X"B0",X"00",
		X"00",X"99",X"05",X"00",X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"00",X"00",X"90",X"05",X"00",
		X"0B",X"00",X"B5",X"00",X"B0",X"00",X"B0",X"00",X"00",X"BB",X"05",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"22",X"99",X"99",X"00",X"99",X"97",X"99",X"00",
		X"99",X"92",X"99",X"00",X"99",X"22",X"99",X"00",X"92",X"72",X"99",X"00",X"29",X"72",X"99",X"00",
		X"69",X"72",X"99",X"00",X"69",X"72",X"90",X"00",X"69",X"72",X"90",X"00",X"69",X"72",X"00",X"00",
		X"69",X"72",X"00",X"00",X"69",X"72",X"00",X"00",X"69",X"72",X"90",X"00",X"69",X"72",X"90",X"00",
		X"29",X"72",X"99",X"00",X"92",X"77",X"99",X"00",X"99",X"22",X"99",X"00",X"22",X"22",X"99",X"00",
		X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",
		X"67",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",
		X"66",X"29",X"00",X"00",X"69",X"29",X"00",X"00",X"69",X"29",X"09",X"00",X"69",X"92",X"99",X"00",
		X"99",X"92",X"99",X"00",X"99",X"92",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"27",X"99",X"00",
		X"29",X"27",X"99",X"00",X"29",X"79",X"00",X"00",X"22",X"79",X"00",X"00",X"99",X"79",X"00",X"00",
		X"99",X"79",X"00",X"00",X"99",X"79",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"69",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"26",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"77",X"90",X"00",
		X"22",X"77",X"90",X"00",X"29",X"99",X"90",X"00",X"90",X"99",X"00",X"00",X"29",X"99",X"00",X"00",
		X"29",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"90",X"00",X"00",X"97",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"97",X"90",X"00",X"00",
		X"22",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"79",X"00",X"00",X"22",X"70",X"00",X"00",
		X"22",X"70",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"66",X"69",X"00",X"00",X"26",X"69",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"72",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"27",X"00",
		X"00",X"29",X"72",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"97",X"00",X"00",X"22",X"99",X"00",
		X"00",X"22",X"99",X"00",X"00",X"22",X"27",X"00",X"00",X"27",X"22",X"00",X"00",X"77",X"22",X"00",
		X"00",X"99",X"29",X"00",X"00",X"99",X"76",X"00",X"00",X"99",X"77",X"00",X"00",X"79",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"99",X"99",X"00",X"9E",X"99",X"22",X"00",X"9E",X"99",X"99",
		X"00",X"9E",X"66",X"99",X"00",X"9E",X"22",X"29",X"00",X"9E",X"22",X"92",X"00",X"99",X"22",X"96",
		X"00",X"99",X"22",X"96",X"00",X"92",X"77",X"96",X"00",X"92",X"66",X"96",X"00",X"22",X"22",X"96",
		X"00",X"22",X"22",X"96",X"00",X"92",X"66",X"96",X"00",X"92",X"77",X"96",X"00",X"99",X"22",X"96",
		X"00",X"99",X"22",X"96",X"00",X"9E",X"22",X"92",X"00",X"9E",X"22",X"29",X"00",X"9E",X"66",X"99",
		X"00",X"0E",X"92",X"99",X"00",X"0E",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",
		X"00",X"09",X"62",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"29",X"99",X"00",X"99",X"22",X"29",
		X"00",X"99",X"72",X"22",X"00",X"99",X"77",X"99",X"00",X"99",X"62",X"29",X"00",X"99",X"22",X"92",
		X"00",X"99",X"22",X"92",X"00",X"99",X"22",X"99",X"00",X"9E",X"22",X"99",X"00",X"9E",X"22",X"92",
		X"00",X"EE",X"97",X"96",X"00",X"EE",X"27",X"96",X"00",X"E3",X"22",X"26",X"00",X"33",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"90",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",X"09",X"22",X"29",X"00",X"09",X"22",X"29",
		X"00",X"09",X"22",X"99",X"00",X"09",X"76",X"92",X"00",X"09",X"77",X"29",X"00",X"09",X"27",X"99",
		X"00",X"09",X"22",X"99",X"00",X"09",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"99",
		X"00",X"00",X"62",X"96",X"00",X"00",X"22",X"96",X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"EE",
		X"00",X"00",X"99",X"EE",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",
		X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"72",X"00",X"00",X"97",X"72",
		X"00",X"00",X"27",X"72",X"00",X"00",X"22",X"27",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"92",X"97",X"00",X"00",X"26",X"62",X"00",X"00",X"96",X"69",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"09",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"37",X"EE",X"00",X"00",X"32",X"EE",X"00",X"00",X"76",X"99",X"00",X"00",X"76",X"22",X"00",
		X"00",X"76",X"22",X"00",X"00",X"26",X"22",X"00",X"00",X"27",X"99",X"00",X"00",X"27",X"99",X"00",
		X"00",X"27",X"29",X"00",X"00",X"27",X"29",X"00",X"00",X"27",X"22",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"99",X"27",X"00",X"00",X"92",X"92",X"00",X"00",X"29",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"66",X"99",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"EE",X"99",X"22",X"00",X"EE",X"99",X"99",
		X"00",X"EE",X"66",X"99",X"00",X"EE",X"22",X"29",X"00",X"EE",X"22",X"92",X"00",X"99",X"22",X"96",
		X"00",X"99",X"22",X"96",X"00",X"92",X"77",X"96",X"00",X"92",X"66",X"96",X"00",X"22",X"22",X"96",
		X"00",X"22",X"22",X"96",X"00",X"92",X"66",X"96",X"00",X"92",X"77",X"96",X"00",X"99",X"22",X"96",
		X"00",X"99",X"22",X"96",X"00",X"9E",X"22",X"92",X"00",X"EE",X"22",X"29",X"00",X"9E",X"66",X"99",
		X"00",X"3E",X"92",X"99",X"00",X"03",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"67",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",
		X"00",X"09",X"62",X"00",X"00",X"99",X"29",X"90",X"00",X"99",X"29",X"99",X"00",X"99",X"22",X"29",
		X"00",X"99",X"72",X"22",X"00",X"99",X"77",X"99",X"00",X"99",X"62",X"29",X"00",X"99",X"22",X"92",
		X"00",X"99",X"22",X"92",X"00",X"99",X"22",X"99",X"00",X"9E",X"22",X"99",X"00",X"9E",X"22",X"92",
		X"00",X"EE",X"97",X"96",X"00",X"EE",X"27",X"96",X"00",X"EE",X"22",X"26",X"00",X"9E",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",X"09",X"22",X"29",X"00",X"09",X"22",X"29",
		X"00",X"09",X"22",X"99",X"00",X"09",X"76",X"92",X"00",X"09",X"77",X"29",X"00",X"09",X"27",X"99",
		X"00",X"09",X"22",X"99",X"00",X"09",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"99",
		X"00",X"00",X"62",X"96",X"00",X"00",X"22",X"96",X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"09",X"EE",
		X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",
		X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"72",X"00",X"00",X"97",X"72",
		X"00",X"00",X"27",X"72",X"00",X"00",X"22",X"27",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"92",X"97",X"00",X"00",X"26",X"62",X"00",X"00",X"96",X"69",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"09",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"97",X"EE",X"00",X"00",X"32",X"EE",X"00",X"00",X"36",X"99",X"00",X"00",X"76",X"22",X"00",
		X"00",X"76",X"22",X"00",X"00",X"26",X"22",X"00",X"00",X"27",X"99",X"00",X"00",X"27",X"99",X"00",
		X"09",X"27",X"29",X"00",X"09",X"27",X"29",X"00",X"09",X"27",X"22",X"00",X"09",X"22",X"29",X"00",
		X"09",X"22",X"29",X"00",X"09",X"99",X"27",X"00",X"09",X"92",X"92",X"00",X"09",X"29",X"99",X"00",
		X"09",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"66",X"99",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"22",X"99",X"99",X"00",X"99",X"97",X"99",X"00",
		X"99",X"92",X"99",X"00",X"99",X"22",X"99",X"00",X"92",X"72",X"99",X"00",X"29",X"72",X"99",X"00",
		X"69",X"72",X"99",X"00",X"69",X"72",X"90",X"00",X"69",X"72",X"90",X"00",X"69",X"72",X"00",X"00",
		X"69",X"72",X"00",X"00",X"69",X"72",X"00",X"00",X"69",X"72",X"90",X"00",X"69",X"72",X"90",X"00",
		X"29",X"72",X"99",X"00",X"92",X"77",X"99",X"00",X"99",X"22",X"99",X"00",X"22",X"22",X"99",X"00",
		X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"29",X"00",X"00",X"69",X"29",X"00",X"00",X"69",X"29",X"09",X"00",X"69",X"92",X"99",X"00",
		X"99",X"92",X"99",X"00",X"99",X"92",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"27",X"99",X"00",
		X"29",X"27",X"99",X"00",X"29",X"79",X"00",X"00",X"22",X"79",X"00",X"00",X"99",X"79",X"00",X"00",
		X"99",X"79",X"00",X"00",X"09",X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"62",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"96",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"69",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"26",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"77",X"90",X"00",
		X"22",X"77",X"90",X"00",X"29",X"99",X"90",X"00",X"90",X"99",X"00",X"00",X"29",X"99",X"00",X"00",
		X"29",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"90",X"00",X"00",X"97",X"90",X"00",X"00",
		X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"99",X"00",X"00",
		X"22",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"79",X"00",X"00",X"22",X"70",X"00",X"00",
		X"22",X"70",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"72",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"27",X"00",
		X"00",X"29",X"72",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"97",X"00",X"00",X"22",X"99",X"00",
		X"00",X"22",X"99",X"00",X"00",X"22",X"27",X"00",X"00",X"27",X"22",X"00",X"00",X"77",X"22",X"00",
		X"00",X"99",X"29",X"00",X"00",X"99",X"76",X"00",X"00",X"99",X"77",X"00",X"00",X"79",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"02",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"29",X"00",X"00",
		X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"02",X"06",X"90",
		X"00",X"26",X"22",X"90",X"00",X"62",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"20",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"22",X"22",X"99",
		X"00",X"22",X"22",X"00",X"02",X"22",X"00",X"00",X"29",X"22",X"99",X"00",X"00",X"22",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"03",X"99",X"99",X"00",X"03",X"11",X"55",X"00",X"03",X"44",X"15",
		X"00",X"09",X"44",X"55",X"00",X"09",X"55",X"49",X"00",X"95",X"55",X"95",X"00",X"90",X"44",X"95",
		X"00",X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"41",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"14",X"99",X"00",X"09",X"41",X"99",
		X"00",X"09",X"14",X"99",X"00",X"90",X"55",X"99",X"00",X"93",X"55",X"91",X"00",X"09",X"55",X"19",
		X"00",X"09",X"11",X"59",X"00",X"03",X"11",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"99",X"19",X"00",X"55",X"11",X"59",X"00",X"51",X"55",X"90",X"00",
		X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"59",X"95",X"59",X"00",X"41",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",
		X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"59",X"00",X"44",X"44",X"59",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"90",X"00",
		X"95",X"99",X"90",X"00",X"55",X"55",X"90",X"00",X"99",X"99",X"19",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"34",X"90",
		X"00",X"00",X"44",X"99",X"00",X"00",X"55",X"19",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"44",
		X"00",X"00",X"14",X"95",X"00",X"00",X"54",X"59",X"00",X"00",X"14",X"59",X"00",X"00",X"54",X"99",
		X"00",X"00",X"59",X"99",X"00",X"00",X"41",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"99",
		X"00",X"0E",X"44",X"95",X"00",X"9E",X"14",X"91",X"00",X"9E",X"51",X"94",X"00",X"95",X"95",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"45",X"51",X"00",X"00",X"44",X"55",X"90",X"00",
		X"44",X"99",X"99",X"00",X"44",X"99",X"55",X"00",X"44",X"59",X"59",X"00",X"44",X"44",X"59",X"00",
		X"00",X"95",X"45",X"54",X"00",X"09",X"11",X"14",X"00",X"00",X"51",X"54",X"00",X"00",X"95",X"55",
		X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",
		X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",X"54",X"44",X"00",X"00",X"99",X"44",X"00",X"00",
		X"99",X"49",X"00",X"00",X"59",X"49",X"00",X"00",X"51",X"19",X"00",X"00",X"51",X"19",X"00",X"00",
		X"99",X"91",X"00",X"00",X"09",X"55",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"95",X"99",X"00",X"00",X"54",X"59",X"00",X"00",X"49",X"19",X"00",X"00",X"95",X"15",
		X"00",X"00",X"51",X"41",X"00",X"00",X"51",X"44",X"00",X"09",X"99",X"94",X"00",X"09",X"99",X"59",
		X"00",X"09",X"15",X"45",X"00",X"09",X"44",X"44",X"00",X"9E",X"44",X"59",X"00",X"9E",X"44",X"99",
		X"00",X"99",X"14",X"95",X"00",X"95",X"14",X"99",X"00",X"09",X"54",X"99",X"00",X"00",X"51",X"95",
		X"00",X"00",X"95",X"91",X"00",X"00",X"19",X"14",X"00",X"00",X"45",X"11",X"00",X"00",X"14",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"45",X"90",X"00",X"00",
		X"00",X"00",X"54",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"15",X"00",X"00",X"44",X"51",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"14",X"59",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"95",X"00",X"00",X"94",X"51",X"00",X"00",X"99",X"45",X"00",X"00",
		X"99",X"59",X"00",X"00",X"95",X"90",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"19",X"00",X"00",X"99",X"95",
		X"00",X"00",X"99",X"51",X"00",X"00",X"EE",X"15",X"00",X"00",X"EE",X"55",X"00",X"00",X"53",X"11",
		X"00",X"00",X"14",X"54",X"00",X"00",X"14",X"54",X"00",X"00",X"14",X"91",X"00",X"00",X"54",X"55",
		X"00",X"00",X"51",X"19",X"00",X"00",X"95",X"49",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"59",
		X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"19",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"51",X"00",X"00",
		X"44",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"54",X"00",X"00",
		X"49",X"55",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"59",X"00",X"00",X"09",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"59",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"14",X"EE",X"00",X"09",X"99",X"EE",X"00",
		X"09",X"55",X"33",X"00",X"00",X"15",X"91",X"00",X"00",X"49",X"91",X"00",X"00",X"41",X"91",X"00",
		X"00",X"41",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"14",X"55",X"00",X"00",X"44",X"55",X"00",
		X"00",X"41",X"55",X"00",X"00",X"41",X"15",X"00",X"00",X"44",X"15",X"00",X"00",X"99",X"19",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"59",X"00",
		X"00",X"11",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"44",X"59",X"00",
		X"00",X"44",X"59",X"00",X"00",X"14",X"59",X"00",X"00",X"44",X"99",X"00",X"00",X"14",X"59",X"00",
		X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"54",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",
		X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",
		X"00",X"44",X"59",X"00",X"00",X"11",X"59",X"00",X"00",X"99",X"49",X"00",X"00",X"99",X"91",X"00",
		X"00",X"55",X"55",X"00",X"00",X"15",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"39",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"93",X"05",X"00",X"99",X"39",X"50",X"00",
		X"99",X"93",X"05",X"00",X"99",X"99",X"50",X"00",X"99",X"99",X"05",X"00",X"99",X"99",X"50",X"00",
		X"09",X"90",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"9D",X"00",X"00",X"93",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",X"00",X"00",
		X"39",X"59",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"05",X"00",X"99",X"99",X"50",X"00",
		X"99",X"90",X"05",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",
		X"09",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"99",X"59",X"00",X"55",X"11",X"59",X"00",X"11",X"55",X"90",X"00",
		X"99",X"99",X"90",X"00",X"99",X"59",X"90",X"00",X"59",X"95",X"59",X"00",X"41",X"45",X"99",X"00",
		X"44",X"49",X"99",X"00",X"44",X"19",X"90",X"00",X"44",X"49",X"90",X"00",X"44",X"59",X"90",X"00",
		X"44",X"59",X"90",X"00",X"44",X"59",X"90",X"00",X"44",X"59",X"90",X"00",X"44",X"55",X"90",X"00",
		X"44",X"49",X"90",X"00",X"44",X"41",X"90",X"00",X"99",X"95",X"90",X"00",X"99",X"99",X"90",X"00",
		X"95",X"55",X"90",X"00",X"51",X"51",X"50",X"00",X"99",X"99",X"59",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"45",X"51",X"00",X"00",X"44",X"55",X"90",X"00",
		X"44",X"99",X"99",X"00",X"44",X"99",X"55",X"00",X"44",X"59",X"59",X"00",X"44",X"41",X"59",X"00",
		X"44",X"95",X"99",X"00",X"44",X"99",X"90",X"00",X"44",X"99",X"90",X"00",X"44",X"99",X"90",X"00",
		X"44",X"99",X"90",X"00",X"44",X"99",X"90",X"00",X"54",X"99",X"00",X"00",X"99",X"55",X"00",X"00",
		X"99",X"99",X"00",X"00",X"59",X"55",X"00",X"00",X"51",X"55",X"00",X"00",X"51",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"09",X"59",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"15",X"00",X"00",X"44",X"51",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"51",X"00",X"00",
		X"44",X"95",X"00",X"00",X"54",X"99",X"00",X"00",X"15",X"99",X"00",X"00",X"55",X"99",X"00",X"00",
		X"45",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"19",X"55",X"00",X"00",X"49",X"45",X"00",X"00",
		X"45",X"59",X"00",X"00",X"45",X"90",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"19",X"00",X"00",X"54",X"19",X"00",X"00",X"45",X"55",X"00",X"00",X"55",X"51",X"00",X"00",
		X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"51",X"00",X"00",X"99",X"54",X"00",X"00",
		X"99",X"55",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"59",X"00",X"00",X"14",X"59",X"00",X"00",X"44",X"99",X"00",X"00",X"14",X"59",X"00",
		X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"54",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",
		X"00",X"45",X"59",X"00",X"00",X"55",X"59",X"00",X"00",X"59",X"59",X"00",X"00",X"99",X"19",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"54",X"00",X"00",X"55",X"94",X"00",X"00",X"55",X"95",X"00",
		X"00",X"59",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"55",X"00",X"09",X"44",X"15",
		X"00",X"09",X"44",X"55",X"00",X"09",X"55",X"49",X"00",X"95",X"55",X"95",X"00",X"90",X"99",X"95",
		X"00",X"09",X"D9",X"99",X"00",X"09",X"DD",X"99",X"00",X"09",X"9D",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"9D",X"99",X"00",X"09",X"DD",X"99",X"00",X"99",X"D9",X"99",
		X"00",X"99",X"99",X"99",X"00",X"90",X"99",X"99",X"00",X"95",X"55",X"91",X"00",X"09",X"55",X"19",
		X"00",X"09",X"11",X"59",X"00",X"00",X"11",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"E5",X"90",X"00",X"00",X"35",X"99",X"00",X"00",X"34",X"99",
		X"00",X"00",X"34",X"99",X"00",X"00",X"55",X"19",X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"44",
		X"00",X"00",X"DD",X"15",X"00",X"00",X"9D",X"59",X"00",X"00",X"DD",X"59",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"DD",X"99",
		X"00",X"09",X"99",X"95",X"00",X"9E",X"99",X"91",X"00",X"9E",X"59",X"94",X"00",X"95",X"95",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"54",X"59",X"00",X"00",X"4D",X"19",X"00",X"00",X"DD",X"15",
		X"00",X"00",X"D9",X"41",X"00",X"00",X"99",X"44",X"00",X"09",X"9D",X"54",X"00",X"09",X"DD",X"55",
		X"00",X"09",X"D9",X"55",X"00",X"09",X"9D",X"11",X"00",X"9E",X"D9",X"59",X"00",X"9E",X"DD",X"99",
		X"00",X"99",X"9D",X"95",X"00",X"95",X"99",X"99",X"00",X"09",X"59",X"99",X"00",X"00",X"55",X"95",
		X"00",X"00",X"95",X"91",X"00",X"00",X"19",X"14",X"00",X"00",X"45",X"11",X"00",X"00",X"14",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"DD",X"00",X"00",X"99",X"D9",
		X"00",X"00",X"99",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"DD",X"00",X"00",X"53",X"DD",
		X"00",X"00",X"33",X"D9",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"D9",X"00",X"00",X"54",X"9D",
		X"00",X"00",X"51",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"59",
		X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"59",X"95",X"00",X"00",X"09",X"99",X"00",X"00",X"1D",X"EE",X"00",X"09",X"DD",X"EE",X"00",
		X"09",X"59",X"33",X"00",X"00",X"DD",X"51",X"00",X"00",X"DD",X"51",X"00",X"00",X"DD",X"51",X"00",
		X"00",X"DD",X"55",X"00",X"00",X"DD",X"55",X"00",X"00",X"DD",X"55",X"00",X"00",X"DD",X"55",X"00",
		X"00",X"99",X"55",X"00",X"00",X"99",X"95",X"00",X"00",X"11",X"15",X"00",X"00",X"99",X"11",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"59",X"00",
		X"00",X"11",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"44",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"55",X"00",X"09",X"44",X"15",
		X"00",X"09",X"44",X"55",X"00",X"09",X"55",X"49",X"00",X"95",X"55",X"95",X"00",X"90",X"99",X"95",
		X"00",X"09",X"D9",X"99",X"00",X"09",X"DD",X"99",X"00",X"09",X"9D",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"9D",X"99",X"00",X"09",X"DD",X"99",X"00",X"99",X"D9",X"99",
		X"00",X"99",X"99",X"99",X"00",X"90",X"99",X"99",X"00",X"95",X"55",X"91",X"00",X"09",X"55",X"19",
		X"00",X"09",X"11",X"59",X"00",X"00",X"11",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"45",X"51",X"00",X"00",X"44",X"55",X"90",X"00",
		X"44",X"99",X"99",X"00",X"44",X"99",X"55",X"00",X"44",X"59",X"59",X"00",X"44",X"41",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"34",X"90",
		X"00",X"00",X"44",X"99",X"00",X"00",X"55",X"19",X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"44",
		X"00",X"00",X"DD",X"15",X"00",X"00",X"9D",X"59",X"00",X"00",X"DD",X"59",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"DD",X"99",
		X"00",X"09",X"99",X"95",X"00",X"9E",X"99",X"91",X"00",X"9E",X"59",X"94",X"00",X"95",X"95",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"95",X"90",X"00",X"00",X"54",X"59",X"00",X"00",X"4D",X"19",X"00",X"00",X"DD",X"15",
		X"00",X"00",X"D9",X"41",X"00",X"00",X"99",X"44",X"00",X"09",X"9D",X"54",X"00",X"09",X"DD",X"55",
		X"00",X"09",X"D9",X"55",X"00",X"09",X"9D",X"11",X"00",X"9E",X"D9",X"59",X"00",X"9E",X"DD",X"99",
		X"00",X"99",X"9D",X"95",X"00",X"95",X"99",X"99",X"00",X"09",X"59",X"99",X"00",X"00",X"55",X"95",
		X"00",X"00",X"95",X"91",X"00",X"00",X"19",X"14",X"00",X"00",X"45",X"11",X"00",X"00",X"14",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"DD",X"00",X"00",X"99",X"D9",
		X"00",X"00",X"99",X"99",X"00",X"00",X"91",X"99",X"00",X"00",X"EE",X"DD",X"00",X"00",X"E3",X"DD",
		X"00",X"00",X"33",X"D9",X"00",X"00",X"34",X"99",X"00",X"00",X"14",X"D9",X"00",X"00",X"54",X"9D",
		X"00",X"00",X"51",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"59",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"09",X"95",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"59",X"95",X"00",X"00",X"09",X"99",X"00",X"00",X"1D",X"1E",X"00",X"09",X"DD",X"EE",X"00",
		X"09",X"59",X"31",X"00",X"00",X"DD",X"53",X"00",X"00",X"DD",X"51",X"00",X"00",X"DD",X"51",X"00",
		X"09",X"DD",X"55",X"00",X"09",X"DD",X"55",X"00",X"99",X"DD",X"55",X"00",X"09",X"DD",X"55",X"00",
		X"99",X"99",X"55",X"00",X"09",X"99",X"95",X"00",X"99",X"11",X"15",X"00",X"00",X"99",X"11",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"59",X"00",
		X"00",X"11",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"44",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"99",X"59",X"00",X"55",X"11",X"59",X"00",X"11",X"55",X"90",X"00",
		X"99",X"99",X"90",X"00",X"99",X"59",X"90",X"00",X"59",X"95",X"59",X"00",X"41",X"45",X"99",X"00",
		X"44",X"49",X"99",X"00",X"44",X"19",X"90",X"00",X"44",X"49",X"90",X"00",X"44",X"59",X"90",X"00",
		X"44",X"59",X"90",X"00",X"44",X"59",X"90",X"00",X"44",X"59",X"90",X"00",X"44",X"55",X"90",X"00",
		X"44",X"49",X"90",X"00",X"44",X"41",X"90",X"00",X"99",X"95",X"90",X"00",X"99",X"99",X"90",X"00",
		X"95",X"55",X"90",X"00",X"51",X"51",X"50",X"00",X"99",X"99",X"59",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"95",X"99",X"00",X"44",X"99",X"90",X"00",X"44",X"99",X"90",X"00",X"44",X"99",X"90",X"00",
		X"44",X"99",X"90",X"00",X"44",X"99",X"90",X"00",X"54",X"99",X"00",X"00",X"99",X"55",X"00",X"00",
		X"99",X"99",X"00",X"00",X"59",X"55",X"00",X"00",X"51",X"55",X"00",X"00",X"51",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"11",X"00",X"00",X"09",X"14",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"45",X"54",X"00",X"09",X"11",X"14",X"00",X"00",X"51",X"54",X"00",X"00",X"95",X"55",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"19",X"00",X"00",X"90",X"55",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"15",X"00",X"00",X"44",X"51",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"51",X"00",X"00",
		X"44",X"95",X"00",X"00",X"54",X"99",X"00",X"00",X"15",X"99",X"00",X"00",X"55",X"99",X"00",X"00",
		X"45",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"19",X"55",X"00",X"00",X"49",X"45",X"00",X"00",
		X"45",X"59",X"00",X"00",X"45",X"90",X"00",X"00",X"51",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"19",X"00",X"00",X"54",X"19",X"00",X"00",X"45",X"55",X"00",X"00",X"55",X"51",X"00",X"00",
		X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"51",X"00",X"00",X"99",X"54",X"00",X"00",
		X"99",X"55",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"59",X"00",X"00",X"14",X"59",X"00",X"00",X"44",X"99",X"00",X"00",X"14",X"59",X"00",
		X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"54",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"59",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"59",X"00",
		X"09",X"45",X"59",X"00",X"09",X"55",X"59",X"00",X"99",X"59",X"59",X"00",X"09",X"99",X"19",X"00",
		X"99",X"99",X"44",X"00",X"09",X"99",X"54",X"00",X"99",X"55",X"94",X"00",X"00",X"55",X"95",X"00",
		X"00",X"59",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"92",X"09",X"09",X"00",X"92",X"99",X"99",X"90",X"92",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",
		X"99",X"92",X"92",X"90",X"00",X"92",X"92",X"90",X"00",X"92",X"92",X"90",X"99",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"99",X"99",X"99",X"90",X"99",X"09",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"90",X"90",X"90",X"90",X"99",X"99",X"99",X"90",X"29",X"29",X"29",X"90",X"22",X"22",X"22",
		X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",
		X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",
		X"90",X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"99",X"29",X"29",X"29",X"29",X"99",X"99",X"99",
		X"99",X"90",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"22",X"29",X"29",X"29",X"99",X"92",X"92",X"92",X"99",X"92",X"92",X"92",
		X"00",X"92",X"92",X"92",X"99",X"92",X"92",X"92",X"22",X"92",X"92",X"92",X"22",X"92",X"92",X"92",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"22",X"29",X"29",X"29",
		X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"99",X"90",X"90",X"29",X"29",X"99",X"99",X"22",X"99",X"29",X"29",X"22",X"00",X"22",X"22",
		X"22",X"00",X"22",X"22",X"22",X"99",X"22",X"22",X"29",X"99",X"22",X"22",X"99",X"29",X"22",X"22",
		X"99",X"29",X"22",X"22",X"90",X"29",X"22",X"22",X"90",X"29",X"22",X"22",X"00",X"29",X"22",X"22",
		X"00",X"29",X"22",X"22",X"00",X"29",X"22",X"22",X"99",X"29",X"29",X"29",X"22",X"99",X"99",X"99",
		X"99",X"90",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"90",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"9A",X"99",X"99",X"00",X"A9",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"90",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"90",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"90",X"00",X"00",X"93",X"90",X"00",X"00",X"93",X"00",X"05",X"00",X"99",X"00",X"50",X"00",
		X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"09",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"99",X"00",X"00",X"09",X"99",X"99",X"00",X"05",X"55",X"59",X"00",X"05",X"11",X"95",
		X"00",X"5E",X"44",X"55",X"00",X"9E",X"41",X"15",X"00",X"95",X"99",X"95",X"00",X"59",X"55",X"91",
		X"00",X"95",X"11",X"54",X"00",X"95",X"44",X"54",X"00",X"55",X"44",X"54",X"00",X"55",X"44",X"14",
		X"00",X"55",X"55",X"54",X"00",X"55",X"41",X"14",X"00",X"55",X"11",X"14",X"00",X"55",X"11",X"54",
		X"00",X"59",X"51",X"94",X"00",X"95",X"95",X"91",X"00",X"9E",X"59",X"55",X"00",X"5E",X"11",X"15",
		X"00",X"55",X"14",X"55",X"00",X"05",X"41",X"91",X"00",X"09",X"99",X"59",X"00",X"09",X"99",X"99",
		X"00",X"01",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"50",X"00",X"00",X"99",X"95",X"00",X"99",X"41",X"59",X"00",X"15",X"14",X"59",X"00",
		X"94",X"59",X"59",X"00",X"55",X"99",X"59",X"00",X"49",X"41",X"59",X"00",X"44",X"44",X"59",X"00",
		X"44",X"44",X"59",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"59",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"59",X"00",
		X"44",X"44",X"59",X"00",X"41",X"44",X"59",X"00",X"49",X"45",X"59",X"00",X"51",X"99",X"59",X"00",
		X"94",X"99",X"59",X"00",X"51",X"44",X"55",X"00",X"99",X"44",X"55",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"E3",X"90",
		X"00",X"00",X"E3",X"95",X"00",X"00",X"34",X"55",X"00",X"00",X"44",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"55",X"00",X"00",X"51",X"49",X"00",X"00",X"44",X"99",
		X"00",X"00",X"55",X"99",X"00",X"00",X"14",X"99",X"00",X"59",X"41",X"99",X"00",X"09",X"14",X"99",
		X"00",X"09",X"54",X"99",X"00",X"55",X"91",X"95",X"00",X"95",X"95",X"91",X"00",X"95",X"49",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"99",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"41",X"54",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"49",X"00",X"44",X"94",X"59",X"00",
		X"00",X"95",X"11",X"94",X"00",X"09",X"14",X"91",X"00",X"00",X"14",X"54",X"00",X"00",X"91",X"91",
		X"00",X"00",X"99",X"55",X"00",X"00",X"09",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"54",X"59",X"00",X"44",X"14",X"54",X"00",X"44",X"44",X"51",X"00",X"44",X"44",X"15",X"00",
		X"44",X"44",X"45",X"00",X"44",X"44",X"15",X"00",X"14",X"44",X"59",X"00",X"99",X"44",X"55",X"00",
		X"99",X"44",X"50",X"00",X"19",X"45",X"50",X"00",X"59",X"49",X"50",X"00",X"94",X"95",X"00",X"00",
		X"99",X"95",X"00",X"00",X"09",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"99",X"95",
		X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"59",X"00",X"00",X"99",X"45",X"00",X"00",X"55",X"14",
		X"00",X"00",X"14",X"44",X"00",X"00",X"99",X"54",X"00",X"00",X"95",X"99",X"00",X"09",X"54",X"55",
		X"00",X"09",X"11",X"11",X"00",X"95",X"14",X"41",X"00",X"95",X"54",X"59",X"00",X"99",X"51",X"99",
		X"00",X"99",X"91",X"99",X"00",X"09",X"95",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"19",X"91",
		X"00",X"00",X"49",X"51",X"00",X"00",X"49",X"41",X"00",X"00",X"44",X"44",X"00",X"00",X"54",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"95",X"00",X"00",
		X"00",X"00",X"95",X"44",X"00",X"00",X"99",X"14",X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"54",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"54",X"00",X"00",
		X"44",X"94",X"00",X"00",X"14",X"95",X"00",X"00",X"45",X"99",X"00",X"00",X"59",X"59",X"00",X"00",
		X"99",X"55",X"00",X"00",X"99",X"95",X"50",X"00",X"99",X"51",X"50",X"00",X"95",X"55",X"00",X"00",
		X"54",X"15",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"15",X"00",X"00",X"95",X"55",X"00",X"00",
		X"55",X"95",X"00",X"00",X"15",X"95",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"59",X"00",X"00",
		X"54",X"90",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",
		X"00",X"00",X"91",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"55",X"99",X"00",X"00",X"EE",X"19",
		X"00",X"00",X"EE",X"11",X"00",X"00",X"E3",X"44",X"00",X"00",X"34",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"14",X"00",X"00",X"14",X"54",X"00",X"00",X"11",X"54",
		X"00",X"00",X"54",X"44",X"00",X"00",X"94",X"49",X"00",X"00",X"91",X"99",X"00",X"00",X"91",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"51",X"00",X"00",X"09",X"11",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"45",
		X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"55",X"95",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"49",X"00",X"00",X"54",X"45",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"55",X"45",X"00",X"00",
		X"55",X"59",X"00",X"00",X"51",X"41",X"00",X"00",X"15",X"55",X"00",X"00",X"55",X"59",X"00",X"00",
		X"55",X"90",X"00",X"00",X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"99",X"59",X"00",X"00",X"55",X"5E",X"00",
		X"00",X"99",X"EE",X"00",X"00",X"99",X"9E",X"00",X"00",X"59",X"53",X"00",X"00",X"99",X"11",X"00",
		X"00",X"95",X"44",X"00",X"00",X"91",X"11",X"00",X"00",X"54",X"14",X"00",X"00",X"54",X"51",X"00",
		X"00",X"14",X"94",X"00",X"00",X"14",X"91",X"00",X"00",X"44",X"95",X"00",X"00",X"14",X"59",X"00",
		X"00",X"14",X"19",X"00",X"00",X"45",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"41",X"19",X"00",X"00",X"11",X"55",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",
		X"00",X"44",X"14",X"00",X"00",X"44",X"95",X"00",X"00",X"14",X"99",X"00",X"00",X"41",X"59",X"00",
		X"00",X"44",X"49",X"00",X"00",X"59",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"11",X"41",X"00",X"00",X"41",X"49",X"00",X"00",X"44",X"15",X"00",X"00",X"41",X"99",X"00",
		X"00",X"44",X"95",X"00",X"00",X"59",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"51",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"95",X"95",X"00",X"00",X"11",X"14",X"00",X"00",X"55",X"51",X"00",
		X"00",X"55",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"39",X"00",X"00",X"09",X"39",X"00",X"00",X"09",X"39",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9A",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"39",X"99",X"00",X"00",
		X"93",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"05",X"00",X"99",X"90",X"50",X"00",
		X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",
		X"00",X"39",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"00",
		X"00",X"99",X"55",X"00",X"00",X"99",X"50",X"00",X"00",X"99",X"05",X"00",X"00",X"90",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"50",X"00",X"00",X"99",X"95",X"00",X"99",X"41",X"59",X"00",X"15",X"14",X"59",X"00",
		X"94",X"59",X"99",X"00",X"55",X"99",X"99",X"00",X"49",X"41",X"59",X"00",X"44",X"44",X"59",X"00",
		X"44",X"44",X"99",X"00",X"44",X"45",X"99",X"00",X"44",X"45",X"90",X"00",X"44",X"45",X"00",X"00",
		X"44",X"44",X"90",X"00",X"44",X"45",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",
		X"44",X"44",X"09",X"00",X"41",X"44",X"99",X"00",X"49",X"45",X"59",X"00",X"51",X"99",X"99",X"00",
		X"94",X"99",X"99",X"00",X"51",X"44",X"99",X"00",X"99",X"45",X"99",X"00",X"00",X"99",X"09",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"99",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"41",X"54",X"90",X"00",
		X"44",X"59",X"99",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"49",X"00",X"44",X"94",X"59",X"00",
		X"44",X"54",X"59",X"00",X"44",X"14",X"59",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"90",X"00",X"14",X"45",X"50",X"00",X"99",X"44",X"55",X"00",
		X"99",X"45",X"00",X"00",X"19",X"41",X"00",X"00",X"59",X"41",X"00",X"00",X"94",X"95",X"00",X"00",
		X"99",X"95",X"00",X"00",X"09",X"45",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"45",X"00",X"00",
		X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"54",X"00",X"00",
		X"44",X"94",X"00",X"00",X"14",X"95",X"00",X"00",X"45",X"99",X"00",X"00",X"59",X"59",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"99",X"50",X"00",X"99",X"99",X"50",X"00",X"95",X"95",X"00",X"00",
		X"54",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"95",X"99",X"00",X"00",
		X"55",X"99",X"00",X"00",X"15",X"95",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",
		X"54",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"49",X"00",X"00",X"54",X"45",X"00",X"00",X"44",X"54",X"00",X"00",
		X"44",X"45",X"00",X"00",X"54",X"59",X"00",X"00",X"55",X"49",X"00",X"00",X"59",X"95",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"59",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"45",
		X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",
		X"00",X"44",X"14",X"00",X"00",X"44",X"95",X"00",X"00",X"14",X"99",X"00",X"00",X"41",X"59",X"00",
		X"00",X"44",X"49",X"00",X"00",X"59",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"11",X"41",X"00",X"00",X"41",X"49",X"00",X"00",X"44",X"15",X"00",X"00",X"11",X"99",X"00",
		X"00",X"15",X"95",X"00",X"00",X"59",X"55",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"55",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"05",X"99",X"00",X"00",X"09",X"99",X"99",X"00",X"05",X"55",X"59",X"00",X"05",X"11",X"95",
		X"00",X"59",X"44",X"55",X"00",X"93",X"41",X"15",X"00",X"95",X"99",X"95",X"00",X"59",X"99",X"91",
		X"00",X"05",X"99",X"54",X"00",X"05",X"DD",X"54",X"00",X"05",X"D9",X"54",X"00",X"05",X"9D",X"14",
		X"00",X"00",X"99",X"54",X"00",X"00",X"9D",X"14",X"00",X"00",X"D9",X"14",X"00",X"05",X"DD",X"54",
		X"00",X"09",X"99",X"94",X"00",X"95",X"99",X"91",X"00",X"95",X"59",X"55",X"00",X"59",X"11",X"15",
		X"00",X"55",X"14",X"55",X"00",X"05",X"41",X"91",X"00",X"09",X"99",X"59",X"00",X"09",X"99",X"99",
		X"00",X"01",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"E3",X"99",X"00",X"00",X"E3",X"99",
		X"00",X"00",X"35",X"95",X"00",X"00",X"34",X"55",X"00",X"00",X"34",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"51",X"00",X"00",X"9D",X"49",X"00",X"00",X"99",X"99",
		X"00",X"00",X"9D",X"99",X"00",X"00",X"9D",X"99",X"00",X"05",X"9D",X"99",X"00",X"05",X"DD",X"99",
		X"00",X"59",X"9D",X"99",X"00",X"55",X"99",X"95",X"00",X"95",X"99",X"91",X"00",X"95",X"49",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"59",X"00",X"00",X"99",X"45",X"00",X"00",X"5D",X"14",
		X"00",X"00",X"D9",X"44",X"00",X"00",X"99",X"54",X"00",X"00",X"9D",X"99",X"00",X"09",X"9D",X"99",
		X"00",X"09",X"9D",X"91",X"00",X"95",X"D9",X"41",X"00",X"95",X"9D",X"59",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"19",X"91",
		X"00",X"00",X"49",X"51",X"00",X"00",X"49",X"41",X"00",X"00",X"44",X"44",X"00",X"00",X"54",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",
		X"00",X"00",X"01",X"DE",X"00",X"00",X"59",X"95",X"00",X"00",X"55",X"99",X"00",X"00",X"EE",X"D9",
		X"00",X"00",X"EE",X"D9",X"00",X"00",X"3E",X"9D",X"00",X"00",X"33",X"9D",X"00",X"00",X"44",X"DD",
		X"00",X"00",X"54",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"11",X"99",
		X"00",X"00",X"54",X"14",X"00",X"00",X"94",X"49",X"00",X"00",X"91",X"99",X"00",X"00",X"91",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"51",X"00",X"00",X"09",X"11",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"99",X"59",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"EE",X"00",X"00",X"99",X"EE",X"00",X"00",X"59",X"33",X"00",X"00",X"99",X"11",X"00",
		X"00",X"95",X"44",X"00",X"00",X"99",X"11",X"00",X"00",X"59",X"14",X"00",X"00",X"59",X"51",X"00",
		X"00",X"99",X"94",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"11",X"99",X"00",X"00",X"45",X"49",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"41",X"19",X"00",X"00",X"11",X"55",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"09",X"00",X"00",X"09",X"99",X"99",X"00",X"05",X"55",X"59",X"00",X"05",X"11",X"95",
		X"00",X"5E",X"44",X"55",X"00",X"91",X"41",X"15",X"00",X"95",X"99",X"95",X"00",X"59",X"99",X"91",
		X"00",X"05",X"99",X"54",X"00",X"05",X"DD",X"54",X"00",X"05",X"D9",X"54",X"00",X"05",X"9D",X"14",
		X"00",X"00",X"99",X"54",X"00",X"00",X"9D",X"14",X"00",X"00",X"D9",X"14",X"00",X"05",X"DD",X"54",
		X"00",X"09",X"99",X"94",X"00",X"95",X"99",X"91",X"00",X"95",X"59",X"55",X"00",X"59",X"11",X"15",
		X"00",X"55",X"14",X"55",X"00",X"05",X"41",X"91",X"00",X"09",X"99",X"59",X"00",X"09",X"99",X"99",
		X"00",X"01",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"41",X"54",X"00",X"00",
		X"44",X"59",X"99",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"49",X"00",X"44",X"94",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"E3",X"99",
		X"00",X"00",X"EE",X"95",X"00",X"00",X"E3",X"55",X"00",X"00",X"E3",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"51",X"00",X"00",X"9D",X"49",X"00",X"00",X"99",X"99",
		X"00",X"00",X"9D",X"99",X"00",X"00",X"9D",X"99",X"00",X"05",X"9D",X"99",X"00",X"05",X"DD",X"99",
		X"00",X"59",X"9D",X"99",X"00",X"55",X"99",X"95",X"00",X"95",X"99",X"91",X"00",X"95",X"49",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"59",X"00",X"00",X"99",X"45",X"00",X"00",X"5D",X"14",
		X"00",X"00",X"D9",X"44",X"00",X"00",X"99",X"54",X"00",X"00",X"9D",X"99",X"00",X"09",X"9D",X"99",
		X"00",X"09",X"9D",X"91",X"00",X"95",X"D9",X"41",X"00",X"95",X"9D",X"59",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"19",X"91",
		X"00",X"09",X"49",X"51",X"00",X"09",X"49",X"41",X"00",X"00",X"44",X"44",X"00",X"00",X"54",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",
		X"00",X"00",X"01",X"D9",X"00",X"00",X"59",X"95",X"00",X"00",X"55",X"99",X"00",X"00",X"EE",X"D9",
		X"00",X"00",X"EE",X"D9",X"00",X"00",X"3E",X"9D",X"00",X"00",X"53",X"9D",X"00",X"00",X"44",X"DD",
		X"00",X"00",X"54",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"11",X"99",
		X"00",X"00",X"54",X"14",X"00",X"00",X"94",X"49",X"00",X"00",X"91",X"99",X"00",X"00",X"91",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"51",X"00",X"00",X"09",X"11",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"99",X"59",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"5E",X"00",X"00",X"99",X"EE",X"00",X"00",X"59",X"EE",X"00",X"99",X"99",X"33",X"00",
		X"09",X"95",X"44",X"00",X"99",X"99",X"11",X"00",X"09",X"59",X"14",X"00",X"99",X"59",X"51",X"00",
		X"09",X"99",X"94",X"00",X"99",X"99",X"91",X"00",X"09",X"99",X"95",X"00",X"09",X"99",X"59",X"00",
		X"09",X"11",X"99",X"00",X"09",X"45",X"49",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"41",X"19",X"00",X"00",X"11",X"55",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"50",X"00",X"00",X"99",X"95",X"00",X"99",X"41",X"59",X"00",X"15",X"14",X"59",X"00",
		X"94",X"59",X"99",X"00",X"55",X"99",X"99",X"00",X"49",X"41",X"59",X"00",X"44",X"44",X"59",X"00",
		X"44",X"44",X"99",X"00",X"44",X"45",X"99",X"00",X"44",X"45",X"90",X"00",X"44",X"45",X"00",X"00",
		X"44",X"44",X"90",X"00",X"44",X"45",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"90",X"00",
		X"44",X"44",X"09",X"00",X"41",X"44",X"99",X"00",X"49",X"45",X"59",X"00",X"51",X"99",X"99",X"00",
		X"94",X"99",X"99",X"00",X"51",X"44",X"99",X"00",X"99",X"45",X"99",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"54",X"59",X"00",X"44",X"14",X"59",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"90",X"00",X"14",X"45",X"50",X"00",X"99",X"44",X"55",X"00",
		X"99",X"45",X"00",X"00",X"19",X"41",X"00",X"00",X"59",X"41",X"00",X"00",X"94",X"95",X"00",X"00",
		X"99",X"95",X"00",X"00",X"99",X"45",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"45",X"00",X"00",
		X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"11",X"94",X"00",X"09",X"14",X"91",X"00",X"00",X"14",X"54",X"00",X"09",X"91",X"91",
		X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"19",X"00",X"00",X"99",X"19",X"00",X"00",X"09",X"95",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"19",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"54",X"00",X"00",
		X"44",X"94",X"00",X"00",X"14",X"95",X"00",X"00",X"45",X"99",X"00",X"00",X"59",X"59",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"99",X"50",X"00",X"99",X"99",X"50",X"00",X"95",X"95",X"00",X"00",
		X"54",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"95",X"99",X"00",X"00",
		X"55",X"99",X"00",X"00",X"15",X"95",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",
		X"54",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"49",X"00",X"00",X"54",X"45",X"00",X"00",X"44",X"54",X"00",X"00",
		X"44",X"45",X"00",X"00",X"54",X"59",X"00",X"00",X"55",X"49",X"00",X"00",X"59",X"95",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"59",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"45",
		X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",
		X"00",X"44",X"14",X"00",X"00",X"44",X"95",X"00",X"00",X"14",X"99",X"00",X"00",X"41",X"59",X"00",
		X"00",X"44",X"49",X"00",X"00",X"59",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"99",X"11",X"41",X"00",X"09",X"41",X"49",X"00",X"99",X"44",X"15",X"00",X"99",X"11",X"99",X"00",
		X"99",X"15",X"95",X"00",X"99",X"59",X"55",X"00",X"09",X"99",X"95",X"00",X"99",X"99",X"59",X"00",
		X"99",X"99",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"55",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"D9",X"99",X"00",
		X"00",X"99",X"99",X"00",X"C0",X"99",X"99",X"00",X"0C",X"99",X"99",X"C0",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"CC",X"99",X"99",X"00",X"0C",X"99",X"99",X"00",
		X"00",X"99",X"95",X"00",X"00",X"99",X"50",X"00",X"0C",X"99",X"00",X"00",X"00",X"05",X"50",X"00",
		X"00",X"05",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"CC",X"C0",X"00",X"00",X"CC",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"07",X"77",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"74",X"00",X"00",X"77",X"74",
		X"00",X"00",X"77",X"74",X"00",X"00",X"77",X"12",X"00",X"00",X"77",X"23",X"00",X"00",X"77",X"33",
		X"00",X"00",X"77",X"33",X"00",X"00",X"77",X"32",X"00",X"00",X"77",X"33",X"00",X"00",X"77",X"33",
		X"00",X"00",X"77",X"23",X"00",X"00",X"77",X"33",X"00",X"00",X"77",X"23",X"00",X"00",X"77",X"22",
		X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"12",X"00",X"00",X"74",X"12",X"00",X"00",X"77",X"12",
		X"00",X"00",X"47",X"22",X"00",X"00",X"07",X"22",X"00",X"00",X"07",X"22",X"00",X"00",X"07",X"22",
		X"00",X"00",X"07",X"22",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"23",X"00",X"00",X"77",X"12",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"70",X"00",
		X"77",X"77",X"70",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"07",X"00",
		X"77",X"77",X"70",X"00",X"77",X"77",X"77",X"00",X"47",X"77",X"77",X"00",X"44",X"77",X"77",X"00",
		X"44",X"77",X"77",X"00",X"11",X"77",X"77",X"00",X"11",X"77",X"77",X"00",X"11",X"77",X"77",X"00",
		X"11",X"77",X"77",X"70",X"22",X"77",X"77",X"07",X"44",X"77",X"77",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"17",X"77",X"77",X"70",X"67",X"77",X"77",X"70",X"17",X"77",X"77",X"77",
		X"14",X"77",X"77",X"77",X"22",X"77",X"77",X"77",X"33",X"77",X"77",X"77",X"23",X"77",X"77",X"77",
		X"33",X"77",X"77",X"77",X"22",X"77",X"77",X"47",X"22",X"77",X"77",X"77",X"11",X"77",X"77",X"74",
		X"00",X"00",X"77",X"11",X"00",X"00",X"77",X"21",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"11",
		X"00",X"00",X"77",X"14",X"00",X"00",X"07",X"14",X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"42",
		X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"74",X"00",X"00",X"00",X"74",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"74",
		X"00",X"00",X"0B",X"44",X"00",X"99",X"BC",X"42",X"00",X"9B",X"CB",X"12",X"00",X"A9",X"BB",X"21",
		X"04",X"BB",X"B9",X"22",X"09",X"AB",X"B7",X"22",X"99",X"BA",X"B7",X"12",X"99",X"BA",X"B7",X"12",
		X"AC",X"AA",X"B7",X"12",X"AB",X"AA",X"97",X"11",X"AB",X"AA",X"B7",X"11",X"AB",X"AA",X"B7",X"11",
		X"11",X"77",X"77",X"77",X"11",X"77",X"77",X"77",X"41",X"77",X"77",X"77",X"41",X"77",X"77",X"77",
		X"42",X"77",X"77",X"77",X"11",X"77",X"77",X"77",X"11",X"77",X"77",X"77",X"12",X"77",X"77",X"77",
		X"21",X"77",X"77",X"77",X"14",X"77",X"77",X"77",X"14",X"79",X"77",X"77",X"47",X"47",X"77",X"77",
		X"47",X"77",X"77",X"77",X"77",X"47",X"77",X"77",X"74",X"44",X"77",X"77",X"11",X"41",X"77",X"77",
		X"11",X"41",X"77",X"77",X"11",X"42",X"A7",X"77",X"11",X"41",X"A7",X"77",X"21",X"41",X"AA",X"77",
		X"22",X"41",X"AA",X"77",X"22",X"41",X"BA",X"74",X"22",X"21",X"BA",X"99",X"22",X"11",X"BA",X"99",
		X"22",X"12",X"BB",X"99",X"22",X"22",X"BB",X"99",X"23",X"21",X"BB",X"99",X"32",X"24",X"BB",X"99",
		X"22",X"19",X"9A",X"A9",X"22",X"49",X"77",X"AA",X"22",X"9A",X"79",X"AA",X"22",X"99",X"77",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"CB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"B7",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"02",X"22",X"00",X"00",X"02",X"21",X"00",X"00",X"22",X"21",X"00",X"00",X"23",X"21",
		X"BB",X"BA",X"B7",X"11",X"BB",X"AA",X"B7",X"11",X"BB",X"BA",X"79",X"11",X"BB",X"AA",X"79",X"11",
		X"BB",X"AA",X"99",X"11",X"BA",X"9A",X"99",X"11",X"BA",X"AA",X"9A",X"11",X"AA",X"AA",X"AA",X"11",
		X"9B",X"AA",X"AA",X"41",X"9A",X"BA",X"A9",X"41",X"9A",X"AA",X"99",X"41",X"99",X"AA",X"A9",X"41",
		X"A9",X"AA",X"99",X"41",X"BA",X"BA",X"99",X"41",X"A7",X"AA",X"99",X"44",X"A4",X"BA",X"99",X"A4",
		X"A4",X"AA",X"99",X"A4",X"94",X"AA",X"99",X"A4",X"99",X"AA",X"99",X"94",X"79",X"AA",X"99",X"A4",
		X"79",X"AA",X"99",X"94",X"99",X"AA",X"97",X"97",X"9B",X"AA",X"99",X"97",X"9B",X"9B",X"99",X"97",
		X"9B",X"9A",X"99",X"77",X"9B",X"AB",X"99",X"79",X"BB",X"BB",X"99",X"74",X"AB",X"BB",X"A9",X"49",
		X"AB",X"BB",X"99",X"77",X"AB",X"BB",X"A9",X"79",X"AA",X"BB",X"A9",X"49",X"AA",X"BB",X"99",X"94",
		X"22",X"AB",X"99",X"BA",X"22",X"BB",X"99",X"BB",X"22",X"BB",X"A9",X"CC",X"22",X"BA",X"99",X"CC",
		X"22",X"A9",X"99",X"CC",X"22",X"A9",X"9A",X"CB",X"22",X"99",X"BB",X"BB",X"22",X"9A",X"9B",X"BB",
		X"22",X"AA",X"BB",X"BB",X"32",X"AA",X"BA",X"BB",X"22",X"AA",X"BB",X"BB",X"24",X"AA",X"BB",X"BA",
		X"4B",X"AA",X"AB",X"BB",X"AB",X"AA",X"BB",X"A7",X"AB",X"BA",X"AA",X"AA",X"9B",X"AA",X"BB",X"AB",
		X"AA",X"AA",X"BB",X"AA",X"AA",X"AA",X"BB",X"AA",X"BA",X"BA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"BA",X"BA",X"AA",X"99",X"BA",X"AA",X"AA",X"77",X"BB",
		X"BA",X"AA",X"77",X"BB",X"AB",X"BA",X"77",X"BB",X"BB",X"BA",X"77",X"BB",X"BB",X"BB",X"97",X"1A",
		X"BB",X"BB",X"77",X"77",X"BB",X"BB",X"77",X"17",X"BB",X"BB",X"97",X"22",X"BB",X"BB",X"77",X"22",
		X"00",X"00",X"23",X"11",X"00",X"00",X"32",X"11",X"00",X"00",X"22",X"14",X"00",X"00",X"22",X"11",
		X"00",X"00",X"22",X"41",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"21",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"21",X"00",
		X"00",X"01",X"21",X"00",X"00",X"01",X"22",X"00",X"00",X"02",X"22",X"00",X"00",X"01",X"22",X"00",
		X"00",X"01",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"AA",X"CB",X"99",X"97",X"AA",X"BB",X"99",X"99",X"BA",X"BA",X"99",X"97",X"0A",X"BA",X"99",X"99",
		X"0B",X"AA",X"99",X"97",X"09",X"AA",X"99",X"9B",X"00",X"AA",X"79",X"7B",X"09",X"9A",X"99",X"B6",
		X"09",X"99",X"99",X"6D",X"99",X"99",X"AA",X"79",X"BB",X"9A",X"AA",X"A7",X"B9",X"99",X"A9",X"99",
		X"99",X"99",X"AB",X"99",X"44",X"A9",X"AB",X"99",X"77",X"AB",X"AB",X"99",X"07",X"99",X"AA",X"A9",
		X"00",X"49",X"9A",X"BA",X"00",X"77",X"9A",X"BD",X"00",X"11",X"99",X"96",X"00",X"21",X"B9",X"97",
		X"00",X"12",X"BB",X"99",X"00",X"22",X"9B",X"9B",X"00",X"22",X"99",X"9B",X"00",X"22",X"79",X"AB",
		X"00",X"22",X"7B",X"BB",X"00",X"22",X"7B",X"AA",X"00",X"22",X"7B",X"77",X"00",X"22",X"BB",X"14",
		X"00",X"22",X"79",X"22",X"00",X"22",X"47",X"22",X"00",X"22",X"47",X"22",X"00",X"22",X"72",X"A2",
		X"BC",X"BB",X"77",X"22",X"CC",X"BB",X"77",X"42",X"CC",X"BA",X"97",X"42",X"CC",X"BA",X"97",X"42",
		X"CC",X"BB",X"97",X"44",X"CC",X"BB",X"77",X"44",X"BC",X"BB",X"77",X"44",X"BB",X"BA",X"77",X"44",
		X"BB",X"BB",X"97",X"44",X"AB",X"BA",X"77",X"44",X"AA",X"BA",X"77",X"44",X"AA",X"AA",X"77",X"41",
		X"AA",X"BA",X"77",X"41",X"AA",X"A9",X"77",X"12",X"AA",X"99",X"77",X"11",X"AA",X"99",X"79",X"42",
		X"BB",X"97",X"97",X"12",X"B9",X"79",X"70",X"12",X"99",X"97",X"90",X"22",X"9A",X"77",X"00",X"C1",
		X"AA",X"77",X"00",X"22",X"AA",X"77",X"00",X"12",X"BB",X"77",X"00",X"22",X"A9",X"77",X"00",X"22",
		X"99",X"77",X"00",X"22",X"77",X"77",X"00",X"22",X"79",X"77",X"00",X"22",X"77",X"97",X"00",X"22",
		X"21",X"49",X"00",X"22",X"12",X"41",X"00",X"22",X"22",X"41",X"00",X"22",X"21",X"12",X"00",X"21",
		X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"27",X"00",X"00",X"22",X"22",X"00",X"00",X"12",X"12",
		X"00",X"00",X"12",X"11",X"00",X"00",X"11",X"21",X"00",X"00",X"01",X"11",X"00",X"00",X"01",X"21",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"12",X"92",X"00",X"12",X"22",X"9A",X"00",X"21",X"22",X"7B",X"00",X"11",X"22",X"27",
		X"00",X"12",X"22",X"22",X"00",X"21",X"22",X"23",X"00",X"12",X"12",X"22",X"00",X"21",X"11",X"23",
		X"00",X"12",X"24",X"32",X"00",X"42",X"42",X"23",X"00",X"12",X"22",X"22",X"00",X"11",X"32",X"22",
		X"00",X"41",X"22",X"22",X"00",X"14",X"22",X"22",X"00",X"41",X"22",X"22",X"00",X"12",X"22",X"22",
		X"00",X"14",X"22",X"22",X"00",X"44",X"22",X"22",X"22",X"11",X"12",X"2C",X"22",X"22",X"22",X"22",
		X"21",X"12",X"21",X"22",X"22",X"11",X"12",X"11",X"22",X"22",X"41",X"22",X"22",X"22",X"44",X"55",
		X"21",X"22",X"44",X"5E",X"21",X"11",X"77",X"EE",X"22",X"14",X"47",X"57",X"21",X"14",X"44",X"55",
		X"12",X"21",X"55",X"55",X"44",X"11",X"5E",X"55",X"01",X"11",X"E7",X"55",X"00",X"41",X"5E",X"65",
		X"22",X"44",X"00",X"22",X"22",X"44",X"00",X"22",X"22",X"14",X"00",X"22",X"22",X"14",X"00",X"22",
		X"22",X"14",X"00",X"22",X"22",X"14",X"00",X"22",X"22",X"44",X"00",X"22",X"22",X"47",X"00",X"22",
		X"22",X"47",X"00",X"22",X"32",X"75",X"E0",X"12",X"32",X"75",X"E0",X"12",X"22",X"55",X"7E",X"12",
		X"22",X"55",X"55",X"41",X"22",X"57",X"77",X"01",X"22",X"75",X"75",X"04",X"22",X"55",X"75",X"00",
		X"22",X"E5",X"77",X"00",X"27",X"E5",X"57",X"00",X"2E",X"E5",X"57",X"00",X"EE",X"E5",X"77",X"00",
		X"E5",X"E5",X"55",X"00",X"E5",X"55",X"55",X"00",X"5E",X"E7",X"55",X"00",X"E5",X"55",X"55",X"00",
		X"E5",X"75",X"55",X"00",X"EE",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"57",X"55",X"55",X"00",X"55",X"55",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"01",X"22",
		X"00",X"00",X"02",X"22",X"00",X"00",X"12",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",
		X"00",X"41",X"55",X"55",X"00",X"71",X"75",X"55",X"00",X"71",X"55",X"55",X"00",X"71",X"75",X"55",
		X"00",X"74",X"57",X"55",X"00",X"77",X"75",X"55",X"05",X"47",X"57",X"55",X"55",X"55",X"55",X"55",
		X"EE",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"77",X"55",X"EE",X"45",X"22",X"55",X"77",X"57",
		X"22",X"55",X"55",X"75",X"23",X"55",X"55",X"77",X"32",X"55",X"EE",X"77",X"25",X"55",X"EE",X"77",
		X"22",X"55",X"EE",X"57",X"22",X"5E",X"E5",X"77",X"22",X"75",X"55",X"75",X"22",X"17",X"55",X"77",
		X"22",X"21",X"55",X"57",X"22",X"22",X"55",X"77",X"22",X"22",X"E5",X"77",X"22",X"21",X"75",X"77",
		X"22",X"22",X"77",X"77",X"22",X"22",X"17",X"75",X"22",X"22",X"71",X"75",X"22",X"22",X"17",X"50",
		X"22",X"22",X"71",X"20",X"22",X"11",X"17",X"00",X"22",X"21",X"77",X"00",X"11",X"11",X"74",X"00",
		X"57",X"55",X"55",X"50",X"55",X"EE",X"55",X"50",X"55",X"5E",X"55",X"50",X"75",X"EE",X"55",X"50",
		X"57",X"EE",X"55",X"50",X"75",X"EE",X"55",X"50",X"57",X"55",X"55",X"50",X"55",X"EE",X"55",X"50",
		X"57",X"5E",X"55",X"50",X"55",X"EE",X"55",X"50",X"55",X"EE",X"55",X"50",X"55",X"E5",X"55",X"50",
		X"55",X"EE",X"55",X"50",X"55",X"5E",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"77",X"55",X"50",
		X"55",X"11",X"77",X"50",X"51",X"22",X"11",X"50",X"77",X"22",X"12",X"50",X"12",X"22",X"21",X"50",
		X"21",X"22",X"22",X"50",X"12",X"22",X"22",X"00",X"21",X"22",X"22",X"00",X"12",X"22",X"22",X"00",
		X"22",X"22",X"21",X"00",X"22",X"22",X"22",X"00",X"12",X"22",X"22",X"00",X"12",X"22",X"21",X"00",
		X"12",X"22",X"22",X"00",X"12",X"22",X"21",X"00",X"12",X"22",X"12",X"00",X"12",X"22",X"21",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"04",X"00",X"77",X"44",X"4C",X"00",
		X"74",X"FD",X"4C",X"00",X"CC",X"FF",X"CC",X"00",X"77",X"FD",X"CC",X"00",X"7C",X"6C",X"CB",X"00",
		X"77",X"F6",X"D7",X"00",X"7C",X"F6",X"C7",X"00",X"77",X"F6",X"C7",X"00",X"7B",X"F6",X"C7",X"00",
		X"77",X"FD",X"C7",X"00",X"7C",X"FD",X"77",X"00",X"00",X"FD",X"77",X"00",X"C7",X"6D",X"74",X"00",
		X"D7",X"FD",X"74",X"00",X"D0",X"6D",X"7D",X"00",X"7B",X"FD",X"7D",X"00",X"7D",X"6D",X"DD",X"00",
		X"7D",X"CD",X"D9",X"00",X"77",X"CC",X"C7",X"00",X"07",X"DC",X"77",X"00",X"07",X"DC",X"77",X"00",
		X"07",X"DC",X"70",X"00",X"00",X"CD",X"70",X"00",X"00",X"CD",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"CF",X"00",X"00",
		X"00",X"CF",X"00",X"00",X"00",X"C6",X"00",X"00",X"00",X"DF",X"00",X"00",X"00",X"CF",X"00",X"00",
		X"00",X"CF",X"00",X"00",X"00",X"C6",X"00",X"00",X"00",X"FF",X"70",X"00",X"00",X"FF",X"70",X"00",
		X"00",X"FF",X"77",X"00",X"07",X"CC",X"77",X"00",X"07",X"77",X"77",X"00",X"07",X"77",X"77",X"00",
		X"07",X"F7",X"57",X"00",X"07",X"F7",X"77",X"00",X"07",X"F7",X"77",X"00",X"07",X"F7",X"77",X"00",
		X"07",X"F7",X"77",X"00",X"07",X"F7",X"77",X"00",X"07",X"77",X"77",X"00",X"07",X"67",X"57",X"00",
		X"07",X"77",X"77",X"00",X"07",X"77",X"57",X"00",X"77",X"77",X"77",X"00",X"77",X"F7",X"77",X"00",
		X"77",X"77",X"77",X"00",X"07",X"77",X"77",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"BA",X"B7",X"11",X"BB",X"AA",X"B7",X"11",X"BB",X"BA",X"79",X"11",X"BB",X"AA",X"79",X"11",
		X"BB",X"AA",X"99",X"11",X"BA",X"9A",X"99",X"11",X"BA",X"AA",X"9A",X"11",X"AA",X"AA",X"AA",X"11",
		X"9B",X"AA",X"AA",X"41",X"9A",X"BA",X"A9",X"41",X"9A",X"AA",X"99",X"41",X"99",X"AA",X"A9",X"41",
		X"A9",X"AA",X"99",X"41",X"BA",X"BA",X"99",X"41",X"A7",X"AA",X"99",X"44",X"A4",X"BA",X"99",X"A4",
		X"A4",X"AA",X"99",X"A4",X"94",X"AA",X"99",X"A4",X"99",X"AA",X"99",X"94",X"79",X"AA",X"99",X"A4",
		X"79",X"AA",X"99",X"94",X"99",X"AA",X"97",X"97",X"9B",X"AA",X"99",X"97",X"9B",X"9B",X"99",X"97",
		X"9B",X"BA",X"99",X"77",X"9B",X"BB",X"99",X"79",X"BB",X"BB",X"99",X"74",X"AB",X"BB",X"A9",X"49",
		X"AB",X"BB",X"99",X"77",X"AB",X"BB",X"A9",X"79",X"AA",X"BB",X"A9",X"49",X"AA",X"BB",X"99",X"94",
		X"BC",X"BB",X"77",X"22",X"CC",X"BB",X"77",X"42",X"CC",X"BB",X"97",X"42",X"CC",X"BB",X"97",X"42",
		X"CC",X"BB",X"97",X"44",X"CC",X"BB",X"77",X"44",X"BC",X"BB",X"77",X"44",X"BB",X"BA",X"77",X"44",
		X"BB",X"BB",X"97",X"44",X"AB",X"BA",X"77",X"44",X"AA",X"BA",X"77",X"44",X"AA",X"AA",X"77",X"41",
		X"AA",X"BA",X"77",X"41",X"AA",X"A9",X"77",X"12",X"AA",X"99",X"77",X"11",X"AA",X"99",X"79",X"42",
		X"BB",X"97",X"97",X"12",X"B9",X"79",X"70",X"12",X"99",X"97",X"90",X"22",X"9A",X"77",X"00",X"C1",
		X"AA",X"77",X"00",X"22",X"AA",X"77",X"00",X"12",X"BB",X"77",X"00",X"22",X"A9",X"77",X"00",X"22",
		X"99",X"77",X"00",X"22",X"77",X"77",X"00",X"22",X"79",X"77",X"00",X"22",X"77",X"97",X"00",X"22",
		X"21",X"49",X"00",X"22",X"12",X"41",X"00",X"22",X"22",X"41",X"00",X"22",X"21",X"12",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"22",X"77",X"00",
		X"00",X"23",X"77",X"00",X"00",X"23",X"77",X"70",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"70",
		X"00",X"72",X"77",X"70",X"00",X"71",X"47",X"77",X"00",X"12",X"47",X"77",X"00",X"22",X"47",X"77",
		X"00",X"22",X"77",X"77",X"00",X"21",X"77",X"77",X"00",X"22",X"77",X"77",X"00",X"12",X"77",X"77",
		X"00",X"21",X"77",X"77",X"00",X"12",X"77",X"77",X"00",X"72",X"77",X"77",X"00",X"71",X"77",X"77",
		X"00",X"74",X"47",X"77",X"00",X"07",X"44",X"77",X"00",X"B7",X"44",X"77",X"00",X"97",X"14",X"77",
		X"00",X"94",X"14",X"47",X"99",X"71",X"22",X"99",X"9B",X"71",X"11",X"99",X"AB",X"71",X"22",X"A9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",
		X"BB",X"74",X"12",X"AA",X"9A",X"7A",X"2A",X"BA",X"AB",X"9A",X"4B",X"AB",X"9B",X"9A",X"AB",X"AC",
		X"BA",X"9A",X"BA",X"BB",X"AA",X"99",X"AA",X"BB",X"9A",X"96",X"BA",X"BA",X"A9",X"99",X"AA",X"AA",
		X"9A",X"99",X"AA",X"99",X"9A",X"99",X"AA",X"97",X"AA",X"99",X"AA",X"97",X"AB",X"A9",X"AA",X"77",
		X"BA",X"AA",X"AB",X"77",X"BB",X"9A",X"AA",X"79",X"AA",X"A9",X"BB",X"77",X"AA",X"AA",X"BB",X"74",
		X"AA",X"AA",X"CB",X"71",X"9A",X"AA",X"BB",X"71",X"99",X"79",X"BC",X"71",X"99",X"9A",X"AB",X"71",
		X"79",X"AA",X"AA",X"71",X"99",X"A9",X"AA",X"71",X"9A",X"A9",X"99",X"11",X"49",X"97",X"79",X"11",
		X"44",X"99",X"99",X"11",X"21",X"9A",X"99",X"11",X"11",X"B9",X"97",X"11",X"11",X"B9",X"97",X"11",
		X"12",X"AA",X"77",X"11",X"02",X"77",X"77",X"12",X"01",X"7A",X"14",X"12",X"01",X"9B",X"44",X"12",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"01",X"19",X"11",X"12",X"01",X"12",X"22",X"41",X"01",X"22",X"22",X"01",X"01",X"22",X"11",X"01",
		X"01",X"22",X"11",X"04",X"01",X"22",X"17",X"00",X"01",X"22",X"75",X"00",X"04",X"22",X"55",X"00",
		X"04",X"22",X"E7",X"00",X"22",X"22",X"5E",X"E0",X"22",X"77",X"E5",X"55",X"12",X"55",X"E5",X"55",
		X"21",X"55",X"75",X"55",X"12",X"4E",X"5E",X"55",X"21",X"E5",X"EE",X"75",X"21",X"56",X"5E",X"75",
		X"41",X"56",X"55",X"55",X"71",X"57",X"55",X"55",X"77",X"55",X"55",X"55",X"57",X"55",X"55",X"57",
		X"E5",X"77",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"5E",X"55",X"55",X"57",X"55",X"57",
		X"47",X"E5",X"55",X"55",X"22",X"57",X"75",X"05",X"21",X"77",X"21",X"17",X"11",X"57",X"22",X"14",
		X"12",X"77",X"22",X"14",X"22",X"77",X"22",X"14",X"22",X"11",X"22",X"14",X"22",X"14",X"22",X"14",
		X"00",X"FF",X"0D",X"D0",X"6F",X"06",X"0D",X"0D",X"F0",X"00",X"DD",X"0D",X"00",X"00",X"0D",X"0D",
		X"00",X"00",X"0D",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",X"0D",X"0D",X"06",X"00",X"0D",X"0D",
		X"06",X"00",X"0D",X"DD",X"06",X"00",X"0D",X"D0",X"06",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"DD",X"F0",X"06",X"00",X"0D",
		X"FF",X"FF",X"DD",X"0D",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"DD",X"0D",X"00",X"00",X"DD",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"0D",X"00",X"D0",X"D0",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"0D",X"00",X"00",X"D0",X"0D",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"D0",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"D0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"0D",X"00",X"00",X"D0",X"0D",X"00",X"00",X"D0",X"0D",X"00",X"00",
		X"D0",X"D0",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"DD",X"D0",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"0D",X"0D",X"00",X"00",
		X"0D",X"0D",X"00",X"00",X"D0",X"DD",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"31",X"31",X"00",
		X"00",X"11",X"11",X"00",X"00",X"13",X"13",X"00",X"03",X"13",X"13",X"00",X"03",X"13",X"13",X"00",
		X"03",X"13",X"13",X"00",X"00",X"13",X"13",X"00",X"00",X"13",X"13",X"00",X"00",X"13",X"13",X"00",
		X"03",X"11",X"11",X"00",X"03",X"31",X"31",X"00",X"03",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"00",X"33",X"31",X"03",X"00",
		X"31",X"31",X"33",X"00",X"31",X"31",X"31",X"00",X"33",X"31",X"31",X"00",X"03",X"31",X"31",X"00",
		X"00",X"33",X"31",X"00",X"00",X"00",X"31",X"00",X"03",X"33",X"31",X"00",X"33",X"31",X"31",X"00",
		X"31",X"31",X"33",X"00",X"31",X"33",X"03",X"00",X"33",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"31",X"03",X"03",X"00",
		X"31",X"33",X"33",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",
		X"33",X"31",X"31",X"00",X"00",X"31",X"31",X"00",X"33",X"31",X"31",X"00",X"31",X"31",X"31",X"00",
		X"31",X"33",X"33",X"00",X"33",X"03",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"00",X"31",X"31",X"03",X"00",
		X"31",X"31",X"33",X"00",X"31",X"31",X"31",X"00",X"03",X"31",X"31",X"00",X"00",X"31",X"31",X"00",
		X"00",X"33",X"31",X"00",X"00",X"00",X"31",X"00",X"03",X"33",X"31",X"00",X"03",X"31",X"31",X"00",
		X"03",X"31",X"33",X"00",X"03",X"33",X"03",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"13",X"30",X"30",X"30",
		X"13",X"33",X"33",X"33",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"33",X"33",X"33",X"11",X"30",X"30",X"30",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"30",X"13",X"13",X"13",X"33",
		X"13",X"11",X"33",X"13",X"13",X"11",X"30",X"11",X"13",X"11",X"33",X"11",X"13",X"11",X"13",X"11",
		X"13",X"13",X"11",X"11",X"13",X"33",X"11",X"11",X"13",X"33",X"11",X"11",X"13",X"33",X"11",X"11",
		X"13",X"33",X"13",X"13",X"11",X"11",X"33",X"33",X"33",X"33",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"30",X"30",X"13",X"13",X"33",X"33",
		X"13",X"13",X"13",X"13",X"13",X"30",X"11",X"11",X"13",X"33",X"11",X"11",X"13",X"13",X"11",X"11",
		X"13",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"13",X"11",X"11",X"11",
		X"13",X"13",X"13",X"13",X"11",X"33",X"33",X"33",X"33",X"30",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"32",X"32",X"00",
		X"00",X"22",X"22",X"00",X"00",X"23",X"23",X"00",X"03",X"23",X"23",X"00",X"03",X"23",X"23",X"00",
		X"03",X"23",X"23",X"00",X"00",X"23",X"23",X"00",X"00",X"23",X"23",X"00",X"00",X"23",X"23",X"00",
		X"03",X"22",X"22",X"00",X"03",X"32",X"32",X"00",X"03",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"00",X"33",X"32",X"03",X"00",
		X"32",X"32",X"33",X"00",X"32",X"32",X"32",X"00",X"33",X"32",X"32",X"00",X"03",X"32",X"32",X"00",
		X"00",X"33",X"32",X"00",X"00",X"00",X"32",X"00",X"03",X"33",X"32",X"00",X"33",X"32",X"32",X"00",
		X"32",X"32",X"33",X"00",X"32",X"33",X"03",X"00",X"33",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"03",X"03",X"00",
		X"32",X"33",X"33",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",
		X"33",X"32",X"32",X"00",X"00",X"32",X"32",X"00",X"33",X"32",X"32",X"00",X"32",X"32",X"32",X"00",
		X"32",X"33",X"33",X"00",X"33",X"03",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"00",X"32",X"32",X"03",X"00",
		X"32",X"32",X"33",X"00",X"32",X"32",X"32",X"00",X"03",X"32",X"32",X"00",X"00",X"32",X"32",X"00",
		X"00",X"33",X"32",X"00",X"00",X"00",X"32",X"00",X"03",X"33",X"32",X"00",X"03",X"32",X"32",X"00",
		X"03",X"32",X"33",X"00",X"03",X"33",X"03",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"30",X"30",X"30",
		X"23",X"33",X"33",X"33",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",
		X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",X"23",
		X"23",X"33",X"33",X"33",X"22",X"30",X"30",X"30",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"30",X"23",X"23",X"23",X"33",
		X"23",X"22",X"33",X"23",X"23",X"22",X"30",X"22",X"23",X"22",X"33",X"22",X"23",X"22",X"23",X"22",
		X"23",X"23",X"22",X"22",X"23",X"33",X"22",X"22",X"23",X"33",X"22",X"22",X"23",X"33",X"22",X"22",
		X"23",X"33",X"23",X"23",X"22",X"22",X"33",X"33",X"33",X"33",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"30",X"30",X"23",X"23",X"33",X"33",
		X"23",X"23",X"23",X"23",X"23",X"30",X"22",X"22",X"23",X"33",X"22",X"22",X"23",X"23",X"22",X"22",
		X"23",X"22",X"22",X"22",X"23",X"22",X"22",X"22",X"23",X"22",X"22",X"22",X"23",X"22",X"22",X"22",
		X"23",X"23",X"23",X"23",X"22",X"33",X"33",X"33",X"33",X"30",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
