library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity domino_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of domino_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",
		X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",
		X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"EA",X"C0",X"FA",X"C0",X"3E",X"C0",X"0F",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"C0",X"0F",X"C0",X"3E",X"C0",X"FA",X"FF",X"EA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"BC",X"00",X"AF",X"00",X"AB",X"C0",X"AA",X"F0",
		X"AA",X"B0",X"AA",X"B0",X"AA",X"BC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",
		X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"BC",X"AA",X"B0",X"AA",X"B0",
		X"AA",X"F0",X"AB",X"C0",X"AF",X"00",X"BC",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"FE",X"00",X"EA",X"03",X"EA",X"0F",X"AA",
		X"0E",X"AA",X"0E",X"AA",X"3E",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",
		X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3A",X"AA",X"3E",X"AA",X"0E",X"AA",X"0E",X"AA",
		X"0F",X"AA",X"03",X"EA",X"00",X"EA",X"00",X"FE",X"00",X"0F",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FC",X"FA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"FA",X"BC",X"3E",X"F0",X"0F",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"F0",X"0F",X"BC",X"3E",X"AF",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AF",X"3F",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"BF",X"00",X"AB",X"00",X"AB",X"C0",X"AA",X"F0",
		X"AA",X"B0",X"AA",X"B0",X"AA",X"BC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",
		X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"BC",X"AA",X"B0",X"AA",X"B0",
		X"AA",X"F0",X"AB",X"C0",X"AB",X"00",X"BF",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"03",X"C0",X"03",X"F0",X"0F",X"B0",X"0E",X"B0",X"0E",X"BC",X"3E",X"AC",X"3A",
		X"AF",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FE",X"BF",X"CE",X"B3",X"CE",X"B3",X"CF",X"F3",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",
		X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",
		X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"AA",X"AC",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"03",X"FF",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"FF",
		X"03",X"FF",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AB",
		X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",
		X"EA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"FF",X"C0",
		X"FF",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"FF",X"C0",X"00",X"00",
		X"00",X"00",X"C0",X"03",X"C0",X"03",X"F0",X"03",X"B0",X"03",X"BC",X"03",X"AC",X"03",X"AF",X"03",
		X"AB",X"03",X"AB",X"C3",X"AA",X"C3",X"AA",X"F3",X"AA",X"B3",X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"CE",X"AA",X"CF",X"AA",X"C3",X"AA",X"C3",X"EA",X"C0",X"EA",
		X"C0",X"FA",X"C0",X"3A",X"C0",X"3E",X"C0",X"0E",X"C0",X"0F",X"C0",X"03",X"C0",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0E",
		X"00",X"0E",X"00",X"0E",X"00",X"3E",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"FA",X"00",X"EA",
		X"00",X"EA",X"00",X"EA",X"03",X"EA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"0F",X"AA",
		X"0E",X"AA",X"3E",X"AB",X"3A",X"AB",X"3A",X"AF",X"3A",X"AC",X"3A",X"AC",X"3F",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"EA",X"AB",X"EA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"EA",X"AF",X"FA",X"AC",X"3A",X"AC",X"3A",X"BC",X"3E",X"B0",X"0E",X"B0",X"0E",X"BF",X"FE",
		X"00",X"00",X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",
		X"00",X"00",X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",
		X"00",X"00",X"2A",X"A0",X"20",X"A0",X"00",X"A0",X"2A",X"A0",X"28",X"00",X"28",X"20",X"2A",X"A0",
		X"00",X"00",X"2A",X"A0",X"20",X"A0",X"00",X"A0",X"0A",X"80",X"00",X"A0",X"20",X"A0",X"2A",X"A0",
		X"00",X"00",X"00",X"A0",X"28",X"A0",X"28",X"A0",X"2A",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",
		X"00",X"00",X"2A",X"A0",X"28",X"20",X"28",X"00",X"2A",X"A0",X"00",X"A0",X"20",X"A0",X"2A",X"A0",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A0",X"28",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"0A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"00",X"28",X"28",X"28",X"2A",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FE",X"B0",X"0E",X"F0",X"0F",
		X"C0",X"03",X"C0",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"B0",X"00",
		X"B0",X"00",X"B0",X"00",X"BC",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AF",X"00",X"AB",X"00",
		X"AB",X"00",X"AB",X"00",X"AB",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"F0",
		X"AA",X"B0",X"EA",X"BC",X"EA",X"AC",X"FA",X"AC",X"3A",X"AC",X"3A",X"AC",X"3F",X"FC",X"00",X"00",
		X"02",X"A0",X"0A",X"A8",X"08",X"88",X"28",X"0A",X"2A",X"AA",X"0A",X"A8",X"0A",X"28",X"15",X"15",
		X"00",X"00",X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"28",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A0",X"28",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"A8",X"2A",X"A0",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",X"28",X"00",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"28",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",
		X"00",X"00",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",
		X"00",X"00",X"02",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A0",X"28",X"A0",X"2A",X"A0",
		X"00",X"00",X"28",X"20",X"28",X"A0",X"2A",X"A0",X"2A",X"00",X"2A",X"A0",X"28",X"A0",X"28",X"A0",
		X"00",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"A8",X"A8",X"AA",X"A8",X"A2",X"28",X"A2",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"00",X"00",X"A0",X"28",X"A8",X"28",X"AA",X"28",X"AA",X"A8",X"A2",X"A8",X"A0",X"A8",X"A0",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"00",X"28",X"00",X"28",X"00",
		X"00",X"00",X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A2",X"A0",X"A2",X"A8",X"AA",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"A8",X"00",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"2A",X"A8",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"28",X"08",X"28",X"08",X"28",X"08",X"28",X"28",X"28",X"A0",X"2A",X"80",X"2A",X"00",
		X"00",X"00",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A2",X"28",X"A2",X"28",X"AA",X"A8",X"A8",X"A8",
		X"00",X"00",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",
		X"00",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"00",X"A0",X"02",X"80",X"0A",X"00",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F5",X"FF",X"D5",X"FF",X"54",X"FD",X"50",X"F5",X"40",X"D5",X"00",X"54",X"00",X"50",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"02",X"AA",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"AA",X"02",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",
		X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"8A",X"AA",X"80",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",
		X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",
		X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"00",X"02",X"AA",X"AA",
		X"00",X"00",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",
		X"55",X"55",X"D5",X"55",X"F5",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"F5",X"FF",X"FD",
		X"80",X"08",X"80",X"08",X"80",X"28",X"A8",X"20",X"88",X"28",X"A0",X"08",X"88",X"28",X"88",X"20",
		X"80",X"A8",X"80",X"80",X"80",X"80",X"A8",X"A8",X"88",X"88",X"A0",X"A8",X"88",X"88",X"88",X"88",
		X"08",X"0A",X"28",X"02",X"20",X"02",X"A2",X"AA",X"82",X"22",X"A2",X"22",X"22",X"02",X"A2",X"02",
		X"28",X"00",X"08",X"00",X"08",X"00",X"2A",X"A0",X"22",X"20",X"22",X"20",X"20",X"20",X"20",X"20",
		X"28",X"20",X"08",X"20",X"08",X"20",X"28",X"28",X"22",X"08",X"22",X"08",X"22",X"28",X"28",X"20",
		X"20",X"20",X"20",X"20",X"28",X"28",X"08",X"08",X"0A",X"08",X"02",X"08",X"2A",X"28",X"20",X"20",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"95",X"55",
		X"AA",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"54",X"54",X"04",X"40",X"54",X"54",X"40",X"04",X"54",X"54",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"A9",X"55",X"95",X"55",X"55",X"55",
		X"AA",X"A5",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"55",X"AA",
		X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"56",X"AA",X"55",X"6A",
		X"15",X"55",X"05",X"55",X"41",X"55",X"50",X"01",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"40",X"15",X"55",X"01",X"55",X"50",
		X"00",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"00",X"00",X"00",
		X"40",X"01",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"15",X"55",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"95",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"95",X"A9",X"55",X"55",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"AA",X"95",
		X"AA",X"95",X"A9",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AF",X"FA",X"BD",X"7F",X"F5",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"65",X"55",X"69",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"EF",X"FA",X"FD",X"7A",X"55",X"7A",
		X"55",X"7E",X"56",X"5E",X"55",X"7E",X"55",X"7A",X"55",X"7B",X"56",X"7F",X"5A",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"DF",X"EA",X"D5",X"EA",X"55",X"EA",X"57",X"EA",X"5F",X"AA",
		X"5E",X"AA",X"5E",X"AA",X"5E",X"BF",X"5F",X"B5",X"57",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"7A",X"AA",X"7E",X"FE",X"5E",X"DE",X"5F",X"DF",X"55",X"57",
		X"EA",X"AA",X"FE",X"FE",X"5E",X"DE",X"9F",X"DE",X"95",X"5E",X"55",X"7E",X"55",X"7A",X"55",X"7F",
		X"EA",X"BF",X"EA",X"F7",X"EF",X"D7",X"ED",X"55",X"FD",X"59",X"55",X"69",X"55",X"A9",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"7E",X"AA",X"5F",X"AA",X"57",X"AA",X"57",X"AA",
		X"57",X"FA",X"55",X"7A",X"55",X"FA",X"57",X"EA",X"57",X"AA",X"57",X"AA",X"57",X"FE",X"55",X"5F",
		X"EA",X"AA",X"FA",X"AA",X"7E",X"AA",X"5E",X"AA",X"5E",X"AA",X"7E",X"AA",X"7A",X"AA",X"7A",X"AA",
		X"5F",X"FE",X"55",X"5E",X"55",X"7E",X"57",X"FA",X"57",X"AA",X"57",X"EA",X"55",X"FE",X"55",X"5E",
		X"55",X"5F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"5A",X"41",X"6A",X"55",X"69",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"5A",X"41",X"6A",X"55",X"69",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"FF",
		X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AB",X"FF",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AB",X"FF",X"BF",X"FF",
		X"AA",X"AF",X"AA",X"BF",X"AB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"AF",X"FF",X"AF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",
		X"FF",X"FF",X"BF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AA",X"AF",
		X"FF",X"FF",X"AF",X"FF",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"59",X"55",X"59",X"59",X"5A",X"59",X"9A",X"5A",X"9A",X"6A",X"AA",X"6A",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"55",X"FD",X"00",X"FD",X"55",
		X"FF",X"55",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"67",X"FF",X"65",X"FF",
		X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",X"6F",X"FF",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"54",X"00",
		X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A5",X"54",
		X"95",X"50",X"55",X"40",X"55",X"00",X"54",X"00",X"54",X"00",X"54",X"05",X"95",X"56",X"9A",X"AA",
		X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"95",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AB",X"A9",X"FF",
		X"AA",X"7F",X"AA",X"7F",X"AA",X"7F",X"AA",X"5F",X"AA",X"96",X"AA",X"56",X"A9",X"45",X"A9",X"01",
		X"A5",X"01",X"A4",X"01",X"A4",X"01",X"A4",X"01",X"A4",X"01",X"A4",X"00",X"A4",X"00",X"A5",X"00",
		X"A5",X"00",X"A9",X"40",X"A9",X"40",X"AA",X"50",X"AA",X"94",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"15",X"00",X"56",X"05",X"6A",X"56",X"AA",X"6A",X"AA",X"AA",X"A9",X"AA",X"A5",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"B4",X"AA",X"F4",X"FF",X"F4",X"FF",X"F4",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"F9",X"FF",X"E9",X"EA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A5",
		X"5A",X"A9",X"15",X"A9",X"01",X"59",X"00",X"15",X"40",X"0D",X"40",X"15",X"50",X"44",X"15",X"04",
		X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"55",X"00",X"AA",X"AA",X"AA",X"AA",
		X"56",X"AA",X"55",X"AA",X"55",X"6A",X"06",X"6A",X"06",X"5A",X"06",X"9A",X"16",X"9A",X"5A",X"96",
		X"6A",X"A7",X"AA",X"A5",X"AA",X"AD",X"AA",X"AD",X"AA",X"AD",X"AA",X"BD",X"55",X"7D",X"00",X"7F",
		X"00",X"5F",X"00",X"1E",X"15",X"1E",X"55",X"1E",X"55",X"16",X"55",X"06",X"55",X"06",X"15",X"16",
		X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"55",X"05",X"40",X"14",X"00",X"10",X"00",X"50",X"00",
		X"40",X"15",X"40",X"55",X"41",X"55",X"41",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"00",X"55",
		X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"10",X"00",X"A4",X"00",X"A9",X"55",
		X"AA",X"BD",X"AA",X"DF",X"AB",X"F7",X"AD",X"FD",X"AF",X"F7",X"BD",X"DD",X"DF",X"7F",X"FD",X"FD",
		X"FF",X"7D",X"5F",X"DF",X"F7",X"F7",X"DD",X"DD",X"F7",X"F7",X"7D",X"DD",X"7F",X"7F",X"7D",X"FD",
		X"7F",X"7D",X"5F",X"DF",X"77",X"F7",X"5D",X"DD",X"77",X"F7",X"7D",X"DD",X"7F",X"7F",X"7D",X"FD",
		X"77",X"7D",X"5F",X"DF",X"77",X"F7",X"5D",X"DF",X"17",X"F7",X"05",X"00",X"01",X"40",X"00",X"40",
		X"40",X"50",X"40",X"10",X"50",X"10",X"50",X"10",X"50",X"14",X"50",X"04",X"50",X"04",X"50",X"04",
		X"40",X"04",X"00",X"14",X"00",X"10",X"00",X"50",X"00",X"40",X"01",X"40",X"15",X"00",X"50",X"00",
		X"F7",X"7A",X"FF",X"FE",X"DD",X"F7",X"5F",X"7F",X"FF",X"FD",X"FF",X"7F",X"7D",X"F7",X"F7",X"DF",
		X"7F",X"F5",X"DD",X"5F",X"FF",X"F7",X"7D",X"FF",X"D7",X"7D",X"FF",X"DF",X"FD",X"77",X"FD",X"FD",
		X"7F",X"F0",X"DD",X"71",X"FF",X"C0",X"7D",X"D1",X"D7",X"00",X"00",X"14",X"00",X"10",X"00",X"41",
		X"01",X"10",X"00",X"01",X"04",X"40",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"7A",X"AA",X"76",X"AA",X"DF",X"AA",X"7D",X"EA",
		X"DF",X"DA",X"77",X"7C",X"77",X"71",X"FD",X"C0",X"7F",X"10",X"77",X"01",X"DC",X"10",X"71",X"01",
		X"DC",X"10",X"F0",X"40",X"41",X"01",X"C0",X"00",X"C4",X"10",X"C0",X"01",X"D0",X"10",X"01",X"01",
		X"01",X"00",X"10",X"04",X"00",X"40",X"40",X"40",X"10",X"01",X"01",X"10",X"00",X"41",X"44",X"00",
		X"14",X"00",X"00",X"44",X"40",X"00",X"10",X"41",X"01",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"01",X"0A",X"10",X"12",X"00",X"00",X"41",X"10",X"00",X"00",X"04",X"04",X"10",X"40",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"02",X"AA",X"04",X"2A",X"10",X"4A",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"6A",X"AA",X"0A",X"AA",X"02",X"AA",X"10",X"AA",X"41",X"AA",
		X"01",X"04",X"40",X"00",X"00",X"11",X"04",X"00",X"00",X"10",X"10",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"11",X"00",X"04",X"00",X"40",X"40",
		X"41",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"10",X"10",X"00",X"00",X"41",X"10",X"00",X"00",X"04",X"04",X"10",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"AA",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"AA",X"80",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"A2",X"AA",X"A2",X"00",X"02",X"00",X"02",X"00",X"00",
		X"0A",X"A0",X"28",X"28",X"22",X"88",X"22",X"08",X"22",X"08",X"22",X"88",X"28",X"28",X"0A",X"A0",
		X"05",X"54",X"01",X"50",X"05",X"54",X"15",X"54",X"95",X"55",X"95",X"55",X"A5",X"55",X"29",X"54",
		X"05",X"50",X"15",X"54",X"5F",X"F5",X"57",X"F5",X"97",X"76",X"85",X"52",X"29",X"68",X"0A",X"A0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"54",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"54",X"54",X"44",X"44",X"44",X"44",X"44",X"44",X"54",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"54",X"00",X"04",X"00",X"54",X"00",X"40",X"00",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"54",X"00",X"40",X"00",X"54",X"00",X"04",X"00",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A2",X"A2",X"22",X"22",X"82",X"22",X"22",X"22",X"A2",X"A2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A2",X"22",X"22",X"22",X"22",X"22",X"22",X"20",X"22",X"A2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"02",X"AA",X"A2",X"AA",X"20",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",
		X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",
		X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",X"55",X"40",X"55",X"40",
		X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"05",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",
		X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"15",X"FF",X"05",X"7F",X"01",X"5F",X"00",X"57",
		X"00",X"15",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"15",X"FF",X"05",X"7F",X"01",X"5F",X"00",X"57",
		X"00",X"15",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"50",X"00",X"D4",X"00",X"F5",X"00",X"FD",X"40",X"FF",X"50",X"FF",X"D4",X"FF",X"F5",
		X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"54",X"FD",X"50",X"F5",X"40",X"D5",X"00",
		X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"54",X"FD",X"50",X"F5",X"40",X"D5",X"00",
		X"54",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"05",X"00",X"17",X"00",X"5F",X"01",X"7F",X"05",X"FF",X"17",X"FF",X"5F",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"15",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"54",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"50",X"00",X"10",X"00",X"14",X"00",X"04",X"00",X"05",X"00",X"01",
		X"40",X"00",X"40",X"00",X"50",X"00",X"10",X"00",X"14",X"00",X"04",X"00",X"05",X"00",X"01",X"00",
		X"01",X"40",X"00",X"40",X"00",X"50",X"00",X"10",X"00",X"14",X"00",X"04",X"00",X"05",X"00",X"01",
		X"55",X"55",X"55",X"55",X"50",X"00",X"10",X"00",X"14",X"00",X"04",X"00",X"05",X"00",X"01",X"00",
		X"00",X"00",X"15",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"05",X"00",X"04",X"00",X"14",X"00",X"10",X"00",X"50",
		X"00",X"40",X"55",X"55",X"55",X"55",X"05",X"00",X"04",X"00",X"14",X"00",X"10",X"00",X"50",X"00",
		X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"01",X"40",X"01",X"00",X"05",X"00",X"04",X"00",X"14",X"00",X"10",X"00",X"50",X"00",
		X"55",X"55",X"55",X"55",X"00",X"01",X"00",X"05",X"00",X"04",X"00",X"14",X"00",X"10",X"00",X"50",
		X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"FF",X"FF",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
