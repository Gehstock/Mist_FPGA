library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sound_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sound_prog is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"48",X"8A",X"48",X"98",X"48",X"AD",X"00",X"A0",X"48",X"F0",X"66",X"29",X"C0",X"D0",X"28",X"68",
		X"29",X"1F",X"F0",X"52",X"C5",X"13",X"90",X"4E",X"85",X"13",X"A8",X"0A",X"AA",X"B9",X"7C",X"F2",
		X"85",X"03",X"BD",X"F1",X"F2",X"85",X"05",X"E8",X"BD",X"F1",X"F2",X"85",X"06",X"A9",X"00",X"85",
		X"01",X"A2",X"FF",X"9A",X"4C",X"A6",X"F0",X"68",X"30",X"32",X"29",X"0F",X"85",X"14",X"AA",X"BD",
		X"8D",X"F2",X"85",X"04",X"BD",X"95",X"F2",X"85",X"15",X"A9",X"00",X"85",X"02",X"85",X"0E",X"85",
		X"1C",X"85",X"1A",X"A5",X"14",X"C9",X"01",X"F0",X"09",X"38",X"E9",X"06",X"B0",X"04",X"A9",X"01",
		X"85",X"1C",X"A9",X"01",X"85",X"19",X"68",X"A8",X"68",X"AA",X"68",X"40",X"E6",X"1B",X"4C",X"66",
		X"F0",X"78",X"D8",X"A2",X"FF",X"9A",X"A2",X"40",X"A9",X"00",X"95",X"01",X"CA",X"10",X"FB",X"A2",
		X"0B",X"A0",X"00",X"B9",X"9D",X"F2",X"8D",X"00",X"40",X"8D",X"00",X"80",X"C8",X"B9",X"9D",X"F2",
		X"8D",X"00",X"20",X"8D",X"00",X"60",X"C8",X"CA",X"10",X"E9",X"AD",X"00",X"A0",X"A9",X"FF",X"8D",
		X"00",X"C0",X"58",X"4C",X"A3",X"F0",X"A9",X"07",X"8D",X"00",X"40",X"A5",X"03",X"8D",X"00",X"20",
		X"A4",X"01",X"B1",X"05",X"C9",X"80",X"F0",X"1F",X"85",X"0B",X"C8",X"B1",X"05",X"85",X"0C",X"C8",
		X"B1",X"05",X"85",X"0D",X"A5",X"0B",X"8D",X"00",X"40",X"A5",X"0C",X"8D",X"00",X"20",X"C8",X"84",
		X"01",X"20",X"72",X"F2",X"4C",X"B0",X"F0",X"A2",X"00",X"86",X"13",X"BD",X"B5",X"F2",X"8D",X"00",
		X"40",X"E8",X"BD",X"B5",X"F2",X"8D",X"00",X"20",X"E8",X"E0",X"08",X"D0",X"EE",X"4C",X"A2",X"F0",
		X"48",X"8A",X"48",X"98",X"48",X"A5",X"1B",X"F0",X"06",X"20",X"54",X"F2",X"4C",X"41",X"F1",X"A5",
		X"19",X"F0",X"3E",X"A5",X"1C",X"D0",X"40",X"A5",X"1A",X"D0",X"31",X"E6",X"1A",X"A2",X"00",X"A4",
		X"15",X"B9",X"13",X"F3",X"95",X"07",X"C8",X"E8",X"E0",X"04",X"D0",X"F5",X"A9",X"07",X"8D",X"00",
		X"80",X"A5",X"04",X"8D",X"00",X"60",X"A0",X"00",X"A9",X"09",X"8D",X"00",X"80",X"B1",X"07",X"8D",
		X"00",X"60",X"A9",X"0A",X"8D",X"00",X"80",X"B1",X"09",X"8D",X"00",X"60",X"20",X"7A",X"F1",X"C6",
		X"0E",X"68",X"A8",X"68",X"AA",X"68",X"40",X"A5",X"1A",X"D0",X"27",X"E6",X"1A",X"A6",X"15",X"BD",
		X"13",X"F3",X"85",X"07",X"E8",X"BD",X"13",X"F3",X"85",X"08",X"A9",X"07",X"8D",X"00",X"80",X"A5",
		X"04",X"8D",X"00",X"60",X"A0",X"00",X"A9",X"08",X"8D",X"00",X"80",X"B1",X"07",X"85",X"17",X"8D",
		X"00",X"60",X"20",X"D0",X"F1",X"C6",X"0E",X"4C",X"41",X"F1",X"A4",X"02",X"A5",X"0E",X"D0",X"46",
		X"A6",X"14",X"BD",X"DB",X"F2",X"85",X"0E",X"C8",X"A9",X"03",X"8D",X"00",X"80",X"B1",X"07",X"C9",
		X"80",X"F0",X"39",X"C9",X"81",X"F0",X"30",X"48",X"4A",X"4A",X"4A",X"4A",X"8D",X"00",X"60",X"A9",
		X"02",X"8D",X"00",X"80",X"68",X"29",X"0F",X"AA",X"BD",X"BD",X"F2",X"8D",X"00",X"60",X"A9",X"00",
		X"8D",X"00",X"80",X"B1",X"09",X"85",X"10",X"8D",X"00",X"60",X"A9",X"04",X"8D",X"00",X"80",X"A5",
		X"10",X"8D",X"00",X"60",X"84",X"02",X"60",X"A9",X"00",X"85",X"02",X"60",X"20",X"54",X"F2",X"60",
		X"A4",X"02",X"A5",X"0E",X"D0",X"40",X"A6",X"14",X"BD",X"DB",X"F2",X"85",X"0E",X"A5",X"02",X"29",
		X"03",X"D0",X"3D",X"A9",X"08",X"8D",X"00",X"80",X"A5",X"17",X"8D",X"00",X"60",X"C8",X"A9",X"01",
		X"8D",X"00",X"80",X"B1",X"07",X"C9",X"80",X"F0",X"23",X"C9",X"81",X"F0",X"1A",X"48",X"4A",X"4A",
		X"4A",X"4A",X"8D",X"00",X"60",X"A9",X"00",X"8D",X"00",X"80",X"68",X"29",X"0F",X"AA",X"BD",X"BD",
		X"F2",X"8D",X"00",X"60",X"84",X"02",X"60",X"A9",X"00",X"85",X"02",X"60",X"20",X"54",X"F2",X"60",
		X"4A",X"B0",X"09",X"4A",X"B0",X"1A",X"4A",X"B0",X"21",X"4C",X"ED",X"F1",X"A5",X"17",X"38",X"E9",
		X"01",X"85",X"18",X"A9",X"08",X"8D",X"00",X"80",X"A5",X"18",X"8D",X"00",X"60",X"4C",X"ED",X"F1",
		X"A5",X"17",X"38",X"E9",X"02",X"85",X"18",X"4C",X"33",X"F2",X"A5",X"17",X"38",X"E9",X"04",X"85",
		X"18",X"4C",X"33",X"F2",X"A2",X"00",X"BD",X"B5",X"F2",X"8D",X"00",X"80",X"E8",X"BD",X"B5",X"F2",
		X"8D",X"00",X"60",X"E8",X"E0",X"08",X"D0",X"EE",X"A9",X"00",X"A2",X"04",X"95",X"19",X"CA",X"10",
		X"FB",X"60",X"A2",X"80",X"CA",X"D0",X"FD",X"C6",X"0D",X"D0",X"F7",X"60",X"00",X"FE",X"FE",X"FE",
		X"F7",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"F7",X"FD",X"FB",X"FB",X"00",X"F9",X"FE",
		X"FE",X"FE",X"FE",X"F9",X"FF",X"00",X"02",X"06",X"08",X"0A",X"0C",X"0E",X"12",X"00",X"00",X"01",
		X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"07",X"FF",X"08",X"00",X"09",X"00",X"0A",
		X"00",X"0E",X"00",X"0F",X"00",X"07",X"FF",X"08",X"00",X"09",X"00",X"0A",X"00",X"00",X"F5",X"BC",
		X"86",X"BC",X"24",X"F7",X"CC",X"A4",X"7E",X"5A",X"38",X"18",X"FA",X"68",X"43",X"00",X"00",X"01",
		X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"07",X"FF",X"00",X"60",X"30",X"28",X"20",
		X"18",X"40",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"07",
		X"FF",X"00",X"00",X"33",X"F3",X"67",X"F3",X"86",X"F3",X"A5",X"F3",X"3C",X"F4",X"6D",X"F4",X"9E",
		X"F4",X"CF",X"F4",X"00",X"F5",X"6A",X"F5",X"98",X"F5",X"CF",X"F5",X"F4",X"F5",X"61",X"F6",X"5B",
		X"F7",X"98",X"F7",X"00",X"00",X"C3",X"F7",X"F9",X"F7",X"2E",X"F8",X"D0",X"F8",X"72",X"F9",X"14",
		X"FA",X"B6",X"FA",X"38",X"FB",X"B9",X"FB",X"B9",X"FB",X"B9",X"FB",X"B9",X"FB",X"B9",X"FB",X"B9",
		X"FB",X"B9",X"FB",X"01",X"00",X"01",X"08",X"0F",X"01",X"00",X"2C",X"10",X"00",X"3B",X"10",X"00",
		X"2C",X"10",X"00",X"3B",X"10",X"00",X"2C",X"10",X"00",X"3B",X"10",X"00",X"37",X"10",X"00",X"3B",
		X"10",X"00",X"37",X"10",X"00",X"3B",X"10",X"00",X"37",X"10",X"00",X"3B",X"10",X"00",X"2C",X"10",
		X"00",X"3B",X"10",X"00",X"2C",X"10",X"80",X"01",X"00",X"01",X"08",X"0D",X"01",X"00",X"59",X"08",
		X"00",X"4F",X"08",X"00",X"47",X"08",X"00",X"43",X"08",X"00",X"3B",X"08",X"00",X"35",X"08",X"00",
		X"2F",X"08",X"00",X"2C",X"08",X"80",X"01",X"00",X"01",X"08",X"0D",X"01",X"00",X"2C",X"08",X"00",
		X"2F",X"08",X"00",X"35",X"08",X"00",X"3B",X"08",X"00",X"43",X"08",X"00",X"47",X"08",X"00",X"4F",
		X"08",X"00",X"59",X"08",X"80",X"06",X"09",X"08",X"08",X"0B",X"02",X"08",X"0C",X"02",X"08",X"0D",
		X"02",X"08",X"0E",X"02",X"08",X"0F",X"02",X"08",X"0E",X"02",X"08",X"0D",X"02",X"08",X"0C",X"02",
		X"08",X"0B",X"02",X"08",X"0A",X"02",X"08",X"0A",X"02",X"08",X"08",X"02",X"08",X"07",X"02",X"08",
		X"06",X"02",X"08",X"05",X"02",X"08",X"06",X"02",X"08",X"07",X"02",X"08",X"08",X"02",X"08",X"09",
		X"02",X"08",X"0A",X"02",X"08",X"0B",X"02",X"08",X"0C",X"02",X"08",X"0D",X"02",X"08",X"0E",X"02",
		X"08",X"0F",X"02",X"06",X"0C",X"08",X"08",X"0E",X"02",X"06",X"0B",X"08",X"08",X"0D",X"02",X"06",
		X"0A",X"08",X"08",X"0C",X"02",X"06",X"09",X"08",X"08",X"0B",X"02",X"06",X"08",X"08",X"08",X"0A",
		X"02",X"06",X"07",X"08",X"08",X"09",X"02",X"06",X"06",X"08",X"08",X"08",X"02",X"06",X"05",X"08",
		X"08",X"07",X"02",X"06",X"04",X"08",X"08",X"06",X"02",X"06",X"03",X"08",X"08",X"05",X"02",X"06",
		X"02",X"08",X"08",X"04",X"02",X"06",X"08",X"08",X"08",X"03",X"02",X"80",X"09",X"10",X"01",X"0C",
		X"08",X"01",X"0D",X"09",X"01",X"03",X"01",X"01",X"02",X"FA",X"20",X"02",X"F8",X"02",X"02",X"FA",
		X"20",X"02",X"FC",X"02",X"02",X"FA",X"20",X"02",X"F8",X"02",X"02",X"FA",X"20",X"02",X"FC",X"02",
		X"02",X"FF",X"02",X"02",X"FF",X"02",X"02",X"FF",X"02",X"02",X"FF",X"02",X"80",X"09",X"10",X"01",
		X"0C",X"08",X"01",X"0D",X"09",X"01",X"03",X"01",X"01",X"02",X"92",X"20",X"02",X"90",X"02",X"02",
		X"92",X"20",X"02",X"94",X"02",X"02",X"92",X"20",X"02",X"9C",X"02",X"02",X"92",X"20",X"02",X"9F",
		X"02",X"02",X"98",X"02",X"02",X"9C",X"02",X"02",X"98",X"02",X"02",X"9C",X"02",X"80",X"09",X"10",
		X"01",X"0C",X"08",X"01",X"0D",X"09",X"01",X"03",X"01",X"01",X"02",X"66",X"20",X"02",X"68",X"02",
		X"02",X"66",X"20",X"02",X"6C",X"02",X"02",X"66",X"20",X"02",X"68",X"02",X"02",X"66",X"20",X"02",
		X"6C",X"02",X"02",X"66",X"02",X"02",X"6F",X"02",X"02",X"66",X"02",X"02",X"6F",X"02",X"80",X"09",
		X"10",X"01",X"0C",X"08",X"01",X"0D",X"09",X"01",X"03",X"00",X"01",X"02",X"FA",X"20",X"02",X"F8",
		X"02",X"02",X"FA",X"20",X"02",X"FC",X"02",X"02",X"FA",X"20",X"02",X"F8",X"02",X"02",X"FA",X"20",
		X"02",X"FC",X"02",X"02",X"FF",X"02",X"02",X"FF",X"02",X"02",X"FF",X"02",X"02",X"FF",X"02",X"80",
		X"03",X"00",X"01",X"09",X"10",X"01",X"0C",X"08",X"01",X"0D",X"09",X"01",X"02",X"70",X"01",X"02",
		X"6F",X"01",X"02",X"6E",X"01",X"02",X"6D",X"01",X"02",X"6C",X"01",X"02",X"6B",X"01",X"02",X"6A",
		X"01",X"02",X"69",X"01",X"02",X"68",X"04",X"02",X"67",X"04",X"02",X"66",X"04",X"02",X"65",X"04",
		X"02",X"64",X"04",X"02",X"63",X"08",X"02",X"62",X"08",X"02",X"61",X"08",X"02",X"60",X"08",X"02",
		X"5F",X"08",X"02",X"5E",X"08",X"02",X"5D",X"08",X"02",X"5C",X"08",X"02",X"5B",X"08",X"02",X"5A",
		X"08",X"02",X"59",X"08",X"02",X"58",X"08",X"02",X"57",X"08",X"02",X"56",X"08",X"02",X"55",X"08",
		X"02",X"54",X"10",X"02",X"53",X"10",X"02",X"52",X"10",X"80",X"09",X"10",X"01",X"0C",X"08",X"01",
		X"0D",X"09",X"01",X"03",X"0F",X"01",X"02",X"FF",X"08",X"03",X"00",X"01",X"02",X"F0",X"08",X"03",
		X"0E",X"01",X"02",X"FF",X"08",X"03",X"00",X"01",X"02",X"A0",X"08",X"03",X"0D",X"01",X"02",X"FF",
		X"08",X"03",X"00",X"01",X"02",X"60",X"20",X"80",X"03",X"00",X"01",X"09",X"10",X"01",X"0C",X"08",
		X"01",X"0D",X"09",X"01",X"02",X"11",X"10",X"02",X"77",X"10",X"02",X"D5",X"10",X"02",X"49",X"10",
		X"03",X"04",X"01",X"02",X"6A",X"10",X"03",X"01",X"01",X"02",X"49",X"10",X"02",X"D5",X"10",X"02",
		X"77",X"10",X"02",X"19",X"10",X"02",X"00",X"10",X"03",X"00",X"01",X"02",X"EA",X"10",X"80",X"08",
		X"10",X"01",X"09",X"10",X"01",X"0C",X"08",X"01",X"0D",X"09",X"01",X"01",X"03",X"01",X"00",X"F5",
		X"10",X"03",X"01",X"01",X"02",X"FA",X"10",X"00",X"24",X"10",X"02",X"92",X"10",X"00",X"A4",X"10",
		X"02",X"52",X"10",X"80",X"06",X"03",X"10",X"08",X"0F",X"02",X"08",X"0E",X"02",X"08",X"0D",X"02",
		X"08",X"0C",X"02",X"08",X"0B",X"02",X"08",X"0A",X"02",X"08",X"09",X"02",X"08",X"07",X"02",X"08",
		X"06",X"02",X"08",X"07",X"02",X"08",X"08",X"02",X"06",X"0A",X"10",X"08",X"09",X"02",X"08",X"0A",
		X"10",X"08",X"0B",X"10",X"08",X"0C",X"02",X"08",X"0D",X"02",X"06",X"07",X"10",X"08",X"0C",X"02",
		X"06",X"06",X"10",X"08",X"0B",X"02",X"06",X"05",X"10",X"08",X"0A",X"02",X"06",X"04",X"10",X"08",
		X"09",X"02",X"06",X"03",X"10",X"08",X"08",X"02",X"06",X"02",X"10",X"08",X"07",X"02",X"06",X"01",
		X"02",X"08",X"06",X"02",X"08",X"05",X"02",X"08",X"04",X"02",X"08",X"03",X"02",X"08",X"02",X"02",
		X"80",X"09",X"10",X"01",X"03",X"00",X"01",X"0C",X"80",X"01",X"0D",X"09",X"01",X"02",X"3F",X"10",
		X"02",X"3D",X"10",X"02",X"3B",X"10",X"02",X"39",X"10",X"02",X"37",X"10",X"02",X"35",X"10",X"02",
		X"33",X"10",X"02",X"31",X"10",X"02",X"2F",X"10",X"02",X"2D",X"10",X"02",X"2B",X"10",X"02",X"29",
		X"10",X"02",X"27",X"10",X"02",X"25",X"10",X"02",X"23",X"10",X"02",X"21",X"10",X"02",X"1F",X"10",
		X"02",X"20",X"10",X"02",X"22",X"10",X"02",X"24",X"10",X"02",X"26",X"10",X"02",X"28",X"10",X"02",
		X"2A",X"10",X"02",X"2C",X"10",X"02",X"2E",X"10",X"02",X"30",X"10",X"02",X"32",X"10",X"02",X"34",
		X"10",X"02",X"36",X"10",X"02",X"38",X"10",X"02",X"3A",X"10",X"02",X"3C",X"10",X"02",X"3E",X"10",
		X"02",X"40",X"08",X"02",X"42",X"08",X"02",X"44",X"08",X"02",X"46",X"08",X"02",X"48",X"08",X"02",
		X"4A",X"08",X"02",X"4C",X"08",X"02",X"50",X"08",X"02",X"52",X"08",X"02",X"54",X"08",X"02",X"56",
		X"08",X"02",X"58",X"08",X"02",X"5A",X"08",X"02",X"5C",X"08",X"02",X"5E",X"08",X"02",X"60",X"04",
		X"02",X"64",X"04",X"02",X"68",X"04",X"02",X"6C",X"04",X"02",X"70",X"04",X"02",X"74",X"04",X"02",
		X"78",X"04",X"02",X"7C",X"04",X"02",X"80",X"04",X"02",X"84",X"04",X"02",X"88",X"04",X"02",X"8C",
		X"04",X"02",X"90",X"04",X"02",X"94",X"04",X"02",X"98",X"04",X"02",X"9C",X"04",X"02",X"A0",X"04",
		X"02",X"A4",X"04",X"02",X"A4",X"04",X"02",X"A8",X"04",X"02",X"AC",X"04",X"02",X"B0",X"04",X"02",
		X"B4",X"04",X"02",X"B8",X"04",X"02",X"BC",X"04",X"02",X"C0",X"04",X"02",X"C4",X"04",X"02",X"C8",
		X"04",X"02",X"CC",X"04",X"02",X"D0",X"04",X"02",X"D4",X"04",X"80",X"0A",X"0F",X"01",X"04",X"40",
		X"20",X"04",X"80",X"20",X"04",X"40",X"20",X"04",X"80",X"20",X"04",X"40",X"20",X"04",X"80",X"20",
		X"04",X"40",X"20",X"04",X"80",X"20",X"04",X"40",X"20",X"04",X"80",X"20",X"04",X"40",X"20",X"04",
		X"80",X"20",X"04",X"40",X"20",X"04",X"80",X"20",X"04",X"40",X"20",X"04",X"80",X"20",X"04",X"40",
		X"20",X"04",X"80",X"20",X"04",X"40",X"20",X"80",X"0A",X"10",X"01",X"0C",X"08",X"01",X"0D",X"09",
		X"01",X"04",X"32",X"10",X"04",X"2A",X"10",X"04",X"32",X"10",X"04",X"2A",X"10",X"04",X"32",X"10",
		X"04",X"2A",X"10",X"04",X"32",X"10",X"04",X"2A",X"10",X"04",X"32",X"10",X"04",X"2A",X"10",X"04",
		X"32",X"10",X"80",X"08",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"35",X"35",X"35",X"35",
		X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"00",X"1D",X"1D",X"2C",X"2C",X"2A",X"2A",X"28",X"28",
		X"26",X"26",X"35",X"35",X"33",X"33",X"31",X"31",X"81",X"0A",X"A9",X"C9",X"FD",X"A9",X"C9",X"FD",
		X"A9",X"C9",X"FD",X"A9",X"C9",X"FD",X"96",X"BD",X"E1",X"96",X"BD",X"E1",X"96",X"BD",X"E1",X"96",
		X"BD",X"E1",X"86",X"A9",X"C9",X"86",X"A9",X"C9",X"86",X"A9",X"C9",X"86",X"A9",X"C9",X"7E",X"7E",
		X"86",X"86",X"96",X"96",X"A9",X"A9",X"BC",X"BC",X"C9",X"C9",X"E1",X"E1",X"FD",X"FD",X"07",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"81",
		X"08",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"81",X"09",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"81",X"0A",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"21",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"81",X"08",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"00",X"00",X"26",X"26",X"00",X"00",X"35",
		X"35",X"00",X"00",X"33",X"33",X"00",X"00",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"00",X"00",X"26",X"26",X"00",X"00",X"35",
		X"35",X"00",X"00",X"33",X"33",X"00",X"00",X"81",X"08",X"7E",X"7E",X"00",X"00",X"96",X"00",X"7E",
		X"7E",X"00",X"00",X"96",X"00",X"7E",X"00",X"96",X"00",X"86",X"86",X"00",X"00",X"A9",X"00",X"86",
		X"86",X"00",X"00",X"A9",X"00",X"86",X"00",X"A9",X"00",X"96",X"96",X"00",X"00",X"BD",X"00",X"96",
		X"96",X"00",X"00",X"BD",X"00",X"96",X"00",X"BD",X"00",X"A9",X"A9",X"00",X"00",X"BD",X"BD",X"00",
		X"00",X"C9",X"C9",X"00",X"00",X"E1",X"E1",X"00",X"00",X"7E",X"7E",X"00",X"00",X"96",X"00",X"7E",
		X"7E",X"00",X"00",X"96",X"00",X"7E",X"00",X"96",X"00",X"86",X"86",X"00",X"00",X"A9",X"00",X"86",
		X"86",X"00",X"00",X"A9",X"00",X"86",X"00",X"A9",X"00",X"96",X"96",X"00",X"00",X"BD",X"00",X"96",
		X"96",X"00",X"00",X"BD",X"00",X"96",X"00",X"BD",X"00",X"A9",X"A9",X"00",X"00",X"BD",X"BD",X"00",
		X"00",X"C9",X"C9",X"00",X"00",X"E1",X"E1",X"00",X"00",X"4C",X"71",X"FC",X"78",X"D8",X"A2",X"FF",
		X"9A",X"AD",X"00",X"A0",X"A9",X"00",X"8D",X"00",X"C0",X"A0",X"00",X"A2",X"00",X"B9",X"00",X"F0",
		X"95",X"00",X"C8",X"E8",X"D0",X"F7",X"B9",X"00",X"F0",X"9D",X"00",X"01",X"C8",X"E8",X"D0",X"F6",
		X"B5",X"00",X"D9",X"00",X"F0",X"D0",X"D2",X"C8",X"E8",X"D0",X"F5",X"BD",X"00",X"01",X"D9",X"00",
		X"F0",X"D0",X"7E",X"C8",X"E8",X"D0",X"F4",X"C8",X"C0",X"20",X"D0",X"CF",X"A2",X"00",X"A0",X"00",
		X"98",X"85",X"1D",X"A9",X"02",X"85",X"1E",X"BD",X"00",X"F0",X"91",X"1D",X"E8",X"C8",X"D0",X"F7",
		X"E6",X"1E",X"A5",X"1E",X"C9",X"04",X"90",X"EF",X"A9",X"00",X"85",X"1D",X"A9",X"02",X"85",X"1E",
		X"B1",X"1D",X"DD",X"00",X"F0",X"D0",X"4A",X"E8",X"C8",X"D0",X"F5",X"E6",X"1E",X"A5",X"1E",X"C9",
		X"04",X"90",X"ED",X"E8",X"E0",X"20",X"D0",X"C6",X"A2",X"00",X"BD",X"59",X"FC",X"8D",X"00",X"40",
		X"E8",X"BD",X"59",X"FC",X"8D",X"00",X"20",X"E8",X"E0",X"18",X"D0",X"EE",X"A2",X"80",X"A0",X"00",
		X"88",X"D0",X"FD",X"CA",X"D0",X"FA",X"4C",X"71",X"F0",X"00",X"66",X"01",X"01",X"02",X"1C",X"03",
		X"01",X"04",X"EF",X"05",X"00",X"07",X"F8",X"08",X"10",X"09",X"10",X"0A",X"10",X"0C",X"30",X"0D",
		X"09",X"A0",X"00",X"B9",X"92",X"FC",X"8D",X"00",X"40",X"C8",X"B9",X"92",X"FC",X"8D",X"00",X"20",
		X"C8",X"C0",X"18",X"D0",X"EE",X"A2",X"A0",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"FA",X"4C",
		X"71",X"FC",X"00",X"CC",X"01",X"02",X"02",X"A4",X"03",X"02",X"04",X"7E",X"05",X"02",X"07",X"38",
		X"08",X"10",X"09",X"10",X"0A",X"10",X"0C",X"30",X"0D",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"BC",X"FB",X"00",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
