library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_big_sprite_tile_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_big_sprite_tile_bit2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"03",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F8",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A3",X"F8",X"F0",X"E0",X"C0",X"80",X"80",X"80",
		X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",
		X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",
		X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"80",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A0",X"80",
		X"A3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",
		X"A3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",X"A3",
		X"00",X"80",X"E0",X"F8",X"FA",X"FA",X"FA",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"1A",X"0A",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"00",X"80",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"0A",X"00",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"A3",X"A0",X"7F",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"20",X"20",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"F0",X"78",X"3C",X"3E",X"3F",X"3E",X"20",
		X"A0",X"A0",X"A3",X"A3",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"A2",X"A3",X"23",
		X"A0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"A3",X"A3",X"A3",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"01",X"FF",X"FF",X"1F",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"F8",X"FA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"7A",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"00",X"00",X"00",X"00",X"0E",X"1F",X"1F",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"FF",X"FF",X"FE",X"FC",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A2",X"A3",X"A3",X"03",X"00",X"A0",X"A2",X"A3",X"03",X"00",X"00",X"00",X"00",
		X"03",X"03",X"01",X"00",X"00",X"20",X"A0",X"A0",X"A0",X"A2",X"A3",X"A3",X"23",X"23",X"03",X"03",
		X"03",X"03",X"01",X"00",X"00",X"20",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"A0",X"23",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"00",X"80",X"E0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"1F",X"3F",X"3F",X"3F",X"1F",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"00",X"01",X"03",X"03",X"03",X"23",X"A3",X"A3",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"21",X"23",X"03",X"00",X"00",X"01",X"01",X"03",X"07",X"03",X"01",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"01",X"01",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"01",X"03",X"3F",X"0F",X"03",X"01",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A3",X"BF",X"BF",X"81",X"BF",X"BF",X"BF",X"A3",X"81",X"83",X"A3",X"A3",X"A3",X"83",X"81",X"A3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"01",X"00",X"00",X"00",X"E0",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"F8",X"FC",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"3F",X"1F",X"10",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"04",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"7E",X"40",X"40",X"40",X"00",X"7E",X"30",X"18",X"0C",X"18",X"30",X"7E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"9F",X"8F",X"87",X"C3",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"00",X"00",X"20",X"20",X"23",X"37",X"1F",X"1F",
		X"1F",X"19",X"18",X"08",X"08",X"00",X"00",X"00",X"1F",X"1F",X"0F",X"07",X"03",X"07",X"07",X"0F",
		X"01",X"03",X"47",X"6F",X"7F",X"3F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"23",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"37",
		X"47",X"6F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"E0",X"E0",X"C0",X"80",X"C0",X"71",X"10",X"F1",X"C0",X"80",X"00",X"80",X"C0",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"07",X"03",X"01",X"01",X"00",X"07",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"F9",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",
		X"83",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0C",X"0E",X"07",X"07",
		X"FF",X"FF",X"F9",X"78",X"70",X"FC",X"FC",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"E0",X"E0",X"C0",X"80",X"C0",X"FF",X"FF",
		X"FF",X"F3",X"31",X"70",X"FC",X"FC",X"F0",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"F0",X"FC",X"FC",X"70",X"31",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"00",X"00",X"00",X"00",X"00",X"F1",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"E0",X"E0",X"00",X"00",X"00",X"00",X"73",X"FB",X"FB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"03",X"03",X"03",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F0",X"E0",X"E0",X"E0",X"E0",X"00",X"03",X"03",X"07",X"7F",X"FF",X"FF",X"FF",
		X"FB",X"F3",X"C3",X"00",X"00",X"00",X"00",X"00",X"80",X"C7",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"C7",X"80",X"00",X"00",X"00",X"00",X"00",X"C3",X"F3",X"FB",
		X"8F",X"87",X"83",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"7F",X"FF",X"9F",X"9F",
		X"9F",X"9F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"83",X"87",X"8F",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"5F",X"CF",X"87",X"C0",X"40",
		X"5F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"3F",X"00",X"00",X"18",X"30",X"60",X"C7",X"8F",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"BF",X"BF",X"9F",X"CF",X"67",X"23",
		X"3F",X"3F",X"3F",X"1F",X"3F",X"7F",X"7F",X"7F",X"03",X"06",X"04",X"05",X"07",X"0F",X"1F",X"3F",
		X"FF",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"FF",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F9",X"01",
		X"81",X"81",X"81",X"FB",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"E3",X"C1",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"F1",X"01",X"F1",X"39",X"3C",X"FC",X"01",X"01",
		X"00",X"00",X"00",X"F8",X"1C",X"1C",X"1C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E8",X"F5",X"F2",X"DF",X"60",X"00",X"00",X"00",X"FF",X"F8",X"F9",X"F8",X"F9",X"F1",X"E1",X"FF",
		X"07",X"E7",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FC",X"00",X"7C",X"FE",X"FF",X"FF",X"8F",X"07",
		X"BF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"BF",
		X"91",X"51",X"F1",X"D0",X"F0",X"F3",X"E7",X"C7",X"E1",X"E1",X"FF",X"FF",X"1F",X"FF",X"37",X"51",
		X"FF",X"8F",X"03",X"01",X"01",X"81",X"C1",X"E1",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"91",X"51",X"F0",X"D0",X"F0",X"F3",X"E7",X"C7",X"C0",X"E0",X"FE",X"FF",X"1F",X"FF",X"36",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"5F",X"4F",X"87",X"01",X"03",X"0F",X"0F",X"C3",X"C7",X"C7",X"EF",X"FF",X"FF",X"BF",X"9F",
		X"FF",X"0F",X"03",X"01",X"01",X"01",X"81",X"C3",X"00",X"00",X"3C",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"FE",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",
		X"F8",X"C0",X"0C",X"3C",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"E0",X"00",X"FE",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"16",X"17",X"17",X"0F",X"07",X"03",X"00",
		X"00",X"03",X"04",X"08",X"09",X"0B",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"02",X"02",
		X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"06",X"03",X"00",X"00",X"1E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"07",X"07",X"0F",X"1F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"01",
		X"08",X"0C",X"04",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"30",X"19",X"0B",X"E7",X"3F",X"03",X"71",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"EA",X"F4",X"DF",X"60",X"00",X"00",X"00",X"0F",X"18",X"19",X"98",X"B9",X"B1",X"21",X"7F",
		X"00",X"E0",X"70",X"F0",X"F0",X"E7",X"C7",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7C",X"3C",X"18",X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"7F",X"7F",X"3F",X"7F",
		X"7F",X"3F",X"7F",X"FF",X"FF",X"7F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"18",X"3C",X"7C",X"7F",
		X"3F",X"3F",X"1F",X"1F",X"0E",X"FC",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FE",X"FE",X"FF",X"3F",X"3F",X"7F",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"1F",X"8F",X"FE",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"3F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",
		X"D1",X"43",X"43",X"80",X"00",X"03",X"0F",X"0F",X"C0",X"C0",X"C0",X"EC",X"FC",X"FC",X"B8",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C7",X"03",X"03",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"C7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0C",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"0F",X"03",X"C7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0C",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"8F",X"81",X"C1",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"F0",X"80",X"1C",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"1F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7B",X"30",X"00",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"03",X"33",X"7B",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"CE",X"8C",X"00",X"10",X"F0",X"E7",X"C3",X"83",X"82",X"82",X"C0",X"C0",X"E6",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"FE",X"FF",X"FF",X"EE",X"CC",X"80",X"00",X"E0",X"E7",X"C3",X"83",X"82",X"82",X"C0",X"C0",X"E6",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"47",X"63",X"21",X"30",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",X"4F",X"4F",
		X"67",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"60",X"C0",X"80",X"81",X"C3",
		X"43",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"9F",X"8F",X"87",X"C3",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"00",X"00",X"20",X"20",X"23",X"37",X"1F",X"1F",
		X"23",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"37",
		X"47",X"6F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"41",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"DF",X"CF",X"8F",X"87",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"10",X"30",X"30",X"3B",X"3F",
		X"FF",X"FF",X"FE",X"7C",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"66",X"FF",X"FF",
		X"F1",X"E0",X"E0",X"C0",X"80",X"C0",X"71",X"10",X"F1",X"C0",X"80",X"00",X"80",X"C0",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",
		X"C7",X"03",X"01",X"00",X"00",X"01",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"EF",X"C3",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"7C",X"FF",X"FF",X"FF",
		X"F1",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"F9",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",
		X"83",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0C",X"0E",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"E0",X"F8",X"E0",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3C",X"7E",X"7E",X"32",X"38",X"F1",X"FF",X"FF",
		X"FB",X"E3",X"C3",X"00",X"00",X"00",X"00",X"00",X"80",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"80",X"00",X"00",X"00",X"00",X"00",X"C3",X"E3",X"FB",
		X"F1",X"00",X"00",X"00",X"00",X"00",X"F1",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"E0",X"E0",X"00",X"00",X"00",X"00",X"73",X"FB",X"FB",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"03",X"03",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F8",X"F0",X"E0",X"E0",X"E0",X"00",X"03",X"03",X"07",X"7F",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
