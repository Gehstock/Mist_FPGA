library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity romf is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of romf is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7E",X"A7",X"CA",X"0E",X"10",X"C6",X"99",X"27",X"77",X"C2",X"0E",X"10",X"06",X"01",X"21",X"22",
		X"20",X"CD",X"32",X"10",X"21",X"23",X"20",X"CD",X"32",X"10",X"23",X"CD",X"32",X"10",X"23",X"CD",
		X"32",X"10",X"23",X"CD",X"32",X"10",X"23",X"CD",X"32",X"10",X"23",X"CD",X"32",X"10",X"32",X"4B",
		X"20",X"C9",X"7E",X"A7",X"CA",X"3C",X"10",X"35",X"C2",X"3C",X"10",X"37",X"78",X"17",X"47",X"C9",
		X"21",X"86",X"20",X"11",X"0B",X"00",X"19",X"E5",X"E5",X"CD",X"A6",X"10",X"E1",X"7D",X"FE",X"B2",
		X"C2",X"43",X"10",X"E1",X"CD",X"0D",X"12",X"E1",X"CD",X"0D",X"12",X"E1",X"CD",X"0D",X"12",X"E1",
		X"C3",X"0D",X"12",X"11",X"54",X"20",X"1A",X"3C",X"FE",X"03",X"C2",X"6E",X"10",X"AF",X"12",X"21",
		X"49",X"20",X"11",X"12",X"00",X"19",X"3D",X"F2",X"75",X"10",X"C9",X"7E",X"E6",X"20",X"C8",X"7E",
		X"E6",X"9F",X"77",X"01",X"06",X"00",X"09",X"11",X"33",X"20",X"CD",X"91",X"10",X"23",X"23",X"23",
		X"23",X"1A",X"13",X"77",X"23",X"1A",X"13",X"77",X"23",X"13",X"13",X"13",X"1A",X"13",X"3C",X"77",
		X"23",X"1A",X"13",X"77",X"23",X"C9",X"3A",X"0B",X"20",X"AE",X"E6",X"10",X"C0",X"7E",X"E6",X"20",
		X"C8",X"7E",X"E6",X"40",X"C2",X"B9",X"10",X"36",X"00",X"01",X"05",X"00",X"09",X"5E",X"23",X"56",
		X"23",X"EB",X"CD",X"C8",X"10",X"0E",X"1F",X"09",X"1A",X"13",X"77",X"23",X"1A",X"13",X"77",X"C9",
		X"7E",X"E6",X"20",X"C8",X"23",X"01",X"05",X"00",X"09",X"5E",X"23",X"56",X"23",X"7B",X"B2",X"C8",
		X"D5",X"5E",X"23",X"56",X"09",X"E3",X"CD",X"F6",X"10",X"E1",X"5E",X"23",X"56",X"23",X"7B",X"B2",
		X"C8",X"D5",X"5E",X"23",X"56",X"E1",X"01",X"20",X"00",X"E5",X"7B",X"36",X"00",X"23",X"3D",X"C2",
		X"FB",X"10",X"E1",X"09",X"15",X"C2",X"F9",X"10",X"C9",X"21",X"33",X"20",X"5E",X"23",X"56",X"23",
		X"7A",X"B3",X"C8",X"D5",X"7E",X"23",X"D3",X"01",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",
		X"E3",X"E6",X"08",X"CC",X"94",X"11",X"C4",X"EB",X"11",X"E1",X"C3",X"0C",X"11",X"7E",X"E6",X"40",
		X"C8",X"7E",X"E6",X"BF",X"F6",X"20",X"77",X"E6",X"08",X"47",X"23",X"23",X"5E",X"23",X"7B",X"E6",
		X"07",X"05",X"FA",X"46",X"11",X"2F",X"32",X"35",X"20",X"32",X"3C",X"20",X"56",X"23",X"CD",X"D9",
		X"11",X"EB",X"22",X"33",X"20",X"EB",X"D5",X"CD",X"B3",X"11",X"23",X"23",X"23",X"23",X"E5",X"21",
		X"36",X"20",X"CD",X"87",X"11",X"E1",X"C1",X"5E",X"23",X"7B",X"A7",X"C8",X"16",X"00",X"3E",X"05",
		X"EB",X"29",X"3D",X"C2",X"71",X"11",X"09",X"EB",X"7E",X"23",X"83",X"5F",X"EB",X"22",X"3A",X"20",
		X"EB",X"CD",X"B3",X"11",X"21",X"3D",X"20",X"73",X"23",X"72",X"23",X"71",X"23",X"70",X"23",X"AF",
		X"77",X"23",X"77",X"C9",X"C5",X"E5",X"1A",X"13",X"D3",X"02",X"DB",X"03",X"77",X"23",X"0D",X"C2",
		X"96",X"11",X"AF",X"D3",X"02",X"DB",X"03",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",
		X"94",X"11",X"C9",X"5E",X"23",X"E5",X"16",X"00",X"21",X"01",X"03",X"19",X"19",X"5E",X"23",X"56",
		X"EB",X"E3",X"5E",X"23",X"E3",X"16",X"00",X"19",X"19",X"5E",X"23",X"56",X"E1",X"EB",X"4E",X"23",
		X"46",X"23",X"EB",X"C9",X"7B",X"E6",X"07",X"D3",X"01",X"06",X"03",X"AF",X"7A",X"1F",X"57",X"7B",
		X"1F",X"5F",X"05",X"C2",X"DB",X"11",X"7A",X"C6",X"24",X"57",X"C9",X"79",X"85",X"6F",X"C5",X"E5",
		X"1A",X"13",X"D3",X"02",X"DB",X"03",X"77",X"2B",X"0D",X"C2",X"F0",X"11",X"AF",X"D3",X"02",X"DB",
		X"03",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"EE",X"11",X"C9",X"3A",X"0B",X"20",
		X"AE",X"E6",X"10",X"C0",X"7E",X"E6",X"40",X"C8",X"7E",X"F6",X"20",X"77",X"23",X"23",X"5E",X"23",
		X"23",X"56",X"23",X"CD",X"D4",X"11",X"73",X"23",X"72",X"23",X"EB",X"CD",X"32",X"12",X"01",X"1F",
		X"00",X"09",X"7E",X"12",X"13",X"3E",X"03",X"D3",X"02",X"DB",X"03",X"B6",X"77",X"23",X"7E",X"12",
		X"13",X"AF",X"D3",X"02",X"DB",X"03",X"B6",X"77",X"C9",X"F3",X"E1",X"01",X"00",X"00",X"11",X"00",
		X"00",X"31",X"20",X"40",X"3E",X"10",X"C5",X"13",X"BA",X"C2",X"56",X"12",X"31",X"00",X"24",X"E9",
		X"7E",X"A7",X"F0",X"E6",X"04",X"01",X"00",X"00",X"11",X"04",X"FC",X"CA",X"71",X"12",X"11",X"06",
		X"FA",X"23",X"7E",X"E6",X"0F",X"CA",X"A9",X"12",X"1F",X"D2",X"7D",X"12",X"42",X"1F",X"D2",X"82",
		X"12",X"43",X"1F",X"D2",X"87",X"12",X"4A",X"1F",X"D2",X"8C",X"12",X"4B",X"79",X"0E",X"00",X"23",
		X"A7",X"C4",X"D0",X"12",X"23",X"78",X"A7",X"C4",X"C6",X"12",X"2B",X"2B",X"79",X"A7",X"CA",X"A9",
		X"12",X"2B",X"7E",X"E6",X"ED",X"F6",X"60",X"77",X"C9",X"2B",X"7E",X"E6",X"02",X"C2",X"A2",X"12",
		X"54",X"5D",X"01",X"0C",X"00",X"09",X"7E",X"FE",X"08",X"C8",X"36",X"08",X"EB",X"7E",X"E6",X"10",
		X"C0",X"7E",X"F6",X"70",X"77",X"C9",X"86",X"FE",X"11",X"D8",X"FE",X"B4",X"D0",X"77",X"0C",X"C9",
		X"86",X"E5",X"F5",X"23",X"23",X"23",X"5E",X"16",X"00",X"7D",X"FE",X"60",X"21",X"60",X"1A",X"CA",
		X"E5",X"12",X"21",X"6A",X"1A",X"19",X"19",X"5E",X"23",X"56",X"F1",X"E1",X"BB",X"D8",X"BA",X"D0",
		X"77",X"0C",X"C9",X"21",X"5B",X"20",X"7E",X"A7",X"F2",X"10",X"13",X"CD",X"39",X"13",X"11",X"46",
		X"1A",X"3A",X"5C",X"20",X"CD",X"50",X"13",X"21",X"98",X"19",X"CD",X"99",X"13",X"22",X"65",X"20",
		X"21",X"6D",X"20",X"7E",X"A7",X"F2",X"2D",X"13",X"CD",X"39",X"13",X"11",X"53",X"1A",X"3A",X"6E",
		X"20",X"CD",X"50",X"13",X"21",X"A4",X"19",X"CD",X"99",X"13",X"22",X"77",X"20",X"21",X"7F",X"20",
		X"7E",X"A7",X"F0",X"CD",X"39",X"13",X"23",X"71",X"C9",X"23",X"23",X"22",X"50",X"20",X"23",X"7E",
		X"23",X"EB",X"21",X"73",X"19",X"01",X"FF",X"00",X"0C",X"BE",X"23",X"DA",X"48",X"13",X"EB",X"C9",
		X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",X"C2",X"5B",X"13",X"3E",X"01",X"77",X"23",X"F5",X"E5",X"46",
		X"71",X"CD",X"7A",X"13",X"E1",X"F1",X"11",X"08",X"00",X"42",X"19",X"71",X"FE",X"0B",X"FA",X"73",
		X"13",X"0E",X"05",X"2B",X"7E",X"A7",X"C0",X"36",X"08",X"C9",X"21",X"2C",X"1A",X"78",X"BE",X"C2",
		X"8F",X"13",X"23",X"79",X"BE",X"C2",X"90",X"13",X"1A",X"2A",X"50",X"20",X"86",X"77",X"C9",X"23",
		X"23",X"13",X"7D",X"FE",X"06",X"C2",X"7D",X"13",X"C9",X"09",X"09",X"5E",X"23",X"56",X"EB",X"C9",
		X"3A",X"43",X"20",X"A7",X"C0",X"21",X"91",X"20",X"CD",X"BD",X"13",X"21",X"9C",X"20",X"CD",X"BD",
		X"13",X"21",X"A7",X"20",X"CD",X"F0",X"13",X"21",X"B2",X"20",X"C3",X"F0",X"13",X"7E",X"A7",X"F0",
		X"CD",X"95",X"14",X"C8",X"CD",X"6C",X"14",X"FE",X"07",X"F8",X"CD",X"5A",X"14",X"FE",X"0A",X"F8",
		X"D6",X"09",X"21",X"90",X"19",X"FE",X"04",X"FA",X"A0",X"14",X"21",X"6E",X"20",X"3E",X"30",X"77",
		X"32",X"5C",X"20",X"23",X"7E",X"FE",X"DE",X"DA",X"EC",X"13",X"36",X"DE",X"AF",X"C3",X"1F",X"14",
		X"7E",X"A7",X"F0",X"CD",X"95",X"14",X"C8",X"CD",X"6C",X"14",X"FE",X"0A",X"F0",X"CD",X"5A",X"14",
		X"FE",X"07",X"F0",X"D6",X"03",X"FE",X"01",X"21",X"8A",X"19",X"F2",X"A0",X"14",X"21",X"5C",X"20",
		X"3E",X"30",X"77",X"32",X"6E",X"20",X"23",X"7E",X"FE",X"30",X"DA",X"1F",X"14",X"36",X"30",X"32",
		X"55",X"20",X"AF",X"32",X"25",X"20",X"32",X"27",X"20",X"32",X"28",X"20",X"32",X"57",X"20",X"32",
		X"58",X"20",X"32",X"22",X"20",X"3C",X"32",X"49",X"20",X"32",X"45",X"20",X"32",X"24",X"20",X"32",
		X"43",X"20",X"3A",X"0A",X"20",X"A7",X"C8",X"3E",X"04",X"32",X"26",X"20",X"3A",X"55",X"20",X"A7",
		X"3E",X"48",X"CA",X"57",X"14",X"3E",X"88",X"D3",X"03",X"C9",X"7E",X"E6",X"BF",X"77",X"11",X"07",
		X"00",X"19",X"AF",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"78",X"C9",X"E5",X"23",X"23",X"7E",
		X"E5",X"21",X"81",X"19",X"06",X"01",X"04",X"04",X"04",X"BE",X"23",X"D2",X"76",X"14",X"E1",X"23",
		X"23",X"7E",X"21",X"85",X"19",X"11",X"88",X"19",X"05",X"13",X"23",X"BE",X"DA",X"88",X"14",X"EB",
		X"96",X"4F",X"78",X"E1",X"C9",X"E5",X"11",X"07",X"00",X"19",X"7E",X"23",X"23",X"B6",X"E1",X"C9",
		X"23",X"23",X"3D",X"C2",X"A0",X"14",X"5E",X"23",X"56",X"2E",X"01",X"61",X"EB",X"C3",X"F6",X"10",
		X"21",X"86",X"20",X"11",X"0B",X"00",X"19",X"E5",X"CD",X"C3",X"14",X"E1",X"7D",X"FE",X"B2",X"C2",
		X"B3",X"14",X"C9",X"7E",X"A7",X"F0",X"23",X"23",X"7E",X"FE",X"08",X"DA",X"E4",X"14",X"FE",X"F8",
		X"D2",X"E4",X"14",X"23",X"23",X"7E",X"FE",X"10",X"DA",X"DE",X"14",X"FE",X"CC",X"D8",X"2B",X"7E",
		X"2F",X"3C",X"77",X"C9",X"2B",X"2B",X"7E",X"E6",X"BF",X"77",X"C9",X"21",X"6D",X"20",X"11",X"0D",
		X"20",X"CD",X"FA",X"14",X"21",X"5B",X"20",X"11",X"0E",X"20",X"7E",X"A7",X"F0",X"E6",X"01",X"C8",
		X"23",X"23",X"23",X"7E",X"FE",X"17",X"D0",X"AF",X"32",X"45",X"20",X"2B",X"2B",X"7E",X"E6",X"0F",
		X"F6",X"E0",X"77",X"2B",X"7E",X"E6",X"FE",X"77",X"3E",X"02",X"32",X"22",X"20",X"3A",X"0A",X"20",
		X"A7",X"C8",X"1A",X"3C",X"27",X"12",X"C3",X"24",X"1C",X"3A",X"09",X"20",X"D6",X"05",X"F8",X"C2",
		X"2C",X"15",X"2A",X"4C",X"20",X"7D",X"FE",X"20",X"D2",X"3E",X"15",X"21",X"23",X"1A",X"46",X"2B",
		X"22",X"4C",X"20",X"3A",X"5C",X"20",X"E6",X"0F",X"CA",X"4F",X"15",X"78",X"32",X"67",X"20",X"3A",
		X"6E",X"20",X"E6",X"0F",X"C8",X"78",X"32",X"79",X"20",X"C9",X"3A",X"57",X"20",X"A7",X"CA",X"70",
		X"15",X"DB",X"00",X"47",X"DB",X"00",X"21",X"20",X"20",X"11",X"B0",X"19",X"B8",X"CC",X"82",X"15",
		X"3A",X"58",X"20",X"A7",X"C8",X"DB",X"01",X"47",X"DB",X"01",X"21",X"21",X"20",X"11",X"C0",X"19",
		X"B8",X"C0",X"E5",X"2F",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"4F",X"06",X"00",X"21",X"B4",
		X"15",X"09",X"F1",X"E6",X"8F",X"B6",X"E1",X"AE",X"C8",X"4F",X"06",X"01",X"79",X"0F",X"DA",X"AA",
		X"15",X"4F",X"78",X"07",X"47",X"13",X"13",X"C3",X"9C",X"15",X"78",X"AE",X"77",X"A0",X"EB",X"4E",
		X"23",X"66",X"69",X"E9",X"30",X"70",X"40",X"50",X"20",X"50",X"60",X"10",X"21",X"5B",X"20",X"11",
		X"20",X"20",X"C3",X"CB",X"15",X"21",X"6D",X"20",X"11",X"21",X"20",X"7E",X"F6",X"02",X"77",X"1A",
		X"E6",X"7F",X"23",X"77",X"C9",X"C8",X"21",X"91",X"20",X"7E",X"A7",X"F2",X"E4",X"15",X"21",X"9C",
		X"20",X"7E",X"A7",X"F8",X"11",X"59",X"20",X"1A",X"FE",X"07",X"F0",X"D5",X"3C",X"12",X"11",X"04",
		X"00",X"19",X"E5",X"21",X"28",X"1E",X"11",X"A2",X"3E",X"CD",X"30",X"01",X"21",X"5F",X"20",X"5E",
		X"16",X"00",X"2B",X"E5",X"21",X"CC",X"19",X"06",X"18",X"3A",X"0A",X"20",X"A7",X"CA",X"18",X"16",
		X"78",X"D3",X"03",X"3E",X"04",X"32",X"26",X"20",X"19",X"19",X"19",X"19",X"5E",X"23",X"56",X"23",
		X"4E",X"23",X"46",X"E1",X"7E",X"80",X"47",X"2B",X"7E",X"81",X"4F",X"E1",X"70",X"2B",X"72",X"2B",
		X"71",X"2B",X"73",X"2B",X"36",X"C0",X"D1",X"1A",X"FE",X"06",X"C0",X"3C",X"12",X"13",X"7B",X"FE",
		X"5A",X"CA",X"46",X"16",X"1B",X"1B",X"06",X"0A",X"3A",X"11",X"20",X"A7",X"CA",X"51",X"16",X"06",
		X"05",X"1A",X"FE",X"06",X"FA",X"59",X"16",X"06",X"02",X"78",X"32",X"25",X"20",X"32",X"4A",X"20",
		X"C9",X"C8",X"21",X"A7",X"20",X"7E",X"A7",X"F2",X"70",X"16",X"21",X"B2",X"20",X"7E",X"A7",X"F8",
		X"11",X"5A",X"20",X"1A",X"FE",X"07",X"F0",X"D5",X"3C",X"12",X"11",X"04",X"00",X"19",X"E5",X"21",
		X"28",X"1E",X"11",X"B8",X"3E",X"CD",X"30",X"01",X"21",X"71",X"20",X"5E",X"16",X"00",X"2B",X"E5",
		X"21",X"E8",X"19",X"06",X"28",X"C3",X"09",X"16",X"21",X"0C",X"20",X"DB",X"02",X"2F",X"47",X"DB",
		X"02",X"2F",X"B8",X"C0",X"E6",X"40",X"47",X"AE",X"C8",X"70",X"78",X"A7",X"C8",X"3E",X"0C",X"D3",
		X"03",X"01",X"64",X"00",X"D3",X"04",X"05",X"C2",X"B4",X"16",X"0D",X"C2",X"B4",X"16",X"3E",X"08",
		X"D3",X"03",X"21",X"12",X"20",X"34",X"21",X"BA",X"1D",X"CD",X"87",X"1C",X"3A",X"0A",X"20",X"A7",
		X"C0",X"21",X"E7",X"1A",X"22",X"06",X"20",X"31",X"00",X"24",X"C3",X"7E",X"0F",X"3A",X"44",X"20",
		X"A7",X"C8",X"11",X"08",X"20",X"01",X"29",X"20",X"CD",X"44",X"1C",X"21",X"29",X"20",X"11",X"0F",
		X"24",X"3E",X"02",X"C3",X"30",X"01",X"21",X"7F",X"20",X"7E",X"A7",X"F0",X"23",X"23",X"23",X"7E",
		X"FE",X"17",X"D2",X"08",X"17",X"3E",X"B6",X"77",X"EB",X"21",X"72",X"19",X"01",X"77",X"19",X"23",
		X"03",X"BE",X"DA",X"0F",X"17",X"EB",X"0A",X"2B",X"77",X"C9",X"21",X"4B",X"20",X"7E",X"A7",X"C8",
		X"36",X"00",X"1F",X"F5",X"DC",X"54",X"17",X"F1",X"1F",X"F5",X"DC",X"A8",X"17",X"F1",X"1F",X"F5",
		X"DC",X"4F",X"17",X"F1",X"1F",X"F5",X"DC",X"49",X"18",X"F1",X"1F",X"F5",X"DC",X"8A",X"18",X"F1",
		X"1F",X"DC",X"1B",X"19",X"1F",X"F5",X"DC",X"10",X"19",X"F1",X"1F",X"DC",X"23",X"19",X"C9",X"3E",
		X"08",X"D3",X"03",X"C9",X"21",X"13",X"20",X"06",X"08",X"7E",X"07",X"07",X"07",X"AE",X"17",X"17",
		X"21",X"13",X"20",X"7E",X"17",X"77",X"23",X"7E",X"17",X"77",X"05",X"C2",X"59",X"17",X"F6",X"02",
		X"E6",X"1F",X"32",X"28",X"20",X"E6",X"07",X"4F",X"06",X"00",X"21",X"74",X"1A",X"09",X"46",X"21",
		X"5E",X"20",X"7E",X"FE",X"A0",X"DA",X"8A",X"17",X"06",X"01",X"FE",X"18",X"D2",X"91",X"17",X"06",
		X"02",X"2B",X"7E",X"FE",X"38",X"DA",X"9A",X"17",X"06",X"04",X"FE",X"10",X"D2",X"A1",X"17",X"06",
		X"08",X"2B",X"7E",X"E6",X"F0",X"B0",X"77",X"C9",X"3A",X"09",X"20",X"F6",X"20",X"32",X"27",X"20",
		X"AF",X"CD",X"C2",X"17",X"32",X"5F",X"20",X"21",X"5C",X"20",X"7E",X"E6",X"0F",X"B0",X"77",X"C3",
		X"D5",X"15",X"F5",X"21",X"5D",X"20",X"4E",X"23",X"5E",X"21",X"6F",X"20",X"46",X"23",X"56",X"CD",
		X"EF",X"17",X"C6",X"14",X"21",X"7A",X"1A",X"23",X"23",X"BE",X"23",X"DA",X"D7",X"17",X"F1",X"A7",
		X"CA",X"E4",X"17",X"23",X"7E",X"4F",X"17",X"17",X"17",X"17",X"E6",X"F0",X"47",X"79",X"C9",X"7A",
		X"93",X"C8",X"5F",X"9F",X"57",X"21",X"00",X"00",X"3E",X"06",X"19",X"3D",X"C2",X"FA",X"17",X"7C");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
