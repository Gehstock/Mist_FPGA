library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"05",X"00",X"22",X"00",X"40",X"C3",X"0B",X"02",X"D3",X"80",X"78",X"D3",X"40",X"CA",X"FF",X"FF",
		X"C3",X"B7",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"7C",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"C7",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"3C",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"60",X"01",X"3D",X"FF",X"CA",X"FF",X"FF",X"08",X"DA",X"22",X"6E",X"00",X"E6",X"3D",X"0D",
		X"CE",X"C2",X"01",X"B7",X"28",X"2B",X"57",X"FD",X"FF",X"20",X"02",X"C7",X"E5",X"0F",X"4F",X"79",
		X"AA",X"28",X"07",X"7A",X"B7",X"28",X"03",X"79",X"18",X"3E",X"79",X"E5",X"0F",X"20",X"38",X"79",
		X"C5",X"11",X"07",X"07",X"07",X"CB",X"7F",X"28",X"2D",X"CB",X"BF",X"18",X"13",X"DA",X"08",X"FB",
		X"CA",X"05",X"05",X"22",X"40",X"40",X"77",X"23",X"10",X"FC",X"3D",X"07",X"05",X"3F",X"CF",X"CA",
		X"CE",X"E5",X"00",X"D0",X"CE",X"8C",X"00",X"AF",X"77",X"23",X"77",X"CA",X"47",X"22",X"3D",X"40",
		X"12",X"01",X"00",X"1A",X"10",X"FE",X"CA",X"31",X"45",X"40",X"CE",X"E5",X"00",X"D8",X"CE",X"E5",
		X"00",X"38",X"38",X"39",X"40",X"40",X"CE",X"01",X"02",X"47",X"39",X"41",X"40",X"CE",X"01",X"02",
		X"4F",X"39",X"44",X"40",X"CE",X"01",X"02",X"31",X"4A",X"40",X"39",X"45",X"40",X"CE",X"01",X"02",
		X"5F",X"22",X"4A",X"40",X"55",X"78",X"BA",X"38",X"02",X"7A",X"B9",X"38",X"02",X"79",X"BB",X"D0",
		X"1D",X"02",X"B8",X"28",X"06",X"1C",X"BA",X"28",X"02",X"1C",X"7B",X"CE",X"8C",X"00",X"39",X"45",
		X"40",X"77",X"23",X"35",X"00",X"CA",X"0D",X"02",X"22",X"40",X"40",X"BD",X"28",X"0D",X"0C",X"23",
		X"23",X"BD",X"28",X"08",X"0C",X"23",X"23",X"BD",X"28",X"01",X"AF",X"CA",X"23",X"35",X"00",X"7A",
		X"37",X"CA",X"22",X"83",X"01",X"5F",X"15",X"00",X"1A",X"7D",X"CA",X"70",X"23",X"7C",X"D5",X"44",
		X"20",X"FA",X"FA",X"3E",X"31",X"80",X"41",X"EE",X"55",X"12",X"3F",X"00",X"CE",X"6E",X"01",X"3D",
		X"08",X"05",X"00",X"CF",X"3D",X"0A",X"CF",X"3D",X"09",X"CF",X"3D",X"07",X"05",X"3F",X"CF",X"22",
		X"00",X"60",X"21",X"4D",X"40",X"77",X"FB",X"22",X"3F",X"40",X"34",X"3D",X"0F",X"CE",X"C2",X"01",
		X"E5",X"08",X"20",X"F7",X"3D",X"0F",X"CE",X"C2",X"01",X"E5",X"08",X"28",X"F7",X"F3",X"3D",X"02",
		X"31",X"4B",X"40",X"22",X"42",X"40",X"7D",X"2B",X"B7",X"28",X"30",X"7D",X"CE",X"E8",X"02",X"FB",
		X"00",X"00",X"00",X"F3",X"22",X"4B",X"40",X"34",X"22",X"43",X"40",X"7D",X"2B",X"B7",X"28",X"22",
		X"7D",X"CE",X"E8",X"02",X"FB",X"00",X"00",X"00",X"F3",X"22",X"4B",X"40",X"34",X"22",X"46",X"40",
		X"7D",X"2B",X"B7",X"28",X"11",X"7D",X"CE",X"E8",X"02",X"18",X"AB",X"7D",X"CE",X"DA",X"02",X"18",
		X"CD",X"7D",X"CE",X"DA",X"02",X"18",X"DE",X"7D",X"CE",X"DA",X"02",X"18",X"9A",X"87",X"5F",X"15",
		X"00",X"1A",X"5D",X"23",X"55",X"EB",X"EA",X"9C",X"01",X"0F",X"03",X"BE",X"03",X"5E",X"04",X"81",
		X"14",X"66",X"14",X"9E",X"0B",X"8E",X"04",X"67",X"0B",X"7F",X"07",X"8B",X"07",X"8D",X"07",X"B0",
		X"09",X"C4",X"09",X"8C",X"0B",X"16",X"10",X"EB",X"05",X"3B",X"0B",X"53",X"0B",X"5E",X"0B",X"00",
		X"00",X"06",X"06",X"23",X"10",X"C3",X"06",X"3E",X"05",X"22",X"A7",X"02",X"CE",X"9E",X"02",X"39",
		X"4B",X"40",X"CE",X"8C",X"00",X"23",X"77",X"CA",X"B7",X"C8",X"22",X"26",X"01",X"E6",X"22",X"F3",
		X"02",X"18",X"A9",X"33",X"00",X"33",X"03",X"D1",X"03",X"76",X"04",X"8C",X"14",X"71",X"14",X"A7",
		X"0B",X"A9",X"04",X"8F",X"0B",X"92",X"07",X"97",X"07",X"9E",X"07",X"BE",X"09",X"C7",X"09",X"95",
		X"0B",X"25",X"10",X"0D",X"07",X"4C",X"0B",X"55",X"0B",X"60",X"0B",X"00",X"00",X"1C",X"06",X"2E",
		X"10",X"E6",X"06",X"62",X"05",X"B7",X"C8",X"CE",X"9C",X"01",X"39",X"4B",X"40",X"C3",X"84",X"00",
		X"39",X"4B",X"40",X"E5",X"03",X"C8",X"C5",X"07",X"05",X"00",X"CF",X"CA",X"39",X"4B",X"40",X"3E",
		X"87",X"47",X"CE",X"0A",X"03",X"04",X"78",X"D3",X"80",X"7C",X"D3",X"40",X"CA",X"39",X"4B",X"40",
		X"3E",X"87",X"47",X"D3",X"80",X"DB",X"40",X"6F",X"04",X"78",X"D3",X"80",X"DB",X"40",X"67",X"CA",
		X"12",X"04",X"7F",X"39",X"4B",X"40",X"47",X"CB",X"01",X"CB",X"03",X"10",X"F9",X"3D",X"07",X"D3",
		X"80",X"39",X"4C",X"40",X"A1",X"B3",X"31",X"4C",X"40",X"D3",X"40",X"CA",X"39",X"4B",X"40",X"C5",
		X"07",X"CF",X"CA",X"00",X"06",X"09",X"0E",X"18",X"07",X"0D",X"0C",X"05",X"16",X"14",X"13",X"10",
		X"0F",X"04",X"15",X"03",X"11",X"12",X"01",X"0A",X"08",X"02",X"15",X"17",X"39",X"4B",X"40",X"47",
		X"3D",X"84",X"07",X"10",X"FE",X"5F",X"15",X"FF",X"CE",X"6E",X"01",X"CE",X"30",X"01",X"18",X"17",
		X"12",X"80",X"FB",X"18",X"AD",X"CF",X"CA",X"39",X"4B",X"40",X"E5",X"03",X"C8",X"C5",X"07",X"18",
		X"00",X"D3",X"80",X"DB",X"40",X"47",X"CA",X"02",X"00",X"00",X"12",X"FF",X"FC",X"39",X"4B",X"40",
		X"FD",X"01",X"28",X"16",X"38",X"08",X"15",X"F3",X"CB",X"00",X"CB",X"00",X"18",X"0B",X"12",X"3F",
		X"FF",X"CB",X"38",X"CB",X"1A",X"CB",X"38",X"CB",X"1A",X"29",X"4D",X"40",X"7C",X"A1",X"B0",X"67",
		X"7E",X"A3",X"B2",X"6F",X"21",X"4D",X"40",X"77",X"CA",X"02",X"00",X"03",X"C3",X"C9",X"01",X"02",
		X"00",X"02",X"18",X"C5",X"02",X"00",X"01",X"18",X"C2",X"D3",X"80",X"7E",X"D3",X"40",X"CA",X"E7",
		X"3D",X"20",X"22",X"60",X"40",X"77",X"3D",X"03",X"23",X"77",X"3D",X"14",X"23",X"77",X"3D",X"02",
		X"23",X"77",X"AF",X"23",X"77",X"22",X"10",X"00",X"21",X"66",X"40",X"2D",X"20",X"EF",X"F7",X"05",
		X"0A",X"DF",X"CA",X"39",X"64",X"40",X"A7",X"28",X"0E",X"FD",X"02",X"28",X"1F",X"FD",X"03",X"38",
		X"2B",X"28",X"4A",X"C3",X"72",X"05",X"22",X"60",X"40",X"36",X"20",X"6F",X"35",X"20",X"D7",X"3E",
		X"28",X"04",X"47",X"DF",X"18",X"66",X"22",X"64",X"40",X"34",X"18",X"F5",X"22",X"00",X"03",X"21",
		X"67",X"40",X"EF",X"05",X"08",X"DF",X"22",X"64",X"40",X"34",X"18",X"4F",X"22",X"62",X"40",X"36",
		X"20",X"4A",X"35",X"03",X"CE",X"4E",X"01",X"B7",X"12",X"08",X"00",X"EE",X"51",X"EF",X"22",X"61",
		X"40",X"36",X"20",X"37",X"35",X"14",X"22",X"64",X"40",X"34",X"18",X"2F",X"22",X"63",X"40",X"36",
		X"20",X"1E",X"35",X"02",X"B7",X"29",X"67",X"40",X"12",X"20",X"00",X"EE",X"51",X"21",X"67",X"40",
		X"EF",X"29",X"66",X"40",X"2B",X"7E",X"B4",X"20",X"0B",X"22",X"64",X"40",X"34",X"18",X"0C",X"29",
		X"67",X"40",X"18",X"EC",X"21",X"66",X"40",X"22",X"64",X"40",X"36",X"AF",X"CA",X"3D",X"80",X"31",
		X"5E",X"40",X"05",X"0D",X"CE",X"7C",X"01",X"22",X"70",X"00",X"CE",X"3C",X"01",X"F7",X"CE",X"04",
		X"03",X"CA",X"39",X"5E",X"40",X"3E",X"31",X"5E",X"40",X"28",X"26",X"FD",X"FF",X"28",X"39",X"FD",
		X"20",X"38",X"09",X"FD",X"30",X"38",X"0C",X"FD",X"70",X"38",X"01",X"AF",X"CA",X"05",X"00",X"CE",
		X"7C",X"01",X"CA",X"22",X"3C",X"00",X"CE",X"3C",X"01",X"05",X"0B",X"CE",X"7C",X"01",X"AF",X"CA",
		X"CE",X"04",X"03",X"3D",X"80",X"31",X"5D",X"40",X"05",X"09",X"CE",X"7C",X"01",X"22",X"FC",X"00",
		X"CE",X"3C",X"01",X"F7",X"AF",X"31",X"5E",X"40",X"CA",X"39",X"5D",X"40",X"3E",X"31",X"5D",X"40",
		X"FD",X"42",X"38",X"0B",X"CE",X"4E",X"01",X"2E",X"2E",X"EF",X"AF",X"31",X"5E",X"40",X"CA",X"FD",
		X"40",X"28",X"0D",X"B7",X"28",X"12",X"CE",X"4E",X"01",X"2C",X"2C",X"EF",X"AF",X"31",X"5E",X"40",
		X"CA",X"D7",X"06",X"DF",X"C3",X"33",X"04",X"D7",X"06",X"28",X"0F",X"DF",X"22",X"00",X"00",X"CE",
		X"3C",X"01",X"3D",X"80",X"31",X"5D",X"40",X"C3",X"1A",X"04",X"3D",X"FF",X"CA",X"CE",X"C7",X"01",
		X"CE",X"60",X"01",X"22",X"00",X"02",X"CE",X"3C",X"01",X"05",X"09",X"CE",X"7C",X"01",X"22",X"90",
		X"01",X"21",X"30",X"42",X"CA",X"29",X"30",X"42",X"2B",X"21",X"30",X"42",X"7C",X"B6",X"3D",X"FF",
		X"C8",X"CE",X"4E",X"01",X"12",X"03",X"00",X"1A",X"CE",X"3C",X"01",X"AF",X"CA",X"E7",X"3D",X"08",
		X"31",X"70",X"42",X"3D",X"0C",X"31",X"72",X"42",X"3D",X"10",X"31",X"71",X"42",X"AF",X"31",X"73",
		X"42",X"22",X"50",X"00",X"EF",X"F7",X"05",X"00",X"DF",X"CA",X"39",X"73",X"42",X"A7",X"28",X"17",
		X"FD",X"02",X"28",X"22",X"FD",X"03",X"38",X"21",X"28",X"2C",X"22",X"71",X"42",X"36",X"3D",X"FF",
		X"C8",X"AF",X"31",X"73",X"42",X"AF",X"CA",X"D7",X"3C",X"FD",X"0E",X"20",X"04",X"22",X"73",X"42",
		X"34",X"47",X"DF",X"18",X"F0",X"CE",X"EB",X"04",X"18",X"EB",X"D7",X"3E",X"20",X"04",X"22",X"73",
		X"42",X"34",X"47",X"DF",X"18",X"DF",X"CE",X"F8",X"04",X"18",X"D9",X"22",X"70",X"42",X"36",X"C0",
		X"3D",X"08",X"77",X"22",X"73",X"42",X"34",X"CA",X"22",X"72",X"42",X"36",X"C0",X"3D",X"0C",X"77",
		X"22",X"73",X"42",X"34",X"CA",X"CE",X"04",X"03",X"22",X"00",X"02",X"21",X"75",X"42",X"F7",X"05",
		X"05",X"DF",X"3D",X"08",X"31",X"76",X"42",X"AF",X"31",X"78",X"42",X"CA",X"39",X"78",X"42",X"FD",
		X"02",X"28",X"34",X"FD",X"01",X"28",X"48",X"FD",X"03",X"28",X"6A",X"FD",X"04",X"28",X"75",X"22",
		X"76",X"42",X"36",X"20",X"15",X"35",X"08",X"12",X"F0",X"FF",X"29",X"75",X"42",X"1A",X"21",X"75",
		X"42",X"7C",X"A7",X"20",X"06",X"7E",X"FD",X"38",X"38",X"03",X"EF",X"AF",X"CA",X"3D",X"20",X"31",
		X"76",X"42",X"44",X"3D",X"02",X"18",X"11",X"22",X"76",X"42",X"36",X"20",X"ED",X"35",X"06",X"3D",
		X"03",X"22",X"60",X"00",X"05",X"01",X"21",X"75",X"42",X"31",X"78",X"42",X"DF",X"AF",X"CA",X"22",
		X"76",X"42",X"36",X"20",X"D5",X"35",X"05",X"12",X"FC",X"FF",X"29",X"75",X"42",X"1A",X"21",X"75",
		X"42",X"7C",X"A7",X"20",X"C6",X"7E",X"FD",X"30",X"30",X"C0",X"3D",X"30",X"31",X"76",X"42",X"44",
		X"3D",X"03",X"18",X"D6",X"22",X"76",X"42",X"36",X"20",X"B2",X"35",X"04",X"3D",X"04",X"22",X"60",
		X"00",X"05",X"04",X"18",X"C2",X"22",X"76",X"42",X"36",X"20",X"A0",X"35",X"04",X"12",X"10",X"00",
		X"29",X"75",X"42",X"1A",X"21",X"75",X"42",X"7C",X"A7",X"28",X"8F",X"7E",X"FD",X"80",X"38",X"89",
		X"C3",X"06",X"06",X"AF",X"22",X"10",X"42",X"77",X"23",X"35",X"04",X"23",X"35",X"04",X"23",X"35",
		X"04",X"23",X"35",X"68",X"CE",X"B0",X"01",X"3D",X"05",X"05",X"18",X"CF",X"05",X"04",X"CE",X"7C",
		X"01",X"CE",X"C7",X"01",X"CA",X"CE",X"1C",X"05",X"CE",X"EE",X"06",X"AF",X"CA",X"39",X"10",X"42",
		X"CB",X"47",X"28",X"10",X"22",X"11",X"42",X"36",X"C0",X"35",X"04",X"05",X"00",X"CE",X"7C",X"01",
		X"0D",X"02",X"18",X"10",X"22",X"12",X"42",X"36",X"C0",X"35",X"04",X"39",X"13",X"42",X"47",X"CE",
		X"7C",X"01",X"0D",X"02",X"39",X"10",X"42",X"AA",X"31",X"10",X"42",X"CA",X"22",X"14",X"42",X"36",
		X"C0",X"35",X"68",X"22",X"13",X"42",X"39",X"10",X"42",X"CB",X"4F",X"20",X"0A",X"34",X"3D",X"07",
		X"BD",X"0D",X"01",X"28",X"DF",X"CA",X"36",X"7D",X"3C",X"C0",X"E2",X"3E",X"CA",X"E7",X"3D",X"20",
		X"22",X"E0",X"42",X"77",X"3D",X"03",X"23",X"77",X"3D",X"14",X"23",X"77",X"3D",X"02",X"23",X"77",
		X"23",X"35",X"00",X"22",X"10",X"00",X"21",X"E6",X"42",X"2D",X"20",X"EF",X"F7",X"05",X"0A",X"DF",
		X"CA",X"39",X"E4",X"42",X"A7",X"28",X"1C",X"FD",X"02",X"28",X"1F",X"FD",X"03",X"38",X"2B",X"28",
		X"4A",X"D7",X"3E",X"28",X"04",X"47",X"DF",X"AF",X"CA",X"AF",X"31",X"A6",X"41",X"3E",X"CA",X"47",
		X"DF",X"18",X"65",X"22",X"E4",X"42",X"34",X"AF",X"18",X"F6",X"22",X"00",X"03",X"21",X"E7",X"42",
		X"EF",X"05",X"08",X"DF",X"22",X"E4",X"42",X"34",X"18",X"4F",X"22",X"E2",X"42",X"36",X"20",X"4A",
		X"35",X"03",X"CE",X"4E",X"01",X"B7",X"12",X"08",X"00",X"EE",X"51",X"EF",X"22",X"E1",X"42",X"36",
		X"20",X"37",X"35",X"14",X"22",X"E4",X"42",X"34",X"18",X"2F",X"22",X"E3",X"42",X"36",X"20",X"1E",
		X"35",X"02",X"B7",X"29",X"E7",X"42",X"12",X"20",X"00",X"EE",X"51",X"21",X"E7",X"42",X"EF",X"29",
		X"E6",X"42",X"2B",X"7E",X"B4",X"20",X"0B",X"22",X"E4",X"42",X"34",X"18",X"0C",X"29",X"E7",X"42",
		X"18",X"EC",X"21",X"E6",X"42",X"22",X"E4",X"42",X"36",X"AF",X"CA",X"22",X"50",X"00",X"21",X"80",
		X"42",X"22",X"24",X"0A",X"21",X"81",X"42",X"3D",X"00",X"31",X"84",X"42",X"05",X"0E",X"CE",X"7C",
		X"01",X"22",X"50",X"00",X"CE",X"3C",X"01",X"CE",X"60",X"01",X"CE",X"C7",X"01",X"CA",X"29",X"80",
		X"42",X"2B",X"21",X"80",X"42",X"7C",X"B6",X"3D",X"00",X"28",X"47",X"39",X"84",X"42",X"CB",X"47",
		X"3D",X"00",X"28",X"0D",X"22",X"81",X"42",X"36",X"C0",X"35",X"24",X"05",X"0E",X"CE",X"7C",X"01",
		X"18",X"26",X"CE",X"4E",X"01",X"12",X"09",X"00",X"39",X"84",X"42",X"CB",X"4F",X"28",X"04",X"AF",
		X"EE",X"51",X"3D",X"1A",X"CE",X"3C",X"01",X"0D",X"01",X"CE",X"5A",X"07",X"22",X"83",X"42",X"36",
		X"C0",X"35",X"0A",X"47",X"CE",X"7C",X"01",X"0D",X"02",X"39",X"84",X"42",X"AA",X"31",X"84",X"42",
		X"AF",X"CA",X"22",X"84",X"42",X"CB",X"55",X"20",X"0D",X"CE",X"EB",X"05",X"05",X"00",X"CE",X"7C",
		X"01",X"22",X"84",X"42",X"CB",X"D5",X"CA",X"05",X"00",X"CE",X"7C",X"01",X"3D",X"FF",X"CA",X"E7",
		X"AF",X"31",X"C8",X"41",X"31",X"A3",X"41",X"F7",X"C3",X"62",X"0A",X"E7",X"F7",X"CA",X"E7",X"F7",
		X"CA",X"DE",X"22",X"80",X"41",X"18",X"09",X"DE",X"22",X"88",X"41",X"18",X"04",X"DE",X"22",X"90",
		X"41",X"DE",X"7D",X"00",X"FD",X"FF",X"28",X"06",X"CE",X"B7",X"07",X"AF",X"CA",X"AF",X"31",X"A6",
		X"41",X"31",X"A5",X"41",X"3D",X"FF",X"CA",X"DE",X"36",X"02",X"C0",X"39",X"A1",X"41",X"DE",X"77",
		X"02",X"DE",X"CB",X"00",X"45",X"C1",X"D6",X"07",X"DE",X"7D",X"07",X"D5",X"02",X"F9",X"D6",X"07",
		X"DE",X"77",X"07",X"47",X"DF",X"DE",X"36",X"00",X"C0",X"DE",X"6D",X"01",X"DE",X"65",X"03",X"7D",
		X"47",X"E5",X"1F",X"C9",X"69",X"08",X"FD",X"1F",X"C1",X"84",X"08",X"23",X"DE",X"76",X"01",X"DE",
		X"74",X"03",X"78",X"E5",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",X"05",X"00",X"22",X"06",X"08",X"0A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
