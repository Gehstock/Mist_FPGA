library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity terrain_2b is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of terrain_2b is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"19",X"1C",X"1F",X"20",X"19",X"1A",X"1B",X"1C",X"1E",X"10",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"08",X"00",X"07",X"00",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"0A",X"0B",
		X"0A",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",
		X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",
		X"07",X"08",X"0A",X"11",X"0A",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",
		X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",
		X"07",X"08",X"07",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"14",X"1A",X"1D",X"19",X"1C",X"1F",X"19",
		X"1A",X"1D",X"20",X"1B",X"1C",X"1D",X"1E",X"19",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"11",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"2B",X"09",X"00",X"00",X"15",X"1B",X"1E",X"1A",X"1D",X"20",X"1A",
		X"1B",X"1E",X"1A",X"1C",X"1D",X"1E",X"1F",X"1D",X"2D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0E",X"0B",
		X"0E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"0E",X"11",X"0E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"64",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"64",X"09",X"00",X"00",X"15",X"1C",X"1F",X"1B",X"1E",X"19",X"1B",
		X"1C",X"1F",X"1B",X"20",X"19",X"1A",X"19",X"10",X"02",X"02",X"02",X"02",X"02",X"02",X"0C",X"04",
		X"0F",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"10",X"0B",
		X"10",X"02",X"04",X"63",X"0C",X"04",X"0F",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"10",X"11",X"10",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"63",X"2C",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"61",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"15",X"1D",X"20",X"1C",X"1F",X"1A",X"1C",
		X"1D",X"20",X"1C",X"1A",X"1B",X"1E",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"0A",X"00",X"09",X"13",X"00",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"28",X"11",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"22",X"1E",X"19",X"1D",X"20",X"1B",X"1D",
		X"1E",X"19",X"1D",X"1C",X"19",X"1C",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"0A",X"00",X"09",X"13",X"00",X"00",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"03",X"21",X"1F",X"1A",X"1E",X"19",X"1C",X"1E",
		X"1F",X"1A",X"1E",X"1B",X"20",X"1F",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"0A",X"00",X"09",X"13",X"00",X"00",X"00",X"03",X"04",X"03",X"13",X"16",X"1C",X"1C",X"1B",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"09",X"03",X"03",X"11",X"20",X"1B",X"1F",X"1A",X"1D",X"1F",
		X"20",X"1B",X"1F",X"19",X"1A",X"1C",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"0A",X"00",X"09",X"13",X"00",X"00",X"00",X"00",X"03",X"04",X"03",X"12",X"1F",X"1A",X"1C",X"1E",
		X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"64",X"04",X"03",X"00",X"13",X"19",X"1C",X"20",X"1B",X"1E",X"20",
		X"19",X"1C",X"20",X"1E",X"1C",X"1D",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"0A",X"00",X"09",X"63",X"14",X"14",X"14",X"14",X"14",X"0F",X"04",X"17",X"12",X"19",X"1B",X"1D",
		X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"23",X"24",X"00",X"5F",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"5E",X"01",
		X"01",X"01",X"01",X"01",X"2B",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"5E",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"64",X"04",X"03",X"00",X"00",X"19",X"1A",X"1D",X"19",X"1C",X"1F",X"19",
		X"1A",X"1D",X"1C",X"1D",X"1E",X"1B",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"02",
		X"02",X"02",X"02",X"02",X"0F",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0E",X"0B",
		X"0E",X"01",X"04",X"13",X"00",X"00",X"00",X"03",X"04",X"04",X"04",X"16",X"00",X"1B",X"1C",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"26",X"26",X"01",X"04",X"01",X"01",X"01",X"01",X"04",X"01",X"01",X"04",X"04",X"04",
		X"5E",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"0C",
		X"01",X"01",X"01",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"15",X"1B",X"1E",X"1A",X"1D",X"20",X"1A",
		X"1B",X"1E",X"1D",X"1C",X"1F",X"1E",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"01",
		X"01",X"01",X"01",X"01",X"01",X"04",X"2C",X"02",X"02",X"02",X"02",X"02",X"0F",X"0C",X"10",X"0B",
		X"10",X"02",X"04",X"13",X"00",X"00",X"03",X"04",X"03",X"00",X"16",X"04",X"17",X"08",X"00",X"00",
		X"00",X"00",X"00",X"61",X"5E",X"01",X"01",X"04",X"0C",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"63",X"02",X"25",X"25",X"02",X"5F",X"00",X"00",X"00",X"00",X"5F",X"67",X"5F",X"5F",X"5E",X"04",
		X"5E",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"1C",X"1F",X"1B",X"1E",X"19",X"1B",
		X"1C",X"1F",X"1E",X"1D",X"20",X"1F",X"11",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"0A",X"0B",
		X"28",X"00",X"09",X"63",X"02",X"0C",X"04",X"03",X"00",X"00",X"17",X"04",X"16",X"07",X"00",X"00",
		X"00",X"00",X"61",X"64",X"64",X"02",X"02",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"00",X"24",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"67",X"61",X"5F",
		X"5E",X"04",X"5E",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"17",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"1D",X"20",X"1C",X"1F",X"1A",X"1C",
		X"1D",X"20",X"1F",X"19",X"1E",X"20",X"11",X"00",X"00",X"00",X"00",X"03",X"04",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"20",X"0B",
		X"21",X"00",X"09",X"04",X"01",X"01",X"04",X"5E",X"5F",X"00",X"00",X"16",X"04",X"17",X"00",X"00",
		X"00",X"61",X"64",X"64",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"00",X"0B",X"2B",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"1C",X"12",X"1B",X"1F",X"65",
		X"61",X"5F",X"5E",X"04",X"5E",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"19",X"1D",X"20",X"1B",X"1D",
		X"1E",X"19",X"20",X"1F",X"1A",X"1D",X"14",X"00",X"00",X"00",X"03",X"04",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"21",
		X"11",X"00",X"09",X"09",X"00",X"00",X"5F",X"5E",X"04",X"04",X"04",X"04",X"04",X"16",X"00",X"00",
		X"5F",X"64",X"64",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"27",X"11",X"28",X"00",X"00",X"00",X"00",X"1B",X"16",X"1D",X"19",X"1B",X"1D",X"1F",X"1E",
		X"65",X"5F",X"00",X"5F",X"5E",X"04",X"5E",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"63",X"02",X"02",X"02",X"02",X"02",X"02",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"1E",X"19",X"1C",X"1E",
		X"1F",X"1A",X"1D",X"1E",X"1B",X"20",X"24",X"01",X"01",X"01",X"04",X"04",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"04",X"09",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"28",
		X"11",X"0A",X"09",X"09",X"00",X"00",X"00",X"00",X"5F",X"02",X"02",X"02",X"64",X"04",X"0C",X"5E",
		X"04",X"64",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"61",
		X"13",X"28",X"11",X"27",X"00",X"00",X"00",X"12",X"19",X"1D",X"19",X"1F",X"1D",X"1A",X"20",X"1F",
		X"1D",X"1F",X"67",X"5F",X"00",X"5F",X"5E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"5E",X"5F",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"1F",X"1A",X"1D",X"1F",
		X"20",X"1B",X"1E",X"1F",X"1C",X"1E",X"23",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"04",X"09",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"0A",
		X"11",X"0A",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"04",X"04",X"04",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"61",X"23",X"21",X"00",X"00",X"00",X"19",X"1D",X"20",X"1C",X"20",X"1E",X"1C",X"19",X"1F",X"1E",
		X"1C",X"1D",X"1A",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"5E",X"04",X"5E",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"1D",X"20",X"1B",X"1E",X"20",
		X"1F",X"1C",X"1D",X"1E",X"19",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"01",X"01",X"01",X"01",X"01",X"2B",X"01",X"01",X"0E",
		X"11",X"0E",X"04",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"04",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"18",
		X"00",X"24",X"28",X"00",X"00",X"17",X"16",X"1C",X"1F",X"1B",X"1F",X"1D",X"1B",X"20",X"1E",X"1D",
		X"1B",X"1C",X"20",X"16",X"1F",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"5E",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"7F",X"19",X"1C",X"1F",X"19",
		X"1E",X"1D",X"1A",X"1C",X"1A",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"64",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"63",X"10",
		X"11",X"10",X"63",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"04",X"64",
		X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"61",
		X"27",X"11",X"27",X"00",X"00",X"10",X"1E",X"1B",X"1E",X"1A",X"1E",X"1C",X"1A",X"1F",X"1D",X"1C",
		X"1A",X"1B",X"1F",X"1A",X"1C",X"1E",X"67",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"1A",X"1D",X"20",X"1A",
		X"1D",X"1E",X"19",X"1F",X"1B",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"64",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",
		X"28",X"34",X"12",X"16",X"16",X"1B",X"1D",X"1A",X"1D",X"19",X"1D",X"1B",X"20",X"1E",X"1C",X"1B",
		X"19",X"1A",X"1E",X"19",X"1B",X"1E",X"12",X"68",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",
		X"14",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"1B",X"1E",X"19",X"1B",
		X"1C",X"1F",X"1A",X"1E",X"1C",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"04",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"00",
		X"21",X"35",X"1D",X"20",X"1D",X"1A",X"1C",X"19",X"1C",X"20",X"1C",X"1A",X"1F",X"1D",X"1B",X"1A",
		X"20",X"19",X"1D",X"20",X"1A",X"1D",X"1B",X"10",X"1F",X"68",X"00",X"00",X"00",X"5F",X"67",X"1F",
		X"1C",X"1F",X"67",X"67",X"67",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"20",X"1C",X"1F",X"1A",X"1C",
		X"1B",X"20",X"1C",X"1B",X"1D",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"17",X"04",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"22",
		X"11",X"36",X"1C",X"1F",X"1C",X"19",X"1B",X"20",X"1B",X"1F",X"1B",X"19",X"1E",X"82",X"86",X"88",
		X"8A",X"20",X"1C",X"1F",X"19",X"1C",X"1A",X"1F",X"19",X"1E",X"14",X"67",X"67",X"5F",X"12",X"1D",
		X"20",X"1B",X"10",X"1B",X"1C",X"1F",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"19",X"1D",X"20",X"1B",X"1D",
		X"1A",X"1E",X"1D",X"19",X"1E",X"12",X"00",X"00",X"12",X"04",X"04",X"64",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"16",X"04",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"18",X"61",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"19",X"1B",X"56",X"57",X"21",
		X"34",X"19",X"1B",X"1E",X"1B",X"20",X"1A",X"1F",X"1A",X"1E",X"1A",X"20",X"1D",X"83",X"04",X"04",
		X"8B",X"1F",X"8A",X"88",X"86",X"82",X"19",X"1E",X"1D",X"1C",X"10",X"1B",X"1C",X"16",X"1D",X"1C",
		X"1F",X"1A",X"1C",X"1B",X"1F",X"1A",X"1E",X"14",X"14",X"67",X"14",X"5F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"1A",X"1E",X"19",X"1C",X"1E",
		X"19",X"1D",X"1F",X"1B",X"1F",X"10",X"00",X"00",X"16",X"04",X"04",X"04",X"17",X"00",X"00",X"00",
		X"00",X"00",X"17",X"04",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"04",X"0C",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"0C",
		X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"17",X"1C",X"16",X"1A",X"20",X"75",X"53",X"37",X"11",
		X"35",X"20",X"1A",X"1D",X"1A",X"1F",X"19",X"1E",X"19",X"1D",X"19",X"1F",X"1C",X"84",X"04",X"04",
		X"8C",X"1E",X"8B",X"04",X"04",X"83",X"20",X"1D",X"1C",X"20",X"1D",X"1B",X"1A",X"1E",X"1C",X"1B",
		X"1E",X"19",X"1B",X"1A",X"1E",X"19",X"1B",X"19",X"1C",X"16",X"1C",X"1F",X"14",X"67",X"62",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1B",X"1F",X"1A",X"1D",X"1F",
		X"20",X"1C",X"19",X"1A",X"20",X"15",X"00",X"00",X"04",X"04",X"04",X"04",X"12",X"00",X"00",X"00",
		X"00",X"00",X"18",X"04",X"01",X"01",X"04",X"01",X"01",X"01",X"17",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"04",X"2B",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"64",X"0C",X"04",X"64",X"17",X"1C",X"1C",X"16",X"1C",X"75",X"53",X"04",X"04",X"55",X"36",X"11",
		X"36",X"1F",X"19",X"1C",X"19",X"1E",X"20",X"1D",X"20",X"1C",X"20",X"1E",X"1B",X"85",X"87",X"89",
		X"8D",X"1D",X"8C",X"04",X"04",X"84",X"1F",X"1C",X"85",X"87",X"89",X"8D",X"20",X"1D",X"1B",X"1A",
		X"1D",X"20",X"1A",X"19",X"1D",X"20",X"1A",X"20",X"82",X"86",X"88",X"8A",X"1D",X"19",X"1F",X"65",
		X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"20",X"1B",X"1E",X"20",
		X"1F",X"1B",X"1C",X"1D",X"19",X"10",X"00",X"00",X"64",X"04",X"04",X"04",X"12",X"00",X"00",X"00",
		X"00",X"03",X"04",X"03",X"00",X"00",X"62",X"02",X"02",X"64",X"16",X"00",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"2C",X"61",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",X"07",X"08",
		X"00",X"00",X"51",X"52",X"16",X"20",X"1C",X"1F",X"1B",X"7C",X"04",X"04",X"04",X"7C",X"36",X"11",
		X"37",X"1E",X"20",X"1B",X"20",X"1D",X"1F",X"1C",X"1F",X"1B",X"1F",X"1D",X"1A",X"20",X"1E",X"1D",
		X"1B",X"1C",X"8D",X"89",X"87",X"85",X"1E",X"1B",X"84",X"04",X"04",X"8C",X"1F",X"1C",X"1A",X"19",
		X"1C",X"1F",X"19",X"20",X"1C",X"1F",X"19",X"1F",X"83",X"04",X"04",X"8B",X"1C",X"20",X"1D",X"12",
		X"1F",X"67",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"1F",X"19",
		X"1E",X"1A",X"19",X"1C",X"1A",X"16",X"17",X"00",X"13",X"04",X"04",X"04",X"64",X"14",X"14",X"14",
		X"0C",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"04",X"03",X"00",X"00",X"0D",X"0A",
		X"11",X"0A",X"13",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",
		X"1C",X"1C",X"16",X"19",X"1C",X"1F",X"1B",X"1E",X"1A",X"7C",X"04",X"04",X"53",X"75",X"37",X"34",
		X"19",X"1D",X"1F",X"1A",X"1F",X"1C",X"1E",X"1B",X"1E",X"1A",X"1E",X"1C",X"19",X"1F",X"1D",X"1C",
		X"1A",X"1B",X"1F",X"1A",X"1C",X"1F",X"1D",X"1A",X"83",X"04",X"04",X"8B",X"1E",X"1B",X"19",X"20",
		X"1B",X"1E",X"20",X"1F",X"1B",X"1E",X"20",X"1E",X"84",X"04",X"04",X"8C",X"1B",X"1F",X"1C",X"20",
		X"16",X"17",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"1D",X"20",X"1A",
		X"1D",X"20",X"1E",X"19",X"1B",X"1F",X"16",X"17",X"61",X"02",X"02",X"5F",X"08",X"08",X"07",X"18",
		X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"0C",X"02",X"63",X"10",
		X"11",X"10",X"63",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"16",X"1E",
		X"1A",X"1C",X"1E",X"20",X"1B",X"1E",X"1A",X"1D",X"20",X"54",X"53",X"73",X"75",X"1C",X"32",X"34",
		X"1F",X"1C",X"1E",X"19",X"70",X"73",X"73",X"73",X"74",X"74",X"73",X"70",X"20",X"1E",X"1C",X"1B",
		X"19",X"1A",X"1E",X"19",X"1B",X"1E",X"1C",X"19",X"82",X"86",X"88",X"8A",X"1D",X"1A",X"20",X"1F",
		X"1A",X"1D",X"1F",X"1E",X"1A",X"1D",X"1F",X"1D",X"85",X"87",X"89",X"8D",X"1A",X"1E",X"1B",X"1F",
		X"1A",X"1C",X"16",X"1F",X"65",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"1E",X"1F",X"1B",
		X"1C",X"1F",X"1A",X"20",X"1C",X"19",X"1D",X"12",X"00",X"00",X"07",X"08",X"07",X"07",X"61",X"64",
		X"16",X"00",X"00",X"17",X"1C",X"17",X"1B",X"1C",X"1B",X"00",X"00",X"03",X"01",X"01",X"01",X"0E",
		X"11",X"0E",X"2B",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"16",X"20",X"1D",X"1F",
		X"19",X"1B",X"1D",X"1F",X"1A",X"1D",X"19",X"77",X"7B",X"73",X"75",X"1A",X"19",X"32",X"46",X"45",
		X"33",X"31",X"30",X"30",X"46",X"45",X"5A",X"5D",X"5A",X"5A",X"5D",X"5B",X"74",X"70",X"1B",X"1A",
		X"20",X"19",X"50",X"70",X"73",X"73",X"73",X"73",X"70",X"50",X"20",X"1E",X"1C",X"19",X"1F",X"1E",
		X"19",X"1C",X"1E",X"1D",X"19",X"1C",X"1E",X"1C",X"1F",X"1D",X"20",X"1C",X"19",X"1D",X"1A",X"1E",
		X"19",X"1B",X"1D",X"1E",X"1E",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"1E",X"1C",
		X"1B",X"1E",X"19",X"1B",X"1D",X"1A",X"1B",X"1C",X"28",X"64",X"02",X"02",X"02",X"02",X"64",X"64",
		X"61",X"00",X"00",X"15",X"1C",X"19",X"1E",X"1C",X"1A",X"12",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"11",X"0A",X"13",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"1C",X"19",X"1D",X"19",X"1D",
		X"1D",X"20",X"1A",X"77",X"75",X"75",X"76",X"73",X"75",X"19",X"1C",X"20",X"59",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"5A",X"5B",X"5C",X"5C",
		X"5C",X"5B",X"5D",X"5A",X"5A",X"5B",X"5C",X"5B",X"5D",X"5B",X"74",X"70",X"1B",X"1F",X"1E",X"1C",
		X"20",X"1A",X"19",X"1B",X"20",X"1B",X"20",X"1D",X"1C",X"19",X"1C",X"1E",X"1D",X"1C",X"20",X"1D",
		X"1D",X"19",X"20",X"1C",X"13",X"17",X"17",X"00",X"00",X"00",X"00",X"00",X"19",X"20",X"1D",X"1D",
		X"1A",X"1D",X"1F",X"1A",X"1E",X"19",X"20",X"1F",X"27",X"5E",X"01",X"01",X"01",X"04",X"5E",X"61",
		X"00",X"00",X"00",X"1A",X"1B",X"20",X"1D",X"1B",X"19",X"1E",X"1C",X"1C",X"17",X"00",X"00",X"0A",
		X"11",X"0A",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"1D",X"1B",X"20",X"1C",X"20",X"1C",
		X"1B",X"1C",X"78",X"75",X"77",X"77",X"1D",X"20",X"1E",X"1F",X"1B",X"59",X"52",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"5A",X"5D",X"5B",X"74",X"70",X"1B",
		X"1F",X"1C",X"1D",X"20",X"1F",X"1A",X"19",X"1B",X"1F",X"1E",X"1B",X"1D",X"20",X"1D",X"1F",X"1C",
		X"1E",X"1A",X"1D",X"1B",X"11",X"00",X"6B",X"00",X"00",X"00",X"00",X"00",X"12",X"19",X"1C",X"1E",
		X"19",X"1C",X"1A",X"19",X"1F",X"1A",X"1B",X"1C",X"15",X"00",X"00",X"00",X"61",X"16",X"00",X"00",
		X"00",X"00",X"00",X"10",X"1A",X"1F",X"1C",X"1A",X"20",X"1D",X"1B",X"19",X"1D",X"12",X"00",X"27",
		X"11",X"0A",X"0D",X"00",X"00",X"00",X"00",X"00",X"18",X"1F",X"1C",X"1A",X"1F",X"1B",X"1F",X"1B",
		X"1F",X"1E",X"79",X"1B",X"19",X"1F",X"1C",X"19",X"1D",X"59",X"53",X"54",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"5A",X"5D",X"5B",
		X"74",X"73",X"74",X"01",X"74",X"73",X"70",X"1A",X"19",X"1F",X"1A",X"1F",X"1C",X"19",X"1E",X"1B",
		X"1F",X"1B",X"1E",X"10",X"00",X"00",X"17",X"03",X"00",X"00",X"00",X"11",X"1F",X"1A",X"1B",X"1F",
		X"1A",X"20",X"1B",X"1E",X"20",X"1F",X"1D",X"1E",X"10",X"00",X"00",X"5F",X"6A",X"61",X"00",X"00",
		X"00",X"00",X"00",X"15",X"19",X"1E",X"1B",X"19",X"1F",X"1C",X"1A",X"20",X"1C",X"1A",X"00",X"00",
		X"24",X"28",X"12",X"17",X"00",X"00",X"00",X"00",X"10",X"1E",X"1B",X"19",X"1E",X"1A",X"1E",X"1A",
		X"19",X"75",X"7A",X"1E",X"1D",X"20",X"1B",X"57",X"58",X"52",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"5A",X"5D",X"5D",X"5D",X"5A",X"5A",X"5B",X"74",X"73",X"70",X"19",X"20",X"1B",X"20",X"1D",X"1A",
		X"20",X"1C",X"16",X"17",X"00",X"00",X"00",X"03",X"17",X"00",X"00",X"12",X"20",X"1B",X"1A",X"20",
		X"1B",X"1E",X"1F",X"1D",X"19",X"1E",X"1C",X"1F",X"2A",X"14",X"5E",X"5E",X"61",X"00",X"00",X"00",
		X"00",X"00",X"00",X"17",X"16",X"1D",X"1A",X"20",X"1E",X"1B",X"19",X"1F",X"1B",X"16",X"00",X"00",
		X"23",X"21",X"2E",X"65",X"5F",X"00",X"00",X"19",X"1A",X"1D",X"1A",X"20",X"1D",X"75",X"73",X"71",
		X"75",X"7A",X"75",X"20",X"1F",X"1C",X"59",X"4F",X"51",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"5A",X"5D",X"5B",X"74",X"70",X"1B",X"1C",X"19",
		X"70",X"71",X"51",X"00",X"00",X"5F",X"14",X"14",X"16",X"00",X"14",X"1B",X"1A",X"1C",X"19",X"19",
		X"1C",X"1F",X"20",X"1C",X"1A",X"1D",X"20",X"19",X"29",X"14",X"5F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1B",X"16",X"1F",X"1D",X"1A",X"20",X"1E",X"1A",X"1E",X"10",X"00",
		X"22",X"11",X"29",X"00",X"5F",X"67",X"02",X"5F",X"19",X"1C",X"19",X"1F",X"75",X"7B",X"75",X"19",
		X"77",X"75",X"1D",X"19",X"57",X"58",X"4F",X"4F",X"4E",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"5A",X"5B",X"74",X"73",X"72",
		X"5F",X"00",X"5F",X"14",X"14",X"5F",X"00",X"00",X"5F",X"5E",X"25",X"1F",X"1B",X"1D",X"20",X"1A",
		X"1D",X"20",X"1A",X"19",X"1B",X"1C",X"1E",X"1A",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"16",X"19",X"1F",X"1D",X"19",X"1D",X"1F",X"11",
		X"00",X"29",X"11",X"29",X"00",X"00",X"5F",X"5E",X"7D",X"1B",X"20",X"1E",X"7C",X"75",X"1D",X"20",
		X"1A",X"1B",X"57",X"58",X"50",X"50",X"50",X"50",X"4D",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"4F",X"60",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1B",X"20",X"1C",X"1E",X"1F",X"1B",
		X"1E",X"19",X"1B",X"20",X"1C",X"19",X"1B",X"1F",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"1B",X"12",X"20",X"1C",X"1E",X"12",
		X"00",X"00",X"29",X"11",X"29",X"00",X"14",X"1B",X"7D",X"7D",X"1E",X"1D",X"79",X"20",X"1C",X"1F",
		X"20",X"56",X"47",X"47",X"47",X"47",X"47",X"47",X"48",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"52",X"4F",X"60",
		X"5E",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",X"19",X"1D",X"1F",X"1E",X"1B",
		X"1F",X"1A",X"1C",X"1B",X"1D",X"20",X"1A",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"32",X"32",X"32",X"32",X"32",X"32",X"3A",X"37",X"18",X"1F",X"1B",X"1D",X"1A",
		X"12",X"1B",X"17",X"29",X"11",X"22",X"15",X"1A",X"1F",X"70",X"76",X"76",X"75",X"1F",X"1B",X"1E",
		X"55",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"4C",X"49",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"49",X"49",X"49",X"4C",X"50",X"50",
		X"50",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1A",X"1E",X"20",X"1D",X"1A",
		X"20",X"1B",X"1D",X"1A",X"1E",X"1F",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"40",X"34",X"34",X"35",X"35",X"35",X"39",X"36",X"11",X"1E",X"1A",X"1C",X"20",
		X"1A",X"1F",X"1C",X"10",X"29",X"21",X"14",X"19",X"1E",X"1A",X"1D",X"20",X"1B",X"1E",X"1A",X"56",
		X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"4B",X"49",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"47",X"47",X"47",X"47",X"47",X"47",
		X"47",X"04",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"1B",X"1F",X"19",X"1C",X"19",
		X"19",X"1C",X"1E",X"19",X"1F",X"1E",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"3D",X"3F",X"44",X"35",X"35",X"35",X"34",X"36",X"13",X"1D",X"19",X"1B",X"1F",
		X"19",X"1E",X"1B",X"1A",X"00",X"29",X"29",X"14",X"1D",X"19",X"1C",X"1F",X"1A",X"1D",X"19",X"47",
		X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"48",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"49",X"49",X"47",X"47",X"47",X"47",X"47",X"47",
		X"47",X"04",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"1A",X"1B",X"20",
		X"1A",X"1D",X"1F",X"1D",X"20",X"1D",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"3B",X"3C",X"35",X"35",X"35",X"34",X"36",X"19",X"1C",X"20",X"1A",X"1E",
		X"20",X"1D",X"1A",X"15",X"00",X"00",X"21",X"29",X"12",X"20",X"1B",X"10",X"10",X"1C",X"56",X"47",
		X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"4C",X"49",X"49",X"49",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"4A",X"4A",X"47",X"47",X"47",X"47",X"47",X"47",
		X"47",X"04",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"26",X"19",X"1B",X"1A",X"1F",
		X"1B",X"1E",X"20",X"1C",X"19",X"1C",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"3D",X"3C",X"3B",X"35",X"35",X"35",X"38",X"36",X"15",X"1B",X"1F",X"19",X"1D",
		X"1F",X"1C",X"19",X"19",X"00",X"00",X"22",X"11",X"29",X"1B",X"1B",X"48",X"59",X"58",X"47",X"47",
		X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"4A",X"4A",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"49",X"47",X"47",X"47",X"47",X"47",X"47",
		X"47",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"5E",X"03",X"15",X"1A",X"1C",X"19",X"1E",
		X"1C",X"1F",X"19",X"1F",X"1A",X"1B",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"33",X"34",X"35",X"35",X"35",X"39",X"36",X"19",X"1A",X"1E",X"20",X"1C",
		X"1E",X"1B",X"20",X"00",X"00",X"00",X"00",X"29",X"2A",X"44",X"44",X"2A",X"5A",X"5B",X"5C",X"47",
		X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"48",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"49",X"49",X"47",X"47",X"47",X"47",X"47",X"47",X"47",
		X"47",X"16",X"00",X"00",X"00",X"00",X"5F",X"5E",X"5E",X"5F",X"00",X"15",X"1B",X"1D",X"20",X"1D",
		X"1D",X"20",X"1A",X"1E",X"1B",X"1F",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"33",X"34",X"35",X"35",X"35",X"39",X"36",X"00",X"1A",X"1D",X"1F",X"1B",
		X"1D",X"16",X"1B",X"00",X"00",X"00",X"00",X"00",X"45",X"45",X"48",X"40",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"45",X"46",X"45",X"46",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",
		X"2F",X"17",X"00",X"00",X"5F",X"5E",X"5E",X"5F",X"00",X"00",X"00",X"15",X"1C",X"1E",X"1F",X"1C",
		X"1E",X"19",X"1C",X"1B",X"1C",X"19",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"33",X"34",X"35",X"35",X"35",X"39",X"36",X"00",X"17",X"16",X"19",X"1A",
		X"1B",X"00",X"00",X"00",X"A5",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"40",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"46",X"45",X"46",X"45",X"46",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"47",X"47",X"47",X"47",X"47",X"2F",
		X"04",X"5E",X"5E",X"5E",X"02",X"5F",X"00",X"00",X"00",X"00",X"13",X"1D",X"1D",X"1F",X"1E",X"1B",
		X"1F",X"1A",X"1D",X"1A",X"1D",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"33",X"34",X"35",X"35",X"35",X"39",X"36",X"00",X"00",X"00",X"1B",X"1C",
		X"00",X"00",X"A5",X"A6",X"A0",X"A0",X"A6",X"A7",X"A5",X"00",X"00",X"00",X"00",X"00",X"48",X"48",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"52",X"4F",X"4F",X"60",X"04",
		X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1C",X"1E",X"20",X"1D",X"1A",
		X"20",X"1B",X"1F",X"19",X"1E",X"1C",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"33",X"34",X"35",X"35",X"35",X"39",X"36",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A4",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A7",X"A5",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"52",X"4F",X"4F",X"60",X"03",X"03",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1B",X"1D",X"1F",X"1C",X"19",
		X"19",X"1C",X"19",X"20",X"1F",X"1D",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"3D",X"3F",X"35",X"35",X"35",X"38",X"36",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A5",X"00",X"00",
		X"00",X"00",X"00",X"45",X"47",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"45",X"45",X"54",X"53",X"4F",X"4F",X"60",X"03",X"00",X"00",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"1A",X"1C",X"1E",X"1B",X"20",
		X"1A",X"1D",X"1A",X"1E",X"20",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"42",X"34",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"00",X"00",
		X"A1",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A8",
		X"A9",X"00",X"00",X"00",X"00",X"00",X"40",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",
		X"46",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",
		X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"52",X"4F",X"6C",X"6D",X"6E",X"5F",X"00",X"00",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1E",X"19",X"1B",X"1D",X"1A",X"1F",
		X"1B",X"1E",X"1B",X"1D",X"19",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"3B",X"43",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"00",X"A2",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A6",X"A5",X"00",X"00",X"00",X"00",X"41",X"42",X"46",X"44",X"43",X"45",X"48",X"48",X"45",
		X"47",X"45",X"48",X"45",X"49",X"4A",X"48",X"45",X"47",X"43",X"44",X"46",X"45",X"46",X"45",X"46",
		X"45",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"47",X"43",X"43",X"47",X"43",
		X"43",X"47",X"47",X"43",X"43",X"47",X"6F",X"6E",X"14",X"5F",X"00",X"1B",X"16",X"10",X"1B",X"1B",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"1D",X"20",X"1A",X"1C",X"19",X"1E",
		X"1C",X"1F",X"1D",X"1C",X"1A",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"34",X"3B",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"00",X"A3",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A6",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4B",X"4C",X"00",X"00",X"00",X"00",X"00",X"45",X"47",X"43",X"44",X"44",
		X"44",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"47",X"45",X"00",X"00",X"00",X"17",X"16",X"1C",
		X"13",X"00",X"07",X"07",X"08",X"03",X"16",X"00",X"17",X"1C",X"16",X"1F",X"1D",X"1A",X"20",X"1E",
		X"17",X"00",X"16",X"03",X"00",X"00",X"00",X"00",X"00",X"15",X"1C",X"1F",X"19",X"1B",X"20",X"1D",
		X"1D",X"20",X"1E",X"19",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"33",X"34",X"34",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"00",X"A1",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"C3",X"DF",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"BA",X"A0",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4E",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"48",X"45",X"43",X"43",X"47",X"45",X"00",X"00",X"00",X"03",X"64",X"02",X"1F",X"1C",X"1B",
		X"5F",X"02",X"5E",X"5E",X"0C",X"64",X"61",X"00",X"15",X"1A",X"1F",X"1D",X"1C",X"19",X"1F",X"1D",
		X"20",X"17",X"17",X"04",X"03",X"00",X"00",X"00",X"00",X"14",X"1B",X"1E",X"20",X"1A",X"1F",X"1C",
		X"1E",X"1A",X"1C",X"20",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"3E",X"3B",X"34",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"A2",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"C1",X"CF",X"D3",X"A0",X"A0",X"A0",X"A0",X"F7",X"FD",X"01",X"03",
		X"07",X"A0",X"A0",X"BB",X"BA",X"A0",X"A6",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"4D",X"47",X"46",X"46",X"45",X"46",X"45",X"45",X"4D",X"00",X"62",X"02",X"5E",X"04",X"5E",
		X"02",X"02",X"5F",X"5F",X"62",X"00",X"00",X"03",X"0C",X"5E",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"18",X"00",X"00",X"15",X"20",X"1E",X"1C",X"1B",X"20",X"1E",X"1C",
		X"1F",X"17",X"00",X"09",X"03",X"03",X"00",X"00",X"00",X"11",X"1A",X"1D",X"1F",X"19",X"1E",X"1B",
		X"1F",X"1B",X"20",X"1F",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"3E",X"3C",X"3B",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"A3",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"C1",X"CD",X"D5",X"C3",X"DF",X"ED",X"EF",X"F5",X"FB",X"FF",X"06",
		X"02",X"A0",X"BB",X"BA",X"BB",X"BA",X"A0",X"A0",X"A6",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"4B",X"45",X"46",X"45",X"46",X"45",X"46",X"45",X"49",X"00",X"09",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"0C",X"0C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"00",X"14",X"1F",X"1D",X"1B",X"1A",X"1F",X"1D",X"1B",
		X"1E",X"1C",X"11",X"16",X"00",X"03",X"03",X"00",X"00",X"13",X"19",X"1C",X"1E",X"20",X"1D",X"1A",
		X"20",X"1C",X"19",X"1D",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"3E",X"3B",X"3C",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"00",X"A1",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"C1",X"CD",X"D5",X"C1",X"CF",X"E9",X"EB",X"F3",X"F9",X"05",X"FE",
		X"00",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A5",X"00",X"00",X"00",X"00",
		X"00",X"4B",X"46",X"45",X"46",X"45",X"46",X"45",X"46",X"4E",X"17",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"11",X"1E",X"1C",X"1A",X"20",X"1E",X"1C",X"1A",
		X"1D",X"1B",X"11",X"13",X"17",X"00",X"03",X"03",X"00",X"19",X"20",X"1B",X"1D",X"1F",X"1C",X"19",
		X"19",X"1D",X"1A",X"1C",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"3E",X"34",X"3B",X"35",X"35",X"35",X"34",X"36",X"00",X"00",X"A2",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"BF",X"C9",X"D5",X"C1",X"CD",X"E5",X"E7",X"F1",X"04",X"F8",X"FA",
		X"FC",X"A0",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A5",X"00",X"00",
		X"00",X"4D",X"46",X"46",X"45",X"46",X"45",X"46",X"45",X"4B",X"13",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"17",X"12",X"1B",X"19",X"1F",X"1D",X"1B",X"19",
		X"1C",X"1A",X"17",X"17",X"13",X"00",X"00",X"03",X"03",X"14",X"1F",X"1A",X"1C",X"1E",X"1B",X"20",
		X"1A",X"1E",X"1D",X"1B",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"41",X"32",X"32",X"32",X"32",X"32",X"32",X"37",X"00",X"00",X"A3",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"BB",X"BD",X"CB",X"D7",X"CD",X"E5",X"E3",X"A0",X"F0",X"F2",X"F4",
		X"F6",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"0B",X"A0",X"A0",X"A0",X"A0",X"A6",X"A5",
		X"00",X"00",X"00",X"40",X"46",X"45",X"46",X"45",X"49",X"4D",X"15",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"64",X"11",X"1A",X"20",X"1E",X"1C",X"1A",X"20",
		X"1B",X"19",X"12",X"00",X"13",X"00",X"00",X"00",X"03",X"03",X"1E",X"19",X"1B",X"1D",X"1A",X"1F",
		X"1B",X"19",X"1C",X"20",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"BB",X"BA",X"C6",X"C7",X"E1",X"A0",X"E2",X"E6",X"EA",X"EE",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"0A",X"0C",X"0B",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A4",X"00",X"00",X"00",X"45",X"45",X"45",X"45",X"00",X"00",X"15",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"09",X"11",X"19",X"1F",X"1D",X"1B",X"19",X"1F",
		X"1A",X"20",X"1E",X"11",X"0D",X"00",X"00",X"00",X"00",X"7E",X"1D",X"20",X"1A",X"1C",X"19",X"1E",
		X"1C",X"20",X"1B",X"1F",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"E0",X"E4",X"E4",X"E8",X"EC",
		X"A0",X"A0",X"D8",X"D9",X"A0",X"A0",X"0B",X"08",X"09",X"0D",X"0F",X"0B",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"09",X"19",X"20",X"1E",X"1C",X"1A",X"20",X"1E",
		X"19",X"1F",X"1D",X"13",X"16",X"00",X"00",X"00",X"00",X"15",X"1C",X"1F",X"19",X"1B",X"20",X"1D",
		X"1D",X"1F",X"19",X"1E",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A3",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"B9",X"A0",X"A0",X"C5",X"CC",X"CC",X"CE",X"DE",
		X"A0",X"A0",X"DB",X"DA",X"DA",X"A0",X"A0",X"0E",X"0D",X"0E",X"EF",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A6",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"02",X"02",X"62",X"03",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"09",X"15",X"1F",X"1D",X"1B",X"19",X"1F",X"1D",
		X"20",X"1E",X"1C",X"11",X"16",X"61",X"00",X"00",X"17",X"1A",X"1B",X"1E",X"20",X"1A",X"1F",X"1C",
		X"1E",X"1E",X"20",X"1D",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"B7",X"B3",X"B8",X"BA",X"C4",X"D6",X"C0",X"C0",X"C2",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"0E",X"A0",X"A0",X"A0",X"A0",X"A0",X"B0",X"B4",
		X"A0",X"A0",X"A0",X"A0",X"AA",X"AB",X"A8",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"02",X"0C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"15",X"1E",X"1C",X"1A",X"20",X"1E",X"1C",
		X"1F",X"1D",X"1B",X"11",X"13",X"16",X"00",X"00",X"15",X"20",X"1A",X"1D",X"1F",X"19",X"1E",X"1B",
		X"1F",X"1D",X"19",X"1B",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"B5",X"B2",X"B6",X"A0",X"BB",X"BA",X"CA",X"D4",X"D4",X"D4",
		X"D2",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"BB",X"A0",X"A0",X"A0",X"A0",X"BB",X"BA",X"B5",X"B1",
		X"B4",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A8",X"A9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"62",X"02",X"0C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"16",X"00",X"12",X"1D",X"1B",X"19",X"1F",X"1D",X"1B",
		X"1E",X"1C",X"1A",X"19",X"17",X"04",X"5E",X"5F",X"1A",X"1F",X"19",X"1C",X"1E",X"20",X"1D",X"1A",
		X"20",X"1C",X"20",X"1A",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A3",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"B5",X"B1",X"B4",X"A0",X"A0",X"A0",X"BB",X"BC",X"C8",X"CC",X"CC",
		X"CE",X"DE",X"A0",X"A0",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"B5",
		X"B2",X"DD",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A8",X"A9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"0C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"17",X"19",X"1B",X"1C",X"1A",X"20",X"1E",X"1C",X"1A",
		X"1D",X"1B",X"19",X"10",X"00",X"16",X"61",X"81",X"19",X"1E",X"20",X"1B",X"1D",X"1F",X"1C",X"19",
		X"19",X"20",X"1E",X"19",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"B0",X"B4",X"A0",X"A0",X"A0",X"A0",X"A0",X"BB",X"BE",X"C0",X"C0",
		X"C0",X"C2",X"A0",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"A0",X"BB",X"BA",X"A0",X"A0",X"A0",X"A0",
		X"B7",X"DC",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A6",X"A8",
		X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"5E",X"5F",X"17",X"16",X"1A",X"1B",X"19",X"1F",X"1D",X"1B",X"19",
		X"1C",X"1A",X"20",X"1E",X"11",X"0D",X"13",X"19",X"20",X"1D",X"1F",X"1A",X"1C",X"1E",X"1B",X"20",
		X"AC",X"AD",X"AE",X"AF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"BA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"01",X"01",X"01",X"04",X"04",X"04",
		X"04",X"04",X"04",X"64",X"62",X"00",X"17",X"16",X"1A",X"19",X"1A",X"20",X"1E",X"1C",X"1A",X"20",
		X"1B",X"19",X"1F",X"1D",X"11",X"13",X"17",X"10",X"1F",X"1C",X"1E",X"19",X"1B",X"1D",X"1A",X"1F");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
