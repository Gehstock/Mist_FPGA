-------------------------------------------------------------------------------
--
-- i8244 Video Display Controller
--
-- $Id: i8244_minor-c.vhd,v 1.2 2007/02/05 21:57:37 arnim Exp $
--
-------------------------------------------------------------------------------

configuration i8244_minor_rtl_c0 of i8244_minor is

  for rtl
  end for;

end i8244_minor_rtl_c0;
