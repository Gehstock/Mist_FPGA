library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"13",X"60",X"B9",X"11",X"60",X"AA",X"A9",X"00",X"85",X"D4",X"A0",X"E2",X"A5",X"CE",X"4C",X"F6",
		X"6A",X"1D",X"B0",X"A5",X"93",X"D0",X"03",X"20",X"96",X"5F",X"F8",X"A5",X"D1",X"18",X"79",X"D6",
		X"01",X"99",X"D6",X"01",X"85",X"D1",X"B9",X"D8",X"01",X"65",X"D2",X"99",X"D8",X"01",X"85",X"D2",
		X"B9",X"DA",X"01",X"65",X"D3",X"99",X"DA",X"01",X"85",X"D3",X"A9",X"FF",X"85",X"D4",X"D8",X"60",
		X"A5",X"F4",X"29",X"70",X"4A",X"4A",X"4A",X"4A",X"A8",X"B9",X"7B",X"60",X"85",X"99",X"F0",X"EF",
		X"A6",X"B9",X"BD",X"D8",X"01",X"4A",X"4A",X"4A",X"4A",X"85",X"98",X"BD",X"DA",X"01",X"0A",X"0A",
		X"0A",X"0A",X"05",X"98",X"F8",X"38",X"F5",X"C3",X"38",X"E5",X"99",X"90",X"D1",X"F6",X"C0",X"48",
		X"B5",X"C3",X"18",X"65",X"99",X"95",X"C3",X"68",X"4C",X"68",X"60",X"10",X"12",X"14",X"15",X"18",
		X"20",X"08",X"00",X"01",X"20",X"01",X"40",X"01",X"50",X"01",X"80",X"01",X"00",X"02",X"80",X"00",
		X"0C",X"0F",X"12",X"0C",X"10",X"0E",X"11",X"0A",X"0D",X"10",X"13",X"0C",X"0E",X"10",X"12",X"0E",
		X"11",X"13",X"16",X"D0",X"E0",X"C0",X"08",X"A0",X"60",X"40",X"20",X"10",X"0A",X"06",X"04",X"02",
		X"01",X"00",X"04",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"03",X"04",X"04",X"05",X"05",X"06",X"06",
		X"07",X"07",X"07",X"07",X"80",X"60",X"40",X"30",X"20",X"20",X"10",X"F0",X"A0",X"80",X"80",X"60",
		X"40",X"20",X"5F",X"B4",X"94",X"2C",X"47",X"D0",X"14",X"7B",X"F0",X"10",X"15",X"12",X"12",X"11",
		X"11",X"16",X"16",X"16",X"18",X"18",X"18",X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"A5",
		X"8D",X"F0",X"42",X"AD",X"6D",X"01",X"D0",X"3D",X"A4",X"A7",X"C0",X"02",X"90",X"37",X"A5",X"E3",
		X"C5",X"E2",X"90",X"31",X"A2",X"00",X"86",X"C7",X"86",X"C9",X"AD",X"0A",X"40",X"10",X"01",X"CA",
		X"86",X"C8",X"8E",X"38",X"01",X"29",X"01",X"85",X"D6",X"AD",X"0A",X"40",X"4A",X"4A",X"4A",X"69",
		X"64",X"C0",X"06",X"B0",X"02",X"69",X"20",X"C0",X"04",X"B0",X"02",X"69",X"10",X"8D",X"6D",X"01",
		X"20",X"DC",X"7A",X"C6",X"DE",X"60",X"E6",X"E3",X"D0",X"02",X"C6",X"E3",X"AD",X"6D",X"01",X"F0",
		X"29",X"85",X"B1",X"C6",X"C7",X"10",X"23",X"E6",X"C9",X"A4",X"D6",X"B9",X"7B",X"61",X"85",X"C7",
		X"AD",X"38",X"01",X"20",X"7D",X"61",X"D0",X"0F",X"A9",X"00",X"8D",X"6D",X"01",X"85",X"C9",X"85",
		X"E3",X"20",X"F8",X"7A",X"B8",X"50",X"03",X"8D",X"38",X"01",X"60",X"01",X"02",X"84",X"AB",X"84",
		X"99",X"85",X"B0",X"A5",X"C8",X"30",X"05",X"E6",X"B0",X"B8",X"50",X"02",X"C6",X"B0",X"B9",X"ED",
		X"61",X"85",X"99",X"A6",X"99",X"BD",X"F5",X"61",X"85",X"98",X"BD",X"FB",X"61",X"85",X"B6",X"BC",
		X"EF",X"61",X"A6",X"99",X"B9",X"63",X"62",X"18",X"65",X"B1",X"49",X"FF",X"85",X"07",X"B9",X"13",
		X"62",X"45",X"C8",X"10",X"0A",X"18",X"65",X"B0",X"C5",X"B0",X"B0",X"1C",X"B8",X"50",X"07",X"18",
		X"65",X"B0",X"C5",X"B0",X"90",X"12",X"DD",X"01",X"62",X"90",X"0D",X"DD",X"07",X"62",X"B0",X"08",
		X"85",X"06",X"A2",X"00",X"A5",X"B6",X"81",X"06",X"C8",X"C6",X"98",X"10",X"C5",X"A4",X"99",X"C6",
		X"99",X"B9",X"0D",X"62",X"10",X"AD",X"A5",X"B0",X"F0",X"02",X"C9",X"FF",X"60",X"03",X"05",X"00",
		X"17",X"2C",X"30",X"36",X"43",X"16",X"14",X"03",X"05",X"0C",X"0C",X"40",X"00",X"80",X"E0",X"40",
		X"00",X"08",X"08",X"08",X"08",X"09",X"09",X"F8",X"F8",X"F8",X"F8",X"F7",X"F7",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"03",X"03",X"04",X"04",X"04",X"03",X"03",X"01",X"01",X"05",X"04",X"04",X"05",
		X"FB",X"FC",X"FC",X"FB",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"05",X"04",X"03",X"03",X"04",X"05",
		X"FE",X"FE",X"F9",X"FA",X"FB",X"FC",X"FC",X"FB",X"FB",X"FB",X"FC",X"FC",X"FB",X"FA",X"F9",X"06",
		X"06",X"FA",X"FA",X"02",X"02",X"02",X"FE",X"FE",X"FE",X"07",X"05",X"03",X"FF",X"FE",X"FD",X"00",
		X"FF",X"FE",X"FD",X"FC",X"F9",X"FA",X"FB",X"FC",X"FC",X"F8",X"F8",X"F8",X"F7",X"FA",X"FB",X"FB",
		X"FA",X"FA",X"F9",X"03",X"02",X"01",X"00",X"FF",X"FE",X"FD",X"04",X"FC",X"05",X"04",X"FC",X"FB",
		X"05",X"04",X"FC",X"FB",X"01",X"00",X"FF",X"01",X"00",X"FF",X"06",X"05",X"04",X"FC",X"FB",X"FA",
		X"04",X"FC",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"FF",X"FE",X"FD",X"FC",X"FB",X"FA",X"06",
		X"FA",X"06",X"FA",X"01",X"00",X"FF",X"01",X"00",X"FF",X"00",X"01",X"02",X"03",X"04",X"05",X"FF",
		X"FE",X"FD",X"FC",X"FB",X"04",X"03",X"05",X"04",X"03",X"04",X"03",X"02",X"01",X"00",X"FF",X"FE",
		X"FD",X"FC",X"FB",X"A2",X"13",X"A9",X"00",X"85",X"9A",X"BD",X"6E",X"01",X"F0",X"06",X"BD",X"C2",
		X"01",X"20",X"F1",X"62",X"A9",X"FC",X"85",X"EC",X"AD",X"0A",X"40",X"29",X"07",X"09",X"04",X"9D",
		X"C2",X"01",X"85",X"9A",X"AD",X"0A",X"40",X"9D",X"39",X"01",X"AD",X"0A",X"40",X"C9",X"D0",X"B0",
		X"F9",X"C9",X"38",X"90",X"F5",X"9D",X"6E",X"01",X"A9",X"00",X"20",X"F1",X"62",X"CA",X"10",X"C5",
		X"60",X"85",X"B5",X"BD",X"6E",X"01",X"85",X"9C",X"BD",X"39",X"01",X"85",X"9B",X"4C",X"71",X"5E",
		X"A5",X"A7",X"C9",X"28",X"90",X"02",X"A9",X"14",X"85",X"A7",X"4C",X"86",X"69",X"20",X"4D",X"63",
		X"A5",X"D5",X"D0",X"06",X"20",X"11",X"54",X"B8",X"50",X"32",X"C9",X"FF",X"D0",X"06",X"20",X"11",
		X"54",X"B8",X"50",X"28",X"20",X"8C",X"63",X"A5",X"D5",X"A4",X"A7",X"C0",X"09",X"B0",X"02",X"09",
		X"01",X"85",X"D5",X"20",X"00",X"64",X"D0",X"06",X"20",X"5D",X"64",X"B8",X"50",X"0E",X"20",X"2D",
		X"64",X"D0",X"06",X"20",X"5D",X"64",X"B8",X"50",X"03",X"20",X"11",X"54",X"60",X"A9",X"00",X"85",
		X"D5",X"86",X"AC",X"A0",X"07",X"A6",X"97",X"BD",X"5D",X"01",X"18",X"79",X"82",X"63",X"49",X"FF",
		X"85",X"B1",X"BD",X"28",X"01",X"18",X"79",X"84",X"63",X"85",X"B0",X"A2",X"00",X"A1",X"B0",X"29",
		X"C0",X"C9",X"80",X"D0",X"07",X"A5",X"D5",X"19",X"F8",X"63",X"85",X"D5",X"88",X"10",X"D6",X"A6",
		X"AC",X"60",X"08",X"06",X"00",X"FA",X"F8",X"FA",X"00",X"06",X"08",X"06",X"A4",X"97",X"20",X"F6",
		X"58",X"A4",X"B0",X"A5",X"B1",X"D0",X"05",X"A9",X"04",X"B8",X"50",X"16",X"20",X"BB",X"59",X"A0",
		X"04",X"A5",X"A9",X"D9",X"DE",X"63",X"D0",X"05",X"A5",X"AA",X"D9",X"E3",X"63",X"88",X"90",X"F1",
		X"C8",X"98",X"85",X"98",X"A6",X"97",X"BD",X"10",X"06",X"5D",X"30",X"06",X"10",X"07",X"A9",X"04",
		X"38",X"E5",X"98",X"85",X"98",X"BD",X"10",X"06",X"2A",X"BD",X"30",X"06",X"2A",X"2A",X"29",X"03",
		X"A8",X"B9",X"DA",X"63",X"18",X"65",X"98",X"85",X"D0",X"60",X"0C",X"08",X"00",X"04",X"00",X"00",
		X"00",X"01",X"05",X"00",X"32",X"AB",X"7F",X"06",X"83",X"87",X"07",X"0F",X"0E",X"1E",X"1C",X"3C",
		X"38",X"78",X"70",X"F0",X"E0",X"E1",X"C1",X"C3",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",
		X"A4",X"D0",X"A6",X"D0",X"A9",X"08",X"85",X"98",X"A5",X"D5",X"39",X"E8",X"63",X"D0",X"01",X"60",
		X"A5",X"D5",X"3D",X"E8",X"63",X"D0",X"05",X"8A",X"A8",X"A9",X"00",X"60",X"88",X"10",X"02",X"A0",
		X"0F",X"E8",X"E0",X"10",X"90",X"02",X"A2",X"00",X"C6",X"98",X"10",X"DC",X"60",X"A5",X"D0",X"4A",
		X"A8",X"AA",X"A9",X"04",X"85",X"98",X"A5",X"D5",X"39",X"F8",X"63",X"F0",X"09",X"A5",X"D5",X"3D",
		X"F8",X"63",X"D0",X"08",X"8A",X"A8",X"98",X"0A",X"A8",X"A9",X"00",X"60",X"88",X"10",X"02",X"A0",
		X"07",X"E8",X"E0",X"08",X"90",X"02",X"A2",X"00",X"C6",X"98",X"10",X"DA",X"60",X"A6",X"97",X"BD",
		X"28",X"01",X"C9",X"F7",X"B0",X"19",X"C9",X"08",X"90",X"15",X"BD",X"5D",X"01",X"C9",X"CE",X"B0",
		X"0E",X"C9",X"2D",X"90",X"0A",X"20",X"82",X"64",X"A4",X"97",X"20",X"F6",X"58",X"18",X"60",X"4C",
		X"11",X"54",X"A6",X"97",X"B9",X"AF",X"64",X"18",X"7D",X"18",X"01",X"9D",X"18",X"01",X"B9",X"C3",
		X"64",X"7D",X"28",X"01",X"9D",X"28",X"01",X"B9",X"AB",X"64",X"18",X"7D",X"4D",X"01",X"9D",X"4D",
		X"01",X"B9",X"BF",X"64",X"7D",X"5D",X"01",X"9D",X"5D",X"01",X"60",X"00",X"EC",X"B4",X"62",X"00",
		X"9E",X"4C",X"14",X"00",X"14",X"4C",X"9E",X"00",X"62",X"B4",X"EC",X"00",X"EC",X"B4",X"62",X"01",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"A9",X"E0",X"4C",X"DA",X"64",X"A9",X"00",X"85",X"98",X"A5",X"0A",X"C9",X"18",
		X"90",X"78",X"18",X"69",X"03",X"49",X"FF",X"85",X"07",X"A5",X"09",X"85",X"06",X"38",X"E9",X"03",
		X"85",X"03",X"A5",X"0A",X"49",X"FF",X"85",X"04",X"A5",X"A6",X"C9",X"18",X"90",X"5C",X"85",X"0A",
		X"18",X"69",X"03",X"49",X"FF",X"85",X"01",X"A5",X"A5",X"85",X"09",X"85",X"00",X"38",X"E9",X"03",
		X"85",X"0D",X"A5",X"A6",X"49",X"FF",X"85",X"0E",X"A0",X"06",X"A2",X"00",X"A1",X"03",X"29",X"E0",
		X"C9",X"E0",X"D0",X"05",X"B9",X"16",X"00",X"81",X"03",X"A1",X"06",X"29",X"E0",X"C9",X"E0",X"D0",
		X"05",X"B9",X"0F",X"00",X"81",X"06",X"E6",X"03",X"E6",X"07",X"88",X"10",X"DF",X"A0",X"06",X"A2",
		X"00",X"A1",X"00",X"99",X"0F",X"00",X"A5",X"98",X"81",X"00",X"E6",X"01",X"A1",X"0D",X"99",X"16",
		X"00",X"A5",X"98",X"81",X"0D",X"E6",X"0D",X"88",X"10",X"E7",X"60",X"16",X"A9",X"80",X"85",X"09",
		X"85",X"A5",X"A9",X"50",X"85",X"0A",X"85",X"A6",X"A9",X"00",X"A2",X"0D",X"95",X"0F",X"CA",X"10",
		X"FB",X"60",X"20",X"D8",X"64",X"A9",X"00",X"85",X"A6",X"85",X"0A",X"60",X"86",X"23",X"A9",X"80",
		X"85",X"0B",X"A5",X"A6",X"49",X"FF",X"38",X"E9",X"02",X"85",X"07",X"85",X"01",X"A5",X"A5",X"4C",
		X"A9",X"65",X"86",X"23",X"A9",X"00",X"85",X"0B",X"A6",X"97",X"BD",X"B2",X"01",X"49",X"FF",X"38",
		X"E9",X"02",X"85",X"07",X"85",X"01",X"BD",X"A2",X"01",X"18",X"69",X"02",X"85",X"06",X"38",X"E9",
		X"04",X"85",X"00",X"A2",X"00",X"A9",X"04",X"85",X"98",X"A5",X"0B",X"81",X"06",X"81",X"00",X"E6",
		X"07",X"C6",X"06",X"E6",X"01",X"E6",X"00",X"C6",X"98",X"10",X"F0",X"A6",X"23",X"60",X"A0",X"E0",
		X"A5",X"B9",X"20",X"DB",X"65",X"A0",X"00",X"A5",X"B9",X"49",X"01",X"84",X"0B",X"AA",X"BD",X"EC",
		X"65",X"48",X"BD",X"EE",X"65",X"AA",X"A0",X"E2",X"68",X"4C",X"00",X"66",X"21",X"22",X"4D",X"A8",
		X"A5",X"D7",X"D0",X"06",X"20",X"CE",X"65",X"B8",X"50",X"05",X"A0",X"00",X"20",X"D0",X"65",X"60",
		X"85",X"0D",X"86",X"00",X"84",X"01",X"A9",X"00",X"85",X"0E",X"A9",X"FF",X"85",X"08",X"06",X"0D",
		X"26",X"0E",X"06",X"0D",X"26",X"0E",X"06",X"0D",X"26",X"0E",X"A9",X"62",X"18",X"65",X"0D",X"85",
		X"0D",X"A9",X"73",X"65",X"0E",X"85",X"0E",X"A9",X"01",X"85",X"22",X"85",X"21",X"A0",X"07",X"A5",
		X"01",X"18",X"69",X"04",X"49",X"FF",X"85",X"07",X"A5",X"21",X"85",X"04",X"A5",X"00",X"38",X"E9",
		X"04",X"24",X"FC",X"50",X"02",X"49",X"FF",X"85",X"06",X"A2",X"00",X"A9",X"07",X"85",X"98",X"B1",
		X"0D",X"0A",X"48",X"A5",X"22",X"85",X"03",X"A5",X"0B",X"B0",X"0B",X"A5",X"08",X"10",X"05",X"A1",
		X"06",X"B8",X"50",X"02",X"A5",X"0C",X"81",X"06",X"24",X"FC",X"50",X"05",X"C6",X"06",X"B8",X"50",
		X"02",X"E6",X"06",X"C6",X"03",X"D0",X"EF",X"68",X"C6",X"98",X"10",X"D5",X"E6",X"07",X"C6",X"04",
		X"D0",X"BA",X"88",X"10",X"B3",X"60",X"86",X"23",X"84",X"24",X"A4",X"97",X"A9",X"00",X"85",X"98",
		X"A9",X"FF",X"85",X"99",X"B9",X"92",X"01",X"49",X"FF",X"85",X"07",X"B9",X"82",X"01",X"85",X"06",
		X"B9",X"00",X"06",X"85",X"03",X"B9",X"20",X"06",X"85",X"04",X"B9",X"10",X"06",X"85",X"00",X"B9",
		X"30",X"06",X"85",X"01",X"B9",X"5D",X"01",X"49",X"FF",X"85",X"02",X"C5",X"07",X"F0",X"2C",X"A2",
		X"00",X"A9",X"00",X"81",X"06",X"A5",X"98",X"18",X"65",X"03",X"85",X"98",X"A5",X"06",X"65",X"00",
		X"85",X"06",X"A5",X"99",X"38",X"E5",X"04",X"85",X"99",X"A5",X"07",X"E5",X"01",X"85",X"07",X"C9",
		X"18",X"90",X"08",X"C5",X"02",X"D0",X"DA",X"A9",X"00",X"81",X"06",X"A6",X"23",X"A4",X"24",X"60",
		X"A4",X"97",X"A9",X"80",X"4C",X"01",X"67",X"A9",X"E0",X"A4",X"97",X"C0",X"08",X"90",X"02",X"A9",
		X"40",X"85",X"0B",X"86",X"98",X"B9",X"28",X"01",X"85",X"06",X"B9",X"5D",X"01",X"49",X"FF",X"85",
		X"07",X"A5",X"0B",X"A2",X"00",X"81",X"06",X"A6",X"98",X"60",X"A2",X"07",X"A9",X"0E",X"95",X"E4",
		X"CA",X"10",X"FB",X"20",X"00",X"63",X"20",X"7C",X"68",X"20",X"5E",X"67",X"20",X"21",X"69",X"A5",
		X"F3",X"4A",X"4A",X"4A",X"4A",X"29",X"06",X"A8",X"B9",X"95",X"6A",X"85",X"2A",X"B9",X"96",X"6A",
		X"85",X"2B",X"A9",X"00",X"A4",X"F4",X"10",X"08",X"09",X"80",X"A4",X"B9",X"F0",X"02",X"09",X"7F",
		X"85",X"FC",X"60",X"BE",X"E2",X"60",X"B9",X"EB",X"60",X"A8",X"A9",X"00",X"F0",X"21",X"A0",X"05",
		X"84",X"99",X"A4",X"B9",X"B9",X"C5",X"00",X"A4",X"99",X"39",X"F7",X"60",X"F0",X"0C",X"BE",X"E2",
		X"60",X"B9",X"EB",X"60",X"A8",X"A9",X"E6",X"20",X"7F",X"67",X"C6",X"99",X"10",X"E4",X"60",X"48",
		X"A5",X"FC",X"29",X"BF",X"85",X"FC",X"68",X"20",X"95",X"67",X"A5",X"FC",X"29",X"3F",X"F0",X"04",
		X"09",X"C0",X"85",X"FC",X"60",X"86",X"1D",X"84",X"1E",X"85",X"1F",X"0A",X"0A",X"0A",X"0A",X"85",
		X"20",X"A2",X"03",X"86",X"05",X"A6",X"05",X"BC",X"C5",X"67",X"B9",X"1F",X"00",X"85",X"0B",X"A4",
		X"1E",X"BD",X"C9",X"67",X"48",X"A5",X"1D",X"18",X"7D",X"CD",X"67",X"AA",X"68",X"20",X"00",X"66",
		X"C6",X"05",X"10",X"E1",X"60",X"01",X"00",X"01",X"00",X"1E",X"1D",X"20",X"1F",X"FC",X"FC",X"04",
		X"04",X"BE",X"A0",X"00",X"E8",X"A9",X"20",X"18",X"48",X"B9",X"E8",X"60",X"7D",X"19",X"68",X"85",
		X"06",X"18",X"B9",X"F1",X"60",X"7D",X"0F",X"68",X"49",X"FF",X"85",X"07",X"68",X"A2",X"00",X"81",
		X"06",X"E6",X"07",X"81",X"06",X"E6",X"07",X"81",X"06",X"E6",X"07",X"81",X"06",X"C6",X"06",X"81",
		X"06",X"E6",X"07",X"81",X"06",X"E6",X"06",X"E6",X"06",X"81",X"06",X"C6",X"07",X"81",X"06",X"60",
		X"02",X"FF",X"FF",X"FC",X"FC",X"FC",X"F9",X"F9",X"F9",X"F9",X"00",X"FD",X"03",X"FA",X"00",X"06",
		X"FD",X"03",X"F7",X"09",X"86",X"23",X"84",X"24",X"AA",X"BD",X"61",X"68",X"24",X"FC",X"50",X"03",
		X"BD",X"67",X"68",X"4C",X"56",X"68",X"85",X"02",X"86",X"23",X"84",X"24",X"AA",X"BD",X"61",X"68",
		X"24",X"FC",X"50",X"03",X"BD",X"67",X"68",X"20",X"4D",X"6A",X"A6",X"02",X"BD",X"5E",X"68",X"24",
		X"FC",X"50",X"03",X"BD",X"64",X"68",X"20",X"55",X"6A",X"A6",X"23",X"A4",X"24",X"60",X"0F",X"10",
		X"11",X"16",X"17",X"18",X"11",X"10",X"0F",X"18",X"17",X"16",X"BE",X"A0",X"00",X"F0",X"0C",X"86",
		X"02",X"A9",X"E0",X"20",X"D7",X"67",X"A6",X"02",X"CA",X"D0",X"F4",X"60",X"A2",X"00",X"A0",X"00",
		X"A9",X"E6",X"85",X"07",X"B9",X"AB",X"68",X"85",X"06",X"C8",X"A9",X"20",X"81",X"06",X"A5",X"06",
		X"D9",X"AB",X"68",X"E6",X"06",X"90",X"F3",X"C8",X"B9",X"AB",X"68",X"C9",X"FF",X"D0",X"09",X"C8",
		X"C0",X"74",X"90",X"02",X"A0",X"73",X"E6",X"07",X"D0",X"DA",X"60",X"0C",X"0D",X"1D",X"1E",X"75",
		X"76",X"81",X"82",X"E9",X"EA",X"FA",X"FB",X"FF",X"0B",X"0E",X"1C",X"1F",X"75",X"77",X"80",X"83",
		X"E7",X"EA",X"F9",X"FC",X"FF",X"0A",X"20",X"74",X"84",X"E6",X"FD",X"FF",X"09",X"21",X"73",X"84",
		X"E6",X"FE",X"FF",X"08",X"22",X"73",X"85",X"E5",X"FE",X"FF",X"06",X"23",X"72",X"85",X"E4",X"FE",
		X"FF",X"05",X"23",X"71",X"86",X"AC",X"BB",X"E3",X"FE",X"FF",X"04",X"24",X"38",X"39",X"70",X"87",
		X"AB",X"BC",X"E2",X"FE",X"FF",X"03",X"25",X"37",X"3A",X"6F",X"87",X"AA",X"BD",X"E1",X"FF",X"FF",
		X"01",X"26",X"32",X"3B",X"6B",X"98",X"A8",X"BD",X"DF",X"FF",X"FF",X"00",X"3C",X"49",X"58",X"67",
		X"C0",X"DE",X"FE",X"FF",X"00",X"5A",X"65",X"FF",X"FF",X"00",X"5C",X"64",X"FF",X"FF",X"00",X"FF",
		X"FF",X"A5",X"A7",X"38",X"E9",X"01",X"4A",X"C9",X"0A",X"90",X"03",X"38",X"E9",X"0A",X"C9",X"0A",
		X"B0",X"F5",X"AA",X"BC",X"4E",X"69",X"A2",X"06",X"B9",X"4E",X"69",X"29",X"0F",X"95",X"E5",X"B9",
		X"4E",X"69",X"4A",X"4A",X"4A",X"4A",X"95",X"E4",X"88",X"CA",X"CA",X"10",X"EB",X"60",X"19",X"1D",
		X"21",X"15",X"25",X"2D",X"31",X"0D",X"11",X"29",X"2A",X"E0",X"E2",X"66",X"06",X"42",X"40",X"AA",
		X"E6",X"22",X"0A",X"CC",X"E2",X"68",X"6E",X"CC",X"E2",X"A8",X"AE",X"CC",X"EC",X"62",X"64",X"AA",
		X"C2",X"64",X"6C",X"EE",X"62",X"EA",X"E6",X"CC",X"82",X"6E",X"68",X"CC",X"4A",X"EE",X"48",X"22",
		X"A9",X"06",X"A2",X"28",X"D0",X"04",X"A2",X"3D",X"A9",X"02",X"85",X"07",X"A0",X"00",X"84",X"06",
		X"A9",X"00",X"91",X"06",X"C8",X"D0",X"FB",X"E6",X"07",X"CA",X"10",X"F6",X"60",X"29",X"7F",X"C9",
		X"41",X"90",X"07",X"29",X"3F",X"A2",X"02",X"B8",X"50",X"18",X"C9",X"3A",X"90",X"06",X"20",X"D3",
		X"69",X"B8",X"50",X"0E",X"C9",X"30",X"B0",X"06",X"20",X"D3",X"69",X"B8",X"50",X"04",X"29",X"0F",
		X"A2",X"00",X"0A",X"0A",X"0A",X"18",X"7D",X"1E",X"6A",X"85",X"0D",X"BD",X"1F",X"6A",X"69",X"00",
		X"85",X"0E",X"60",X"A2",X"06",X"DD",X"E8",X"69",X"D0",X"06",X"BD",X"EF",X"69",X"A2",X"06",X"60",
		X"CA",X"10",X"F2",X"A9",X"00",X"A2",X"04",X"60",X"20",X"40",X"3A",X"3F",X"23",X"24",X"25",X"00",
		X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"A0",X"00",X"B1",X"1D",X"85",X"05",X"20",X"9D",X"69",X"A5",
		X"1F",X"85",X"00",X"A5",X"20",X"85",X"01",X"98",X"48",X"20",X"2D",X"66",X"A5",X"22",X"0A",X"0A",
		X"0A",X"18",X"65",X"1F",X"85",X"1F",X"68",X"A8",X"C8",X"A5",X"05",X"10",X"DB",X"60",X"1A",X"73",
		X"62",X"73",X"12",X"73",X"3A",X"74",X"B1",X"2A",X"C0",X"54",X"90",X"10",X"B9",X"12",X"6E",X"85",
		X"1F",X"B9",X"13",X"6E",X"85",X"1D",X"B9",X"14",X"6E",X"B8",X"50",X"0A",X"85",X"1F",X"C8",X"B1",
		X"2A",X"85",X"1D",X"C8",X"B1",X"2A",X"85",X"1E",X"60",X"A0",X"A0",X"30",X"0A",X"A0",X"80",X"30",
		X"06",X"A0",X"00",X"10",X"02",X"A0",X"FF",X"84",X"08",X"A8",X"B9",X"C5",X"6C",X"29",X"0F",X"85",
		X"21",X"B9",X"C5",X"6C",X"4A",X"4A",X"4A",X"4A",X"85",X"22",X"B9",X"ED",X"6C",X"85",X"20",X"98",
		X"85",X"1F",X"0A",X"18",X"65",X"1F",X"A8",X"20",X"26",X"6A",X"A9",X"E0",X"85",X"0B",X"A9",X"00",
		X"85",X"0C",X"A5",X"08",X"C9",X"80",X"D0",X"03",X"4C",X"38",X"6B",X"C9",X"A0",X"D0",X"03",X"4C",
		X"30",X"6B",X"4C",X"F6",X"69",X"12",X"6E",X"16",X"6D",X"6A",X"6D",X"BE",X"6D",X"86",X"1F",X"84",
		X"20",X"86",X"23",X"84",X"24",X"85",X"02",X"C9",X"13",X"B0",X"13",X"C9",X"0A",X"90",X"0A",X"38",
		X"E9",X"0A",X"85",X"02",X"A9",X"01",X"20",X"C8",X"6A",X"A5",X"02",X"B8",X"50",X"02",X"A9",X"FF",
		X"20",X"C8",X"6A",X"A6",X"23",X"A4",X"24",X"60",X"18",X"69",X"01",X"0A",X"0A",X"0A",X"18",X"6D",
		X"22",X"6A",X"85",X"0D",X"AD",X"23",X"6A",X"69",X"00",X"85",X"0E",X"A5",X"1F",X"85",X"00",X"A5",
		X"20",X"85",X"01",X"A9",X"00",X"85",X"0C",X"A9",X"00",X"85",X"08",X"20",X"27",X"66",X"A5",X"1F",
		X"18",X"69",X"08",X"85",X"1F",X"60",X"86",X"1F",X"84",X"20",X"85",X"0B",X"A2",X"02",X"A0",X"00",
		X"84",X"05",X"B5",X"D1",X"4A",X"4A",X"4A",X"4A",X"20",X"1E",X"6B",X"B5",X"D1",X"E0",X"00",X"D0",
		X"04",X"A0",X"FF",X"84",X"05",X"29",X"0F",X"20",X"1E",X"6B",X"CA",X"10",X"E5",X"60",X"F0",X"05",
		X"85",X"05",X"B8",X"50",X"08",X"A9",X"00",X"A4",X"05",X"D0",X"02",X"A9",X"FF",X"4C",X"A1",X"6A",
		X"A9",X"04",X"85",X"1F",X"A0",X"20",X"D0",X"08",X"A0",X"FF",X"C8",X"B1",X"1D",X"10",X"FB",X"C8",
		X"84",X"99",X"06",X"99",X"C6",X"99",X"A5",X"1F",X"38",X"E9",X"04",X"24",X"FC",X"50",X"02",X"49",
		X"FF",X"85",X"1F",X"A5",X"20",X"49",X"FF",X"38",X"E9",X"04",X"85",X"20",X"A9",X"07",X"85",X"98",
		X"46",X"20",X"66",X"1F",X"46",X"20",X"66",X"1F",X"24",X"FC",X"50",X"07",X"A5",X"1F",X"38",X"E5",
		X"99",X"85",X"1F",X"A4",X"99",X"A9",X"00",X"91",X"1F",X"88",X"10",X"F9",X"A5",X"1F",X"18",X"69",
		X"40",X"85",X"1F",X"90",X"02",X"E6",X"20",X"C6",X"98",X"10",X"E8",X"60",X"A9",X"00",X"85",X"B9",
		X"A5",X"FC",X"29",X"80",X"85",X"FC",X"A5",X"66",X"C9",X"28",X"90",X"04",X"A9",X"28",X"85",X"66",
		X"F8",X"85",X"99",X"A9",X"00",X"85",X"98",X"A0",X"07",X"06",X"99",X"A5",X"98",X"65",X"98",X"85",
		X"98",X"88",X"10",X"F5",X"D8",X"A5",X"98",X"C5",X"29",X"F0",X"22",X"85",X"29",X"A5",X"66",X"F0",
		X"05",X"A2",X"00",X"B8",X"50",X"0C",X"A5",X"F3",X"29",X"03",X"AA",X"BD",X"2F",X"6C",X"85",X"28",
		X"A2",X"05",X"86",X"25",X"20",X"B6",X"6C",X"A9",X"00",X"85",X"27",X"85",X"26",X"A5",X"27",X"F0",
		X"05",X"C6",X"27",X"B8",X"50",X"48",X"A6",X"25",X"BD",X"42",X"6C",X"C9",X"00",X"D0",X"09",X"BD",
		X"38",X"6C",X"20",X"7F",X"6C",X"B8",X"50",X"1B",X"BD",X"38",X"6C",X"85",X"06",X"A0",X"00",X"84",
		X"07",X"B1",X"06",X"BC",X"42",X"6C",X"C0",X"02",X"D0",X"06",X"20",X"7F",X"6C",X"B8",X"50",X"03",
		X"20",X"56",X"6C",X"A5",X"27",X"C9",X"FF",X"D0",X"15",X"A6",X"25",X"BD",X"4C",X"6C",X"85",X"27",
		X"E8",X"BD",X"42",X"6C",X"C9",X"03",X"D0",X"04",X"BD",X"38",X"6C",X"AA",X"86",X"25",X"60",X"25",
		X"0A",X"0B",X"0C",X"A9",X"FF",X"85",X"29",X"60",X"03",X"0D",X"29",X"1E",X"00",X"0E",X"04",X"28",
		X"1E",X"05",X"00",X"00",X"01",X"00",X"03",X"00",X"00",X"02",X"00",X"03",X"20",X"08",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"A4",X"26",X"F0",X"0A",X"A0",X"FF",X"84",X"27",X"C8",X"84",
		X"26",X"B8",X"50",X"0E",X"A0",X"07",X"84",X"27",X"E6",X"26",X"4A",X"4A",X"4A",X"4A",X"D0",X"02",
		X"A9",X"FF",X"29",X"0F",X"C9",X"0A",X"B0",X"06",X"18",X"69",X"30",X"20",X"9C",X"6C",X"60",X"85",
		X"1D",X"0A",X"18",X"65",X"1D",X"A8",X"20",X"26",X"6A",X"A4",X"26",X"E6",X"26",X"A9",X"07",X"85",
		X"27",X"B1",X"1D",X"10",X"07",X"A0",X"FF",X"84",X"27",X"C8",X"84",X"26",X"20",X"9D",X"69",X"A9",
		X"FC",X"85",X"00",X"A9",X"03",X"85",X"01",X"A9",X"00",X"85",X"08",X"A9",X"00",X"85",X"0B",X"A9",
		X"20",X"85",X"0C",X"4C",X"27",X"66",X"A0",X"00",X"A9",X"FF",X"99",X"01",X"04",X"99",X"01",X"05",
		X"C8",X"C8",X"D0",X"F6",X"60",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"3A",X"21",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"90",X"D0",X"03",
		X"03",X"03",X"40",X"70",X"A0",X"A0",X"80",X"40",X"40",X"40",X"03",X"A0",X"03",X"03",X"03",X"70",
		X"60",X"50",X"38",X"03",X"03",X"03",X"58",X"58",X"58",X"A0",X"70",X"03",X"70",X"90",X"70",X"90",
		X"80",X"80",X"40",X"34",X"80",X"95",X"60",X"D2",X"6F",X"40",X"BB",X"70",X"06",X"D8",X"6F",X"90",
		X"E5",X"6F",X"78",X"F6",X"6F",X"5C",X"0B",X"70",X"68",X"22",X"70",X"50",X"16",X"70",X"60",X"2A",
		X"70",X"10",X"5F",X"70",X"40",X"2D",X"70",X"40",X"3E",X"70",X"40",X"4E",X"70",X"B0",X"F6",X"6E",
		X"54",X"D8",X"6F",X"04",X"E1",X"70",X"70",X"E1",X"70",X"E4",X"E1",X"70",X"24",X"6E",X"70",X"04",
		X"86",X"70",X"04",X"A1",X"70",X"34",X"CB",X"70",X"0C",X"DE",X"70",X"74",X"DE",X"70",X"E8",X"DE",
		X"70",X"88",X"E5",X"70",X"C8",X"24",X"70",X"28",X"0B",X"70",X"54",X"E6",X"70",X"50",X"D0",X"71",
		X"06",X"ED",X"70",X"90",X"F6",X"70",X"78",X"09",X"71",X"5C",X"17",X"71",X"68",X"2C",X"71",X"58",
		X"21",X"71",X"54",X"34",X"71",X"14",X"6E",X"71",X"40",X"38",X"71",X"40",X"47",X"71",X"40",X"56",
		X"71",X"B0",X"66",X"71",X"58",X"ED",X"70",X"04",X"F7",X"71",X"70",X"F7",X"71",X"E4",X"F7",X"71",
		X"14",X"7C",X"71",X"04",X"98",X"71",X"04",X"B7",X"71",X"30",X"DC",X"71",X"04",X"F2",X"71",X"6C",
		X"F2",X"71",X"DC",X"F2",X"71",X"70",X"FB",X"71",X"C8",X"2E",X"71",X"18",X"17",X"71",X"5C",X"FF",
		X"71",X"64",X"EB",X"72",X"06",X"06",X"72",X"90",X"15",X"72",X"78",X"21",X"72",X"5C",X"2F",X"72",
		X"68",X"51",X"72",X"30",X"3B",X"72",X"60",X"2A",X"70",X"24",X"94",X"72",X"40",X"59",X"72",X"40",
		X"6A",X"72",X"40",X"7A",X"72",X"B0",X"8B",X"72",X"48",X"06",X"72",X"0C",X"0B",X"73",X"74",X"0B",
		X"73",X"E8",X"0B",X"73",X"38",X"A0",X"72",X"04",X"B3",X"72",X"04",X"D3",X"72",X"30",X"F2",X"72",
		X"04",X"07",X"73",X"70",X"07",X"73",X"E4",X"07",X"73",X"70",X"0E",X"73",X"C8",X"53",X"72",X"08",
		X"2F",X"72",X"60",X"8A",X"6E",X"54",X"78",X"6F",X"06",X"90",X"6E",X"90",X"99",X"6E",X"78",X"A4",
		X"6E",X"5C",X"B0",X"6E",X"68",X"22",X"70",X"50",X"BA",X"6E",X"36",X"C6",X"6E",X"2C",X"20",X"6F",
		X"40",X"CD",X"6E",X"40",X"DB",X"6E",X"40",X"E8",X"6E",X"B0",X"F6",X"6E",X"5C",X"90",X"6E",X"0C",
		X"A6",X"6F",X"74",X"A6",X"6F",X"E8",X"A6",X"6F",X"38",X"2B",X"6F",X"04",X"3E",X"6F",X"04",X"59",
		X"6F",X"38",X"83",X"6F",X"0C",X"96",X"6F",X"74",X"96",X"6F",X"E8",X"96",X"6F",X"68",X"C4",X"6F",
		X"C8",X"24",X"70",X"10",X"B0",X"6E",X"20",X"B6",X"6F",X"20",X"BD",X"6F",X"50",X"A9",X"6F",X"5C",
		X"FE",X"6E",X"5C",X"04",X"6F",X"5C",X"0A",X"6F",X"5C",X"11",X"6F",X"5C",X"9F",X"6F",X"5C",X"99",
		X"6F",X"40",X"C9",X"6F",X"50",X"90",X"6F",X"10",X"18",X"6F",X"50",X"4C",X"41",X"59",X"45",X"D2",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"D2",X"50",X"52",X"45",X"53",X"53",X"20",X"53",
		X"54",X"41",X"52",X"D4",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"D3",
		X"42",X"4F",X"4E",X"55",X"53",X"20",X"43",X"49",X"54",X"D9",X"42",X"4F",X"4E",X"55",X"53",X"20",
		X"50",X"4F",X"49",X"4E",X"54",X"D3",X"54",X"48",X"45",X"20",X"45",X"4E",X"C4",X"31",X"20",X"43",
		X"4F",X"49",X"4E",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"D3",X"31",X"20",X"43",X"4F",X"49",
		X"4E",X"20",X"31",X"20",X"50",X"4C",X"41",X"D9",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",
		X"31",X"20",X"50",X"4C",X"41",X"D9",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"BA",X"52",X"41",
		X"4D",X"20",X"4F",X"CB",X"52",X"4F",X"4D",X"20",X"4F",X"CB",X"42",X"41",X"44",X"20",X"52",X"41",
		X"CD",X"42",X"41",X"44",X"20",X"52",X"4F",X"CD",X"42",X"41",X"44",X"20",X"43",X"48",X"49",X"D0",
		X"47",X"52",X"45",X"41",X"54",X"20",X"53",X"43",X"4F",X"52",X"C5",X"45",X"4E",X"54",X"45",X"52",
		X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"D3",X"53",X"50",
		X"49",X"4E",X"20",X"42",X"41",X"4C",X"4C",X"20",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",
		X"45",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"D3",X"50",X"52",X"45",X"53",X"53",X"20",X"41",
		X"4E",X"59",X"20",X"46",X"49",X"52",X"45",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"20",X"54",
		X"4F",X"20",X"53",X"45",X"4C",X"45",X"43",X"D4",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",
		X"52",X"45",X"D3",X"44",X"45",X"46",X"45",X"4E",X"44",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"43",X"49",X"54",X"49",X"45",X"D3",X"4C",X"4F",X"D7",X"4D",X"41",X"50",X"20",X"4F",X"CB",X"42",
		X"41",X"44",X"20",X"4D",X"41",X"D0",X"4F",X"55",X"D4",X"41",X"54",X"41",X"52",X"49",X"20",X"40",
		X"3F",X"20",X"31",X"39",X"38",X"B0",X"4D",X"49",X"53",X"53",X"49",X"4C",X"C5",X"43",X"4F",X"4D",
		X"4D",X"41",X"4E",X"C4",X"45",X"56",X"45",X"52",X"D9",X"46",X"52",X"45",X"45",X"20",X"50",X"4C",
		X"41",X"D9",X"4A",X"4F",X"55",X"45",X"55",X"D2",X"46",X"49",X"4E",X"20",X"44",X"45",X"20",X"50",
		X"41",X"52",X"54",X"49",X"C5",X"41",X"50",X"50",X"55",X"59",X"45",X"5A",X"20",X"53",X"55",X"52",
		X"20",X"53",X"54",X"41",X"52",X"D4",X"49",X"4E",X"54",X"52",X"4F",X"44",X"55",X"49",X"52",X"45");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
