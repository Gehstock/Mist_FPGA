library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GAL_FIR is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GAL_FIR is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AC",X"68",X"72",X"C7",X"93",X"3F",X"80",X"C8",X"5C",X"A1",X"22",X"90",X"B9",X"8A",X"41",X"62",
		X"C2",X"A1",X"40",X"6A",X"C9",X"7F",X"64",X"3C",X"BC",X"AD",X"5B",X"4C",X"D4",X"62",X"3D",X"D3",
		X"7F",X"31",X"A3",X"BE",X"5D",X"49",X"C7",X"7D",X"28",X"C0",X"A1",X"7A",X"7D",X"2B",X"C9",X"91",
		X"80",X"6B",X"39",X"95",X"BA",X"91",X"27",X"C1",X"91",X"7E",X"6D",X"31",X"C0",X"A4",X"7C",X"7B",
		X"37",X"80",X"CB",X"7E",X"88",X"64",X"40",X"8F",X"C3",X"83",X"83",X"68",X"36",X"D0",X"8C",X"29",
		X"B4",X"B1",X"52",X"4B",X"E9",X"3E",X"74",X"C4",X"73",X"81",X"2B",X"AD",X"B9",X"4E",X"4B",X"CB",
		X"91",X"76",X"33",X"B6",X"A5",X"6E",X"4A",X"63",X"D7",X"7C",X"3E",X"7E",X"DE",X"45",X"67",X"C1",
		X"84",X"2D",X"A8",X"A9",X"20",X"AC",X"B5",X"7E",X"47",X"5F",X"DD",X"6E",X"44",X"BD",X"97",X"22",
		X"AE",X"A4",X"25",X"CB",X"93",X"77",X"3C",X"78",X"CB",X"83",X"29",X"B3",X"AB",X"7D",X"5D",X"44",
		X"A4",X"BC",X"79",X"8C",X"3A",X"76",X"CF",X"78",X"44",X"6B",X"D9",X"6B",X"3B",X"9A",X"CC",X"26",
		X"A4",X"A3",X"1D",X"BA",X"A9",X"83",X"71",X"3A",X"8B",X"CC",X"6A",X"3E",X"E5",X"28",X"A4",X"A3",
		X"1E",X"C9",X"9C",X"78",X"32",X"94",X"C4",X"74",X"88",X"2A",X"A2",X"BC",X"1A",X"E2",X"4B",X"86",
		X"B3",X"72",X"48",X"68",X"D2",X"83",X"32",X"A4",X"B2",X"73",X"4E",X"5A",X"C8",X"9C",X"2C",X"90",
		X"C1",X"7B",X"5E",X"41",X"CC",X"99",X"6F",X"3A",X"8B",X"C9",X"7A",X"84",X"23",X"BC",X"9D",X"33",
		X"CC",X"82",X"24",X"D7",X"6C",X"47",X"D1",X"87",X"5C",X"41",X"C5",X"9F",X"71",X"35",X"A8",X"B9",
		X"67",X"4F",X"5F",X"CE",X"8A",X"43",X"C6",X"80",X"54",X"4A",X"B1",X"AE",X"87",X"50",X"4F",X"C6",
		X"9F",X"55",X"45",X"BB",X"AC",X"5C",X"41",X"A9",X"BE",X"5C",X"4C",X"72",X"D4",X"71",X"42",X"DA",
		X"20",X"CF",X"6C",X"3D",X"D5",X"8A",X"78",X"39",X"7B",X"BF",X"99",X"75",X"37",X"99",X"C7",X"28",
		X"7B",X"C3",X"91",X"58",X"46",X"9D",X"BB",X"88",X"60",X"40",X"9A",X"BB",X"8C",X"3B",X"6A",X"BA",
		X"AC",X"31",X"7F",X"C8",X"2F",X"78",X"DC",X"33",X"AE",X"80",X"34",X"EE",X"38",X"74",X"D5",X"1F",
		X"98",X"BA",X"82",X"58",X"4A",X"D6",X"86",X"56",X"49",X"F0",X"34",X"73",X"BD",X"9A",X"43",X"67",
		X"C3",X"8D",X"2E",X"8B",X"B9",X"40",X"C6",X"33",X"B7",X"A5",X"27",X"8A",X"BA",X"42",X"BF",X"8A",
		X"3A",X"6F",X"D1",X"5C",X"41",X"DF",X"6A",X"42",X"C3",X"A4",X"33",X"80",X"CC",X"5C",X"43",X"89",
		X"BE",X"96",X"53",X"4E",X"8D",X"D4",X"2E",X"BD",X"56",X"6C",X"DA",X"53",X"47",X"9C",X"C8",X"2A",
		X"75",X"B3",X"B0",X"2F",X"80",X"CA",X"2B",X"81",X"CD",X"35",X"7E",X"CE",X"32",X"81",X"CD",X"74",
		X"40",X"74",X"D8",X"4E",X"58",X"D3",X"85",X"4D",X"53",X"AE",X"B8",X"61",X"3D",X"9F",X"C3",X"30",
		X"86",X"D0",X"5E",X"47",X"7D",X"C6",X"91",X"4E",X"4E",X"A9",X"B9",X"6D",X"34",X"9F",X"B7",X"3F",
		X"C6",X"7A",X"37",X"81",X"C5",X"8C",X"33",X"88",X"D3",X"44",X"59",X"82",X"C8",X"88",X"42",X"61",
		X"AF",X"A2",X"44",X"D9",X"48",X"52",X"89",X"BC",X"99",X"2E",X"7E",X"B4",X"38",X"B7",X"9E",X"20",
		X"E4",X"56",X"63",X"D9",X"56",X"43",X"B1",X"B8",X"37",X"6B",X"D3",X"6D",X"31",X"C8",X"65",X"8D",
		X"B9",X"0B",X"BA",X"86",X"4D",X"D7",X"4E",X"4B",X"E7",X"3C",X"95",X"AD",X"1D",X"D8",X"72",X"35",
		X"B4",X"A5",X"2F",X"B3",X"B6",X"44",X"57",X"93",X"CB",X"67",X"3F",X"A1",X"C7",X"21",X"89",X"9C",
		X"5A",X"D8",X"20",X"A3",X"BA",X"25",X"89",X"AD",X"37",X"D8",X"5D",X"53",X"DC",X"77",X"43",X"70",
		X"E1",X"46",X"59",X"83",X"CC",X"6E",X"37",X"E7",X"56",X"4E",X"86",X"D3",X"27",X"9E",X"AA",X"44",
		X"C0",X"19",X"E9",X"54",X"63",X"DB",X"51",X"4D",X"88",X"CF",X"30",X"91",X"C5",X"66",X"35",X"C1",
		X"9C",X"33",X"79",X"A7",X"BA",X"53",X"41",X"DD",X"4B",X"73",X"D2",X"25",X"7F",X"BB",X"9D",X"37",
		X"68",X"A9",X"BD",X"3B",X"5C",X"CF",X"61",X"47",X"C9",X"9E",X"47",X"55",X"AF",X"96",X"5D",X"D0",
		X"28",X"7E",X"D3",X"48",X"51",X"C7",X"95",X"21",X"BB",X"A6",X"3A",X"67",X"C3",X"81",X"37",X"DE",
		X"7D",X"3F",X"72",X"AA",X"B4",X"15",X"DC",X"6C",X"47",X"D2",X"71",X"28",X"EB",X"2E",X"9F",X"93",
		X"6C",X"9C",X"37",X"DB",X"43",X"AC",X"37",X"D3",X"4F",X"AC",X"8D",X"1B",X"DF",X"7E",X"46",X"6B",
		X"BA",X"A5",X"35",X"73",X"CB",X"41",X"7E",X"C8",X"1D",X"D3",X"60",X"5F",X"DB",X"44",X"57",X"C2",
		X"A2",X"41",X"5B",X"AE",X"96",X"5E",X"CC",X"10",X"CF",X"83",X"31",X"DF",X"59",X"46",X"CC",X"87",
		X"28",X"D7",X"84",X"3D",X"7A",X"DD",X"3A",X"7B",X"C8",X"36",X"66",X"C8",X"60",X"9A",X"8F",X"29",
		X"A8",X"B3",X"83",X"1F",X"D6",X"81",X"33",X"C4",X"82",X"2A",X"D4",X"6B",X"70",X"CA",X"1B",X"A9",
		X"AB",X"22",X"AE",X"9E",X"49",X"D3",X"45",X"5A",X"A1",X"BB",X"70",X"27",X"E9",X"49",X"72",X"CC",
		X"38",X"67",X"B6",X"AD",X"41",X"57",X"B7",X"8C",X"39",X"E4",X"70",X"4B",X"63",X"C7",X"52",X"AE",
		X"8A",X"36",X"8A",X"BB",X"8E",X"2F",X"87",X"AB",X"B2",X"2D",X"72",X"94",X"CD",X"39",X"67",X"D9",
		X"2B",X"86",X"C8",X"50",X"4D",X"BC",X"A1",X"3F",X"6B",X"BC",X"7C",X"48",X"E0",X"20",X"BA",X"83",
		X"43",X"D4",X"26",X"BD",X"A2",X"3E",X"6C",X"CA",X"8A",X"38",X"7B",X"AF",X"AE",X"23",X"91",X"C0",
		X"37",X"76",X"A3",X"C2",X"39",X"63",X"D9",X"48",X"5A",X"93",X"C9",X"43",X"62",X"90",X"B1",X"37",
		X"D1",X"53",X"74",X"B1",X"37",X"F6",X"23",X"82",X"C3",X"52",X"4A",X"BB",X"75",X"95",X"88",X"3D",
		X"90",X"C3",X"76",X"3B",X"87",X"A9",X"70",X"A6",X"61",X"4F",X"AE",X"B6",X"50",X"4B",X"E2",X"4A",
		X"63",X"DC",X"3E",X"63",X"92",X"CC",X"4F",X"4D",X"E3",X"4A",X"5B",X"89",X"D0",X"47",X"5E",X"90",
		X"D0",X"49",X"5B",X"7E",X"C6",X"76",X"3E",X"8C",X"AA",X"A4",X"15",X"CD",X"89",X"43",X"80",X"BD",
		X"65",X"A8",X"3D",X"8E",X"CF",X"0B",X"C0",X"8E",X"46",X"76",X"C9",X"7A",X"3E",X"88",X"AA",X"A8",
		X"18",X"BF",X"9C",X"2E",X"C3",X"85",X"2B",X"DC",X"6C",X"45",X"DB",X"4B",X"5F",X"92",X"AD",X"3D",
		X"C3",X"4F",X"86",X"A6",X"75",X"81",X"36",X"E7",X"37",X"A6",X"7D",X"A5",X"5A",X"58",X"D8",X"4E",
		X"56",X"AB",X"8E",X"49",X"DD",X"68",X"40",X"8A",X"B0",X"53",X"C3",X"4F",X"60",X"92",X"C6",X"51",
		X"54",X"9A",X"C5",X"55",X"4D",X"93",X"C2",X"70",X"2F",X"E3",X"50",X"5B",X"8D",X"AF",X"48",X"AA",
		X"81",X"98",X"4C",X"65",X"C1",X"66",X"BB",X"23",X"B0",X"9B",X"39",X"83",X"A4",X"B3",X"1A",X"B0",
		X"9D",X"31",X"C3",X"8E",X"2B",X"E2",X"54",X"5A",X"DC",X"32",X"86",X"CA",X"14",X"C9",X"83",X"43",
		X"83",X"AD",X"A6",X"15",X"DA",X"6D",X"4C",X"87",X"AF",X"63",X"B9",X"3A",X"8C",X"C5",X"0D",X"CC",
		X"79",X"58",X"74",X"C9",X"7D",X"42",X"7C",X"B7",X"5C",X"A9",X"7B",X"41",X"93",X"B6",X"81",X"32",
		X"9D",X"92",X"6B",X"87",X"9D",X"94",X"4A",X"6C",X"B7",X"A4",X"1B",X"BD",X"88",X"4D",X"7D",X"BD",
		X"4D",X"99",X"8A",X"51",X"CF",X"1B",X"F2",X"56",X"5A",X"72",X"C3",X"4B",X"BE",X"63",X"52",X"E1",
		X"2F",X"77",X"91",X"93",X"52",X"C0",X"37",X"E1",X"53",X"5A",X"DA",X"35",X"77",X"85",X"D5",X"39",
		X"6D",X"80",X"D3",X"50",X"58",X"D3",X"2D",X"9A",X"B2",X"23",X"BC",X"8C",X"52",X"71",X"C1",X"8D",
		X"3E",X"76",X"B3",X"6F",X"6D",X"A1",X"49",X"C9",X"2E",X"D1",X"38",X"C6",X"55",X"8B",X"7C",X"86",
		X"B2",X"33",X"7E",X"AD",X"99",X"3C",X"80",X"A3",X"6E",X"88",X"98",X"50",X"AA",X"79",X"99",X"27",
		X"FB",X"1D",X"AE",X"63",X"8F",X"94",X"51",X"B0",X"4A",X"AD",X"86",X"8B",X"39",X"EA",X"1B",X"AB",
		X"9A",X"4C",X"73",X"B8",X"9A",X"3A",X"76",X"AC",X"64",X"88",X"8B",X"6D",X"A6",X"71",X"97",X"40",
		X"8C",X"B5",X"4A",X"A0",X"68",X"86",X"8C",X"98",X"69",X"59",X"DE",X"1F",X"AB",X"A0",X"36",X"A8",
		X"A7",X"28",X"E0",X"58",X"59",X"CE",X"37",X"82",X"C8",X"2E",X"A4",X"5A",X"AF",X"62",X"8E",X"C2",
		X"2D",X"79",X"91",X"C2",X"2A",X"96",X"77",X"8A",X"99",X"8E",X"3D",X"C7",X"61",X"57",X"9D",X"A3",
		X"44",X"DE",X"34",X"88",X"B1",X"37",X"89",X"A3",X"B3",X"15",X"CB",X"73",X"43",X"BA",X"8D",X"47",
		X"9D",X"6F",X"C9",X"15",X"D1",X"72",X"53",X"CA",X"48",X"6B",X"9B",X"89",X"6A",X"A0",X"57",X"BE",
		X"45",X"9C",X"A5",X"5E",X"54",X"CA",X"63",X"52",X"E1",X"25",X"AE",X"93",X"35",X"E5",X"2A",X"A5",
		X"97",X"40",X"8A",X"9A",X"73",X"81",X"8E",X"57",X"CC",X"68",X"67",X"5D",X"C5",X"94",X"43",X"6E",
		X"AA",X"A8",X"30",X"9D",X"6E",X"B3",X"6B",X"4B",X"AB",X"79",X"90",X"93",X"50",X"89",X"81",X"8A",
		X"A4",X"42",X"9B",X"7F",X"67",X"9F",X"A8",X"48",X"80",X"BA",X"23",X"C5",X"6A",X"5E",X"91",X"99",
		X"62",X"9A",X"91",X"6A",X"5A",X"D9",X"3D",X"81",X"B2",X"34",X"C5",X"7A",X"3F",X"BB",X"90",X"3D",
		X"D0",X"50",X"65",X"95",X"94",X"63",X"C6",X"2D",X"A6",X"91",X"3D",X"CA",X"5F",X"66",X"91",X"97",
		X"A6",X"35",X"A6",X"97",X"2E",X"D9",X"41",X"8F",X"A4",X"3E",X"A2",X"B0",X"2E",X"B5",X"7A",X"55",
		X"C9",X"3F",X"84",X"C3",X"42",X"8A",X"72",X"9F",X"65",X"95",X"72",X"84",X"8A",X"58",X"C6",X"73",
		X"47",X"D9",X"35",X"90",X"9F",X"4D",X"80",X"A8",X"A1",X"30",X"8F",X"8B",X"C5",X"18",X"B5",X"70",
		X"65",X"B0",X"5D",X"93",X"93",X"7B",X"48",X"CB",X"52",X"7D",X"B0",X"3D",X"98",X"BA",X"2E",X"AD",
		X"86",X"4A",X"BD",X"6E",X"4C",X"DA",X"53",X"78",X"77",X"96",X"75",X"83",X"82",X"82",X"A5",X"3D",
		X"86",X"A2",X"A7",X"31",X"8B",X"8E",X"C3",X"20",X"AA",X"92",X"3A",X"C0",X"87",X"51",X"77",X"AD",
		X"62",X"B9",X"4F",X"7F",X"BC",X"1E",X"BF",X"7E",X"51",X"C3",X"50",X"72",X"C0",X"49",X"8A",X"81",
		X"72",X"AA",X"7B",X"55",X"8C",X"83",X"CA",X"2B",X"97",X"9C",X"4B",X"86",X"9F",X"B0",X"14",X"EA",
		X"3C",X"8A",X"9B",X"51",X"C2",X"25",X"C7",X"70",X"5F",X"AF",X"52",X"C6",X"29",X"B8",X"7F",X"5F",
		X"A3",X"5C",X"CB",X"26",X"AE",X"8B",X"3C",X"D6",X"48",X"8A",X"74",X"A2",X"8D",X"3F",X"D3",X"2A",
		X"B9",X"7B",X"4D",X"A6",X"69",X"B6",X"6E",X"56",X"8A",X"A1",X"64",X"C3",X"28",X"B2",X"7D",X"60",
		X"A6",X"58",X"D4",X"11",X"D1",X"5C",X"7A",X"A8",X"42",X"96",X"C7",X"27",X"A9",X"90",X"44",X"89",
		X"9F",X"69",X"90",X"A7",X"25",X"DB",X"46",X"7C",X"B7",X"42",X"9A",X"6E",X"99",X"8C",X"81",X"41",
		X"C7",X"7A",X"58",X"8D",X"83",X"B2",X"29",X"C1",X"6E",X"52",X"DA",X"44",X"83",X"B6",X"2A",X"C4",
		X"41",X"A6",X"7A",X"76",X"98",X"5B",X"B6",X"86",X"42",X"A2",X"8A",X"4B",X"95",X"97",X"65",X"B7",
		X"56",X"6C",X"D2",X"1E",X"B6",X"94",X"36",X"DD",X"38",X"96",X"7B",X"70",X"9E",X"95",X"59",X"77",
		X"82",X"8D",X"7C",X"78",X"DC",X"01",X"CD",X"70",X"5D",X"76",X"B4",X"91",X"35",X"BD",X"48",X"D3",
		X"36",X"8E",X"B7",X"2C",X"BE",X"49",X"CA",X"4C",X"72",X"CB",X"29",X"B9",X"82",X"3B",X"CC",X"71",
		X"4B",X"D1",X"4F",X"6A",X"8D",X"C9",X"46",X"6A",X"CA",X"28",X"99",X"A9",X"61",X"59",X"AA",X"78",
		X"8F",X"98",X"35",X"CE",X"64",X"58",X"95",X"A7",X"49",X"AC",X"57",X"9B",X"7C",X"70",X"DE",X"14",
		X"A9",X"A3",X"3F",X"7B",X"C9",X"57",X"5F",X"D6",X"17",X"C5",X"7D",X"58",X"9E",X"71",X"B8",X"3D",
		X"72",X"A7",X"6C",X"A7",X"80",X"3A",X"E5",X"22",X"A5",X"61",X"B6",X"86",X"38",X"D9",X"56",X"57",
		X"9A",X"8E",X"64",X"97",X"96",X"7D",X"45",X"CC",X"5D",X"5A",X"A8",X"AA",X"3C",X"7E",X"97",X"C1",
		X"22",X"9B",X"A7",X"45",X"7F",X"A1",X"B4",X"1D",X"BB",X"51",X"B9",X"7A",X"45",X"91",X"A5",X"67",
		X"B8",X"34",X"9E",X"A8",X"35",X"88",X"B0",X"54",X"A8",X"8C",X"31",X"E7",X"41",X"6A",X"C7",X"41",
		X"85",X"BA",X"2D",X"B1",X"A0",X"35",X"90",X"9F",X"75",X"A0",X"5D",X"52",X"CA",X"59",X"84",X"9A",
		X"52",X"B2",X"66",X"AF",X"43",X"6E",X"BC",X"59",X"89",X"95",X"8B",X"74",X"44",X"AE",X"85",X"96",
		X"7B",X"4A",X"8B",X"BD",X"7E",X"2F",X"D2",X"68",X"4D",X"D9",X"41",X"6F",X"CA",X"4D",X"62",X"A0",
		X"B7",X"3C",X"76",X"D1",X"2E",X"98",X"B1",X"2A",X"BB",X"8D",X"2F",X"E2",X"4A",X"6C",X"C4",X"49",
		X"64",X"A5",X"88",X"80",X"9E",X"2A",X"DD",X"59",X"54",X"CE",X"60",X"54",X"9E",X"9D",X"42",X"BF",
		X"92",X"34",X"98",X"B7",X"40",X"77",X"9F",X"BC",X"28",X"93",X"B8",X"44",X"67",X"A7",X"AC",X"41",
		X"6F",X"9F",X"91",X"50",X"C4",X"37",X"B1",X"7A",X"5B",X"DD",X"4C",X"58",X"C6",X"5D",X"51",X"BA",
		X"82",X"47",X"D6",X"6B",X"45",X"AC",X"60",X"C5",X"3D",X"7D",X"CA",X"33",X"8D",X"AE",X"42",X"88",
		X"CB",X"4F",X"5D",X"84",X"C3",X"31",X"B4",X"6B",X"6C",X"AD",X"73",X"AB",X"23",X"D5",X"6B",X"43",
		X"D1",X"6A",X"47",X"CB",X"4B",X"77",X"C4",X"2B",X"BC",X"94",X"35",X"C6",X"77",X"3E",X"9E",X"94",
		X"77",X"A5",X"43",X"7C",X"99",X"BD",X"3A",X"79",X"C8",X"2B",X"B8",X"83",X"37",X"D2",X"77",X"4F",
		X"78",X"BD",X"43",X"AC",X"80",X"66",X"C8",X"28",X"89",X"A3",X"AF",X"2A",X"92",X"B9",X"3D",X"80",
		X"CC",X"27",X"9A",X"B0",X"48",X"66",X"AD",X"8D",X"44",X"D0",X"6A",X"44",X"AA",X"87",X"6B",X"C7",
		X"25",X"A3",X"AB",X"41",X"70",X"AD",X"71",X"9C",X"74",X"45",X"C9",X"91",X"51",X"5D",X"D9",X"4E",
		X"62",X"C7",X"61",X"4C",X"A4",X"97",X"78",X"95",X"3D",X"9E",X"A8",X"30",X"D4",X"4B",X"81",X"B2",
		X"33",X"C5",X"65",X"A4",X"63",X"4E",X"A8",X"98",X"5F",X"C0",X"30",X"96",X"B5",X"3D",X"75",X"B2",
		X"92",X"31",X"B1",X"A5",X"33",X"A4",X"AD",X"43",X"68",X"B4",X"7A",X"51",X"DB",X"45",X"74",X"C9",
		X"2D",X"95",X"AD",X"3B",X"8E",X"A9",X"3D",X"C0",X"70",X"62",X"D5",X"27",X"A7",X"9E",X"3F",X"7C",
		X"BC",X"50",X"A4",X"8E",X"34",X"A3",X"A1",X"4E",X"99",X"BC",X"35",X"7B",X"BD",X"67",X"45",X"AA",
		X"94",X"62",X"C1",X"3E",X"74",X"CB",X"41",X"74",X"A3",X"50",X"B6",X"9F",X"47",X"68",X"A6",X"AF",
		X"4A",X"62",X"94",X"AC",X"3F",X"AD",X"A9",X"3F",X"72",X"8A",X"C7",X"54",X"5E",X"7A",X"C0",X"80",
		X"4D",X"6B",X"B7",X"71",X"86",X"9F",X"2C",X"DC",X"60",X"59",X"79",X"BB",X"7C",X"40",X"A8",X"AC",
		X"63",X"48",X"D4",X"67",X"56",X"79",X"B8",X"8D",X"38",X"BE",X"7E",X"3C",X"B0",X"97",X"54",X"C2",
		X"37",X"98",X"B4",X"32",X"90",X"B9",X"4F",X"5E",X"B2",X"A0",X"34",X"9F",X"A3",X"35",X"AD",X"9B",
		X"38",X"BB",X"97",X"4E",X"64",X"A4",X"94",X"53",X"D0",X"45",X"6A",X"C2",X"6E",X"42",X"CC",X"77",
		X"52",X"73",X"BB",X"61",X"89",X"B2",X"2D",X"9C",X"B4",X"43",X"77",X"C5",X"57",X"59",X"93",X"A6",
		X"5B",X"B6",X"50",X"63",X"BE",X"8D",X"4D",X"6A",X"A2",X"AA",X"6F",X"3F",X"C2",X"86",X"4B",X"75",
		X"BD",X"76",X"4B",X"D2",X"5A",X"5A",X"8A",X"BF",X"5B",X"56",X"B3",X"9F",X"4E",X"66",X"C4",X"5D",
		X"51",X"C0",X"68",X"70",X"C1",X"3E",X"75",X"BB",X"50",X"A6",X"88",X"3A",X"AB",X"A4",X"79",X"3A",
		X"BC",X"8E",X"4A",X"74",X"B7",X"82",X"42",X"D2",X"5F",X"5A",X"7F",X"B4",X"8D",X"41",X"86",X"C0",
		X"55",X"5F",X"C0",X"44",X"96",X"B6",X"5A",X"5A",X"84",X"BD",X"78",X"52",X"6C",X"BA",X"82",X"41",
		X"BD",X"83",X"3E",X"A9",X"91",X"56",X"CA",X"38",X"95",X"AA",X"39",X"8B",X"AE",X"4D",X"8C",X"AC",
		X"35",X"BC",X"79",X"52",X"C1",X"5A",X"80",X"C2",X"41",X"73",X"A8",X"4C",X"B1",X"9C",X"63",X"4F",
		X"BB",X"8B",X"4B",X"70",X"B2",X"7F",X"46",X"D3",X"48",X"A3",X"94",X"3D",X"94",X"B6",X"52",X"61",
		X"BD",X"49",X"91",X"B9",X"58",X"61",X"77",X"BD",X"4D",X"A9",X"84",X"43",X"CF",X"6A",X"58",X"74",
		X"C2",X"57",X"93",X"61",X"84",X"BB",X"2E",X"B6",X"86",X"4B",X"C7",X"71",X"54",X"76",X"AF",X"73",
		X"5D",X"D2",X"40",X"85",X"B7",X"59",X"5A",X"94",X"AF",X"40",X"9D",X"A1",X"32",X"BD",X"71",X"72",
		X"BC",X"51",X"60",X"97",X"AC",X"7F",X"47",X"8D",X"B7",X"57",X"5B",X"C1",X"7B",X"52",X"73",X"AB",
		X"8B",X"44",X"C1",X"82",X"42",X"BD",X"75",X"4B",X"B0",X"9D",X"6A",X"50",X"8A",X"AD",X"8E",X"53",
		X"65",X"9C",X"AE",X"65",X"51",X"AF",X"99",X"43",X"80",X"B4",X"7E",X"3D",X"B9",X"6B",X"66",X"C2",
		X"45",X"B4",X"81",X"50",X"72",X"BC",X"6E",X"4E",X"BA",X"7A",X"4A",X"C1",X"6F",X"5A",X"BB",X"89",
		X"5C",X"5E",X"9B",X"AF",X"5E",X"5C",X"CA",X"43",X"87",X"B0",X"41",X"85",X"BA",X"4D",X"77",X"BA",
		X"76",X"4A",X"A7",X"9D",X"54",X"61",X"AA",X"9C",X"47",X"7B",X"B2",X"8B",X"51",X"6C",X"9A",X"A4",
		X"42",X"A4",X"A6",X"3A",X"A5",X"97",X"3F",X"9E",X"A7",X"78",X"4E",X"7F",X"B1",X"8A",X"58",X"64",
		X"B8",X"88",X"48",X"87",X"B5",X"6E",X"49",X"BE",X"59",X"93",X"A5",X"46",X"74",X"9E",X"A3",X"35",
		X"C2",X"72",X"55",X"C2",X"5B",X"60",X"B9",X"79",X"48",X"C8",X"57",X"84",X"B1",X"4B",X"6C",X"97",
		X"AC",X"3F",X"8C",X"AF",X"47",X"AF",X"89",X"4A",X"7D",X"A4",X"9E",X"4F",X"6A",X"B1",X"8E",X"45",
		X"88",X"B2",X"70",X"4B",X"A7",X"9C",X"41",X"AD",X"96",X"49",X"7B",X"B6",X"77",X"4B",X"B4",X"8D",
		X"56",X"67",X"A2",X"A0",X"3E",X"B2",X"84",X"45",X"AC",X"9A",X"78",X"44",X"B1",X"80",X"52",X"C9",
		X"4B",X"7E",X"B7",X"3C",X"A1",X"99",X"40",X"9F",X"A3",X"7C",X"4C",X"8A",X"B0",X"76",X"4C",X"9D",
		X"A6",X"3F",X"9C",X"A5",X"5E",X"5C",X"B7",X"85",X"4E",X"7E",X"B4",X"6A",X"56",X"CD",X"4B",X"99",
		X"6F",X"69",X"C4",X"45",X"89",X"B2",X"60",X"60",X"7F",X"BB",X"57",X"6E",X"B4",X"84",X"66",X"59",
		X"BD",X"4A",X"9F",X"A0",X"5B",X"5F",X"A1",X"A4",X"65",X"57",X"94",X"A3",X"8E",X"46",X"8A",X"9B",
		X"58",X"B7",X"78",X"4C",X"9B",X"A1",X"40",X"AF",X"87",X"42",X"B4",X"80",X"5E",X"BB",X"4B",X"7D",
		X"BB",X"42",X"95",X"A1",X"42",X"AA",X"98",X"59",X"64",X"A4",X"A0",X"5F",X"5D",X"9C",X"A7",X"66",
		X"57",X"A0",X"A4",X"5E",X"61",X"8A",X"B4",X"4D",X"92",X"A5",X"55",X"68",X"8F",X"B1",X"55",X"6C",
		X"BE",X"51",X"88",X"A6",X"36",X"C2",X"6C",X"60",X"B2",X"84",X"4D",X"84",X"A8",X"4A",X"A5",X"9E",
		X"60",X"5D",X"AD",X"92",X"76",X"4E",X"94",X"A8",X"72",X"4C",X"B0",X"7A",X"57",X"B8",X"85",X"72",
		X"51",X"C2",X"59",X"6C",X"B1",X"86",X"69",X"5A",X"92",X"A9",X"7B",X"50",X"8B",X"B3",X"41",X"AD",
		X"6F",X"61",X"B7",X"82",X"6E",X"55",X"A0",X"9F",X"4B",X"87",X"B1",X"52",X"9B",X"96",X"59",X"68",
		X"B7",X"55",X"85",X"B1",X"64",X"65",X"70",X"BB",X"6A",X"5F",X"B0",X"8A",X"76",X"55",X"82",X"AE",
		X"82",X"5F",X"66",X"A1",X"9C",X"48",X"B7",X"67",X"60",X"B8",X"76",X"4D",X"B7",X"76",X"62",X"B1",
		X"7C",X"55",X"84",X"AD",X"77",X"55",X"8B",X"AC",X"40",X"9A",X"A1",X"75",X"57",X"7D",X"A6",X"91",
		X"75",X"5C",X"74",X"AE",X"7D",X"52",X"C1",X"58",X"74",X"B7",X"45",X"95",X"A1",X"70",X"57",X"89",
		X"AA",X"81",X"5B",X"6D",X"9F",X"9E",X"6F",X"57",X"AB",X"8E",X"63",X"5E",X"B0",X"80",X"4E",X"B1",
		X"88",X"4C",X"9E",X"9A",X"46",X"98",X"A4",X"6C",X"55",X"B0",X"84",X"56",X"B8",X"48",X"92",X"A3",
		X"7D",X"69",X"5C",X"A6",X"98",X"51",X"83",X"B5",X"4C",X"8E",X"A3",X"69",X"5E",X"80",X"AF",X"6B",
		X"5B",X"B3",X"7C",X"52",X"B1",X"88",X"81",X"50",X"88",X"A7",X"83",X"54",X"82",X"AB",X"46",X"9F",
		X"9F",X"4B",X"94",X"9F",X"42",X"A8",X"92",X"84",X"59",X"77",X"B3",X"46",X"A5",X"8C",X"4A",X"AE",
		X"8A",X"59",X"A9",X"82",X"67",X"60",X"99",X"9F",X"81",X"6A",X"5B",X"BF",X"4F",X"9C",X"82",X"54",
		X"BA",X"75",X"55",X"A7",X"8A",X"4B",X"A4",X"96",X"82",X"61",X"67",X"9A",X"9E",X"4D",X"8A",X"A7",
		X"7F",X"73",X"52",X"BB",X"60",X"73",X"AC",X"83",X"73",X"59",X"89",X"A4",X"88",X"50",X"95",X"A2",
		X"67",X"63",X"7D",X"B0",X"72",X"59",X"A9",X"8F",X"50",X"87",X"AC",X"47",X"9C",X"97",X"7B",X"53",
		X"92",X"A0",X"7B",X"5B",X"7F",X"B1",X"49",X"8D",X"A4",X"7B",X"66",X"62",X"B4",X"76",X"66",X"AA",
		X"81",X"62",X"6D",X"AF",X"80",X"6D",X"5C",X"97",X"9C",X"86",X"69",X"60",X"AE",X"80",X"4E",X"B9",
		X"66",X"6D",X"AA",X"83",X"64",X"69",X"AD",X"86",X"6B",X"60",X"8C",X"AA",X"65",X"66",X"AF",X"80",
		X"51",X"9A",X"9B",X"7B",X"72",X"57",X"A5",X"92",X"87",X"67",X"66",X"86",X"B2",X"58",X"8E",X"8B",
		X"5F",X"B0",X"71",X"6B",X"63",X"A7",X"8F",X"85",X"67",X"63",X"B2",X"61",X"6F",X"AE",X"81",X"7F",
		X"4E",X"A4",X"8D",X"51",X"9F",X"99",X"73",X"62",X"75",X"B6",X"66",X"79",X"9F",X"50",X"B7",X"4C",
		X"8E",X"9E",X"7D",X"5C",X"7F",X"AF",X"4B",X"8D",X"A1",X"7D",X"65",X"66",X"AE",X"7B",X"62",X"AD",
		X"7B",X"6C",X"5F",X"A8",X"8D",X"84",X"66",X"65",X"A7",X"8D",X"75",X"58",X"9F",X"97",X"74",X"60",
		X"79",X"A4",X"8E",X"6A",X"5F",X"A7",X"8D",X"53",X"A7",X"87",X"73",X"57",X"B1",X"74",X"68",X"AD",
		X"48",X"A0",X"94",X"81",X"6D",X"5F",X"94",X"9C",X"85",X"6D",X"5F",X"97",X"9D",X"78",X"5B",X"87",
		X"AA",X"5E",X"6C",X"A6",X"8A",X"7A",X"5D",X"7B",X"9E",X"96",X"59",X"7D",X"AB",X"4C",X"98",X"95",
		X"4B",X"A5",X"8B",X"55",X"A5",X"8D",X"71",X"60",X"84",X"A4",X"84",X"7F",X"5A",X"82",X"AB",X"5B",
		X"78",X"B2",X"5B",X"7F",X"A2",X"4D",X"94",X"A2",X"51",X"98",X"93",X"78",X"57",X"9B",X"95",X"7D",
		X"57",X"90",X"9D",X"53",X"A2",X"8D",X"6C",X"65",X"81",X"AD",X"68",X"71",X"A9",X"53",X"A4",X"82",
		X"7A",X"55",X"A4",X"88",X"53",X"A5",X"8D",X"7F",X"6A",X"63",X"A7",X"87",X"59",X"A5",X"8A",X"77",
		X"61",X"7B",X"AD",X"73",X"6B",X"A1",X"7F",X"6F",X"60",X"B2",X"6C",X"66",X"AA",X"82",X"81",X"5E",
		X"75",X"9D",X"92",X"7D",X"6C",X"63",X"B0",X"73",X"60",X"A8",X"86",X"80",X"62",X"71",X"99",X"9A",
		X"50",X"97",X"92",X"51",X"9D",X"96",X"51",X"A5",X"79",X"5D",X"AA",X"85",X"80",X"64",X"6D",X"AB",
		X"77",X"64",X"A9",X"82",X"77",X"5F",X"85",X"A1",X"85",X"7F",X"5B",X"88",X"A4",X"4E",X"95",X"98",
		X"81",X"69",X"69",X"B1",X"55",X"90",X"99",X"4F",X"A7",X"7E",X"59",X"AA",X"7C",X"5B",X"9E",X"92",
		X"7E",X"70",X"5F",X"A1",X"8F",X"85",X"5F",X"78",X"A6",X"7F",X"77",X"5A",X"A0",X"87",X"58",X"A0",
		X"93",X"59",X"97",X"94",X"5B",X"76",X"9F",X"8E",X"63",X"72",X"AC",X"57",X"81",X"A6",X"66",X"68",
		X"A7",X"83",X"5C",X"A7",X"80",X"7A",X"59",X"97",X"9A",X"5D",X"7A",X"AD",X"66",X"72",X"A1",X"80",
		X"70",X"62",X"A7",X"85",X"7B",X"5F",X"7E",X"9D",X"8E",X"73",X"5F",X"93",X"9D",X"63",X"6D",X"AA",
		X"7B",X"89",X"5B",X"7F",X"A0",X"84",X"64",X"78",X"A5",X"7A",X"75",X"5E",X"9C",X"93",X"7F",X"7C",
		X"58",X"A0",X"8D",X"80",X"61",X"77",X"9D",X"91",X"65",X"71",X"A4",X"80",X"76",X"5E",X"A4",X"89",
		X"7C",X"62",X"78",X"9D",X"8D",X"7D",X"6C",X"68",X"B0",X"69",X"78",X"A3",X"54",X"9F",X"8A",X"79",
		X"63",X"7A",X"9E",X"8D",X"64",X"71",X"AD",X"6D",X"6D",X"9D",X"86",X"6F",X"68",X"82",X"A8",X"6A",
		X"74",X"A2",X"7A",X"73",X"61",X"B1",X"66",X"73",X"A8",X"5C",X"7D",X"A7",X"6C",X"6C",X"AA",X"56",
		X"97",X"89",X"55",X"A7",X"85",X"85",X"6E",X"66",X"A6",X"82",X"82",X"5F",X"81",X"A5",X"55",X"8A",
		X"9C",X"7C",X"81",X"5B",X"8A",X"9F",X"5E",X"7E",X"A9",X"5D",X"79",X"9E",X"87",X"61",X"76",X"9E",
		X"8C",X"65",X"72",X"A2",X"83",X"78",X"60",X"A2",X"86",X"7C",X"5E",X"9B",X"8C",X"56",X"AD",X"66",
		X"71",X"A3",X"81",X"82",X"66",X"74",X"AE",X"5E",X"82",X"9B",X"58",X"8E",X"9E",X"63",X"72",X"A1",
		X"84",X"72",X"62",X"9F",X"8B",X"81",X"73",X"65",X"89",X"9D",X"7F",X"84",X"5E",X"84",X"9E",X"7C",
		X"7B",X"5E",X"8B",X"96",X"8C",X"56",X"96",X"90",X"80",X"66",X"74",X"9A",X"92",X"61",X"78",X"9E",
		X"87",X"69",X"72",X"A2",X"7F",X"76",X"63",X"8B",X"9A",X"83",X"5B",X"8F",X"98",X"7B",X"7F",X"5B",
		X"92",X"98",X"5A",X"9D",X"86",X"81",X"62",X"80",X"A0",X"7B",X"76",X"61",X"9A",X"91",X"80",X"7B",
		X"5E",X"91",X"96",X"7F",X"6E",X"69",X"99",X"94",X"64",X"75",X"A6",X"74",X"64",X"8F",X"9D",X"65",
		X"72",X"A1",X"83",X"74",X"62",X"9F",X"89",X"82",X"72",X"67",X"88",X"9D",X"7A",X"62",X"AC",X"5A",
		X"8F",X"90",X"7F",X"6E",X"6B",X"8E",X"9D",X"61",X"86",X"9B",X"56",X"9D",X"88",X"7C",X"64",X"7B",
		X"99",X"8E",X"5E",X"7F",X"9F",X"7F",X"83",X"63",X"7D",X"A5",X"6A",X"6C",X"99",X"8F",X"57",X"A1",
		X"7C",X"68",X"9C",X"86",X"6B",X"72",X"A2",X"7B",X"81",X"5C",X"98",X"90",X"77",X"61",X"A5",X"71",
		X"6B",X"A0",X"87",X"73",X"68",X"A2",X"80",X"80",X"63",X"7D",X"9E",X"81",X"60",X"A2",X"77",X"69",
		X"A8",X"6B",X"6D",X"9D",X"83",X"7E",X"65",X"7C",X"9D",X"86",X"62",X"80",X"A1",X"6F",X"68",X"A0",
		X"83",X"84",X"6C",X"6E",X"92",X"9A",X"5D",X"8C",X"8F",X"5F",X"A1",X"7F",X"7F",X"65",X"7B",X"98",
		X"8C",X"61",X"7C",X"A1",X"78",X"66",X"A3",X"68",X"75",X"A3",X"7A",X"87",X"69",X"70",X"8E",X"97",
		X"7C",X"62",X"93",X"90",X"79",X"6B",X"74",X"A0",X"83",X"63",X"87",X"9E",X"6D",X"70",X"A1",X"60",
		X"8E",X"91",X"7A",X"73",X"68",X"97",X"8E",X"84",X"73",X"68",X"8D",X"9A",X"75",X"66",X"9E",X"7F",
		X"60",X"9A",X"8E",X"61",X"8D",X"92",X"57",X"96",X"8E",X"81",X"79",X"65",X"9C",X"87",X"7A",X"67",
		X"80",X"9E",X"7D",X"85",X"64",X"7B",X"9B",X"85",X"72",X"68",X"98",X"8F",X"74",X"66",X"9A",X"89",
		X"5D",X"8D",X"96",X"7C",X"60",X"A1",X"7C",X"69",X"9D",X"81",X"78",X"65",X"A2",X"78",X"69",X"A8",
		X"62",X"83",X"95",X"7E",X"76",X"67",X"8B",X"97",X"7B",X"61",X"A7",X"6B",X"76",X"9C",X"7F",X"77",
		X"66",X"91",X"95",X"77",X"64",X"98",X"8E",X"64",X"7B",X"9D",X"7F",X"61",X"94",X"8F",X"7C",X"66",
		X"82",X"9D",X"7A",X"87",X"66",X"7A",X"A0",X"6E",X"6D",X"A0",X"7F",X"84",X"71",X"6B",X"9E",X"83",
		X"7E",X"62",X"90",X"92",X"7B",X"79",X"62",X"A4",X"79",X"70",X"99",X"84",X"62",X"8B",X"92",X"7F",
		X"74",X"6B",X"8A",X"99",X"75",X"68",X"99",X"8C",X"68",X"77",X"9D",X"7D",X"83",X"6F",X"6D",X"91",
		X"91",X"83",X"6F",X"6E",X"99",X"8C",X"69",X"76",X"9F",X"79",X"68",X"A1",X"70",X"6D",X"9B",X"86",
		X"60",X"9C",X"7C",X"6A",X"9F",X"7B",X"84",X"65",X"81",X"A0",X"61",X"89",X"91",X"7D",X"7B",X"65",
		X"8D",X"95",X"7E",X"83",X"70",X"6D",X"A3",X"73",X"70",X"A1",X"67",X"7F",X"9C",X"5A",X"98",X"7F",
		X"6B",X"A0",X"78",X"87",X"60",X"8A",X"95",X"7C",X"81",X"61",X"94",X"8E",X"7F",X"7A",X"67",X"88",
		X"93",X"88",X"6F",X"71",X"A0",X"67",X"78",X"98",X"88",X"6D",X"72",X"9E",X"7E",X"83",X"78",X"67",
		X"8D",X"92",X"82",X"63",X"8F",X"8F",X"7D",X"7A",X"66",X"8F",X"93",X"7B",X"66",X"A3",X"6B",X"7B",
		X"97",X"7E",X"74",X"6B",X"9B",X"86",X"7F",X"80",X"66",X"82",X"95",X"87",X"62",X"88",X"95",X"7D",
		X"82",X"6B",X"77",X"99",X"86",X"66",X"91",X"8C",X"74",X"6C",X"98",X"85",X"7B",X"66",X"97",X"87",
		X"80",X"74",X"6D",X"8C",X"96",X"73",X"70",X"A1",X"64",X"7A",X"93",X"8D",X"64",X"80",X"96",X"82",
		X"6F",X"71",X"99",X"87",X"65",X"82",X"98",X"7F",X"82",X"71",X"6F",X"92",X"8D",X"83",X"6E",X"73",
		X"95",X"8C",X"6E",X"74",X"9A",X"7E",X"82",X"69",X"7E",X"9F",X"62",X"88",X"91",X"64",X"8F",X"8F",
		X"65",X"7E",X"96",X"83",X"63",X"8D",X"90",X"7F",X"7D",X"67",X"98",X"85",X"7E",X"66",X"92",X"8B",
		X"7C",X"6C",X"7C",X"9B",X"7C",X"69",X"94",X"86",X"7F",X"72",X"6F",X"8F",X"91",X"78",X"68",X"97",
		X"89",X"7B",X"67",X"97",X"86",X"80",X"74",X"6C",X"94",X"8C",X"7E",X"82",X"6B",X"7C",X"9F",X"67",
		X"82",X"96",X"6A",X"77",X"9A",X"7E",X"83",X"78",X"69",X"98",X"86",X"81",X"74",X"6D",X"8C",X"91",
		X"81",X"7A",X"69",X"99",X"80",X"65",X"90",X"8F",X"7D",X"66",X"96",X"87",X"7F",X"67",X"8D",X"8F",
		X"61",X"98",X"7F",X"67",X"8E",X"90",X"7D",X"82",X"69",X"7D",X"96",X"86",X"6A",X"7D",X"9D",X"6F",
		X"76",X"99",X"6E",X"71",X"99",X"83",X"83",X"71",X"71",X"8F",X"91",X"71",X"72",X"9A",X"7D",X"84",
		X"6A",X"7A",X"8C",X"94",X"6B",X"7D",X"94",X"7F",X"6D",X"79",X"97",X"84",X"67",X"85",X"93",X"81",
		X"73",X"74",X"9B",X"7A",X"84",X"68",X"80",X"97",X"7E",X"83",X"69",X"82",X"99",X"69",X"82",X"97",
		X"65",X"87",X"91",X"63",X"93",X"86",X"7F",X"76",X"6C",X"94",X"89",X"82",X"6D",X"78",X"96",X"86",
		X"69",X"80",X"97",X"79",X"6D",X"97",X"7D",X"6A",X"9A",X"76",X"6D",X"98",X"83",X"81",X"7D",X"6C",
		X"80",X"93",X"87",X"65",X"96",X"83",X"81",X"78",X"6B",X"99",X"82",X"82",X"73",X"70",X"91",X"8D",
		X"7C",X"84",X"69",X"80",X"97",X"7B",X"85",X"6C",X"79",X"92",X"8B",X"73",X"71",X"9B",X"75",X"6E",
		X"91",X"8E",X"70",X"73",X"97",X"84",X"6B",X"80",X"98",X"77",X"70",X"95",X"7F",X"67",X"93",X"89",
		X"7F",X"7E",X"6B",X"83",X"95",X"7F",X"82",X"78",X"6C",X"98",X"83",X"81",X"79",X"6B",X"96",X"84",
		X"67",X"95",X"84",X"68",X"8E",X"8F",X"71",X"72",X"8F",X"8F",X"6B",X"80",X"93",X"7A",X"6B",X"91",
		X"87",X"65",X"90",X"8D",X"74",X"6E",X"93",X"89",X"7D",X"82",X"6B",X"7E",X"93",X"87",X"6B",X"7F",
		X"97",X"7A",X"86",X"6B",X"7E",X"95",X"7D",X"83",X"71",X"74",X"93",X"88",X"7F",X"7E",X"69",X"96",
		X"83",X"81",X"79",X"6C",X"8B",X"90",X"7D",X"83",X"77",X"6E",X"8A",X"92",X"77",X"71",X"98",X"78",
		X"6F",X"9B",X"6E",X"7D",X"94",X"7A",X"83",X"65",X"93",X"88",X"81",X"78",X"6F",X"86",X"96",X"71",
		X"79",X"94",X"7D",X"80",X"6C",X"7E",X"91",X"87",X"7E",X"80",X"6B",X"80",X"8F",X"8B",X"6B",X"7D",
		X"95",X"7D",X"83",X"72",X"73",X"92",X"88",X"80",X"6E",X"7C",X"95",X"80",X"6D",X"7F",X"95",X"7D",
		X"83",X"77",X"6E",X"92",X"88",X"7F",X"6F",X"7A",X"96",X"7F",X"6E",X"80",X"99",X"6B",X"7F",X"90",
		X"80",X"75",X"72",X"94",X"87",X"75",X"72",X"99",X"78",X"6F",X"8C",X"8F",X"6C",X"7C",X"92",X"80",
		X"78",X"6E",X"90",X"8C",X"72",X"73",X"96",X"81",X"81",X"6D",X"7F",X"95",X"7D",X"83",X"7B",X"6E",
		X"83",X"93",X"7E",X"83",X"6A",X"88",X"90",X"66",X"8C",X"8D",X"69",X"86",X"92",X"7B",X"85",X"70",
		X"76",X"8D",X"8E",X"70",X"78",X"96",X"7C",X"85",X"6F",X"79",X"98",X"74",X"71",X"90",X"89",X"7C",
		X"83",X"6B",X"83",X"91",X"80",X"80",X"70",X"79",X"90",X"88",X"7E",X"81",X"6E",X"7D",X"98",X"71",
		X"7B",X"93",X"7A",X"85",X"6B",X"80",X"92",X"81",X"80",X"71",X"79",X"99",X"74",X"78",X"93",X"7C",
		X"83",X"70",X"78",X"8D",X"8B",X"7E",X"80",X"6C",X"82",X"90",X"84",X"6A",X"8B",X"8C",X"7D",X"81",
		X"6B",X"8B",X"8F",X"6D",X"82",X"92",X"6C",X"7F",X"94",X"72",X"74",X"91",X"86",X"6D",X"82",X"93",
		X"69",X"82",X"91",X"80",X"6E",X"81",X"94",X"77",X"73",X"93",X"7C",X"6F",X"97",X"78",X"71",X"8B",
		X"8F",X"6C",X"82",X"8E",X"7D",X"81",X"6F",X"7C",X"8F",X"87",X"7E",X"80",X"6E",X"7E",X"8E",X"8A",
		X"70",X"78",X"95",X"7D",X"84",X"78",X"71",X"87",X"91",X"79",X"70",X"91",X"85",X"7C",X"6F",X"8B",
		X"8C",X"67",X"90",X"82",X"6F",X"91",X"84",X"76",X"72",X"8D",X"8D",X"70",X"7D",X"93",X"6F",X"7D",
		X"95",X"68",X"88",X"8B",X"80",X"78",X"73",X"96",X"7D",X"84",X"73",X"75",X"93",X"83",X"81",X"77",
		X"72",X"8E",X"8A",X"7E",X"80",X"6D",X"8C",X"8C",X"6A",X"83",X"8F",X"81",X"6D",X"85",X"8F",X"7E",
		X"6D",X"88",X"8D",X"7F",X"6F",X"82",X"91",X"7D",X"6F",X"85",X"8F",X"7D",X"7D",X"6D",X"90",X"88",
		X"7C",X"6E",X"94",X"80",X"70",X"8E",X"87",X"76",X"74",X"92",X"81",X"7D",X"6D",X"8F",X"87",X"7F",
		X"71",X"7C",X"92",X"81",X"73",X"7A",X"95",X"7C",X"84",X"7B",X"6F",X"8D",X"8A",X"7B",X"71",X"82",
		X"92",X"79",X"73",X"91",X"7E",X"6D",X"8D",X"89",X"7D",X"83",X"6D",X"84",X"8F",X"7D",X"83",X"70",
		X"7B",X"8B",X"8B",X"7B",X"85",X"71",X"7A",X"93",X"7E",X"82",X"75",X"75",X"89",X"8D",X"7D",X"6D",
		X"90",X"85",X"81",X"79",X"71",X"8D",X"8A",X"79",X"72",X"91",X"83",X"7D",X"6F",X"86",X"8E",X"7D",
		X"70",X"85",X"90",X"7A",X"86",X"74",X"76",X"91",X"82",X"81",X"79",X"72",X"87",X"8D",X"80",X"6D",
		X"86",X"8E",X"7E",X"82",X"76",X"74",X"89",X"8B",X"82",X"72",X"7F",X"94",X"6F",X"80",X"8D",X"7E",
		X"73",X"7B",X"92",X"7F",X"71",X"8A",X"89",X"6A",X"89",X"8B",X"81",X"71",X"7F",X"91",X"7C",X"84",
		X"79",X"72",X"8D",X"89",X"6C",X"8C",X"86",X"7F",X"7C",X"71",X"83",X"8D",X"83",X"7E",X"81",X"6E",
		X"83",X"8D",X"85",X"71",X"7C",X"91",X"7E",X"82",X"7D",X"70",X"88",X"8D",X"7D",X"83",X"6E",X"84",
		X"8F",X"7C",X"83",X"70",X"7E",X"90",X"7F",X"82",X"76",X"76",X"93",X"7E",X"83",X"7A",X"72",X"8D",
		X"89",X"76",X"75",X"92",X"7F",X"83",X"76",X"76",X"92",X"7F",X"6F",X"8A",X"8A",X"7D",X"72",X"83",
		X"90",X"79",X"75",X"8A",X"87",X"6B",X"89",X"89",X"7F",X"7F",X"71",X"81",X"93",X"70",X"7E",X"8E",
		X"80",X"79",X"73",X"8E",X"88",X"79",X"72",X"8E",X"86",X"7B",X"72",X"8E",X"85",X"6E",X"8E",X"84",
		X"6F",X"85",X"8E",X"78",X"74",X"91",X"7C",X"71",X"94",X"7A",X"73",X"8A",X"8C",X"76",X"76",X"8F",
		X"84",X"7D",X"83",X"6E",X"86",X"8B",X"81",X"71",X"83",X"8D",X"7E",X"78",X"75",X"92",X"81",X"81",
		X"7D",X"72",X"82",X"8E",X"80",X"80",X"7E",X"70",X"85",X"8C",X"83",X"70",X"80",X"8E",X"7F",X"72",
		X"81",X"90",X"7A",X"86",X"72",X"7D",X"90",X"77",X"74",X"8C",X"88",X"7D",X"83",X"75",X"78",X"8C",
		X"88",X"7D",X"83",X"74",X"79",X"8F",X"83",X"6F",X"87",X"8C",X"79",X"73",X"8A",X"89",X"7D",X"83",
		X"76",X"76",X"8C",X"87",X"7F",X"7D",X"70",X"8C",X"87",X"80",X"71",X"84",X"8D",X"7C",X"73",X"8C",
		X"83",X"6E",X"89",X"8A",X"7C",X"73",X"90",X"7E",X"83",X"70",X"84",X"8C",X"7E",X"78",X"78",X"93",
		X"7A",X"73",X"8A",X"89",X"7C",X"84",X"77",X"76",X"90",X"81",X"81",X"7A",X"73",X"8B",X"89",X"71",
		X"7E",X"8F",X"7E",X"71",X"8B",X"86",X"7F",X"7E",X"70",X"8D",X"87",X"72",X"7D",X"8E",X"82",X"73",
		X"7E",X"8F",X"7F",X"82",X"7D",X"72",X"88",X"8C",X"6F",X"86",X"89",X"7D",X"81",X"70",X"83",X"8C",
		X"82",X"70",X"83",X"8C",X"81",X"72",X"80",X"8E",X"7D",X"83",X"7A",X"74",X"86",X"8C",X"7C",X"72",
		X"87",X"8B",X"7D",X"83",X"78",X"76",X"8F",X"82",X"71",X"8D",X"82",X"80",X"7E",X"72",X"83",X"8D",
		X"7E",X"83",X"74",X"7E",X"8F",X"7B",X"85",X"74",X"7B",X"8F",X"7F",X"81",X"7B",X"73",X"87",X"8A",
		X"80",X"72",X"8B",X"84",X"7E",X"80",X"70",X"8B",X"87",X"7E",X"82",X"73",X"7D",X"8C",X"86",X"77",
		X"79",X"91",X"79",X"77",X"90",X"7A",X"77",X"90",X"79",X"75",X"8B",X"87",X"77",X"79",X"91",X"74",
		X"7D",X"8C",X"7F",X"72",X"85",X"8B",X"7D",X"72",X"87",X"89",X"7F",X"7B",X"74",X"8D",X"86",X"76",
		X"7A",X"91",X"74",X"7A",X"8B",X"86",X"78",X"77",X"8E",X"82",X"7F",X"81",X"73",X"7E",X"8C",X"84",
		X"76",X"7B",X"91",X"77",X"77",X"8A",X"87",X"76",X"79",X"8B",X"86",X"75",X"7B",X"8B",X"85",X"72",
		X"83",X"89",X"7E",X"7E",X"73",X"8F",X"80",X"73",X"83",X"8D",X"7D",X"84",X"73",X"7E",X"8B",X"84",
		X"74",X"7D",X"8C",X"82",X"74",X"7F",X"8D",X"80",X"7B",X"74",X"8D",X"84",X"79",X"76",X"8F",X"80",
		X"82",X"72",X"85",X"8A",X"7C",X"82",X"71",X"85",X"8A",X"7F",X"81",X"76",X"7B",X"8F",X"7F",X"83",
		X"75",X"7B",X"89",X"89",X"73",X"81",X"8B",X"7C",X"84",X"74",X"7D",X"8C",X"81",X"71",X"89",X"87",
		X"80",X"72",X"88",X"87",X"7F",X"75",X"82",X"8C",X"7B",X"84",X"73",X"7F",X"8E",X"7A",X"76",X"8D",
		X"81",X"7E",X"74",X"8C",X"84",X"71",X"85",X"8A",X"7E",X"74",X"86",X"8A",X"7B",X"75",X"8A",X"85",
		X"71",X"8B",X"83",X"73",X"89",X"85",X"7B",X"75",X"87",X"8A",X"79",X"76",X"8C",X"83",X"7F",X"80",
		X"73",X"81",X"89",X"86",X"73",X"7D",X"8B",X"84",X"7A",X"76",X"8C",X"83",X"7F",X"75",X"81",X"8D",
		X"7D",X"84",X"77",X"7A",X"8E",X"7B",X"75",X"8D",X"80",X"81",X"7B",X"75",X"8C",X"84",X"7F",X"73",
		X"87",X"88",X"7D",X"82",X"75",X"7D",X"8D",X"7F",X"74",X"8D",X"7E",X"75",X"8D",X"7E",X"74",X"88",
		X"88",X"7A",X"78",X"8D",X"7C",X"75",X"87",X"89",X"7A",X"76",X"88",X"89",X"77",X"7A",X"8E",X"7C",
		X"74",X"8A",X"85",X"7E",X"82",X"76",X"7B",X"89",X"87",X"72",X"88",X"85",X"7E",X"81",X"74",X"7F",
		X"88",X"87",X"75",X"7E",X"8E",X"77",X"79",X"8A",X"85",X"77",X"7A",X"8B",X"83",X"76",X"7F",X"8C",
		X"73",X"7E",X"8B",X"82",X"75",X"7E",X"8C",X"7F",X"77",X"7C",X"8D",X"80",X"75",X"86",X"87",X"73",
		X"7F",X"8B",X"80",X"7F",X"74",X"89",X"85",X"72",X"89",X"85",X"73",X"88",X"85",X"7D",X"82",X"71",
		X"8A",X"84",X"83",X"74",X"82",X"89",X"81",X"78",X"7D",X"8C",X"7F",X"7C",X"76",X"8A",X"86",X"7B",
		X"77",X"8C",X"81",X"80",X"7E",X"74",X"86",X"88",X"82",X"7A",X"78",X"8B",X"83",X"7E",X"82",X"77",
		X"7B",X"88",X"87",X"7A",X"77",X"86",X"89",X"78",X"7A",X"8C",X"7F",X"81",X"79",X"78",X"87",X"87",
		X"81",X"76",X"80",X"8D",X"74",X"81",X"89",X"7D",X"83",X"76",X"7D",X"8B",X"81",X"73",X"87",X"88",
		X"7D",X"76",X"8D",X"7D",X"77",X"8A",X"82",X"7A",X"78",X"89",X"86",X"76",X"7C",X"8B",X"81",X"7D",
		X"75",X"8B",X"82",X"74",X"8A",X"82",X"74",X"8B",X"81",X"80",X"7E",X"75",X"85",X"8A",X"77",X"7B",
		X"8A",X"83",X"77",X"7C",X"8B",X"81",X"77",X"7D",X"8D",X"7D",X"83",X"7A",X"78",X"89",X"86",X"7D",
		X"83",X"79",X"79",X"8A",X"84",X"75",X"80",X"8A",X"80",X"7B",X"78",X"8E",X"7C",X"78",X"8B",X"7F",
		X"81",X"7C",X"76",X"86",X"87",X"80",X"74",X"85",X"88",X"7B",X"76",X"8C",X"81",X"82",X"78",X"7C",
		X"8A",X"80",X"7B",X"78",X"8C",X"80",X"7E",X"75",X"87",X"87",X"7D",X"76",X"86",X"88",X"7B",X"77",
		X"87",X"87",X"79",X"7A",X"8C",X"7B",X"78",X"8C",X"80",X"81",X"7D",X"76",X"85",X"88",X"80",X"7E",
		X"76",X"86",X"88",X"7D",X"76",X"84",X"89",X"7B",X"79",X"89",X"81",X"80",X"7B",X"77",X"89",X"84",
		X"80",X"7F",X"75",X"88",X"84",X"7F",X"77",X"7F",X"8B",X"80",X"78",X"7E",X"8C",X"7B",X"79",X"88",
		X"83",X"77",X"7F",X"8C",X"76",X"7F",X"89",X"7F",X"78",X"7C",X"8B",X"81",X"76",X"83",X"8A",X"74",
		X"83",X"88",X"75",X"82",X"89",X"74",X"81",X"89",X"7D",X"83",X"77",X"7C",X"8C",X"7E",X"76",X"88",
		X"86",X"7E",X"83",X"7A",X"79",X"83",X"89",X"7F",X"76",X"88",X"85",X"74",X"84",X"89",X"75",X"82",
		X"88",X"7D",X"83",X"75",X"80",X"88",X"82",X"7A",X"7B",X"8B",X"7E",X"82",X"7B",X"78",X"88",X"86",
		X"76",X"83",X"88",X"74",X"83",X"88",X"7E",X"76",X"85",X"87",X"7E",X"82",X"7C",X"78",X"83",X"87",
		X"83",X"76",X"80",X"89",X"80",X"77",X"81",X"8A",X"7E",X"81",X"7E",X"77",X"81",X"89",X"81",X"78",
		X"7C",X"8B",X"80",X"82",X"74",X"86",X"85",X"80",X"77",X"82",X"88",X"7F",X"7A",X"7B",X"8C",X"7E",
		X"82",X"7B",X"78",X"87",X"86",X"7E",X"82",X"76",X"81",X"8A",X"7A",X"79",X"87",X"86",X"7A",X"79",
		X"89",X"83",X"7F",X"81",X"76",X"83",X"89",X"78",X"7C",X"89",X"82",X"78",X"7C",X"8B",X"7F",X"81",
		X"7C",X"77",X"87",X"85",X"7E",X"81",X"77",X"7E",X"8A",X"80",X"81",X"7F",X"77",X"81",X"89",X"80",
		X"80",X"7F",X"76",X"84",X"88",X"7E",X"82",X"79",X"7B",X"87",X"86",X"7C",X"79",X"88",X"83",X"76",
		X"81",X"88",X"80",X"77",X"81",X"89",X"7D",X"78",X"86",X"84",X"76",X"81",X"88",X"80",X"77",X"85",
		X"86",X"76",X"7E",X"89",X"81",X"78",X"7F",X"8A",X"7E",X"78",X"89",X"81",X"80",X"7E",X"77",X"82",
		X"87",X"82",X"7F",X"81",X"78",X"7D",X"88",X"83",X"7F",X"77",X"86",X"85",X"7E",X"82",X"76",X"80",
		X"88",X"82",X"7E",X"77",X"86",X"85",X"7F",X"77",X"86",X"85",X"7F",X"78",X"81",X"8A",X"75",X"83",
		X"87",X"77",X"7F",X"8A",X"79",X"7B",X"88",X"84",X"76",X"84",X"85",X"7E",X"78",X"82",X"88",X"7F",
		X"78",X"84",X"87",X"76",X"7F",X"88",X"82",X"7E",X"82",X"77",X"7F",X"89",X"7E",X"82",X"7B",X"7A",
		X"87",X"85",X"76",X"81",X"88",X"80",X"77",X"81",X"88",X"7E",X"82",X"7E",X"78",X"82",X"87",X"81",
		X"77",X"80",X"88",X"7F",X"78",X"81",X"89",X"7E",X"82",X"7E",X"78",X"82",X"88",X"81",X"78",X"7F",
		X"89",X"7E",X"82",X"7E",X"78",X"83",X"88",X"7A",X"7B",X"88",X"81",X"7E",X"77",X"87",X"84",X"7F",
		X"78",X"82",X"89",X"75",X"84",X"85",X"7F",X"81",X"78",X"7E",X"8A",X"7E",X"79",X"89",X"80",X"81",
		X"7D",X"78",X"85",X"86",X"81",X"76",X"86",X"84",X"80",X"79",X"7E",X"88",X"81",X"79",X"7D",X"8A",
		X"7E",X"82",X"7E",X"7A",X"7D",X"88",X"82",X"81",X"79",X"7F",X"8A",X"79",X"7B",X"88",X"82",X"7F",
		X"7F",X"77",X"85",X"86",X"7F",X"78",X"82",X"88",X"7F",X"82",X"7B",X"7A",X"86",X"85",X"7F",X"81",
		X"77",X"82",X"87",X"80",X"78",X"83",X"86",X"7D",X"83",X"77",X"81",X"88",X"7F",X"82",X"7B",X"7A",
		X"88",X"83",X"77",X"83",X"87",X"78",X"7E",X"88",X"80",X"80",X"7F",X"79",X"7D",X"87",X"83",X"80",
		X"77",X"83",X"85",X"7F",X"7A",X"7C",X"89",X"81",X"7A",X"7D",X"8A",X"7A",X"7B",X"86",X"84",X"7A",
		X"7C",X"89",X"7F",X"82",X"7C",X"7A",X"88",X"81",X"77",X"85",X"86",X"77",X"84",X"85",X"77",X"81",
		X"88",X"78",X"7D",X"87",X"82",X"78",X"81",X"87",X"7A",X"7C",X"89",X"7D",X"79",X"87",X"83",X"7A",
		X"7C",X"88",X"82",X"7A",X"7D",X"88",X"80",X"78",X"86",X"83",X"76",X"84",X"86",X"7E",X"78",X"86",
		X"83",X"7E",X"81",X"77",X"81",X"86",X"83",X"79",X"7E",X"88",X"7F",X"81",X"7D",X"79",X"86",X"84",
		X"7E",X"82",X"77",X"81",X"86",X"82",X"78",X"82",X"86",X"80",X"7D",X"7A",X"89",X"80",X"7F",X"78",
		X"88",X"81",X"78",X"87",X"81",X"7F",X"81",X"78",X"82",X"88",X"79",X"7F",X"88",X"7B",X"7B",X"85",
		X"85",X"7A",X"7E",X"87",X"7F",X"81",X"7D",X"79",X"84",X"85",X"80",X"80",X"78",X"86",X"84",X"77",
		X"81",X"87",X"7E",X"82",X"7A",X"7D",X"89",X"7E",X"82",X"7D",X"7A",X"82",X"87",X"7F",X"81",X"7F",
		X"79",X"83",X"87",X"7A",X"7C",X"87",X"81",X"7E",X"79",X"85",X"85",X"7E",X"79",X"84",X"86",X"79",
		X"7E",X"88",X"7B",X"7B",X"86",X"83",X"7F",X"82",X"79",X"7E",X"87",X"81",X"7D",X"79",X"86",X"84",
		X"7F",X"79",X"84",X"85",X"77",X"85",X"84",X"7F",X"81",X"7A",X"7D",X"86",X"83",X"7E",X"82",X"7B",
		X"7C",X"87",X"81",X"78",X"81",X"86",X"7F",X"79",X"82",X"86",X"7E",X"79",X"81",X"87",X"7E",X"79",
		X"87",X"82",X"7F",X"80",X"78",X"84",X"85",X"7C",X"7B",X"87",X"81",X"80",X"78",X"86",X"83",X"80",
		X"7B",X"7C",X"88",X"81",X"7C",X"7C",X"89",X"7B",X"7B",X"85",X"84",X"7B",X"7B",X"85",X"84",X"7C",
		X"7A",X"86",X"84",X"7C",X"7B",X"87",X"82",X"7F",X"79",X"85",X"84",X"78",X"84",X"84",X"7A",X"7E",
		X"87",X"81",X"7A",X"81",X"86",X"7A",X"7C",X"87",X"81",X"7F",X"81",X"7A",X"7F",X"88",X"7E",X"7A",
		X"85",X"83",X"7A",X"7E",X"88",X"7B",X"7D",X"88",X"7D",X"7B",X"87",X"80",X"79",X"84",X"84",X"7E",
		X"82",X"79",X"7F",X"87",X"80",X"80",X"79",X"83",X"86",X"7F",X"79",X"83",X"85",X"78",X"80",X"87",
		X"7F",X"81",X"7A",X"7F",X"88",X"7A",X"7E",X"87",X"7F",X"81",X"7D",X"7A",X"84",X"85",X"7F",X"79",
		X"81",X"87",X"7E",X"82",X"7B",X"7E",X"87",X"7E",X"79",X"84",X"85",X"7E",X"82",X"7C",X"7B",X"84",
		X"86",X"78",X"83",X"84",X"80",X"7A",X"7E",X"86",X"82",X"7A",X"7E",X"87",X"81",X"7A",X"7F",X"87",
		X"80",X"7E",X"79",X"86",X"83",X"7F",X"81",X"79",X"81",X"86",X"7E",X"82",X"7B",X"7D",X"87",X"80",
		X"81",X"7F",X"7A",X"81",X"87",X"7C",X"7B",X"86",X"82",X"7C",X"7B",X"86",X"83",X"7D",X"7A",X"88",
		X"7E",X"7B",X"85",X"82",X"7B",X"7D",X"87",X"80",X"7E",X"7A",X"85",X"84",X"7E",X"7A",X"85",X"84",
		X"7E",X"7A",X"84",X"84",X"7E",X"82",X"79",X"80",X"86",X"7E",X"7A",X"85",X"83",X"7F",X"80",X"79",
		X"85",X"84",X"79",X"82",X"86",X"79",X"81",X"86",X"7B",X"7D",X"87",X"7F",X"79",X"86",X"81",X"79",
		X"85",X"83",X"79",X"82",X"85",X"78",X"82",X"85",X"7F",X"81",X"7B",X"7D",X"87",X"80",X"80",X"7F",
		X"7A",X"83",X"86",X"7B",X"7D",X"86",X"81",X"7B",X"7D",X"86",X"82",X"7C",X"7D",X"88",X"7D",X"7B",
		X"83",X"85",X"7E",X"7A",X"83",X"85",X"7C",X"7C",X"86",X"80",X"7F",X"7A",X"85",X"83",X"79",X"85",
		X"83",X"7A",X"81",X"86",X"79",X"80",X"85",X"81",X"7E",X"7B",X"87",X"80",X"81",X"7E",X"7B",X"83",
		X"86",X"79",X"81",X"84",X"80",X"7B",X"80",X"86",X"7F",X"7D",X"7D",X"88",X"7E",X"82",X"7C",X"7C",
		X"85",X"83",X"79",X"81",X"86",X"7F",X"7A",X"82",X"86",X"79",X"80",X"85",X"81",X"7A",X"7F",X"86",
		X"81",X"7B",X"7E",X"87",X"7F",X"80",X"80",X"7B",X"80",X"87",X"7E",X"7A",X"85",X"83",X"7F",X"7A",
		X"84",X"84",X"7F",X"7C",X"7E",X"87",X"7E",X"82",X"7D",X"7B",X"85",X"81",X"7F",X"7A",X"85",X"82",
		X"7F",X"7B",X"80",X"86",X"80",X"7B",X"80",X"86",X"7F",X"80",X"80",X"7A",X"81",X"85",X"7F",X"7A",
		X"82",X"85",X"80",X"7B",X"81",X"86",X"7C",X"7C",X"86",X"81",X"81",X"7C",X"7E",X"86",X"7F",X"80",
		X"79",X"84",X"84",X"7F",X"80",X"7F",X"7A",X"83",X"84",X"7F",X"81",X"7B",X"7E",X"83",X"85",X"7D",
		X"7C",X"86",X"81",X"7A",X"81",X"85",X"7F",X"7B",X"84",X"82",X"7F",X"81",X"7A",X"80",X"85",X"81",
		X"7F",X"81",X"7D",X"7C",X"84",X"84",X"7F",X"7A",X"82",X"85",X"7F",X"81",X"7F",X"7A",X"84",X"83",
		X"7F",X"80",X"7A",X"81",X"85",X"80",X"80",X"7D",X"7C",X"86",X"81",X"80",X"80",X"7A",X"85",X"82",
		X"7F",X"81",X"7B",X"7E",X"85",X"82",X"7F",X"81",X"7B",X"7F",X"84",X"83",X"7C",X"7D",X"85",X"82",
		X"7C",X"7E",X"86",X"7D",X"7C",X"85",X"82",X"7F",X"81",X"7E",X"7B",X"84",X"83",X"81",X"7C",X"7D",
		X"87",X"7C",X"7E",X"86",X"7F",X"7B",X"86",X"80",X"81",X"7C",X"7E",X"86",X"7F",X"7B",X"83",X"84",
		X"7F",X"80",X"7A",X"81",X"85",X"7F",X"82",X"7C",X"7E",X"85",X"80",X"7E",X"7C",X"87",X"7E",X"7C",
		X"85",X"80",X"7B",X"84",X"82",X"79",X"82",X"84",X"81",X"7A",X"81",X"85",X"80",X"7F",X"7B",X"86",
		X"81",X"7A",X"83",X"84",X"7F",X"81",X"7F",X"7B",X"82",X"85",X"7B",X"7D",X"85",X"81",X"7F",X"81",
		X"7D",X"7C",X"85",X"82",X"80",X"7A",X"83",X"83",X"80",X"7D",X"7D",X"86",X"80",X"7F",X"7B",X"84",
		X"83",X"7F",X"81",X"7E",X"7C",X"83",X"84",X"7B",X"81",X"85",X"7C",X"7E",X"86",X"7C",X"7D",X"84",
		X"84",X"7C",X"7E",X"85",X"80",X"7C",X"7D",X"85",X"81",X"7F",X"81",X"7C",X"7F",X"86",X"7F",X"81",
		X"7F",X"7B",X"84",X"83",X"7C",X"7F",X"86",X"7B",X"7E",X"84",X"82",X"7D",X"7D",X"85",X"80",X"7F",
		X"7B",X"86",X"80",X"80",X"7F",X"7B",X"82",X"85",X"7B",X"80",X"84",X"80",X"7D",X"7D",X"85",X"82",
		X"7D",X"7D",X"85",X"81",X"7D",X"7D",X"84",X"82",X"7D",X"7E",X"86",X"7D",X"7C",X"84",X"82",X"7B",
		X"80",X"85",X"7F",X"80",X"80",X"7B",X"81",X"85",X"7F",X"81",X"7D",X"7D",X"82",X"84",X"80",X"7B",
		X"81",X"84",X"7F",X"7B",X"83",X"83",X"7F",X"81",X"7B",X"80",X"83",X"83",X"7D",X"7C",X"85",X"81",
		X"7F",X"81",X"7D",X"7D",X"83",X"83",X"80",X"7B",X"83",X"83",X"80",X"7B",X"81",X"84",X"80",X"7C",
		X"80",X"85",X"7B",X"7E",X"84",X"82",X"7F",X"82",X"7C",X"7E",X"85",X"80",X"80",X"7B",X"83",X"84",
		X"7A",X"83",X"82",X"80",X"7C",X"81",X"85",X"7B",X"7F",X"84",X"80",X"7F",X"81",X"7C",X"7F",X"85",
		X"7E",X"7C",X"83",X"84",X"7F",X"81",X"7B",X"80",X"84",X"7F",X"81",X"7D",X"7C",X"83",X"83",X"80",
		X"7B",X"80",X"84",X"7F",X"7C",X"81",X"84",X"7F",X"81",X"7F",X"7C",X"81",X"85",X"7B",X"7F",X"85",
		X"7F",X"81",X"7D",X"7D",X"82",X"84",X"80",X"80",X"80",X"7B",X"82",X"83",X"7F",X"81",X"7D",X"7D",
		X"85",X"80",X"80",X"80",X"7C",X"80",X"85",X"80",X"80",X"7F",X"7C",X"85",X"81",X"7B",X"82",X"83",
		X"7A",X"82",X"83",X"7F",X"81",X"7B",X"80",X"85",X"7F",X"7C",X"84",X"82",X"7B",X"80",X"84",X"81",
		X"7C",X"7F",X"85",X"7F",X"82",X"7D",X"7E",X"85",X"80",X"7B",X"82",X"83",X"7F",X"80",X"7B",X"85",
		X"81",X"7B",X"81",X"84",X"80",X"7C",X"83",X"82",X"7B",X"80",X"84",X"80",X"81",X"7C",X"81",X"85",
		X"7B",X"7F",X"85",X"7D",X"7D",X"84",X"81",X"80",X"81",X"7E",X"7C",X"83",X"83",X"7F",X"7C",X"81",
		X"84",X"7F",X"81",X"7C",X"7F",X"85",X"7F",X"7C",X"82",X"83",X"7E",X"7C",X"82",X"84",X"7F",X"81",
		X"7F",X"7C",X"81",X"84",X"80",X"80",X"81",X"7C",X"80",X"85",X"7F",X"7C",X"84",X"80",X"81",X"7C",
		X"7F",X"84",X"81",X"7E",X"7D",X"84",X"82",X"7D",X"7D",X"84",X"81",X"7E",X"7C",X"84",X"81",X"7F",
		X"81",X"7D",X"7D",X"82",X"83",X"80",X"7C",X"82",X"83",X"7F",X"7C",X"81",X"84",X"7F",X"81",X"7F",
		X"7C",X"80",X"83",X"82",X"7D",X"7E",X"84",X"81",X"7F",X"81",X"7C",X"80",X"84",X"81",X"7D",X"7E",
		X"84",X"80",X"7F",X"7C",X"83",X"83",X"7E",X"7D",X"84",X"81",X"7B",X"82",X"83",X"7F",X"7C",X"81",
		X"83",X"80",X"7C",X"81",X"84",X"7F",X"80",X"80",X"7C",X"81",X"84",X"7D",X"7D",X"83",X"82",X"7F",
		X"81",X"7D",X"7D",X"82",X"83",X"80",X"80",X"80",X"7B",X"82",X"83",X"80",X"7E",X"7D",X"84",X"81",
		X"7F",X"80",X"7B",X"82",X"83",X"80",X"7E",X"7D",X"85",X"80",X"80",X"7F",X"7C",X"83",X"82",X"7C",
		X"81",X"84",X"7C",X"80",X"84",X"7D",X"7E",X"85",X"7F",X"7C",X"83",X"82",X"7F",X"81",X"7C",X"81",
		X"84",X"80",X"80",X"80",X"7D",X"7F",X"83",X"82",X"7C",X"81",X"83",X"7F",X"81",X"7C",X"7F",X"83",
		X"81",X"7F",X"81",X"7D",X"7E",X"85",X"80",X"80",X"7F",X"7C",X"82",X"83",X"7D",X"7E",X"83",X"82",
		X"7E",X"7D",X"84",X"81",X"80",X"80",X"7C",X"81",X"84",X"80",X"81",X"7E",X"7D",X"84",X"82",X"7C",
		X"82",X"83",X"7C",X"7F",X"84",X"80",X"80",X"81",X"7D",X"7E",X"83",X"82",X"80",X"80",X"7C",X"82",
		X"83",X"7C",X"80",X"84",X"7D",X"7D",X"84",X"80",X"81",X"7C",X"82",X"83",X"7F",X"7E",X"7E",X"84",
		X"80",X"80",X"80",X"7D",X"7E",X"85",X"80",X"7D",X"83",X"81",X"7C",X"81",X"83",X"7F",X"7C",X"82",
		X"83",X"7B",X"80",X"83",X"80",X"7D",X"7E",X"84",X"80",X"80",X"80",X"7D",X"7F",X"84",X"7F",X"7C",
		X"84",X"81",X"80",X"7C",X"83",X"82",X"7C",X"82",X"82",X"7C",X"80",X"84",X"7D",X"7E",X"84",X"80",
		X"80",X"80",X"7C",X"83",X"82",X"80",X"7E",X"7E",X"85",X"7E",X"7D",X"82",X"83",X"7E",X"7D",X"83",
		X"80",X"7C",X"83",X"81",X"7C",X"83",X"81",X"80",X"80",X"7C",X"7F",X"82",X"82",X"7E",X"7D",X"83",
		X"82",X"7E",X"7D",X"83",X"82",X"7E",X"7E",X"84",X"7F",X"7C",X"84",X"80",X"7C",X"83",X"81",X"7F",
		X"80",X"7C",X"81",X"83",X"80",X"7F",X"7D",X"83",X"81",X"7C",X"81",X"83",X"7B",X"82",X"82",X"7F",
		X"80",X"7C",X"82",X"82",X"80",X"7D",X"82",X"83",X"7B",X"82",X"82",X"80",X"7D",X"80",X"83",X"80",
		X"7D",X"80",X"84",X"7F",X"81",X"7F",X"7D",X"82",X"83",X"80",X"7C",X"81",X"83",X"7F",X"7D",X"81",
		X"84",X"7D",X"7F",X"84",X"7F",X"7D",X"84",X"80",X"81",X"7C",X"81",X"83",X"7F",X"81",X"7E",X"7E",
		X"82",X"83",X"7F",X"81",X"7D",X"7F",X"83",X"81",X"7D",X"7F",X"84",X"80",X"7C",X"83",X"81",X"7C",
		X"82",X"82",X"7C",X"80",X"83",X"80",X"80",X"80",X"7D",X"7E",X"83",X"81",X"80",X"80",X"7F",X"7D",
		X"82",X"83",X"80",X"80",X"80",X"7C",X"81",X"83",X"7F",X"81",X"7E",X"7D",X"82",X"82",X"80",X"7E",
		X"7D",X"84",X"81",X"80",X"80",X"7D",X"80",X"84",X"7E",X"7E",X"83",X"81",X"7F",X"7D",X"82",X"82",
		X"7E",X"7E",X"83",X"7F",X"7D",X"82",X"82",X"7F",X"7D",X"82",X"83",X"7F",X"7D",X"83",X"81",X"7C",
		X"82",X"81",X"7F",X"81",X"7D",X"80",X"83",X"7F",X"7D",X"83",X"81",X"7F",X"81",X"7C",X"81",X"83",
		X"7F",X"80",X"7F",X"7D",X"82",X"82",X"80",X"7D",X"80",X"83",X"80",X"7D",X"82",X"82",X"7F",X"81",
		X"7D",X"7F",X"82",X"82",X"7D",X"81",X"83",X"7F",X"81",X"7D",X"7E",X"84",X"7F",X"7D",X"83",X"80",
		X"7D",X"83",X"81",X"80",X"7E",X"7E",X"84",X"7E",X"7E",X"82",X"81",X"7D",X"80",X"83",X"81",X"7E",
		X"7E",X"83",X"81",X"7D",X"80",X"83",X"7E",X"7E",X"83",X"81",X"80",X"80",X"7C",X"82",X"82",X"7E",
		X"7E",X"83",X"81",X"7E",X"7E",X"83",X"80",X"80",X"7F",X"7D",X"83",X"80",X"80",X"7D",X"83",X"81",
		X"80",X"7D",X"80",X"83",X"7F",X"81",X"7E",X"7F",X"83",X"7F",X"7D",X"83",X"80",X"7C",X"83",X"81",
		X"7D",X"82",X"82",X"7C",X"81",X"82",X"80",X"7E",X"7F",X"83",X"81",X"7E",X"7F",X"83",X"80",X"80",
		X"81",X"7D",X"7F",X"83",X"81",X"7D",X"80",X"83",X"80",X"7D",X"81",X"82",X"7F",X"81",X"7D",X"7F",
		X"83",X"80",X"7D",X"83",X"80",X"7F",X"7D",X"83",X"81",X"80",X"80",X"7D",X"81",X"83",X"80",X"7D",
		X"83",X"81",X"80",X"80",X"7D",X"80",X"82",X"81",X"7E",X"7E",X"83",X"81",X"7E",X"7E",X"83",X"81",
		X"80",X"81",X"7E",X"7E",X"82",X"82",X"7F",X"7D",X"82",X"82",X"7C",X"81",X"82",X"81",X"7D",X"81",
		X"82",X"80",X"7E",X"7E",X"83",X"81",X"7E",X"7E",X"83",X"81",X"7F",X"7E",X"83",X"81",X"7E",X"7E",
		X"83",X"81",X"7F",X"7E",X"82",X"82",X"7E",X"7F",X"83",X"7F",X"7D",X"82",X"82",X"7E",X"7E",X"83",
		X"80",X"80",X"7E",X"7E",X"83",X"81",X"7F",X"7E",X"83",X"7F",X"7E",X"83",X"80",X"7D",X"81",X"83",
		X"7F",X"80",X"80",X"7D",X"80",X"83",X"7D",X"7F",X"83",X"80",X"81",X"7E",X"7E",X"83",X"80",X"80",
		X"80",X"7D",X"80",X"82",X"82",X"7D",X"80",X"82",X"80",X"7E",X"7E",X"83",X"81",X"7E",X"7E",X"83",
		X"80",X"80",X"80",X"7D",X"80",X"83",X"7F",X"7D",X"82",X"82",X"7F",X"81",X"7F",X"7E",X"82",X"81",
		X"7D",X"81",X"82",X"7F",X"81",X"7D",X"80",X"82",X"81",X"7E",X"7F",X"83",X"81",X"7E",X"7E",X"83",
		X"80",X"7D",X"81",X"82",X"80",X"80",X"7D",X"81",X"82",X"80",X"80",X"7F",X"7D",X"81",X"83",X"7F",
		X"7E",X"82",X"81",X"7D",X"81",X"82",X"7F",X"81",X"7D",X"81",X"82",X"7F",X"80",X"7E",X"7E",X"82",
		X"82",X"80",X"80",X"7D",X"81",X"83",X"7E",X"7E",X"82",X"82",X"7E",X"7F",X"83",X"7F",X"7D",X"82",
		X"82",X"80",X"80",X"80",X"7D",X"81",X"82",X"81",X"7D",X"80",X"82",X"80",X"7E",X"80",X"83",X"80",
		X"7F",X"7E",X"83",X"81",X"80",X"80",X"7D",X"81",X"82",X"80",X"80",X"80",X"7D",X"80",X"83",X"7F",
		X"7E",X"83",X"80",X"7D",X"81",X"82",X"80",X"7D",X"81",X"82",X"7F",X"80",X"80",X"7D",X"80",X"82",
		X"80",X"7D",X"81",X"82",X"80",X"80",X"80",X"7D",X"80",X"82",X"80",X"7F",X"7E",X"83",X"7F",X"7E",
		X"83",X"80",X"80",X"80",X"7D",X"81",X"82",X"81",X"7D",X"81",X"81",X"80",X"7E",X"7F",X"83",X"80",
		X"7F",X"7E",X"83",X"80",X"80",X"80",X"7F",X"7E",X"82",X"82",X"80",X"80",X"80",X"7D",X"81",X"82",
		X"7D",X"80",X"83",X"7F",X"7E",X"82",X"81",X"7D",X"80",X"82",X"80",X"7D",X"81",X"81",X"80",X"7D",
		X"81",X"82",X"80",X"7E",X"7F",X"83",X"80",X"80",X"80",X"7E",X"7F",X"82",X"82",X"7E",X"7F",X"82",
		X"80",X"7E",X"80",X"82",X"7F",X"81",X"7E",X"7E",X"82",X"82",X"80",X"80",X"80",X"7E",X"80",X"82",
		X"81",X"7E",X"81",X"82",X"7F",X"81",X"7E",X"7F",X"82",X"81",X"80",X"80",X"7D",X"80",X"82",X"81",
		X"7E",X"80",X"82",X"7F",X"81",X"7E",X"7E",X"81",X"82",X"80",X"80",X"80",X"7E",X"80",X"82",X"80",
		X"80",X"80",X"7D",X"82",X"81",X"80",X"80",X"7E",X"7F",X"82",X"81",X"80",X"80",X"7D",X"82",X"81",
		X"7F",X"81",X"7E",X"7F",X"82",X"80",X"7D",X"81",X"82",X"80",X"7D",X"81",X"82",X"7F",X"80",X"7D",
		X"81",X"82",X"7D",X"80",X"82",X"80",X"7E",X"81",X"82",X"7D",X"81",X"81",X"80",X"7D",X"81",X"82",
		X"7F",X"80",X"7E",X"7F",X"82",X"81",X"7F",X"81",X"7D",X"81",X"82",X"7E",X"7F",X"82",X"81",X"7E",
		X"7F",X"83",X"7F",X"7E",X"82",X"81",X"80",X"80",X"7F",X"7E",X"81",X"82",X"80",X"80",X"80",X"7E",
		X"7F",X"82",X"81",X"7E",X"81",X"82",X"7E",X"7F",X"82",X"80",X"80",X"7E",X"81",X"82",X"7F",X"80",
		X"7E",X"80",X"81",X"82",X"7F",X"7E",X"82",X"81",X"7F",X"81",X"7F",X"7E",X"82",X"81",X"7E",X"80",
		X"82",X"7E",X"7F",X"82",X"81",X"7E",X"7F",X"83",X"7F",X"7E",X"82",X"81",X"80",X"80",X"7F",X"7E",
		X"82",X"81",X"80",X"7E",X"7F",X"82",X"81",X"7E",X"7F",X"82",X"80",X"7F",X"7F",X"83",X"7E",X"7F",
		X"82",X"80",X"7F",X"7E",X"82",X"81",X"7F",X"7E",X"82",X"81",X"80",X"7E",X"81",X"81",X"80",X"7E",
		X"80",X"82",X"80",X"7F",X"7E",X"83",X"80",X"80",X"80",X"7E",X"81",X"82",X"80",X"7E",X"7F",X"82",
		X"80",X"7E",X"80",X"82",X"7E",X"7F",X"82",X"81",X"7F",X"7F",X"83",X"7E",X"7F",X"82",X"80",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
