library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_big_sprite_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_big_sprite_tile_bit1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"00",X"1E",X"36",X"60",X"C0",X"CC",X"ED",X"F1",X"1F",X"27",X"47",X"43",X"43",X"43",X"43",X"43",
		X"ED",X"CC",X"C0",X"60",X"36",X"1E",X"0E",X"00",X"43",X"43",X"43",X"43",X"47",X"27",X"1F",X"1F",
		X"00",X"1E",X"36",X"60",X"C0",X"CC",X"ED",X"F1",X"6F",X"F7",X"F7",X"73",X"7B",X"7B",X"7B",X"73",
		X"ED",X"CC",X"C0",X"60",X"36",X"1E",X"0E",X"00",X"7B",X"7B",X"7B",X"73",X"F7",X"F7",X"67",X"0F",
		X"FE",X"47",X"87",X"14",X"85",X"04",X"89",X"F0",X"00",X"00",X"C0",X"C0",X"40",X"C0",X"C0",X"40",
		X"F0",X"89",X"04",X"85",X"14",X"87",X"47",X"FE",X"C0",X"40",X"C0",X"40",X"C0",X"C0",X"00",X"00",
		X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",
		X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"F8",X"F4",X"F0",X"F0",X"28",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"87",X"FF",X"00",X"01",X"02",X"E4",X"F8",X"FA",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FC",X"F8",X"FA",X"FC",X"F8",X"F8",X"30",X"20",
		X"01",X"0F",X"07",X"0F",X"07",X"23",X"13",X"09",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",
		X"51",X"31",X"11",X"01",X"01",X"03",X"01",X"01",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"1F",X"00",X"05",X"02",X"07",X"0F",X"FF",X"FF",X"FF",
		X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"7F",X"FF",
		X"01",X"03",X"07",X"07",X"07",X"03",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EE",X"FF",X"FC",X"F0",X"00",X"C0",X"C0",X"60",X"B0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"CC",
		X"00",X"00",X"01",X"01",X"0F",X"1F",X"3F",X"7F",X"F8",X"FE",X"FD",X"FC",X"F9",X"F8",X"F8",X"F8",
		X"F4",X"F9",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"FC",X"FC",X"32",X"84",X"C3",X"F0",
		X"3F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"F8",X"F0",X"F0",X"A0",X"04",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E6",X"E2",X"E0",X"E0",X"E0",X"E6",X"FC",X"78",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"01",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"78",X"78",X"FC",X"F7",X"E3",X"E1",X"C0",X"FF",X"FF",X"3F",X"9F",X"CF",X"E3",X"C1",X"80",
		X"CC",X"4C",X"00",X"04",X"04",X"00",X"00",X"00",X"08",X"10",X"20",X"20",X"20",X"20",X"20",X"00",
		X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"60",X"F0",X"F8",X"FC",X"FC",X"FE",X"FC",X"EC",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0C",X"08",X"CE",X"CE",X"C0",X"C0",X"E0",X"E0",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"0B",X"FF",X"FF",
		X"07",X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"20",X"5C",X"7F",X"FF",X"7F",X"7F",X"1F",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"FF",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"0F",X"07",X"07",X"0B",X"00",X"00",X"00",X"00",X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"18",X"30",X"F6",X"F7",X"F7",X"F3",X"FB",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"0E",X"00",X"00",X"F9",X"FC",X"E4",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"7F",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"90",X"30",X"70",X"F0",
		X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"80",X"49",X"2A",X"08",X"7E",X"08",X"2A",X"49",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"80",X"00",X"02",X"09",X"80",X"08",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"40",X"61",X"63",X"66",X"6C",X"7A",X"00",X"00",X"81",X"C3",X"E3",X"33",X"1B",X"AF",
		X"7A",X"6C",X"66",X"63",X"61",X"40",X"00",X"00",X"AF",X"1B",X"33",X"E3",X"C3",X"81",X"00",X"00",
		X"00",X"00",X"04",X"06",X"06",X"06",X"06",X"07",X"20",X"70",X"71",X"53",X"DB",X"8B",X"8B",X"FF",
		X"07",X"06",X"06",X"06",X"06",X"04",X"00",X"00",X"FF",X"8B",X"8B",X"DB",X"53",X"71",X"70",X"20",
		X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"CC",
		X"00",X"21",X"00",X"00",X"04",X"00",X"00",X"00",X"FC",X"FC",X"CC",X"78",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"01",X"23",X"03",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"CE",
		X"05",X"01",X"02",X"00",X"10",X"02",X"00",X"00",X"FE",X"FE",X"CC",X"FC",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"06",X"03",X"00",X"00",X"3C",X"FE",X"FE",X"FB",X"F7",X"EF",X"AF",
		X"10",X"0C",X"20",X"10",X"08",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"33",X"61",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"03",X"07",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"F8",X"FC",X"F8",X"FA",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1C",X"38",X"78",X"63",X"E7",X"F3",X"F8",X"CC",X"DE",X"1E",X"3E",X"0E",X"1E",X"1E",X"1E",
		X"F8",X"F3",X"E7",X"E3",X"78",X"78",X"3C",X"1F",X"5E",X"1E",X"1E",X"3E",X"3E",X"1E",X"1E",X"0C",
		X"F0",X"F3",X"E0",X"E0",X"E0",X"E4",X"F0",X"7F",X"3F",X"9F",X"8F",X"73",X"18",X"17",X"15",X"F5",
		X"7C",X"78",X"F0",X"E0",X"E0",X"E0",X"E0",X"F3",X"E3",X"63",X"21",X"31",X"17",X"16",X"A0",X"D9",
		X"E0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"80",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"33",X"7F",X"1F",X"0F",X"07",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"E7",X"CF",X"CF",X"DF",X"DF",X"BE",X"7E",X"A3",X"4F",X"3F",X"FF",X"3F",X"3F",X"3F",X"3F",
		X"FE",X"FC",X"FC",X"78",X"70",X"00",X"00",X"00",X"3F",X"3F",X"1F",X"04",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E4",X"C0",X"C0",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
