library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"24",X"24",X"18",X"00",X"00",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"70",X"F8",X"8D",X"85",X"C0",X"60",X"00",
		X"8E",X"4A",X"2E",X"10",X"E8",X"A4",X"E2",X"00",X"18",X"3C",X"7E",X"FF",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"06",X"06",X"06",X"0E",X"0C",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"3E",X"7E",X"7E",X"3E",X"00",X"00",X"00",X"38",X"6E",X"42",X"42",X"6E",X"38",X"00",
		X"00",X"00",X"1C",X"24",X"24",X"1C",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"00",X"00",
		X"07",X"0F",X"07",X"07",X"04",X"08",X"0F",X"0F",X"E0",X"F0",X"E0",X"E0",X"20",X"10",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"04",X"04",X"07",X"0F",X"07",X"F0",X"F0",X"F0",X"20",X"20",X"E0",X"F0",X"E0",
		X"01",X"0F",X"07",X"07",X"04",X"08",X"0F",X"0F",X"80",X"F0",X"E0",X"E0",X"20",X"10",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"04",X"04",X"07",X"0F",X"07",X"F0",X"F0",X"F0",X"20",X"20",X"E0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"23",X"7D",X"79",X"79",X"00",X"00",X"00",X"00",X"F1",X"FF",X"F3",X"F3",
		X"79",X"79",X"7D",X"23",X"00",X"00",X"00",X"00",X"F3",X"F3",X"FF",X"F1",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"23",X"3D",X"39",X"79",X"00",X"00",X"00",X"00",X"F1",X"FF",X"F3",X"F3",
		X"79",X"39",X"3D",X"23",X"00",X"00",X"00",X"00",X"F3",X"F3",X"FF",X"F1",X"00",X"00",X"00",X"00",
		X"02",X"0E",X"0E",X"0F",X"00",X"00",X"00",X"1F",X"60",X"7F",X"78",X"F8",X"0F",X"0F",X"0E",X"EE",
		X"1F",X"18",X"1F",X"0F",X"00",X"00",X"00",X"00",X"EE",X"6E",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"84",X"84",X"FC",X"FC",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"7E",X"7E",X"42",X"42",X"7E",X"3C",
		X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"7E",X"7E",X"06",X"74",X"74",X"74",X"00",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"3E",X"3E",X"3E",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"21",X"40",X"80",X"80",X"40",X"21",X"1F",X"00",X"49",X"FF",X"49",X"49",X"FF",X"49",X"00",
		X"0F",X"0F",X"03",X"0F",X"0F",X"03",X"0F",X"0F",X"00",X"00",X"0F",X"08",X"0F",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"7E",X"FE",X"FE",X"FE",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"88",X"88",X"88",X"F8",X"F8",X"00",X"00",X"00",X"00",X"F8",X"C8",X"48",X"48",X"48",
		X"0F",X"1F",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"0F",X"09",X"09",X"09",X"0F",X"7F",X"7F",X"41",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"00",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"78",X"78",X"78",X"78",X"58",X"78",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"98",X"98",X"98",X"34",X"34",X"2C",X"2C",X"34",X"34",X"2C",X"2C",
		X"3F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"3F",X"22",X"AA",X"88",X"00",X"00",X"00",X"00",X"00",
		X"22",X"FE",X"C4",X"C6",X"46",X"C6",X"FC",X"AA",X"00",X"00",X"00",X"00",X"00",X"AA",X"88",X"AA",
		X"22",X"AA",X"00",X"FF",X"FF",X"00",X"88",X"AA",X"22",X"AA",X"88",X"0A",X"02",X"02",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"08",X"AA",X"8A",X"A2",X"48",X"48",X"48",X"7E",X"7E",X"00",X"00",X"00",
		X"42",X"42",X"3C",X"18",X"00",X"00",X"60",X"40",X"48",X"7E",X"7E",X"00",X"00",X"18",X"3C",X"42",
		X"40",X"60",X"00",X"00",X"32",X"7E",X"4C",X"48",X"00",X"00",X"60",X"40",X"42",X"7E",X"7E",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"C3",X"C3",X"C3",X"C3",
		X"3F",X"3F",X"3F",X"3F",X"C3",X"C3",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"C3",X"C3",X"C3",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",
		X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"06",X"0C",X"1B",X"33",X"7F",X"FF",X"3C",X"3C",X"3C",X"3C",X"C3",X"C3",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"FC",X"C3",X"C3",X"FF",X"FF",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",
		X"00",X"00",X"08",X"04",X"03",X"0F",X"00",X"0F",X"00",X"00",X"60",X"80",X"01",X"E3",X"06",X"EC",
		X"01",X"03",X"0F",X"00",X"07",X"08",X"07",X"00",X"9E",X"02",X"E2",X"02",X"E2",X"82",X"E2",X"02",
		X"06",X"09",X"09",X"0F",X"00",X"00",X"00",X"00",X"C3",X"23",X"20",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"3F",X"22",X"36",X"36",X"00",X"00",X"00",X"00",X"FF",X"D1",X"DB",X"5B",
		X"36",X"36",X"36",X"3F",X"00",X"00",X"00",X"00",X"1B",X"9B",X"DB",X"FF",X"00",X"00",X"00",X"00",
		X"0F",X"0B",X"08",X"0B",X"0F",X"08",X"0F",X"0E",X"F0",X"F0",X"10",X"F0",X"F0",X"10",X"70",X"F0",
		X"08",X"0F",X"0B",X"08",X"0B",X"0F",X"00",X"00",X"10",X"F0",X"F0",X"10",X"F0",X"F0",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"0C",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"F0",
		X"1F",X"20",X"20",X"20",X"30",X"10",X"00",X"00",X"F8",X"04",X"04",X"04",X"0C",X"08",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"0C",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"F0",
		X"1F",X"20",X"20",X"20",X"30",X"10",X"00",X"00",X"F8",X"04",X"04",X"04",X"0C",X"08",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"0C",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"F0",
		X"1F",X"20",X"20",X"20",X"30",X"10",X"00",X"00",X"F8",X"04",X"04",X"04",X"0C",X"08",X"00",X"00",
		X"0F",X"0E",X"0E",X"0F",X"0F",X"0C",X"0C",X"0F",X"F0",X"70",X"70",X"F0",X"F0",X"30",X"30",X"F0",
		X"1F",X"20",X"20",X"20",X"30",X"10",X"00",X"00",X"F8",X"04",X"04",X"04",X"0C",X"08",X"00",X"00",
		X"02",X"04",X"08",X"10",X"20",X"00",X"34",X"34",X"00",X"00",X"7C",X"00",X"00",X"00",X"2C",X"2C",
		X"37",X"00",X"00",X"00",X"0D",X"05",X"01",X"00",X"EC",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"08",X"08",X"08",X"08",X"08",X"00",X"34",X"34",X"40",X"20",X"10",X"08",X"04",X"00",X"2C",X"2C",
		X"07",X"30",X"00",X"00",X"0D",X"05",X"00",X"01",X"E0",X"0C",X"00",X"00",X"80",X"80",X"00",X"80",
		X"00",X"30",X"20",X"10",X"30",X"00",X"00",X"00",X"00",X"0C",X"04",X"08",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"30",X"10",X"20",X"30",X"0E",X"0E",X"00",X"00",X"0C",X"08",X"04",X"0C",X"70",X"70",
		X"00",X"31",X"11",X"27",X"37",X"07",X"01",X"01",X"00",X"8C",X"88",X"E4",X"EC",X"E0",X"80",X"80",
		X"00",X"00",X"30",X"20",X"10",X"30",X"00",X"00",X"00",X"00",X"0C",X"04",X"08",X"0C",X"00",X"00",
		X"20",X"10",X"08",X"04",X"02",X"00",X"34",X"04",X"10",X"10",X"10",X"10",X"10",X"00",X"2C",X"20",
		X"37",X"30",X"00",X"00",X"01",X"00",X"01",X"01",X"EC",X"0C",X"00",X"00",X"B0",X"20",X"80",X"80",
		X"00",X"00",X"3E",X"00",X"00",X"00",X"04",X"34",X"04",X"08",X"10",X"20",X"40",X"00",X"20",X"2C",
		X"37",X"30",X"00",X"00",X"00",X"01",X"01",X"01",X"EC",X"0C",X"00",X"00",X"30",X"A0",X"80",X"80",
		X"80",X"C0",X"60",X"30",X"D8",X"CC",X"FE",X"FF",X"00",X"00",X"3C",X"3C",X"3C",X"3C",X"00",X"00",
		X"D8",X"D8",X"D8",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"78",
		X"0A",X"3A",X"7A",X"7A",X"7A",X"3A",X"0A",X"04",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"04",
		X"00",X"FF",X"FF",X"81",X"81",X"81",X"81",X"81",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"3C",X"3C",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"FC",X"FC",X"3C",X"FC",X"FC",X"3C",X"FC",X"FC",
		X"81",X"81",X"81",X"81",X"81",X"FF",X"FF",X"00",X"3C",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"18",X"3C",X"18",X"18",X"18",X"18",X"00",X"00",X"18",X"18",X"18",X"18",X"3C",X"18",X"00",
		X"00",X"00",X"20",X"7E",X"7E",X"20",X"00",X"00",X"00",X"00",X"04",X"7E",X"7E",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"04",X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"20",X"00",
		X"02",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"10",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"10",X"02",X"01",X"06",X"00",X"10",X"00",X"02",X"80",X"70",X"50",X"D0",
		X"A3",X"15",X"07",X"02",X"10",X"02",X"00",X"00",X"B0",X"60",X"E2",X"80",X"90",X"02",X"80",X"10",
		X"00",X"00",X"00",X"2C",X"2C",X"03",X"01",X"01",X"00",X"00",X"00",X"16",X"16",X"00",X"FF",X"01",
		X"01",X"01",X"03",X"2C",X"2C",X"00",X"00",X"00",X"01",X"FF",X"00",X"16",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"34",X"34",X"C2",X"C1",X"01",X"00",X"00",X"00",X"1A",X"1A",X"00",X"FE",X"01",
		X"01",X"C1",X"C2",X"34",X"34",X"00",X"00",X"00",X"01",X"FE",X"00",X"1A",X"1A",X"00",X"00",X"00",
		X"06",X"06",X"18",X"18",X"00",X"18",X"04",X"03",X"60",X"60",X"18",X"18",X"00",X"18",X"20",X"C0",
		X"02",X"02",X"02",X"1A",X"1A",X"02",X"1A",X"01",X"40",X"40",X"40",X"58",X"58",X"40",X"58",X"80",
		X"00",X"00",X"18",X"00",X"18",X"18",X"04",X"07",X"00",X"00",X"18",X"00",X"18",X"18",X"20",X"E0",
		X"02",X"02",X"02",X"1A",X"02",X"1A",X"1A",X"03",X"40",X"40",X"40",X"58",X"40",X"58",X"58",X"C0",
		X"80",X"C0",X"60",X"30",X"D8",X"CC",X"C6",X"C3",X"01",X"03",X"06",X"0C",X"1B",X"33",X"63",X"C3",
		X"3C",X"3C",X"3C",X"3C",X"C3",X"C3",X"C3",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
