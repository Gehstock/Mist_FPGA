library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity swimmer_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of swimmer_tile_bit1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"1F",X"1F",X"1E",X"00",X"00",X"00",X"80",X"80",X"30",X"70",X"F8",
		X"3F",X"7F",X"7F",X"7F",X"9F",X"0F",X"3F",X"70",X"F0",X"E0",X"F0",X"F0",X"F0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",
		X"E7",X"F3",X"71",X"00",X"06",X"07",X"07",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"40",X"01",X"03",X"07",X"03",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"7F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"A0",
		X"7F",X"7E",X"3C",X"3B",X"1F",X"0F",X"03",X"00",X"20",X"60",X"E0",X"80",X"80",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"01",X"19",X"3F",X"3E",X"3E",X"00",X"00",X"00",X"E0",X"90",X"38",X"78",X"F8",
		X"1D",X"3F",X"3F",X"3F",X"3F",X"1E",X"00",X"00",X"F8",X"E0",X"E0",X"F0",X"F0",X"E0",X"00",X"00",
		X"03",X"03",X"03",X"04",X"03",X"01",X"00",X"00",X"C0",X"C0",X"A0",X"60",X"C0",X"04",X"0C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"20",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"39",X"39",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"E0",X"F0",X"E8",X"C8",X"98",X"38",
		X"7E",X"FF",X"FF",X"BF",X"BF",X"1F",X"16",X"34",X"E0",X"E0",X"F8",X"F8",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0C",X"1C",X"3D",X"3D",X"3D",X"78",X"78",X"00",X"00",X"00",X"80",X"80",X"80",X"B7",X"37",
		X"30",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"17",X"36",X"F6",X"FC",X"F8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0D",X"1E",X"1E",X"0E",X"00",X"80",X"A0",X"20",X"30",X"78",X"78",X"70",
		X"00",X"00",X"00",X"02",X"13",X"37",X"13",X"12",X"00",X"00",X"00",X"00",X"20",X"40",X"20",X"20",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"01",X"01",X"41",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",
		X"11",X"08",X"00",X"00",X"00",X"F0",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"1F",X"3F",X"7F",X"7F",X"00",X"00",X"E0",X"E0",X"C0",X"EC",X"EC",X"EC",
		X"7F",X"FE",X"F8",X"FF",X"FF",X"FF",X"FF",X"3E",X"9C",X"3C",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"1C",X"1E",X"0E",X"0F",X"0F",X"0F",X"1F",X"1F",X"00",X"78",X"7C",X"F8",X"F2",X"E6",X"CE",X"B8",
		X"7F",X"FF",X"BF",X"6F",X"E7",X"C5",X"08",X"00",X"F8",X"FE",X"FF",X"FF",X"C3",X"80",X"00",X"00",
		X"00",X"00",X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"3C",X"3E",X"7D",X"F9",X"F3",X"E7",X"DC",X"F8",
		X"FF",X"DF",X"37",X"F3",X"E3",X"06",X"FC",X"F8",X"FC",X"FC",X"FC",X"F8",X"F8",X"70",X"60",X"40",
		X"00",X"00",X"00",X"00",X"3C",X"3E",X"3F",X"0F",X"00",X"00",X"00",X"78",X"7C",X"FA",X"F2",X"E6",
		X"1F",X"3F",X"FF",X"FF",X"BF",X"6F",X"E7",X"C7",X"CE",X"B8",X"F0",X"F8",X"FC",X"FC",X"9C",X"1C",
		X"00",X"00",X"00",X"05",X"07",X"07",X"0F",X"1F",X"00",X"00",X"00",X"00",X"B0",X"20",X"70",X"F8",
		X"3F",X"1F",X"0F",X"0F",X"1B",X"1F",X"3E",X"34",X"FC",X"F8",X"F0",X"70",X"30",X"70",X"60",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",
		X"0F",X"3F",X"7F",X"FF",X"F8",X"F0",X"F8",X"78",X"F8",X"FC",X"FE",X"FF",X"1F",X"0F",X"1F",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"0F",X"07",X"0F",X"0F",X"1E",X"3E",X"0F",X"00",X"80",X"80",X"90",X"30",X"38",X"7C",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"0F",X"07",X"0F",X"3F",X"7E",X"7E",X"3F",X"1F",X"80",X"80",X"90",X"3C",X"3E",X"7E",X"FC",X"F8",
		X"01",X"1F",X"3E",X"61",X"7F",X"3F",X"1C",X"39",X"C0",X"C0",X"40",X"C0",X"C0",X"8E",X"30",X"E0",
		X"31",X"03",X"07",X"06",X"00",X"00",X"00",X"00",X"E0",X"84",X"FC",X"F8",X"70",X"00",X"00",X"00",
		X"03",X"07",X"1C",X"3F",X"7F",X"FF",X"E0",X"00",X"C0",X"C0",X"00",X"C0",X"C0",X"80",X"00",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1F",X"1F",X"1E",X"1E",X"3C",X"38",X"30",
		X"03",X"07",X"03",X"07",X"00",X"0F",X"1F",X"1E",X"80",X"C0",X"C0",X"B0",X"60",X"E0",X"C0",X"0C",
		X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"38",X"00",X"F8",X"F0",X"C3",X"F8",X"E0",X"00",X"00",X"00",
		X"00",X"01",X"07",X"0F",X"18",X"1F",X"1E",X"1C",X"00",X"80",X"80",X"80",X"00",X"80",X"80",X"04",
		X"3C",X"3C",X"18",X"00",X"00",X"01",X"01",X"00",X"78",X"38",X"01",X"3F",X"FE",X"FC",X"F8",X"C0",
		X"6D",X"5F",X"78",X"78",X"7C",X"3C",X"1C",X"1C",X"CE",X"DE",X"1E",X"1E",X"3E",X"3C",X"38",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"30",X"38",X"38",X"38",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",
		X"0F",X"3E",X"3E",X"1F",X"07",X"07",X"03",X"00",X"30",X"3C",X"78",X"F8",X"E0",X"E0",X"C0",X"00",
		X"0F",X"0F",X"0F",X"06",X"13",X"37",X"17",X"1E",X"F0",X"F0",X"F0",X"60",X"20",X"40",X"68",X"E8",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"20",X"F0",X"87",X"EF",X"FF",X"77",
		X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"87",X"EF",X"DF",X"07",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"0F",X"3F",X"FF",X"F9",X"00",X"00",X"00",X"00",X"A0",X"F0",X"F8",X"F8",
		X"F8",X"FC",X"3F",X"0F",X"0E",X"02",X"00",X"00",X"F8",X"10",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"30",X"7D",X"7F",X"7F",X"4F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"C7",X"60",X"78",X"7C",X"30",X"20",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3D",X"FE",X"FF",X"F3",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"F0",X"FE",X"FF",X"3F",X"1F",X"00",
		X"00",X"00",X"C1",X"F3",X"7F",X"EF",X"7F",X"3F",X"00",X"00",X"00",X"80",X"C0",X"F8",X"F0",X"F8",
		X"87",X"EF",X"FF",X"3F",X"03",X"C1",X"00",X"00",X"90",X"C0",X"F0",X"D0",X"80",X"00",X"00",X"00",
		X"78",X"FC",X"FE",X"FE",X"DF",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"0F",X"0F",X"0F",X"DF",X"FF",X"FE",X"FC",X"78",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"1F",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"1F",X"1F",X"1F",X"3F",X"00",X"00",X"60",X"70",X"B8",X"D8",X"D8",X"9C",
		X"3F",X"3F",X"3F",X"3E",X"1F",X"1F",X"0F",X"0F",X"DC",X"9C",X"3C",X"7C",X"F8",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",
		X"EF",X"FE",X"7E",X"3F",X"1F",X"0F",X"0F",X"0F",X"37",X"3F",X"7E",X"FC",X"F8",X"F0",X"F0",X"F0",
		X"00",X"03",X"07",X"0F",X"07",X"0F",X"0F",X"1F",X"00",X"80",X"C0",X"80",X"C0",X"D0",X"B0",X"78",
		X"3E",X"7F",X"7F",X"FF",X"FF",X"EF",X"E6",X"C3",X"FC",X"FE",X"FE",X"FF",X"FF",X"F7",X"67",X"23",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",
		X"0F",X"7E",X"FE",X"FF",X"EF",X"0F",X"0F",X"0F",X"30",X"3E",X"7F",X"FF",X"F7",X"F0",X"F0",X"F0",
		X"3E",X"3F",X"3F",X"07",X"01",X"00",X"00",X"00",X"00",X"F0",X"BC",X"C6",X"F0",X"7D",X"3F",X"0E",
		X"00",X"00",X"00",X"01",X"07",X"3F",X"3F",X"3E",X"30",X"3D",X"3B",X"C0",X"F0",X"FC",X"F0",X"00",
		X"03",X"07",X"0F",X"1E",X"FF",X"FF",X"FF",X"F9",X"00",X"00",X"00",X"00",X"A0",X"F0",X"F8",X"F8",
		X"F8",X"FC",X"FF",X"FF",X"1E",X"0F",X"07",X"03",X"F8",X"10",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"1F",X"03",X"01",X"07",X"39",X"FC",X"FF",X"F7",X"FB",
		X"1F",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"F6",X"F8",X"3C",X"00",X"01",X"03",
		X"F8",X"FE",X"7F",X"1F",X"3F",X"7F",X"FF",X"BE",X"00",X"00",X"00",X"80",X"E8",X"FC",X"FE",X"FE",
		X"3E",X"7F",X"FF",X"3F",X"1F",X"7F",X"FE",X"F8",X"7E",X"B4",X"C0",X"E0",X"80",X"00",X"00",X"00",
		X"0F",X"06",X"13",X"37",X"77",X"6E",X"5D",X"7E",X"F0",X"60",X"20",X"44",X"66",X"EE",X"DE",X"7E",
		X"3E",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"7C",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"06",X"13",X"37",X"27",X"6E",X"6E",X"5C",X"78",X"60",X"20",X"44",X"64",X"EE",X"EE",X"1E",X"1E",
		X"78",X"F0",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"1E",X"0F",X"0F",X"07",X"07",X"07",X"00",X"00",
		X"F7",X"A7",X"2E",X"1D",X"1F",X"1F",X"0F",X"0F",X"43",X"61",X"E8",X"D8",X"F8",X"F8",X"F0",X"F0",
		X"07",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",
		X"06",X"13",X"37",X"37",X"6E",X"6E",X"58",X"78",X"60",X"20",X"44",X"64",X"EE",X"EE",X"1E",X"1E",
		X"7C",X"3C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"3E",X"3C",X"38",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"07",X"07",X"00",X"00",X"F0",X"B8",X"DC",X"E1",X"FB",X"BF",X"5D",
		X"00",X"07",X"07",X"01",X"01",X"01",X"00",X"00",X"61",X"FB",X"B7",X"C1",X"E0",X"F8",X"F0",X"00",
		X"00",X"00",X"0F",X"3F",X"FF",X"FF",X"FF",X"F7",X"00",X"00",X"80",X"F0",X"F8",X"FC",X"FC",X"F0",
		X"F3",X"F9",X"FC",X"FF",X"3F",X"0F",X"00",X"00",X"F0",X"6C",X"1C",X"F8",X"F0",X"80",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"BC",X"CE",X"F0",X"3D",X"3F",X"0E",
		X"00",X"00",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"30",X"3D",X"3B",X"C0",X"F0",X"FC",X"F0",X"00",
		X"1C",X"1E",X"1E",X"0E",X"FF",X"FF",X"FF",X"F9",X"00",X"00",X"00",X"00",X"A0",X"F0",X"F8",X"F8",
		X"F8",X"FC",X"FF",X"FF",X"0E",X"1E",X"1E",X"1C",X"F8",X"10",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"0E",X"1C",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"38",X"1C",
		X"1C",X"1C",X"0E",X"0F",X"07",X"01",X"00",X"00",X"1C",X"1C",X"38",X"F8",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"0C",X"1C",X"3F",X"10",X"00",X"60",X"30",X"18",X"18",X"18",X"18",X"98",X"18",
		X"00",X"00",X"3E",X"43",X"00",X"00",X"00",X"00",X"7C",X"0E",X"06",X"07",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"08",X"0C",X"06",X"02",X"00",X"38",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"00",X"00",X"00",X"1C",X"06",X"03",X"03",X"03",X"FC",X"0E",X"07",X"07",X"07",X"07",X"07",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"20",X"20",X"30",X"30",X"30",X"F0",
		X"00",X"44",X"C6",X"FE",X"FE",X"FE",X"7C",X"7C",X"6C",X"6C",X"EE",X"FE",X"EE",X"6C",X"6C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"7C",X"7C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"7C",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"E0",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0E",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"60",X"E0",X"F0",X"F0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"0D",X"09",X"19",X"1F",X"01",X"1D",X"80",X"E0",X"B0",X"90",X"98",X"F8",X"80",X"B8",
		X"01",X"1D",X"01",X"0D",X"01",X"01",X"07",X"1F",X"80",X"B8",X"80",X"B0",X"80",X"80",X"E0",X"F8",
		X"00",X"00",X"00",X"82",X"8A",X"CA",X"C0",X"FF",X"00",X"00",X"00",X"B0",X"BC",X"A6",X"22",X"FF",
		X"FF",X"C0",X"CA",X"8A",X"82",X"00",X"00",X"00",X"FF",X"22",X"A6",X"BC",X"B0",X"00",X"00",X"00",
		X"02",X"03",X"0A",X"0C",X"0E",X"0E",X"0E",X"0C",X"20",X"60",X"28",X"18",X"38",X"38",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"77",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"77",X"F8",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"0C",X"18",X"00",X"00",X"88",X"80",X"80",X"C0",X"E0",X"30",
		X"18",X"0C",X"00",X"00",X"00",X"20",X"00",X"00",X"30",X"60",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"06",X"03",X"00",X"40",X"44",X"40",X"40",X"C0",X"E0",X"30",
		X"03",X"06",X"00",X"00",X"00",X"20",X"00",X"00",X"30",X"60",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"F8",X"F8",X"F0",X"F1",X"E3",X"E3",X"C3",X"00",X"3C",X"7E",X"FF",X"FF",X"E7",X"C3",X"C3",
		X"C3",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"0F",X"1F",X"3F",X"73",X"7B",X"73",X"3E",X"1C",X"E0",X"F0",X"F8",X"9C",X"BC",X"9C",X"F8",X"70",
		X"00",X"1F",X"1F",X"1F",X"9F",X"DF",X"DF",X"DF",X"00",X"3E",X"3E",X"BE",X"BE",X"FE",X"FE",X"FE",
		X"DF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"0E",X"1F",X"3F",X"3F",
		X"04",X"04",X"08",X"08",X"08",X"08",X"07",X"06",X"3F",X"1F",X"0F",X"07",X"03",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"80",X"FF",X"00",X"10",X"10",X"08",X"08",X"08",X"08",X"F0",X"30",
		X"01",X"00",X"08",X"08",X"08",X"00",X"00",X"01",X"FF",X"02",X"02",X"02",X"03",X"00",X"00",X"FF",
		X"FF",X"10",X"10",X"10",X"70",X"00",X"00",X"FF",X"C0",X"00",X"08",X"08",X"08",X"00",X"00",X"C0",
		X"0F",X"FF",X"9F",X"7F",X"5F",X"3F",X"3F",X"04",X"E0",X"FC",X"F4",X"FE",X"F2",X"FF",X"F9",X"28",
		X"20",X"78",X"FC",X"EE",X"E3",X"F1",X"7C",X"1F",X"0E",X"1F",X"3F",X"37",X"67",X"47",X"06",X"0C",
		X"0F",X"3F",X"3F",X"7F",X"5F",X"FF",X"9F",X"88",X"E0",X"FF",X"F1",X"FE",X"F2",X"FC",X"F4",X"48",
		X"20",X"7E",X"FF",X"E3",X"F8",X"7F",X"1F",X"00",X"0E",X"0F",X"9F",X"DF",X"1F",X"DF",X"1E",X"0C",
		X"00",X"03",X"02",X"07",X"04",X"0F",X"08",X"08",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"60",
		X"01",X"01",X"03",X"07",X"07",X"07",X"03",X"00",X"00",X"F0",X"FC",X"0E",X"00",X"80",X"E0",X"F8",
		X"60",X"A0",X"F1",X"97",X"FF",X"1E",X"7C",X"1E",X"00",X"00",X"F0",X"FC",X"9E",X"03",X"01",X"00",
		X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FE",X"78",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"30",X"20",X"28",X"10",X"00",X"06",X"00",X"04",X"04",X"24",X"14",X"08",X"00",X"00",
		X"0F",X"1F",X"13",X"03",X"06",X"0A",X"15",X"0A",X"00",X"48",X"F8",X"78",X"30",X"A8",X"54",X"A8",
		X"00",X"40",X"02",X"0A",X"22",X"02",X"2B",X"82",X"7F",X"04",X"11",X"A4",X"01",X"AA",X"04",X"4A",
		X"2A",X"57",X"22",X"AB",X"14",X"44",X"29",X"0B",X"00",X"4F",X"3F",X"FE",X"DF",X"FF",X"FB",X"FF",
		X"FF",X"00",X"81",X"48",X"02",X"48",X"21",X"52",X"00",X"08",X"25",X"30",X"A5",X"28",X"24",X"29",
		X"02",X"F8",X"FF",X"FF",X"FD",X"BF",X"FF",X"EF",X"B4",X"22",X"20",X"E9",X"94",X"90",X"C8",X"E8",
		X"00",X"03",X"1B",X"37",X"37",X"36",X"05",X"3B",X"00",X"80",X"DC",X"DC",X"E4",X"68",X"BE",X"DE",
		X"7B",X"7F",X"7D",X"33",X"4B",X"3B",X"01",X"00",X"DC",X"D0",X"E8",X"DC",X"DC",X"DC",X"B8",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",
		X"3F",X"7C",X"18",X"1A",X"08",X"00",X"00",X"00",X"FC",X"3E",X"18",X"58",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3C",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"3C",
		X"3E",X"7F",X"1F",X"1C",X"08",X"00",X"00",X"00",X"7C",X"FE",X"F8",X"38",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3C",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"3C",
		X"3E",X"7F",X"0F",X"0C",X"08",X"00",X"00",X"00",X"7C",X"FE",X"F0",X"30",X"10",X"00",X"00",X"00",
		X"00",X"02",X"06",X"06",X"02",X"06",X"06",X"06",X"80",X"A0",X"E0",X"60",X"60",X"60",X"F0",X"B0",
		X"07",X"06",X"07",X"07",X"03",X"03",X"07",X"07",X"F0",X"F0",X"A0",X"A0",X"A0",X"E0",X"A0",X"B0",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FC",X"F8",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"02",X"00",
		X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"40",X"00",X"F0",X"FC",X"FE",X"FE",X"FE",X"CB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"04",X"06",X"02",X"00",X"00",X"00",X"00",X"E6",X"E6",X"37",X"17",X"13",X"33",X"33",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"66",X"66",X"66",X"C6",X"C6",X"E6",X"0C",
		X"00",X"00",X"00",X"01",X"09",X"0D",X"0E",X"11",X"7F",X"FC",X"F0",X"E0",X"C0",X"BC",X"FE",X"E0",
		X"76",X"6F",X"CF",X"DE",X"DC",X"9C",X"9C",X"8C",X"80",X"E0",X"30",X"38",X"78",X"7C",X"FC",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"28",X"FE",X"AA",X"AA",X"AA",X"FE",X"00",X"DF",X"11",X"D1",X"1F",X"12",X"51",X"D1",
		X"06",X"06",X"07",X"07",X"07",X"03",X"0F",X"0F",X"A0",X"A0",X"A0",X"B0",X"B0",X"20",X"20",X"30",
		X"0E",X"06",X"07",X"07",X"07",X"0F",X"1F",X"1F",X"B0",X"A0",X"B0",X"F0",X"F0",X"F8",X"FC",X"FC",
		X"00",X"00",X"03",X"00",X"00",X"01",X"06",X"38",X"00",X"00",X"C0",X"80",X"80",X"40",X"40",X"40",
		X"7C",X"7D",X"7F",X"3B",X"03",X"01",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",
		X"08",X"0F",X"08",X"00",X"01",X"04",X"0F",X"15",X"00",X"E0",X"80",X"00",X"00",X"80",X"00",X"00",
		X"1A",X"32",X"0D",X"12",X"15",X"0A",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"10",X"00",X"00",X"00",X"00",X"00",
		X"40",X"60",X"20",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"84",X"88",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"A0",X"B0",X"F8",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"00",X"F8",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"C0",X"E0",X"E1",X"FF",X"FF",X"FF",X"FF",X"00",X"30",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"07",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"20",X"60",X"F0",X"F0",X"F8",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"00",X"01",X"03",X"07",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"E0",X"F0",X"FC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"1F",X"1F",X"0F",X"0F",X"1F",X"78",X"10",X"10",X"A0",X"D8",X"FC",X"FC",X"F8",
		X"1F",X"0F",X"07",X"0F",X"1F",X"1F",X"0C",X"00",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",
		X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"80",X"08",X"18",
		X"08",X"00",X"08",X"00",X"01",X"07",X"03",X"00",X"1C",X"1C",X"3C",X"78",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"01",X"05",X"08",X"00",X"10",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"9F",X"9F",X"7F",X"7F",X"FB",X"00",X"FF",X"FF",X"33",X"33",X"FF",X"FF",X"FF",
		X"F3",X"E7",X"EF",X"FF",X"FE",X"02",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"11",X"FF",
		X"00",X"0F",X"1F",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"60",X"30",X"10",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
