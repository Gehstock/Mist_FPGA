library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sol_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sol_sp_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"F0",X"00",X"00",X"90",X"00",X"00",X"00",X"FF",X"0B",X"00",
		X"00",X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"0B",X"B6",X"00",
		X"00",X"6B",X"00",X"00",X"00",X"FF",X"B0",X"00",X"00",X"9B",X"0B",X"00",X"00",X"99",X"00",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"BB",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9B",X"00",X"99",X"0F",X"BB",X"00",X"BB",X"BB",X"BB",X"B0",X"B0",X"9B",X"BB",X"B9",
		X"B0",X"BB",X"0B",X"B0",X"B0",X"F9",X"00",X"00",X"00",X"F9",X"F9",X"00",X"00",X"FF",X"F9",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"0F",X"99",X"00",X"00",X"BB",X"9F",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"0B",X"00",X"F9",X"BB",X"0B",X"00",X"99",X"9F",X"BB",
		X"00",X"90",X"90",X"9B",X"00",X"99",X"99",X"90",X"B0",X"FF",X"B9",X"00",X"BB",X"FF",X"BB",X"00",
		X"9B",X"F9",X"BB",X"00",X"9B",X"09",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"99",X"96",X"00",
		X"00",X"99",X"9A",X"00",X"99",X"AA",X"BB",X"00",X"BB",X"AA",X"BB",X"B0",X"B0",X"AA",X"B9",X"B9",
		X"B0",X"AA",X"0B",X"B0",X"B0",X"A9",X"AA",X"00",X"00",X"F9",X"AA",X"00",X"00",X"FF",X"69",X"00",
		X"00",X"AA",X"6A",X"00",X"00",X"0F",X"5A",X"00",X"00",X"BB",X"5A",X"00",X"00",X"A9",X"59",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AB",X"AA",X"0B",X"00",X"A9",X"99",X"0B",X"00",X"A9",X"99",X"BB",
		X"00",X"90",X"99",X"9B",X"00",X"99",X"9A",X"90",X"B0",X"9A",X"9A",X"00",X"BB",X"9A",X"BA",X"00",
		X"9B",X"F9",X"BA",X"00",X"9B",X"09",X"0B",X"00",X"00",X"09",X"0B",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"99",X"44",X"00",X"00",X"B0",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"99",
		X"00",X"99",X"BB",X"99",X"09",X"99",X"BB",X"99",X"04",X"99",X"99",X"09",X"04",X"0B",X"BB",X"09",
		X"44",X"BB",X"0B",X"00",X"49",X"00",X"BB",X"01",X"49",X"0B",X"F0",X"00",X"99",X"0B",X"00",X"B0",
		X"99",X"5B",X"00",X"B0",X"91",X"BB",X"00",X"B0",X"91",X"BB",X"40",X"B0",X"91",X"BB",X"40",X"B9",
		X"49",X"BB",X"40",X"BB",X"99",X"B0",X"00",X"BB",X"49",X"BB",X"B0",X"B0",X"99",X"B0",X"00",X"00",
		X"99",X"BB",X"B0",X"B0",X"99",X"BB",X"BB",X"BB",X"99",X"BB",X"BB",X"1B",X"44",X"1B",X"0B",X"19",
		X"04",X"10",X"00",X"14",X"04",X"11",X"00",X"94",X"04",X"11",X"90",X"94",X"00",X"9F",X"90",X"94",
		X"00",X"99",X"99",X"44",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",
		X"00",X"06",X"66",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F9",X"00",X"00",X"F0",
		X"F9",X"FF",X"FF",X"F0",X"F9",X"99",X"99",X"F0",X"99",X"99",X"99",X"9F",X"99",X"99",X"99",X"9F",
		X"99",X"F9",X"FF",X"9F",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9B",X"99",X"00",X"00",X"BB",X"C9",X"00",X"0F",X"00",X"C9",X"00",X"F9",X"00",X"C0",X"F0",
		X"99",X"99",X"00",X"F0",X"99",X"99",X"00",X"F0",X"99",X"99",X"99",X"F0",X"99",X"9B",X"99",X"F0",
		X"99",X"B0",X"99",X"F0",X"99",X"00",X"99",X"F0",X"99",X"00",X"B9",X"F0",X"BB",X"00",X"0B",X"B0",
		X"BB",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"95",X"00",
		X"00",X"99",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"96",X"00",
		X"00",X"55",X"95",X"00",X"00",X"55",X"65",X"80",X"00",X"55",X"95",X"88",X"99",X"99",X"99",X"88",
		X"99",X"99",X"96",X"99",X"F9",X"55",X"95",X"99",X"06",X"55",X"95",X"99",X"00",X"55",X"95",X"99",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"F9",X"90",X"00",X"00",X"99",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"BB",X"0F",X"90",
		X"00",X"BB",X"9F",X"00",X"00",X"B9",X"FF",X"00",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"F9",X"00",
		X"00",X"99",X"C9",X"99",X"00",X"B9",X"99",X"99",X"00",X"B9",X"99",X"99",X"00",X"B0",X"99",X"09",
		X"00",X"00",X"9B",X"09",X"00",X"00",X"FB",X"00",X"00",X"99",X"BB",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"9F",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"B9",X"00",X"00",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"44",
		X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"04",
		X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",
		X"00",X"04",X"44",X"44",X"00",X"44",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",
		X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"04",X"40",X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",
		X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"69",X"9F",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"69",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"FF",X"BB",X"0F",
		X"00",X"0F",X"BF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"66",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"00",
		X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"FB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"BB",X"00",X"00",X"B9",X"B9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"04",X"40",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"40",X"00",X"00",X"00",
		X"40",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",X"F0",
		X"FB",X"FF",X"FF",X"F0",X"FB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BF",
		X"BB",X"FB",X"FF",X"BF",X"BB",X"FB",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"11",X"1F",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"0F",X"1B",X"11",X"00",X"F1",X"BB",X"B1",X"F0",
		X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",X"BB",X"BF",X"BB",X"F0",
		X"BB",X"F0",X"BB",X"F0",X"BB",X"00",X"BB",X"00",X"FB",X"00",X"FB",X"00",X"0F",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",X"F0",
		X"FB",X"FF",X"FF",X"F0",X"FB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BF",
		X"BB",X"FB",X"FF",X"BF",X"BB",X"FB",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"60",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",
		X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"1B",X"F0",X"00",
		X"00",X"1B",X"F0",X"00",X"00",X"1B",X"F0",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",
		X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",
		X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"F0",X"00",X"00",X"1B",X"F0",X"00",
		X"00",X"1B",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"00",X"00",X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"BF",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"0F",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"BF",X"F0",X"00",X"00",X"FF",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"00",X"6B",X"00",X"00",X"00",X"6B",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"FF",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"BF",X"F0",X"00",X"00",X"FF",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"44",X"40",X"04",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",
		X"00",X"40",X"44",X"44",X"00",X"40",X"44",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"44",
		X"00",X"40",X"00",X"04",X"00",X"04",X"00",X"04",X"44",X"04",X"00",X"04",X"00",X"40",X"00",X"04",
		X"44",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",
		X"00",X"04",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"40",X"04",
		X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",
		X"00",X"44",X"44",X"40",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"50",X"BB",X"00",X"00",X"10",X"FB",X"00",X"00",X"11",X"50",X"00",X"00",X"11",X"00",
		X"00",X"0C",X"11",X"50",X"00",X"00",X"11",X"00",X"00",X"0C",X"10",X"50",X"00",X"00",X"10",X"00",
		X"00",X"0C",X"15",X"00",X"00",X"00",X"10",X"10",X"00",X"CC",X"11",X"11",X"00",X"00",X"10",X"10",
		X"00",X"C0",X"11",X"50",X"00",X"00",X"10",X"00",X"00",X"C0",X"11",X"05",X"00",X"00",X"11",X"00",
		X"00",X"C1",X"11",X"05",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"F5",X"00",X"00",X"10",X"BF",
		X"00",X"00",X"05",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"05",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"40",X"04",
		X"00",X"40",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"40",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",
		X"00",X"04",X"44",X"44",X"00",X"44",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"44",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"40",
		X"00",X"04",X"44",X"44",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"04",X"40",X"04",
		X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"40",X"00",X"44",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"9B",X"B9",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"9B",X"B9",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"F0",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"BB",X"00",
		X"00",X"B6",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"66",X"B0",X"00",X"00",X"66",X"B0",X"00",X"00",X"6F",X"B0",X"00",X"00",X"66",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"06",X"66",X"00",
		X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"6F",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",
		X"00",X"06",X"66",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"00",X"05",X"CC",X"CC",X"00",X"00",X"55",X"CC",X"0C",X"CC",X"55",X"CC",X"00",X"C0",X"55",X"CC",
		X"00",X"05",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"B5",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"C5",X"55",X"00",X"0C",X"CC",X"55",X"00",X"00",X"00",X"55",X"CC",X"00",X"55",X"55",X"CC",
		X"00",X"05",X"CC",X"CC",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"0D",X"00",X"80",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"F0",X"00",X"C0",X"00",X"00",
		X"00",X"0F",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"20",X"00",X"22",X"55",X"22",X"00",X"22",X"55",X"00",X"00",X"25",X"55",X"55",
		X"00",X"50",X"55",X"55",X"00",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"55",X"55",X"F5",X"55",X"00",X"55",X"AF",X"00",X"20",X"55",X"FA",X"20",X"22",X"55",X"FF",X"22",
		X"22",X"55",X"FA",X"22",X"22",X"55",X"FF",X"22",X"20",X"55",X"FA",X"20",X"00",X"55",X"AF",X"00",
		X"55",X"55",X"F5",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"50",X"55",X"55",X"00",X"20",X"00",X"05",X"00",X"22",X"55",X"00",X"00",X"22",X"55",X"22",
		X"00",X"00",X"55",X"20",X"00",X"05",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"60",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"66",X"6B",X"00",X"00",X"66",X"6B",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"FF",X"00",X"00",X"66",X"6B",X"00",X"00",X"66",X"6B",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"B0",X"00",
		X"00",X"B6",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"B0",X"00",X"00",X"66",X"B0",X"00",X"00",X"6F",X"B0",X"00",X"00",X"66",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"4F",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"CB",X"00",X"90",X"00",X"CC",X"99",X"99",X"00",X"0C",X"99",X"99",
		X"00",X"0C",X"99",X"99",X"00",X"CC",X"99",X"99",X"00",X"CB",X"00",X"90",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"00",X"00",X"00",X"00",
		X"0B",X"55",X"05",X"05",X"BB",X"00",X"00",X"00",X"BB",X"50",X"05",X"05",X"00",X"01",X"00",X"00",
		X"05",X"11",X"CC",X"05",X"00",X"11",X"00",X"00",X"05",X"11",X"CC",X"05",X"00",X"01",X"C0",X"00",
		X"00",X"51",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"50",X"10",X"0C",X"00",X"00",X"00",X"00",X"00",X"50",X"11",X"0C",X"50",X"00",X"11",X"00",X"00",
		X"50",X"11",X"11",X"50",X"00",X"01",X"00",X"00",X"50",X"05",X"50",X"50",X"00",X"00",X"00",X"00",
		X"0B",X"55",X"50",X"50",X"0B",X"00",X"00",X"00",X"05",X"50",X"50",X"50",X"00",X"00",X"00",X"00",
		X"00",X"50",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
