library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"80",X"EB",X"C3",X"68",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"B8",X"00",X"47",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"45",X"3A",X"00",X"A0",X"47",X"3A",X"01",X"A0",X"A0",
		X"E6",X"10",X"CA",X"AF",X"56",X"21",X"00",X"E0",X"11",X"01",X"E0",X"01",X"FF",X"0F",X"36",X"00",
		X"ED",X"B0",X"21",X"5B",X"36",X"22",X"7B",X"E0",X"11",X"17",X"E0",X"3E",X"0A",X"21",X"AE",X"00",
		X"01",X"0A",X"00",X"ED",X"B0",X"3D",X"20",X"F5",X"3E",X"03",X"32",X"20",X"E0",X"CD",X"80",X"5A",
		X"3E",X"80",X"32",X"A1",X"E1",X"AF",X"32",X"00",X"98",X"ED",X"56",X"FB",X"18",X"FE",X"01",X"00",
		X"00",X"29",X"29",X"29",X"01",X"01",X"00",X"00",X"C5",X"D5",X"E5",X"F5",X"DD",X"E5",X"FD",X"E5",
		X"FD",X"21",X"00",X"E0",X"FD",X"CB",X"01",X"7E",X"C4",X"6D",X"02",X"FD",X"CB",X"01",X"BE",X"CD",
		X"A6",X"01",X"CD",X"90",X"5A",X"21",X"56",X"01",X"06",X"14",X"FD",X"21",X"97",X"E0",X"3A",X"00",
		X"E0",X"CB",X"67",X"28",X"04",X"FD",X"21",X"1C",X"E1",X"5E",X"23",X"56",X"23",X"D5",X"DD",X"E1",
		X"5E",X"23",X"56",X"23",X"DD",X"CB",X"00",X"7E",X"28",X"0E",X"C5",X"E5",X"FD",X"E5",X"01",X"04",
		X"01",X"C5",X"EB",X"E9",X"FD",X"E1",X"E1",X"C1",X"10",X"DF",X"3A",X"01",X"E0",X"E6",X"20",X"28",
		X"0B",X"21",X"05",X"E0",X"35",X"20",X"05",X"21",X"01",X"E0",X"CB",X"AE",X"3A",X"01",X"E0",X"1F",
		X"38",X"16",X"1F",X"38",X"09",X"1F",X"38",X"19",X"1F",X"38",X"03",X"1F",X"38",X"1F",X"FD",X"E1",
		X"DD",X"E1",X"F1",X"E1",X"D1",X"C1",X"FB",X"C9",X"31",X"80",X"EB",X"FB",X"CD",X"EC",X"54",X"18",
		X"0C",X"31",X"76",X"EB",X"FB",X"CD",X"8E",X"55",X"F1",X"E1",X"D1",X"C1",X"C9",X"31",X"80",X"EB",
		X"FB",X"CD",X"47",X"56",X"18",X"FE",X"1A",X"E2",X"31",X"32",X"2F",X"E2",X"31",X"32",X"44",X"E2",
		X"31",X"32",X"59",X"E2",X"31",X"32",X"6E",X"E2",X"31",X"32",X"83",X"E2",X"31",X"32",X"98",X"E2",
		X"31",X"32",X"AD",X"E2",X"31",X"32",X"C2",X"E2",X"53",X"43",X"D3",X"E2",X"18",X"4B",X"E2",X"E2",
		X"18",X"4B",X"F1",X"E2",X"18",X"4B",X"09",X"E3",X"2B",X"54",X"C5",X"E1",X"B2",X"1F",X"00",X"E3",
		X"02",X"4E",X"D7",X"E1",X"DF",X"28",X"12",X"E2",X"01",X"2F",X"B6",X"E1",X"3C",X"19",X"A9",X"E1",
		X"CE",X"11",X"A1",X"E1",X"2A",X"0D",X"CD",X"DE",X"01",X"3A",X"01",X"A0",X"17",X"38",X"15",X"F5",
		X"3A",X"03",X"E0",X"A7",X"20",X"08",X"3A",X"03",X"A0",X"E6",X"0F",X"CD",X"FA",X"01",X"3E",X"03",
		X"32",X"03",X"E0",X"F1",X"17",X"D8",X"3A",X"04",X"E0",X"A7",X"20",X"0C",X"3A",X"03",X"A0",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"CD",X"FA",X"01",X"3E",X"03",X"32",X"04",X"E0",X"C9",X"21",X"02",
		X"E0",X"7E",X"A7",X"28",X"01",X"35",X"3A",X"00",X"A0",X"17",X"38",X"02",X"36",X"0A",X"23",X"7E",
		X"A7",X"28",X"01",X"35",X"23",X"7E",X"A7",X"C8",X"35",X"C9",X"4F",X"3E",X"14",X"06",X"00",X"CD",
		X"DF",X"02",X"3A",X"02",X"E0",X"A7",X"C0",X"3A",X"03",X"A0",X"47",X"E6",X"F0",X"C8",X"78",X"E6",
		X"0F",X"C8",X"79",X"87",X"5F",X"16",X"00",X"21",X"4D",X"02",X"19",X"EB",X"69",X"01",X"07",X"E0",
		X"09",X"34",X"1A",X"BE",X"C0",X"47",X"3A",X"06",X"E0",X"4F",X"13",X"1A",X"81",X"27",X"38",X"0B",
		X"FE",X"99",X"28",X"07",X"32",X"06",X"E0",X"36",X"00",X"18",X"07",X"3E",X"99",X"32",X"06",X"E0",
		X"05",X"70",X"3A",X"00",X"E0",X"17",X"D8",X"21",X"A1",X"E1",X"CB",X"E6",X"C9",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"01",X"03",X"02",X"03",X"01",X"02",
		X"03",X"02",X"01",X"01",X"05",X"01",X"04",X"01",X"03",X"01",X"02",X"01",X"01",X"21",X"11",X"E3",
		X"11",X"00",X"90",X"06",X"00",X"7E",X"87",X"28",X"08",X"87",X"4F",X"30",X"01",X"04",X"23",X"ED",
		X"B0",X"21",X"11",X"E3",X"3E",X"40",X"96",X"36",X"00",X"C8",X"D8",X"47",X"EB",X"23",X"11",X"04",
		X"00",X"AF",X"77",X"19",X"10",X"FC",X"C9",X"DD",X"56",X"01",X"DD",X"5E",X"03",X"21",X"11",X"E3",
		X"7E",X"87",X"D8",X"87",X"D8",X"D5",X"5F",X"16",X"00",X"23",X"19",X"D1",X"3A",X"00",X"E0",X"1F",
		X"38",X"0A",X"3E",X"08",X"92",X"57",X"7B",X"D6",X"08",X"5F",X"18",X"0C",X"79",X"EE",X"30",X"4F",
		X"7A",X"C6",X"08",X"57",X"3E",X"F8",X"93",X"5F",X"70",X"23",X"72",X"23",X"71",X"23",X"73",X"21",
		X"11",X"E3",X"34",X"21",X"01",X"E0",X"CB",X"FE",X"C9",X"21",X"00",X"E0",X"CB",X"7E",X"C8",X"5F",
		X"16",X"00",X"21",X"00",X"EC",X"19",X"CB",X"C0",X"70",X"C9",X"5F",X"16",X"00",X"21",X"00",X"EC",
		X"19",X"CB",X"D6",X"C9",X"2A",X"7B",X"E0",X"54",X"5D",X"29",X"19",X"7B",X"84",X"67",X"22",X"7B",
		X"E0",X"C9",X"3A",X"00",X"E0",X"17",X"D0",X"FD",X"E5",X"E1",X"01",X"07",X"00",X"09",X"CD",X"18",
		X"03",X"FD",X"E5",X"E1",X"01",X"2F",X"00",X"09",X"37",X"06",X"03",X"7E",X"CE",X"00",X"27",X"FE",
		X"60",X"38",X"01",X"AF",X"77",X"3F",X"2B",X"10",X"F2",X"C9",X"3A",X"00",X"E0",X"17",X"D0",X"FD",
		X"E5",X"E1",X"23",X"23",X"23",X"D5",X"CD",X"74",X"03",X"CD",X"80",X"03",X"FD",X"56",X"18",X"FD",
		X"5E",X"19",X"FD",X"66",X"01",X"FD",X"6E",X"02",X"7A",X"B3",X"20",X"05",X"7C",X"FE",X"90",X"30",
		X"1B",X"A7",X"ED",X"52",X"38",X"16",X"7B",X"C6",X"50",X"27",X"FD",X"77",X"19",X"5F",X"7A",X"CE",
		X"00",X"27",X"FD",X"77",X"18",X"57",X"FD",X"CB",X"1B",X"C6",X"18",X"D6",X"D1",X"FD",X"E5",X"E1",
		X"01",X"2C",X"00",X"09",X"06",X"03",X"AF",X"1A",X"8E",X"27",X"77",X"1B",X"2B",X"10",X"F8",X"C9",
		X"0E",X"09",X"3A",X"00",X"E0",X"CB",X"67",X"20",X"08",X"11",X"BD",X"88",X"21",X"98",X"E0",X"18",
		X"10",X"11",X"BD",X"8A",X"21",X"1D",X"E1",X"18",X"08",X"0E",X"2C",X"11",X"A1",X"8A",X"21",X"17",
		X"E0",X"AF",X"06",X"06",X"EB",X"71",X"C5",X"01",X"00",X"04",X"09",X"C1",X"EB",X"ED",X"6F",X"20",
		X"05",X"F5",X"3E",X"29",X"18",X"05",X"F6",X"80",X"F5",X"E6",X"0F",X"12",X"F1",X"E5",X"21",X"20",
		X"FC",X"19",X"EB",X"E1",X"CB",X"40",X"28",X"03",X"ED",X"6F",X"23",X"CB",X"50",X"20",X"02",X"F6",
		X"80",X"10",X"D1",X"C9",X"5E",X"23",X"56",X"23",X"7E",X"23",X"4E",X"23",X"46",X"23",X"D5",X"D9",
		X"D1",X"D9",X"C5",X"D9",X"21",X"00",X"04",X"19",X"D5",X"D9",X"08",X"7E",X"D9",X"77",X"08",X"12",
		X"13",X"23",X"D9",X"23",X"10",X"F4",X"D9",X"D1",X"21",X"20",X"00",X"19",X"EB",X"D9",X"C1",X"0D",
		X"20",X"E0",X"C9",X"5E",X"23",X"56",X"23",X"7E",X"23",X"46",X"23",X"D5",X"D9",X"D1",X"D9",X"D9",
		X"12",X"21",X"00",X"04",X"19",X"D9",X"08",X"7E",X"D9",X"77",X"21",X"20",X"00",X"19",X"EB",X"D9",
		X"08",X"23",X"10",X"EB",X"C9",X"5E",X"23",X"56",X"23",X"4E",X"23",X"23",X"EB",X"A7",X"28",X"0A",
		X"C5",X"01",X"20",X"00",X"09",X"13",X"3D",X"20",X"FB",X"C1",X"1A",X"71",X"11",X"00",X"04",X"19",
		X"77",X"C9",X"C5",X"D5",X"21",X"00",X"04",X"19",X"12",X"08",X"77",X"3C",X"08",X"13",X"23",X"10",
		X"F7",X"D1",X"21",X"20",X"00",X"19",X"EB",X"C1",X"0D",X"20",X"E7",X"C9",X"C5",X"E5",X"77",X"23",
		X"10",X"FC",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",X"20",X"F1",X"C9",X"AF",X"C5",X"D5",X"21",
		X"00",X"04",X"19",X"12",X"36",X"29",X"13",X"23",X"10",X"F9",X"D1",X"21",X"20",X"00",X"19",X"EB",
		X"C1",X"0D",X"20",X"E9",X"C9",X"11",X"70",X"88",X"21",X"47",X"05",X"3E",X"A5",X"12",X"13",X"06",
		X"04",X"7E",X"12",X"23",X"3A",X"03",X"98",X"E6",X"7E",X"BE",X"C0",X"13",X"23",X"10",X"F2",X"11",
		X"00",X"80",X"01",X"20",X"20",X"CD",X"6C",X"04",X"CD",X"A6",X"01",X"11",X"80",X"88",X"01",X"18",
		X"20",X"CD",X"6C",X"04",X"AF",X"32",X"00",X"F0",X"32",X"00",X"F8",X"32",X"11",X"E3",X"21",X"01",
		X"E0",X"CB",X"FE",X"3A",X"00",X"E0",X"E6",X"10",X"20",X"1F",X"21",X"24",X"05",X"CD",X"03",X"04",
		X"0E",X"09",X"CD",X"89",X"03",X"3A",X"00",X"E0",X"E6",X"20",X"28",X"20",X"21",X"2B",X"05",X"CD",
		X"03",X"04",X"0E",X"08",X"CD",X"91",X"03",X"18",X"13",X"21",X"24",X"05",X"CD",X"03",X"04",X"CD",
		X"03",X"04",X"0E",X"08",X"CD",X"89",X"03",X"0E",X"09",X"CD",X"91",X"03",X"CD",X"4F",X"05",X"CD",
		X"AA",X"05",X"21",X"32",X"05",X"CD",X"03",X"04",X"CD",X"03",X"04",X"FD",X"7E",X"04",X"47",X"E6",
		X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"22",X"8F",X"78",X"E6",X"0F",X"32",X"42",X"8F",
		X"CD",X"99",X"03",X"C9",X"FE",X"88",X"26",X"03",X"01",X"1C",X"1D",X"FE",X"8A",X"26",X"03",X"02",
		X"17",X"0D",X"22",X"8A",X"26",X"0A",X"1C",X"0C",X"0E",X"17",X"0E",X"28",X"28",X"28",X"28",X"29",
		X"21",X"8A",X"2C",X"03",X"1D",X"18",X"19",X"A5",X"40",X"CD",X"16",X"36",X"7A",X"6F",X"3E",X"3E",
		X"2D",X"08",X"3E",X"4C",X"08",X"01",X"0A",X"02",X"11",X"7D",X"89",X"CD",X"42",X"04",X"FD",X"7E",
		X"16",X"06",X"03",X"21",X"9D",X"89",X"87",X"30",X"0E",X"F5",X"C5",X"3E",X"1A",X"01",X"02",X"02",
		X"CD",X"5C",X"04",X"C1",X"F1",X"18",X"04",X"11",X"40",X"00",X"19",X"87",X"30",X"0E",X"F5",X"C5",
		X"3E",X"1A",X"01",X"01",X"02",X"CD",X"5C",X"04",X"C1",X"F1",X"18",X"04",X"11",X"20",X"00",X"19",
		X"10",X"D4",X"C9",X"3A",X"02",X"A0",X"E6",X"C0",X"07",X"07",X"06",X"00",X"4F",X"21",X"A6",X"05",
		X"09",X"7E",X"FD",X"77",X"00",X"C9",X"02",X"05",X"04",X"03",X"11",X"81",X"88",X"FD",X"7E",X"00",
		X"FE",X"07",X"38",X"02",X"3E",X"06",X"4F",X"A7",X"28",X"11",X"47",X"C5",X"08",X"3E",X"2E",X"08",
		X"3E",X"09",X"01",X"02",X"02",X"CD",X"42",X"04",X"C1",X"10",X"F0",X"3E",X"06",X"91",X"C8",X"87",
		X"4F",X"06",X"02",X"CD",X"6C",X"04",X"C9",X"DD",X"7E",X"01",X"FD",X"96",X"01",X"30",X"02",X"ED",
		X"44",X"B8",X"D0",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"30",X"02",X"ED",X"44",X"B9",X"C9",X"7A",
		X"94",X"30",X"02",X"ED",X"44",X"B8",X"D0",X"7B",X"95",X"30",X"02",X"ED",X"44",X"B9",X"C9",X"AF",
		X"32",X"C5",X"E1",X"32",X"C2",X"E2",X"32",X"00",X"E3",X"32",X"D7",X"E1",X"32",X"09",X"E3",X"32",
		X"12",X"E2",X"21",X"1A",X"E2",X"11",X"15",X"00",X"06",X"08",X"CD",X"25",X"06",X"21",X"D3",X"E2",
		X"11",X"0F",X"00",X"06",X"03",X"77",X"19",X"10",X"FC",X"C9",X"21",X"1A",X"E2",X"11",X"15",X"00",
		X"06",X"08",X"7E",X"A7",X"C0",X"19",X"10",X"FA",X"21",X"D3",X"E2",X"11",X"0F",X"00",X"06",X"03",
		X"7E",X"A7",X"C0",X"19",X"10",X"FA",X"3A",X"C2",X"E2",X"A7",X"C0",X"3A",X"09",X"E3",X"A7",X"C0",
		X"3A",X"00",X"E3",X"A7",X"C0",X"3A",X"12",X"E2",X"A7",X"C0",X"3A",X"D7",X"E1",X"A7",X"C0",X"3A",
		X"C5",X"E1",X"A7",X"C9",X"FD",X"E5",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",X"84",X"00",X"ED",
		X"B0",X"CD",X"93",X"05",X"FD",X"36",X"04",X"01",X"CD",X"76",X"1A",X"5F",X"16",X"00",X"21",X"71",
		X"1A",X"19",X"7E",X"FD",X"77",X"0A",X"FD",X"36",X"0B",X"9F",X"FD",X"36",X"19",X"50",X"CD",X"A1",
		X"06",X"CD",X"A6",X"01",X"CD",X"24",X"07",X"CD",X"A6",X"01",X"CD",X"20",X"0B",X"CD",X"E0",X"0B",
		X"C9",X"FD",X"7E",X"04",X"D6",X"01",X"27",X"FE",X"30",X"38",X"05",X"D6",X"30",X"27",X"18",X"F7",
		X"4F",X"E6",X"F0",X"0F",X"47",X"0F",X"0F",X"80",X"47",X"79",X"E6",X"0F",X"80",X"87",X"5F",X"16",
		X"00",X"21",X"E6",X"06",X"19",X"E5",X"7E",X"21",X"83",X"80",X"01",X"18",X"1A",X"CD",X"5C",X"04",
		X"E1",X"23",X"7E",X"21",X"83",X"84",X"01",X"18",X"1A",X"CD",X"5C",X"04",X"01",X"02",X"02",X"11",
		X"CF",X"81",X"CD",X"6C",X"04",X"C9",X"4B",X"0A",X"73",X"01",X"47",X"05",X"47",X"03",X"47",X"04",
		X"47",X"05",X"7E",X"06",X"7E",X"07",X"7E",X"08",X"63",X"09",X"47",X"03",X"47",X"04",X"47",X"05",
		X"7E",X"06",X"7E",X"07",X"7E",X"08",X"73",X"00",X"73",X"01",X"73",X"02",X"4B",X"0A",X"7E",X"06",
		X"7E",X"07",X"7E",X"08",X"73",X"00",X"73",X"01",X"73",X"02",X"47",X"03",X"47",X"04",X"47",X"05",
		X"74",X"0B",X"28",X"0C",X"FD",X"7E",X"04",X"E6",X"0F",X"87",X"5F",X"16",X"00",X"21",X"B7",X"07",
		X"19",X"5E",X"23",X"56",X"D5",X"EB",X"11",X"83",X"88",X"01",X"0D",X"06",X"C5",X"D5",X"C5",X"7E",
		X"E6",X"F0",X"0F",X"0F",X"CD",X"A1",X"07",X"7E",X"E6",X"0F",X"87",X"87",X"CD",X"A1",X"07",X"23",
		X"C1",X"10",X"EB",X"D1",X"13",X"13",X"C1",X"0D",X"20",X"E2",X"21",X"17",X"0B",X"CD",X"D4",X"03",
		X"D1",X"0E",X"0D",X"D9",X"11",X"12",X"E4",X"01",X"1F",X"00",X"D9",X"06",X"06",X"D9",X"62",X"6B",
		X"D9",X"1A",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"D9",X"77",X"23",X"36",X"FF",X"09",X"D9",X"1A",
		X"E6",X"0F",X"D9",X"77",X"23",X"36",X"FF",X"09",X"D9",X"13",X"10",X"E5",X"D9",X"13",X"13",X"D9",
		X"0D",X"20",X"D8",X"21",X"2A",X"E4",X"11",X"20",X"00",X"06",X"0C",X"CB",X"9E",X"19",X"10",X"FB",
		X"C9",X"E5",X"4F",X"06",X"00",X"21",X"D7",X"0A",X"09",X"3E",X"00",X"01",X"02",X"02",X"CD",X"DE",
		X"03",X"D9",X"D5",X"D9",X"D1",X"E1",X"C9",X"CB",X"07",X"19",X"08",X"67",X"08",X"B5",X"08",X"03",
		X"09",X"51",X"09",X"9F",X"09",X"ED",X"09",X"3B",X"0A",X"89",X"0A",X"00",X"C5",X"55",X"55",X"59",
		X"00",X"0C",X"30",X"00",X"00",X"0E",X"90",X"C3",X"00",X"00",X"00",X"C3",X"69",X"A0",X"00",X"00",
		X"0C",X"30",X"0A",X"A0",X"00",X"0C",X"53",X"00",X"0A",X"A0",X"00",X"0A",X"00",X"00",X"0A",X"A0",
		X"00",X"0A",X"00",X"00",X"0A",X"A0",X"00",X"0A",X"00",X"00",X"0A",X"A0",X"00",X"C3",X"00",X"00",
		X"0A",X"A0",X"0C",X"30",X"00",X"00",X"0A",X"69",X"C3",X"00",X"00",X"00",X"C3",X"06",X"B0",X"00",
		X"00",X"0C",X"30",X"00",X"65",X"DD",X"DD",X"53",X"00",X"C5",X"D5",X"5D",X"55",X"59",X"00",X"A0",
		X"A0",X"0A",X"00",X"06",X"90",X"65",X"30",X"0A",X"00",X"00",X"69",X"00",X"00",X"0A",X"00",X"00",
		X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",
		X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",
		X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"C3",X"00",X"00",X"0A",X"00",X"0C",
		X"30",X"00",X"00",X"CF",X"DD",X"53",X"00",X"C5",X"55",X"55",X"55",X"55",X"51",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"06",X"59",X"00",X"00",X"00",X"00",X"00",
		X"06",X"59",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"55",X"90",X"00",X"00",X"02",X"00",X"00",
		X"69",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"80",X"00",X"00",
		X"00",X"00",X"0A",X"69",X"00",X"00",X"00",X"00",X"C3",X"06",X"90",X"00",X"00",X"0C",X"30",X"00",
		X"65",X"DD",X"DD",X"53",X"00",X"0C",X"55",X"55",X"55",X"55",X"90",X"C3",X"00",X"00",X"00",X"00",
		X"69",X"20",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"C3",X"00",X"00",X"4D",X"55",X"55",X"B0",X"00",X"00",X"02",X"00",X"00",X"69",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"80",X"00",X"00",X"00",X"00",
		X"0A",X"69",X"00",X"00",X"00",X"00",X"C3",X"06",X"90",X"00",X"00",X"0C",X"30",X"00",X"65",X"DD",
		X"DD",X"53",X"00",X"00",X"00",X"04",X"55",X"59",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"C5",
		X"55",X"55",X"55",X"5F",X"51",X"A0",X"00",X"00",X"00",X"0A",X"00",X"65",X"90",X"00",X"00",X"0A",
		X"00",X"00",X"E5",X"59",X"00",X"0A",X"00",X"00",X"A0",X"02",X"00",X"0A",X"00",X"00",X"69",X"00",
		X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"06",X"90",X"00",X"0A",X"00",X"00",
		X"00",X"A0",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",X"00",X"ED",X"DD",X"53",
		X"00",X"0C",X"55",X"55",X"55",X"55",X"90",X"C3",X"00",X"00",X"00",X"00",X"69",X"20",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"CD",X"90",X"00",X"0A",X"00",X"00",X"EF",X"B0",X"00",X"C3",X"C5",X"55",X"77",X"75",X"55",
		X"30",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"65",X"55",X"DD",X"DD",X"55",X"51",X"0C",
		X"55",X"55",X"55",X"55",X"90",X"C3",X"00",X"00",X"00",X"00",X"69",X"A0",X"00",X"00",X"00",X"00",
		X"0A",X"A0",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"C3",X"E5",X"55",X"5D",
		X"55",X"55",X"30",X"A0",X"00",X"02",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",
		X"00",X"06",X"90",X"00",X"00",X"00",X"00",X"00",X"65",X"DD",X"DD",X"55",X"51",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"0E",X"90",X"00",
		X"00",X"00",X"00",X"02",X"69",X"00",X"00",X"00",X"00",X"00",X"06",X"90",X"00",X"00",X"00",X"00",
		X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"06",X"90",X"00",X"00",X"00",X"00",X"00",X"69",X"80",
		X"00",X"00",X"00",X"00",X"0A",X"65",X"55",X"DD",X"DD",X"55",X"53",X"0C",X"55",X"55",X"55",X"55",
		X"90",X"C3",X"00",X"00",X"00",X"00",X"69",X"A0",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",
		X"00",X"00",X"0A",X"65",X"90",X"00",X"00",X"0C",X"53",X"00",X"E5",X"5D",X"55",X"5B",X"00",X"0C",
		X"30",X"02",X"00",X"06",X"90",X"C3",X"00",X"00",X"00",X"00",X"69",X"A0",X"00",X"00",X"00",X"00",
		X"0A",X"A0",X"00",X"00",X"00",X"00",X"0A",X"69",X"00",X"00",X"00",X"00",X"C3",X"06",X"90",X"00",
		X"00",X"0C",X"30",X"00",X"65",X"DD",X"DD",X"53",X"00",X"45",X"55",X"55",X"55",X"59",X"00",X"00",
		X"00",X"00",X"00",X"06",X"90",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"0C",X"55",X"5D",X"55",X"55",X"5B",X"C3",X"00",X"02",
		X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"0A",X"69",X"00",X"00",X"00",X"00",X"C3",X"06",X"90",X"00",X"00",X"0C",
		X"30",X"00",X"65",X"DD",X"DD",X"53",X"00",X"77",X"77",X"77",X"77",X"8A",X"88",X"7E",X"7F",X"89",
		X"7C",X"8B",X"7F",X"76",X"88",X"8B",X"7F",X"7D",X"7C",X"8A",X"88",X"8A",X"88",X"8A",X"88",X"89",
		X"7C",X"76",X"88",X"76",X"88",X"76",X"88",X"7D",X"89",X"7E",X"8B",X"8A",X"76",X"7E",X"8B",X"89",
		X"89",X"8B",X"8B",X"76",X"76",X"8B",X"8B",X"7D",X"89",X"8A",X"76",X"8A",X"76",X"8A",X"76",X"89",
		X"89",X"76",X"76",X"76",X"76",X"76",X"76",X"CF",X"89",X"3B",X"02",X"02",X"72",X"73",X"74",X"75",
		X"FD",X"7E",X"04",X"E6",X"0F",X"87",X"47",X"87",X"87",X"80",X"5F",X"16",X"00",X"21",X"75",X"0B",
		X"19",X"06",X"05",X"5E",X"23",X"56",X"23",X"C5",X"E5",X"7A",X"CB",X"BA",X"21",X"00",X"88",X"19",
		X"EB",X"17",X"38",X"0D",X"CD",X"5C",X"0B",X"21",X"7C",X"00",X"19",X"EB",X"CD",X"5C",X"0B",X"18",
		X"06",X"CD",X"5C",X"0B",X"CD",X"5C",X"0B",X"E1",X"C1",X"10",X"D8",X"C9",X"06",X"02",X"C5",X"21",
		X"D9",X"0B",X"E5",X"CD",X"D8",X"03",X"D9",X"E1",X"CD",X"D8",X"03",X"D9",X"21",X"82",X"FF",X"19",
		X"EB",X"C1",X"10",X"EA",X"C9",X"C9",X"00",X"CF",X"00",X"85",X"01",X"13",X"02",X"C9",X"82",X"89",
		X"00",X"93",X"80",X"4F",X"81",X"15",X"02",X"89",X"82",X"8B",X"80",X"15",X"01",X"87",X"01",X"8F",
		X"82",X"05",X"83",X"8D",X"80",X"45",X"81",X"53",X"01",X"47",X"02",X"8F",X"82",X"8D",X"80",X"97",
		X"00",X"C3",X"00",X"4D",X"82",X"11",X"83",X"C7",X"80",X"15",X"01",X"87",X"01",X"93",X"02",X"C7",
		X"82",X"C7",X"00",X"0F",X"81",X"D3",X"01",X"05",X"02",X"0F",X"83",X"89",X"00",X"D1",X"80",X"93",
		X"01",X"45",X"82",X"0B",X"83",X"C7",X"00",X"11",X"81",X"D1",X"81",X"05",X"02",X"91",X"82",X"85",
		X"80",X"0F",X"81",X"D5",X"01",X"07",X"02",X"4F",X"02",X"00",X"02",X"02",X"78",X"79",X"7A",X"7B",
		X"3A",X"00",X"E0",X"E6",X"80",X"28",X"05",X"CD",X"F4",X"02",X"E6",X"06",X"4F",X"87",X"81",X"4F",
		X"FD",X"7E",X"04",X"E6",X"0F",X"87",X"87",X"87",X"47",X"87",X"80",X"81",X"5F",X"16",X"00",X"21",
		X"3A",X"0C",X"19",X"EB",X"FD",X"E5",X"E1",X"01",X"31",X"00",X"09",X"06",X"06",X"36",X"80",X"23",
		X"1A",X"E6",X"F0",X"C6",X"08",X"77",X"23",X"36",X"00",X"23",X"1A",X"E6",X"0F",X"87",X"87",X"87",
		X"87",X"77",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"13",X"23",X"10",X"DE",X"06",
		X"06",X"11",X"07",X"00",X"36",X"00",X"19",X"10",X"FB",X"C9",X"3A",X"57",X"7C",X"7D",X"A9",X"AD",
		X"4A",X"6D",X"85",X"8C",X"AC",X"C9",X"47",X"4B",X"8D",X"9C",X"A8",X"CB",X"4A",X"57",X"85",X"8D",
		X"A8",X"AD",X"3E",X"48",X"5C",X"8D",X"96",X"AA",X"4D",X"4E",X"57",X"95",X"A9",X"CB",X"47",X"49",
		X"6C",X"AD",X"B9",X"C9",X"49",X"4E",X"6C",X"96",X"AA",X"CB",X"49",X"6A",X"6D",X"AC",X"B6",X"BC",
		X"3A",X"5D",X"86",X"9A",X"9B",X"CB",X"3B",X"5A",X"8B",X"8C",X"96",X"AD",X"3A",X"6D",X"86",X"8B",
		X"AD",X"B6",X"4A",X"57",X"7D",X"96",X"9D",X"CB",X"48",X"6D",X"7C",X"9A",X"A6",X"BC",X"3B",X"5C",
		X"69",X"86",X"8C",X"B6",X"3B",X"48",X"7C",X"7D",X"B6",X"CB",X"4B",X"7C",X"89",X"8A",X"AD",X"C7",
		X"3B",X"4E",X"6A",X"87",X"AB",X"C8",X"3E",X"66",X"7D",X"8C",X"9B",X"CD",X"3E",X"66",X"7C",X"89",
		X"AB",X"C8",X"38",X"5D",X"66",X"8C",X"AC",X"CC",X"4D",X"57",X"86",X"8B",X"B8",X"CD",X"3C",X"58",
		X"7D",X"97",X"9C",X"A8",X"3C",X"57",X"8B",X"8C",X"A8",X"CD",X"36",X"5C",X"5D",X"8C",X"95",X"CC",
		X"3B",X"56",X"7D",X"AC",X"B5",X"BB",X"6B",X"6D",X"85",X"9D",X"A6",X"BC",X"36",X"5C",X"85",X"9D",
		X"BB",X"BC",X"4D",X"57",X"6C",X"6D",X"9D",X"A8",X"3D",X"47",X"5B",X"8C",X"AD",X"B6",X"37",X"48",
		X"5C",X"7D",X"A7",X"CA",X"47",X"48",X"4D",X"6C",X"9D",X"B6",X"56",X"5D",X"69",X"9B",X"9C",X"A5",
		X"3B",X"66",X"6C",X"9A",X"AD",X"B5",X"56",X"6B",X"6C",X"8D",X"96",X"9A",X"3B",X"66",X"6D",X"7D",
		X"95",X"9B",X"4C",X"66",X"6C",X"6D",X"AA",X"BC",X"46",X"5C",X"8A",X"9D",X"B6",X"BB",X"3B",X"6A",
		X"8D",X"96",X"AD",X"BA",X"46",X"4C",X"6A",X"96",X"9D",X"AA",X"3A",X"03",X"A0",X"47",X"E6",X"F0",
		X"28",X"05",X"78",X"E6",X"0F",X"20",X"13",X"DD",X"CB",X"00",X"AE",X"3A",X"00",X"A0",X"CB",X"77",
		X"CA",X"72",X"0F",X"CB",X"6F",X"CA",X"9C",X"0F",X"18",X"07",X"3A",X"06",X"E0",X"A7",X"C2",X"DC",
		X"0E",X"3A",X"A9",X"E1",X"17",X"D8",X"DD",X"7E",X"01",X"A7",X"28",X"04",X"DD",X"35",X"01",X"C9",
		X"DD",X"7E",X"02",X"FE",X"03",X"D2",X"4C",X"0E",X"FE",X"02",X"D2",X"D2",X"0D",X"FE",X"01",X"30",
		X"5D",X"DD",X"7E",X"03",X"A7",X"20",X"53",X"DD",X"34",X"03",X"DD",X"36",X"04",X"00",X"CD",X"85",
		X"04",X"CD",X"6E",X"70",X"CD",X"B0",X"11",X"3A",X"03",X"A0",X"47",X"E6",X"F0",X"28",X"34",X"78",
		X"E6",X"0F",X"28",X"2F",X"21",X"2C",X"11",X"CD",X"03",X"04",X"3A",X"03",X"A0",X"E6",X"0F",X"F5",
		X"11",X"2C",X"89",X"CD",X"FB",X"0F",X"F1",X"47",X"3A",X"03",X"A0",X"E6",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"B8",X"C8",X"11",X"29",X"89",X"CD",X"FB",X"0F",X"21",X"3B",X"11",X"CD",X"03",X"04",X"CD",
		X"03",X"04",X"C9",X"21",X"4C",X"11",X"CD",X"03",X"04",X"C9",X"CD",X"01",X"70",X"C9",X"CD",X"A9",
		X"70",X"C9",X"DD",X"7E",X"03",X"A7",X"20",X"47",X"DD",X"34",X"03",X"DD",X"CB",X"00",X"86",X"DD",
		X"36",X"04",X"FF",X"DD",X"36",X"05",X"01",X"CD",X"85",X"04",X"AF",X"FD",X"77",X"08",X"FD",X"77",
		X"09",X"FD",X"36",X"04",X"01",X"FD",X"77",X"0D",X"FD",X"77",X"16",X"FD",X"77",X"17",X"FD",X"77",
		X"1A",X"CD",X"71",X"06",X"CD",X"C3",X"04",X"3E",X"80",X"32",X"C5",X"E1",X"32",X"12",X"E2",X"32",
		X"C2",X"E2",X"32",X"00",X"E3",X"21",X"00",X"E0",X"CB",X"F6",X"DD",X"36",X"01",X"60",X"C9",X"DD",
		X"CB",X"00",X"46",X"20",X"1B",X"DD",X"35",X"05",X"C0",X"DD",X"6E",X"03",X"26",X"00",X"29",X"11",
		X"D2",X"10",X"19",X"7E",X"DD",X"77",X"04",X"23",X"7E",X"DD",X"77",X"05",X"DD",X"34",X"03",X"C9",
		X"DD",X"34",X"02",X"DD",X"36",X"03",X"00",X"FD",X"36",X"00",X"00",X"C9",X"DD",X"7E",X"03",X"A7",
		X"20",X"06",X"CD",X"85",X"04",X"CD",X"86",X"10",X"DD",X"7E",X"03",X"FE",X"0E",X"30",X"57",X"FE",
		X"0D",X"30",X"3F",X"FE",X"08",X"30",X"18",X"21",X"8F",X"15",X"CD",X"25",X"04",X"DD",X"34",X"03",
		X"DD",X"36",X"01",X"02",X"DD",X"7E",X"03",X"FE",X"08",X"D8",X"DD",X"36",X"01",X"10",X"C9",X"D6",
		X"08",X"87",X"5F",X"16",X"00",X"21",X"9B",X"15",X"19",X"5E",X"23",X"56",X"EB",X"CD",X"03",X"04",
		X"DD",X"34",X"03",X"DD",X"36",X"01",X"04",X"DD",X"7E",X"03",X"FE",X"0D",X"D8",X"DD",X"36",X"01",
		X"08",X"C9",X"21",X"CA",X"15",X"06",X"0A",X"C5",X"CD",X"03",X"04",X"C1",X"10",X"F9",X"DD",X"34",
		X"03",X"DD",X"36",X"01",X"10",X"C9",X"06",X"0A",X"11",X"36",X"89",X"21",X"17",X"E0",X"C5",X"D5",
		X"E5",X"CD",X"11",X"16",X"E1",X"01",X"0A",X"00",X"09",X"D1",X"1B",X"1B",X"C1",X"10",X"EF",X"DD",
		X"36",X"01",X"FF",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"00",X"C9",X"FE",X"01",X"20",X"0A",
		X"3A",X"00",X"A0",X"CB",X"6F",X"CA",X"9C",X"0F",X"18",X"0D",X"3A",X"00",X"A0",X"CB",X"77",X"CA",
		X"72",X"0F",X"CB",X"6F",X"CA",X"9C",X"0F",X"3A",X"A9",X"E1",X"17",X"D8",X"DD",X"CB",X"00",X"6E",
		X"20",X"1E",X"DD",X"CB",X"00",X"EE",X"CD",X"FF",X"05",X"CD",X"85",X"04",X"CD",X"6E",X"70",X"21",
		X"59",X"11",X"CD",X"03",X"04",X"CD",X"03",X"04",X"CD",X"03",X"04",X"CD",X"B0",X"11",X"18",X"05",
		X"DD",X"CB",X"00",X"66",X"C8",X"DD",X"CB",X"00",X"A6",X"21",X"75",X"11",X"3A",X"06",X"E0",X"3D",
		X"28",X"03",X"21",X"8D",X"11",X"CD",X"03",X"04",X"21",X"A6",X"11",X"CD",X"03",X"04",X"3A",X"06",
		X"E0",X"FE",X"0A",X"38",X"02",X"3E",X"09",X"32",X"24",X"8F",X"47",X"3E",X"0B",X"32",X"24",X"8B",
		X"11",X"ED",X"88",X"3E",X"09",X"90",X"28",X"09",X"EB",X"11",X"20",X"00",X"19",X"3D",X"20",X"FC",
		X"EB",X"C5",X"08",X"3E",X"32",X"08",X"3E",X"4D",X"01",X"02",X"02",X"CD",X"42",X"04",X"C1",X"10",
		X"F0",X"C9",X"3E",X"E0",X"32",X"00",X"E0",X"3A",X"03",X"A0",X"47",X"E6",X"F0",X"28",X"0E",X"78",
		X"E6",X"0F",X"28",X"09",X"3A",X"06",X"E0",X"D6",X"02",X"27",X"32",X"06",X"E0",X"CD",X"85",X"04",
		X"FD",X"21",X"1C",X"E1",X"CD",X"64",X"06",X"CD",X"A7",X"10",X"18",X"1B",X"3E",X"C0",X"32",X"00",
		X"E0",X"3A",X"03",X"A0",X"47",X"E6",X"F0",X"28",X"0E",X"78",X"E6",X"0F",X"28",X"09",X"3A",X"06",
		X"E0",X"D6",X"01",X"27",X"32",X"06",X"E0",X"CD",X"85",X"04",X"FD",X"21",X"97",X"E0",X"CD",X"64",
		X"06",X"CD",X"C3",X"04",X"CD",X"FF",X"05",X"32",X"A9",X"E1",X"32",X"B6",X"E1",X"DD",X"77",X"00",
		X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"3E",X"80",X"32",X"C5",X"E1",X"32",X"12",
		X"E2",X"32",X"C2",X"E2",X"32",X"00",X"E3",X"32",X"01",X"E0",X"3A",X"00",X"E0",X"32",X"00",X"98",
		X"3E",X"25",X"CD",X"EA",X"02",X"3E",X"21",X"CD",X"EA",X"02",X"C9",X"87",X"F5",X"D9",X"5F",X"16",
		X"00",X"21",X"2A",X"10",X"19",X"5E",X"23",X"56",X"EB",X"06",X"0F",X"3E",X"09",X"CD",X"0F",X"04",
		X"D9",X"21",X"20",X"02",X"19",X"EB",X"F1",X"4F",X"06",X"00",X"21",X"4D",X"02",X"09",X"EB",X"1A",
		X"77",X"01",X"00",X"01",X"09",X"13",X"1A",X"77",X"D9",X"C9",X"4A",X"10",X"4A",X"10",X"4A",X"10",
		X"4A",X"10",X"4A",X"10",X"4A",X"10",X"68",X"10",X"77",X"10",X"68",X"10",X"77",X"10",X"68",X"10",
		X"59",X"10",X"59",X"10",X"59",X"10",X"59",X"10",X"4A",X"10",X"29",X"29",X"0C",X"18",X"12",X"17",
		X"29",X"29",X"29",X"29",X"19",X"15",X"0A",X"22",X"29",X"29",X"29",X"0C",X"18",X"12",X"17",X"29",
		X"29",X"29",X"29",X"19",X"15",X"0A",X"22",X"1C",X"29",X"29",X"0C",X"18",X"12",X"17",X"1C",X"29",
		X"29",X"29",X"19",X"15",X"0A",X"22",X"29",X"29",X"29",X"0C",X"18",X"12",X"17",X"1C",X"29",X"29",
		X"29",X"19",X"15",X"0A",X"22",X"1C",X"3A",X"03",X"A0",X"47",X"E6",X"0F",X"28",X"04",X"78",X"E6",
		X"F0",X"C0",X"21",X"99",X"10",X"CD",X"03",X"04",X"C9",X"22",X"8A",X"09",X"0A",X"0F",X"1B",X"0E",
		X"0E",X"29",X"19",X"15",X"0A",X"22",X"29",X"21",X"83",X"8C",X"11",X"12",X"E6",X"3E",X"18",X"01",
		X"1A",X"00",X"ED",X"B0",X"01",X"06",X"00",X"09",X"3D",X"20",X"F4",X"21",X"12",X"E4",X"11",X"AF",
		X"E8",X"3E",X"0C",X"01",X"0D",X"00",X"ED",X"A0",X"23",X"EA",X"C6",X"10",X"01",X"06",X"00",X"09",
		X"3D",X"20",X"F0",X"C9",X"FB",X"4D",X"FE",X"01",X"EF",X"F0",X"F7",X"43",X"FE",X"48",X"FF",X"3C",
		X"FB",X"30",X"FF",X"96",X"FB",X"0A",X"F7",X"60",X"FE",X"18",X"F7",X"30",X"FE",X"18",X"F7",X"18",
		X"FB",X"48",X"FD",X"18",X"FE",X"43",X"FD",X"48",X"FE",X"36",X"E7",X"01",X"F7",X"3A",X"FE",X"18",
		X"FD",X"48",X"FE",X"18",X"F7",X"4C",X"ED",X"01",X"FE",X"30",X"F7",X"30",X"FE",X"18",X"FD",X"4C",
		X"E7",X"01",X"FB",X"18",X"FD",X"60",X"FE",X"18",X"FD",X"18",X"FB",X"50",X"EE",X"01",X"F7",X"18",
		X"FE",X"18",X"FD",X"57",X"FB",X"8A",X"EE",X"01",X"F7",X"FF",X"FF",X"FF",X"6F",X"89",X"09",X"0B",
		X"12",X"17",X"1C",X"0E",X"1B",X"1D",X"29",X"0C",X"18",X"12",X"17",X"ED",X"88",X"09",X"05",X"1B",
		X"12",X"10",X"11",X"1D",X"EA",X"88",X"09",X"04",X"15",X"0E",X"0F",X"1D",X"8F",X"89",X"09",X"09",
		X"0F",X"1B",X"0E",X"0E",X"29",X"19",X"15",X"0A",X"22",X"B2",X"89",X"09",X"05",X"19",X"1B",X"0E",
		X"1C",X"1C",X"6B",X"89",X"09",X"09",X"19",X"1B",X"0E",X"1C",X"0E",X"17",X"1D",X"0E",X"0D",X"E9",
		X"89",X"09",X"02",X"0B",X"22",X"D0",X"88",X"09",X"14",X"01",X"29",X"19",X"15",X"0A",X"22",X"0E",
		X"1B",X"29",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"29",X"18",X"17",X"15",X"22",X"B0",X"88",X"09",
		X"15",X"01",X"29",X"18",X"1B",X"29",X"02",X"29",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"29",
		X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"44",X"8A",X"0B",X"06",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",
		X"3E",X"36",X"08",X"3E",X"3E",X"01",X"0B",X"02",X"11",X"06",X"89",X"CD",X"42",X"04",X"21",X"C5",
		X"11",X"CD",X"03",X"04",X"C9",X"66",X"8A",X"2C",X"05",X"2A",X"01",X"09",X"08",X"02",X"DD",X"CB",
		X"00",X"76",X"20",X"3B",X"21",X"00",X"E0",X"CB",X"B6",X"CD",X"2A",X"06",X"C0",X"3A",X"00",X"E0",
		X"87",X"D2",X"C0",X"14",X"CD",X"80",X"5A",X"DD",X"CB",X"00",X"F6",X"DD",X"36",X"01",X"40",X"DD",
		X"36",X"03",X"00",X"FD",X"7E",X"00",X"A7",X"20",X"05",X"DD",X"36",X"02",X"00",X"C9",X"CD",X"DE",
		X"14",X"7E",X"A7",X"28",X"05",X"DD",X"36",X"02",X"03",X"C9",X"DD",X"36",X"02",X"05",X"C9",X"DD",
		X"7E",X"01",X"A7",X"28",X"04",X"DD",X"35",X"01",X"C9",X"21",X"01",X"E0",X"CB",X"FE",X"DD",X"7E",
		X"02",X"FE",X"06",X"D2",X"C0",X"14",X"FE",X"05",X"D2",X"A0",X"14",X"FE",X"04",X"D2",X"78",X"14",
		X"FE",X"03",X"D2",X"2C",X"14",X"FE",X"02",X"D2",X"F6",X"13",X"FE",X"01",X"30",X"71",X"DD",X"7E",
		X"03",X"A7",X"20",X"21",X"11",X"51",X"89",X"01",X"0B",X"03",X"CD",X"6C",X"04",X"11",X"51",X"81",
		X"01",X"0B",X"03",X"CD",X"6C",X"04",X"DD",X"36",X"01",X"10",X"DD",X"34",X"03",X"3E",X"21",X"06",
		X"00",X"CD",X"D9",X"02",X"C9",X"DD",X"7E",X"03",X"3D",X"21",X"71",X"15",X"CD",X"25",X"04",X"DD",
		X"36",X"01",X"08",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"0A",X"D8",X"DD",X"36",X"01",X"DC",
		X"DD",X"36",X"03",X"00",X"CD",X"8B",X"16",X"30",X"10",X"DD",X"36",X"02",X"01",X"CD",X"DE",X"14",
		X"7E",X"A7",X"C0",X"21",X"A1",X"E1",X"CB",X"FE",X"C9",X"CD",X"DE",X"14",X"7E",X"A7",X"28",X"05",
		X"DD",X"36",X"02",X"03",X"C9",X"DD",X"36",X"02",X"06",X"21",X"A1",X"E1",X"CB",X"FE",X"C9",X"DD",
		X"7E",X"03",X"A7",X"20",X"03",X"CD",X"85",X"04",X"DD",X"7E",X"03",X"FE",X"13",X"D2",X"CA",X"13",
		X"FE",X"12",X"D2",X"98",X"13",X"FE",X"11",X"D2",X"82",X"13",X"FE",X"10",X"D2",X"6C",X"13",X"FE",
		X"0F",X"D2",X"56",X"13",X"FE",X"0E",X"30",X"57",X"FE",X"0D",X"30",X"3F",X"FE",X"08",X"30",X"18",
		X"21",X"8F",X"15",X"CD",X"25",X"04",X"DD",X"34",X"03",X"DD",X"36",X"01",X"02",X"DD",X"7E",X"03",
		X"FE",X"08",X"D8",X"DD",X"36",X"01",X"10",X"C9",X"D6",X"08",X"87",X"5F",X"16",X"00",X"21",X"9B",
		X"15",X"19",X"5E",X"23",X"56",X"EB",X"CD",X"03",X"04",X"DD",X"34",X"03",X"DD",X"36",X"01",X"04",
		X"DD",X"7E",X"03",X"FE",X"0D",X"D8",X"DD",X"36",X"01",X"08",X"C9",X"21",X"CA",X"15",X"06",X"0A",
		X"C5",X"CD",X"03",X"04",X"C1",X"10",X"F9",X"DD",X"34",X"03",X"DD",X"36",X"01",X"08",X"C9",X"06",
		X"0A",X"11",X"36",X"89",X"21",X"17",X"E0",X"C5",X"D5",X"E5",X"3E",X"0A",X"90",X"DD",X"BE",X"04",
		X"C4",X"11",X"16",X"E1",X"01",X"0A",X"00",X"09",X"D1",X"1B",X"1B",X"C1",X"10",X"E9",X"DD",X"34",
		X"03",X"DD",X"36",X"01",X"08",X"C9",X"11",X"36",X"89",X"21",X"17",X"E0",X"CD",X"2D",X"19",X"0E",
		X"3E",X"CD",X"3B",X"16",X"DD",X"34",X"03",X"DD",X"36",X"01",X"04",X"C9",X"11",X"96",X"8A",X"21",
		X"1D",X"E0",X"CD",X"2D",X"19",X"0E",X"3E",X"CD",X"4F",X"16",X"DD",X"34",X"03",X"DD",X"36",X"01",
		X"04",X"C9",X"11",X"F6",X"8A",X"21",X"1E",X"E0",X"CD",X"2D",X"19",X"0E",X"3E",X"CD",X"64",X"16",
		X"DD",X"34",X"03",X"DD",X"36",X"01",X"04",X"C9",X"DD",X"36",X"05",X"1C",X"DD",X"36",X"06",X"20",
		X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"0A",X"DD",X"36",X"09",X"00",X"DD",X"36",X"0A",X"00",
		X"DD",X"36",X"0B",X"00",X"DD",X"36",X"0C",X"00",X"CD",X"60",X"18",X"DD",X"34",X"03",X"DD",X"36",
		X"01",X"04",X"3E",X"25",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"DD",X"46",X"05",X"DD",X"4E",X"06",
		X"0B",X"DD",X"70",X"05",X"DD",X"71",X"06",X"78",X"B1",X"28",X"09",X"CD",X"2B",X"17",X"DD",X"7E",
		X"07",X"FE",X"03",X"D8",X"DD",X"36",X"02",X"02",X"DD",X"36",X"01",X"08",X"DD",X"36",X"03",X"00",
		X"3E",X"25",X"CD",X"EA",X"02",X"C9",X"DD",X"7E",X"03",X"A7",X"20",X"24",X"11",X"E3",X"81",X"01",
		X"05",X"15",X"CD",X"6C",X"04",X"CD",X"0C",X"18",X"21",X"A1",X"E1",X"CB",X"7E",X"20",X"08",X"DD",
		X"34",X"03",X"DD",X"36",X"01",X"78",X"C9",X"DD",X"36",X"02",X"06",X"DD",X"36",X"01",X"FF",X"C9",
		X"CD",X"85",X"04",X"DD",X"36",X"02",X"03",X"DD",X"36",X"03",X"00",X"C9",X"DD",X"7E",X"03",X"A7",
		X"20",X"1D",X"CD",X"EB",X"14",X"11",X"11",X"89",X"01",X"0F",X"03",X"CD",X"6C",X"04",X"11",X"11",
		X"81",X"01",X"0F",X"03",X"CD",X"6C",X"04",X"DD",X"36",X"01",X"10",X"DD",X"34",X"03",X"C9",X"FE",
		X"0E",X"30",X"19",X"3D",X"21",X"7E",X"15",X"CD",X"25",X"04",X"DD",X"36",X"01",X"08",X"DD",X"34",
		X"03",X"DD",X"7E",X"03",X"FE",X"0E",X"D8",X"DD",X"36",X"01",X"44",X"C9",X"DD",X"36",X"02",X"04",
		X"DD",X"36",X"03",X"00",X"CD",X"05",X"15",X"C9",X"3A",X"00",X"E0",X"E6",X"BF",X"EE",X"10",X"21",
		X"02",X"A0",X"CB",X"6E",X"28",X"05",X"EE",X"01",X"32",X"00",X"98",X"32",X"00",X"E0",X"FD",X"21",
		X"97",X"E0",X"E6",X"10",X"28",X"04",X"FD",X"21",X"1C",X"E1",X"CD",X"1F",X"15",X"CD",X"C3",X"04",
		X"CD",X"A1",X"06",X"21",X"00",X"E0",X"CB",X"9E",X"CB",X"F6",X"23",X"CB",X"B6",X"3E",X"80",X"32",
		X"C5",X"E1",X"32",X"12",X"E2",X"32",X"C2",X"E2",X"32",X"00",X"E3",X"DD",X"36",X"00",X"00",X"C9",
		X"CD",X"FF",X"05",X"21",X"A1",X"E1",X"CB",X"FE",X"CB",X"C6",X"3A",X"00",X"E0",X"E6",X"26",X"32",
		X"00",X"E0",X"32",X"00",X"98",X"AF",X"32",X"01",X"E0",X"DD",X"36",X"00",X"00",X"C9",X"21",X"1C",
		X"E1",X"3A",X"00",X"E0",X"CB",X"67",X"C8",X"21",X"97",X"E0",X"C9",X"21",X"11",X"8D",X"11",X"82",
		X"E8",X"0E",X"0F",X"06",X"03",X"7E",X"12",X"13",X"23",X"10",X"FA",X"79",X"01",X"1D",X"00",X"09",
		X"4F",X"0D",X"20",X"EF",X"C9",X"21",X"11",X"8D",X"11",X"82",X"E8",X"0E",X"0F",X"06",X"03",X"1A",
		X"77",X"13",X"23",X"10",X"FA",X"79",X"01",X"1D",X"00",X"09",X"4F",X"0D",X"20",X"EF",X"C9",X"CD",
		X"A1",X"06",X"21",X"83",X"8C",X"11",X"12",X"E6",X"0E",X"18",X"06",X"1A",X"7E",X"08",X"1A",X"77",
		X"08",X"12",X"13",X"23",X"10",X"F6",X"23",X"23",X"23",X"23",X"23",X"23",X"0D",X"20",X"EB",X"21",
		X"83",X"88",X"01",X"18",X"1A",X"3E",X"00",X"CD",X"5C",X"04",X"21",X"17",X"0B",X"CD",X"D4",X"03",
		X"21",X"12",X"E4",X"11",X"AF",X"E8",X"0E",X"0C",X"06",X"0D",X"7E",X"08",X"1A",X"77",X"08",X"12",
		X"23",X"36",X"FF",X"13",X"23",X"10",X"F3",X"23",X"23",X"23",X"23",X"23",X"23",X"0D",X"20",X"E8",
		X"C9",X"72",X"89",X"2E",X"09",X"10",X"0A",X"16",X"0E",X"29",X"18",X"1F",X"0E",X"1B",X"32",X"89",
		X"3E",X"0D",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"29",X"0C",X"11",X"0A",X"17",X"10",X"0E",X"9B",
		X"89",X"2C",X"08",X"11",X"12",X"2B",X"1C",X"0C",X"18",X"1B",X"0E",X"A5",X"15",X"AC",X"15",X"B4",
		X"15",X"BB",X"15",X"C3",X"15",X"B8",X"88",X"89",X"03",X"00",X"01",X"02",X"58",X"89",X"89",X"04",
		X"03",X"04",X"05",X"FE",X"18",X"8A",X"89",X"03",X"06",X"07",X"08",X"98",X"8A",X"89",X"04",X"09",
		X"0A",X"0B",X"0C",X"38",X"8B",X"89",X"03",X"0D",X"0E",X"0F",X"B6",X"88",X"2C",X"03",X"1D",X"18",
		X"19",X"B4",X"88",X"26",X"03",X"02",X"17",X"0D",X"B2",X"88",X"26",X"03",X"03",X"1B",X"0D",X"B0",
		X"88",X"26",X"03",X"04",X"1D",X"11",X"AE",X"88",X"26",X"03",X"05",X"1D",X"11",X"AC",X"88",X"26",
		X"03",X"06",X"1D",X"11",X"AA",X"88",X"26",X"03",X"07",X"1D",X"11",X"A8",X"88",X"26",X"03",X"08",
		X"1D",X"11",X"A6",X"88",X"26",X"03",X"09",X"1D",X"11",X"84",X"88",X"26",X"04",X"01",X"00",X"1D",
		X"11",X"CD",X"39",X"16",X"D5",X"D9",X"D1",X"21",X"20",X"00",X"19",X"EB",X"D9",X"3E",X"09",X"06",
		X"03",X"CD",X"0F",X"04",X"D9",X"21",X"20",X"00",X"19",X"E5",X"D9",X"D1",X"CD",X"4D",X"16",X"EB",
		X"01",X"20",X"00",X"09",X"EB",X"CD",X"62",X"16",X"C9",X"0E",X"09",X"D5",X"E5",X"11",X"17",X"E0",
		X"A7",X"ED",X"52",X"20",X"02",X"0E",X"2C",X"E1",X"D1",X"CD",X"A1",X"03",X"C9",X"0E",X"09",X"23",
		X"23",X"23",X"CB",X"4E",X"2B",X"2B",X"2B",X"28",X"02",X"0E",X"2C",X"AF",X"06",X"02",X"CD",X"A4",
		X"03",X"C9",X"0E",X"09",X"23",X"23",X"CB",X"46",X"2B",X"2B",X"28",X"02",X"0E",X"2C",X"AF",X"06",
		X"02",X"CD",X"A4",X"03",X"79",X"12",X"E5",X"21",X"00",X"04",X"19",X"36",X"2D",X"21",X"20",X"00",
		X"19",X"EB",X"E1",X"3E",X"80",X"06",X"02",X"CD",X"A4",X"03",X"C9",X"FD",X"E5",X"D1",X"13",X"21",
		X"17",X"E0",X"01",X"00",X"0A",X"D5",X"E5",X"C5",X"CD",X"21",X"17",X"30",X"0C",X"C1",X"E1",X"11",
		X"0A",X"00",X"19",X"D1",X"0C",X"10",X"EE",X"A7",X"C9",X"C1",X"DD",X"71",X"04",X"3E",X"09",X"91",
		X"28",X"0E",X"21",X"70",X"E0",X"11",X"7A",X"E0",X"01",X"0A",X"00",X"ED",X"B8",X"3D",X"20",X"F8",
		X"D1",X"E1",X"01",X"03",X"00",X"ED",X"B0",X"06",X"03",X"3E",X"29",X"12",X"13",X"10",X"FC",X"01",
		X"03",X"00",X"ED",X"B0",X"21",X"20",X"E0",X"11",X"0A",X"00",X"06",X"0A",X"36",X"00",X"19",X"10",
		X"FB",X"11",X"1D",X"E0",X"21",X"27",X"E0",X"06",X"09",X"1A",X"BE",X"30",X"02",X"54",X"5D",X"C5",
		X"01",X"0A",X"00",X"09",X"C1",X"10",X"F2",X"EB",X"23",X"23",X"23",X"CB",X"CE",X"11",X"1E",X"E0",
		X"21",X"28",X"E0",X"06",X"09",X"C5",X"D5",X"E5",X"06",X"02",X"CD",X"23",X"17",X"E1",X"D1",X"30",
		X"02",X"54",X"5D",X"01",X"0A",X"00",X"09",X"C1",X"10",X"EB",X"EB",X"23",X"23",X"CB",X"C6",X"37",
		X"C9",X"06",X"03",X"1A",X"BE",X"C0",X"13",X"23",X"10",X"F9",X"C9",X"DD",X"7E",X"0B",X"A7",X"28",
		X"05",X"DD",X"35",X"0B",X"18",X"3A",X"CD",X"00",X"18",X"CB",X"66",X"20",X"33",X"DD",X"36",X"0B",
		X"20",X"DD",X"7E",X"07",X"57",X"0F",X"0F",X"0F",X"4F",X"06",X"00",X"21",X"16",X"8E",X"09",X"EB",
		X"4C",X"21",X"1A",X"E0",X"09",X"CD",X"2D",X"19",X"DD",X"7E",X"08",X"12",X"77",X"11",X"00",X"FC",
		X"19",X"36",X"3E",X"DD",X"34",X"07",X"DD",X"7E",X"07",X"FE",X"03",X"D0",X"DD",X"36",X"08",X"0A",
		X"DD",X"7E",X"0C",X"A7",X"28",X"05",X"DD",X"35",X"0C",X"18",X"32",X"CD",X"00",X"18",X"7E",X"2F",
		X"E6",X"0F",X"28",X"29",X"DD",X"36",X"0C",X"0F",X"E6",X"06",X"28",X"10",X"DD",X"34",X"08",X"DD",
		X"7E",X"08",X"FE",X"2A",X"38",X"14",X"DD",X"36",X"08",X"0A",X"18",X"0E",X"DD",X"35",X"08",X"DD",
		X"7E",X"08",X"FE",X"0A",X"30",X"04",X"DD",X"36",X"08",X"29",X"CD",X"43",X"18",X"DD",X"34",X"09",
		X"DD",X"7E",X"09",X"E6",X"1F",X"28",X"31",X"FE",X"14",X"20",X"33",X"11",X"36",X"89",X"CD",X"2D",
		X"19",X"01",X"06",X"01",X"CD",X"6C",X"04",X"21",X"A0",X"00",X"19",X"EB",X"01",X"08",X"01",X"CD",
		X"6C",X"04",X"DD",X"7E",X"07",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"16",X"8E",X"19",X"EB",
		X"CD",X"2D",X"19",X"EB",X"36",X"29",X"18",X"06",X"CD",X"0C",X"18",X"CD",X"43",X"18",X"DD",X"34",
		X"0A",X"DD",X"7E",X"0A",X"FE",X"18",X"38",X"04",X"DD",X"36",X"0A",X"00",X"CD",X"60",X"18",X"C9",
		X"21",X"00",X"A0",X"3A",X"00",X"E0",X"1F",X"D0",X"21",X"01",X"A0",X"C9",X"11",X"36",X"89",X"21",
		X"17",X"E0",X"CD",X"2D",X"19",X"0E",X"3E",X"CD",X"3B",X"16",X"D5",X"D9",X"D1",X"21",X"20",X"00",
		X"19",X"EB",X"D9",X"3E",X"3E",X"06",X"03",X"CD",X"0F",X"04",X"D9",X"21",X"20",X"00",X"19",X"E5",
		X"D9",X"D1",X"0E",X"3E",X"CD",X"4F",X"16",X"EB",X"01",X"20",X"00",X"09",X"EB",X"0E",X"3E",X"CD",
		X"64",X"16",X"C9",X"DD",X"7E",X"07",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"16",X"8A",X"19",
		X"EB",X"CD",X"2D",X"19",X"EB",X"36",X"22",X"11",X"00",X"04",X"19",X"DD",X"7E",X"08",X"77",X"C9",
		X"DD",X"7E",X"0A",X"47",X"E6",X"07",X"C0",X"78",X"0F",X"0F",X"0F",X"4F",X"78",X"87",X"91",X"5F",
		X"DD",X"7E",X"07",X"57",X"87",X"87",X"4F",X"87",X"47",X"87",X"87",X"80",X"81",X"82",X"83",X"5F",
		X"16",X"00",X"21",X"A6",X"18",X"19",X"E5",X"11",X"F5",X"81",X"CD",X"2D",X"19",X"E1",X"D5",X"D9",
		X"D1",X"D9",X"3E",X"87",X"01",X"05",X"03",X"CD",X"E2",X"03",X"21",X"21",X"00",X"19",X"EB",X"01",
		X"03",X"01",X"CD",X"6C",X"04",X"C9",X"41",X"44",X"47",X"4B",X"29",X"4C",X"51",X"29",X"52",X"50",
		X"29",X"53",X"56",X"59",X"5C",X"40",X"43",X"46",X"4A",X"29",X"4E",X"50",X"29",X"54",X"4F",X"29",
		X"52",X"55",X"58",X"5B",X"42",X"45",X"48",X"49",X"29",X"4D",X"4F",X"29",X"53",X"51",X"29",X"54",
		X"57",X"5A",X"5D",X"40",X"43",X"46",X"4F",X"29",X"52",X"49",X"29",X"4C",X"4F",X"29",X"52",X"55",
		X"58",X"5B",X"41",X"44",X"47",X"50",X"29",X"53",X"4A",X"29",X"4D",X"50",X"29",X"53",X"56",X"59",
		X"5C",X"42",X"45",X"48",X"51",X"29",X"54",X"4B",X"29",X"4E",X"51",X"29",X"54",X"57",X"5A",X"5D",
		X"42",X"45",X"48",X"51",X"29",X"54",X"50",X"29",X"52",X"4A",X"29",X"4C",X"57",X"5A",X"5D",X"41",
		X"44",X"47",X"50",X"29",X"53",X"4F",X"29",X"54",X"49",X"29",X"4E",X"56",X"59",X"5C",X"40",X"43",
		X"46",X"4F",X"29",X"52",X"51",X"29",X"53",X"4B",X"29",X"4D",X"55",X"58",X"5B",X"DD",X"7E",X"04",
		X"A7",X"C8",X"01",X"0A",X"00",X"09",X"1B",X"1B",X"3D",X"20",X"FA",X"C9",X"AF",X"32",X"A9",X"E1",
		X"DD",X"CB",X"00",X"76",X"20",X"13",X"DD",X"CB",X"00",X"F6",X"DD",X"36",X"01",X"B4",X"CD",X"80",
		X"5A",X"3E",X"22",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"DD",X"7E",X"01",X"A7",X"28",X"04",X"DD",
		X"35",X"01",X"C9",X"3A",X"01",X"E0",X"E6",X"20",X"C0",X"21",X"00",X"E0",X"CB",X"B6",X"CD",X"2A",
		X"06",X"C0",X"3A",X"00",X"E0",X"87",X"38",X"0A",X"21",X"A1",X"E1",X"CB",X"C6",X"DD",X"36",X"00",
		X"00",X"C9",X"DD",X"CB",X"00",X"6E",X"28",X"12",X"DD",X"CB",X"00",X"66",X"20",X"08",X"DD",X"CB",
		X"00",X"E6",X"DD",X"36",X"02",X"00",X"CD",X"A5",X"73",X"C9",X"DD",X"CB",X"00",X"5E",X"28",X"12",
		X"DD",X"CB",X"00",X"56",X"20",X"08",X"DD",X"CB",X"00",X"D6",X"DD",X"36",X"02",X"00",X"CD",X"90",
		X"75",X"C9",X"DD",X"CB",X"00",X"46",X"20",X"27",X"DD",X"CB",X"00",X"C6",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"03",X"00",X"FD",X"7E",X"04",X"E6",X"0F",X"28",X"0F",X"FE",X"03",X"28",X"07",X"FE",
		X"06",X"28",X"03",X"FE",X"09",X"C0",X"DD",X"34",X"02",X"C9",X"DD",X"36",X"02",X"06",X"C9",X"DD",
		X"7E",X"02",X"A7",X"28",X"0C",X"FE",X"06",X"30",X"04",X"CD",X"6A",X"79",X"C9",X"CD",X"E1",X"7A",
		X"C9",X"FD",X"7E",X"04",X"C6",X"01",X"27",X"FD",X"77",X"04",X"21",X"85",X"04",X"06",X"1A",X"AF",
		X"86",X"23",X"10",X"FC",X"21",X"47",X"05",X"06",X"08",X"86",X"23",X"10",X"FC",X"FE",X"4F",X"20",
		X"06",X"FD",X"34",X"08",X"FD",X"34",X"09",X"FD",X"34",X"00",X"CD",X"76",X"1A",X"FE",X"05",X"38",
		X"02",X"3E",X"04",X"5F",X"16",X"00",X"21",X"71",X"1A",X"19",X"7E",X"FD",X"77",X"0A",X"FD",X"36",
		X"0B",X"9F",X"FD",X"E5",X"D1",X"21",X"1C",X"00",X"19",X"EB",X"01",X"23",X"00",X"09",X"01",X"0E",
		X"00",X"ED",X"B0",X"EB",X"36",X"00",X"54",X"5D",X"13",X"01",X"06",X"00",X"ED",X"B0",X"CD",X"85",
		X"04",X"CD",X"8E",X"06",X"21",X"00",X"E0",X"CB",X"9E",X"CB",X"F6",X"23",X"CB",X"B6",X"3E",X"80",
		X"32",X"C5",X"E1",X"32",X"12",X"E2",X"32",X"C2",X"E2",X"32",X"00",X"E3",X"DD",X"36",X"00",X"00",
		X"C9",X"06",X"06",X"08",X"08",X"08",X"FD",X"7E",X"08",X"21",X"00",X"E0",X"CB",X"7E",X"C8",X"FE",
		X"40",X"D0",X"4F",X"3A",X"02",X"A0",X"E6",X"03",X"28",X"09",X"FE",X"03",X"28",X"0B",X"79",X"87",
		X"C6",X"01",X"C9",X"79",X"87",X"87",X"C6",X"03",X"C9",X"79",X"C9",X"DD",X"56",X"01",X"DD",X"5E",
		X"03",X"CD",X"89",X"1D",X"06",X"01",X"CD",X"87",X"1B",X"DD",X"71",X"0B",X"23",X"CD",X"71",X"1B",
		X"DD",X"71",X"0C",X"11",X"E0",X"FF",X"19",X"05",X"CD",X"71",X"1B",X"DD",X"71",X"0A",X"2B",X"CD",
		X"87",X"1B",X"DD",X"71",X"09",X"DD",X"7E",X"07",X"F6",X"04",X"EE",X"08",X"DD",X"77",X"07",X"C9",
		X"DD",X"56",X"01",X"DD",X"5E",X"03",X"CD",X"89",X"1D",X"06",X"04",X"CD",X"87",X"1B",X"DD",X"71",
		X"0C",X"2B",X"CD",X"71",X"1B",X"DD",X"71",X"0B",X"11",X"E0",X"FF",X"19",X"04",X"CD",X"71",X"1B",
		X"DD",X"71",X"09",X"23",X"CD",X"87",X"1B",X"DD",X"71",X"0A",X"DD",X"7E",X"07",X"F6",X"04",X"EE",
		X"08",X"DD",X"77",X"07",X"C9",X"DD",X"56",X"01",X"DD",X"5E",X"03",X"CD",X"89",X"1D",X"06",X"02",
		X"CD",X"87",X"1B",X"DD",X"71",X"0A",X"2B",X"04",X"CD",X"87",X"1B",X"DD",X"71",X"09",X"11",X"20",
		X"00",X"19",X"CD",X"71",X"1B",X"DD",X"71",X"0B",X"23",X"05",X"CD",X"71",X"1B",X"DD",X"71",X"0C",
		X"DD",X"7E",X"07",X"F6",X"04",X"EE",X"08",X"DD",X"77",X"07",X"C9",X"DD",X"56",X"01",X"DD",X"5E",
		X"03",X"CD",X"89",X"1D",X"06",X"07",X"CD",X"87",X"1B",X"DD",X"71",X"0C",X"2B",X"05",X"CD",X"87",
		X"1B",X"DD",X"71",X"0B",X"11",X"E0",X"FF",X"19",X"CD",X"71",X"1B",X"DD",X"71",X"09",X"23",X"04",
		X"CD",X"71",X"1B",X"DD",X"71",X"0A",X"DD",X"7E",X"07",X"F6",X"04",X"EE",X"08",X"DD",X"77",X"07",
		X"C9",X"78",X"87",X"87",X"5F",X"16",X"00",X"E5",X"21",X"C1",X"1B",X"19",X"EB",X"E1",X"0E",X"04",
		X"1A",X"BE",X"C8",X"13",X"0D",X"20",X"F9",X"7E",X"4F",X"D6",X"77",X"D8",X"FE",X"1D",X"30",X"10",
		X"87",X"87",X"87",X"80",X"D9",X"5F",X"16",X"00",X"21",X"E1",X"1B",X"19",X"7E",X"D9",X"77",X"C9",
		X"FE",X"25",X"30",X"0E",X"D6",X"1D",X"D9",X"5F",X"16",X"00",X"21",X"C9",X"1C",X"19",X"7E",X"D9",
		X"77",X"C9",X"D6",X"25",X"1F",X"D9",X"5F",X"16",X"00",X"21",X"D1",X"1C",X"19",X"7E",X"D9",X"77",
		X"C9",X"7C",X"80",X"84",X"88",X"7F",X"83",X"87",X"88",X"7F",X"83",X"87",X"8B",X"7E",X"82",X"86",
		X"8B",X"7E",X"82",X"86",X"8A",X"7D",X"81",X"85",X"8A",X"7D",X"81",X"85",X"89",X"7C",X"80",X"84",
		X"89",X"9D",X"A2",X"A3",X"A0",X"A1",X"9E",X"9F",X"9C",X"98",X"78",X"78",X"96",X"78",X"DE",X"DF",
		X"78",X"DD",X"79",X"9B",X"79",X"79",X"95",X"79",X"DC",X"7A",X"97",X"7A",X"E0",X"E1",X"7A",X"99",
		X"7A",X"7B",X"E2",X"E3",X"7B",X"9A",X"7B",X"7B",X"94",X"A7",X"BC",X"C5",X"AC",X"B3",X"C6",X"BF",
		X"A4",X"C7",X"B0",X"AF",X"C8",X"C1",X"A6",X"A9",X"BE",X"AD",X"CA",X"C3",X"A8",X"AB",X"C0",X"C9",
		X"B2",X"BD",X"AA",X"A5",X"C2",X"CB",X"AE",X"B1",X"C4",X"80",X"EC",X"F5",X"80",X"BB",X"BB",X"80",
		X"E4",X"F7",X"81",X"B7",X"81",X"B7",X"E6",X"81",X"EE",X"B5",X"82",X"82",X"E8",X"B5",X"F0",X"F9",
		X"82",X"83",X"EA",X"83",X"F2",X"FB",X"B9",X"B9",X"83",X"E7",X"84",X"84",X"B4",X"B4",X"F6",X"EF",
		X"84",X"85",X"B8",X"85",X"F8",X"F1",X"B8",X"E9",X"85",X"86",X"FA",X"F3",X"86",X"EB",X"BA",X"86",
		X"BA",X"ED",X"87",X"E5",X"87",X"B6",X"B6",X"87",X"F4",X"D3",X"D2",X"88",X"76",X"D7",X"D6",X"76",
		X"88",X"89",X"76",X"D9",X"D8",X"76",X"89",X"CD",X"CC",X"DB",X"DA",X"76",X"8A",X"CF",X"CE",X"8A",
		X"76",X"76",X"8B",X"D1",X"D0",X"8B",X"76",X"D5",X"D4",X"76",X"8C",X"8C",X"76",X"8C",X"76",X"76",
		X"8C",X"76",X"8D",X"76",X"8D",X"8D",X"76",X"8D",X"76",X"8E",X"76",X"8E",X"76",X"76",X"8E",X"76",
		X"8E",X"8F",X"76",X"76",X"8F",X"76",X"8F",X"8F",X"76",X"FC",X"90",X"90",X"FC",X"90",X"FC",X"FC",
		X"90",X"FD",X"91",X"FD",X"91",X"91",X"FD",X"91",X"FD",X"92",X"FE",X"92",X"FE",X"FE",X"92",X"FE",
		X"92",X"93",X"FF",X"FF",X"93",X"FF",X"93",X"93",X"FF",X"80",X"81",X"82",X"83",X"84",X"85",X"86",
		X"87",X"7C",X"7D",X"7E",X"7F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",
		X"93",X"88",X"89",X"8A",X"8B",X"88",X"89",X"8A",X"8B",X"76",X"76",X"76",X"76",X"76",X"76",X"76",
		X"76",X"7C",X"7D",X"7E",X"7F",X"88",X"89",X"8A",X"8B",X"88",X"89",X"8A",X"8B",X"88",X"89",X"8A",
		X"8B",X"76",X"76",X"DD",X"CB",X"10",X"9E",X"DD",X"7E",X"10",X"E6",X"06",X"28",X"29",X"FE",X"02",
		X"28",X"19",X"FE",X"04",X"28",X"0C",X"DD",X"56",X"01",X"15",X"DD",X"7E",X"03",X"D6",X"08",X"5F",
		X"18",X"1C",X"DD",X"56",X"01",X"15",X"DD",X"5E",X"03",X"18",X"13",X"DD",X"7E",X"01",X"D6",X"08",
		X"57",X"DD",X"5E",X"03",X"1D",X"18",X"07",X"DD",X"56",X"01",X"DD",X"5E",X"03",X"1D",X"CD",X"89",
		X"1D",X"DD",X"7E",X"09",X"CD",X"5C",X"1D",X"23",X"DD",X"7E",X"0A",X"CD",X"5C",X"1D",X"11",X"1F",
		X"00",X"19",X"DD",X"7E",X"0B",X"CD",X"5C",X"1D",X"23",X"DD",X"7E",X"0C",X"FE",X"76",X"D8",X"FE",
		X"94",X"D0",X"47",X"7E",X"FE",X"94",X"D8",X"70",X"C9",X"DD",X"7E",X"07",X"47",X"E6",X"03",X"DD",
		X"77",X"07",X"78",X"E6",X"18",X"FE",X"18",X"C0",X"DD",X"7E",X"00",X"E6",X"03",X"28",X"B8",X"FE",
		X"01",X"28",X"A8",X"FE",X"02",X"28",X"9B",X"18",X"8D",X"7A",X"E6",X"F8",X"6F",X"26",X"00",X"29",
		X"29",X"7B",X"E6",X"F8",X"0F",X"0F",X"0F",X"B5",X"6F",X"11",X"00",X"88",X"19",X"EB",X"21",X"00",
		X"04",X"19",X"C9",X"DD",X"7E",X"01",X"D6",X"20",X"E6",X"F0",X"6F",X"DD",X"7E",X"03",X"D6",X"18",
		X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"B5",X"6F",X"26",X"00",X"29",X"11",X"12",X"E4",X"19",X"C9",
		X"7A",X"D6",X"20",X"E6",X"F0",X"6F",X"7B",X"18",X"E5",X"21",X"01",X"E0",X"CB",X"C6",X"CD",X"A3",
		X"1D",X"CD",X"1E",X"1F",X"7E",X"E6",X"0D",X"C0",X"44",X"4D",X"DD",X"56",X"01",X"DD",X"7E",X"03",
		X"C6",X"03",X"5F",X"CD",X"89",X"1D",X"EB",X"60",X"69",X"1A",X"FE",X"88",X"28",X"0D",X"FE",X"76",
		X"28",X"09",X"FE",X"8B",X"20",X"08",X"CD",X"15",X"1F",X"18",X"03",X"CD",X"27",X"1F",X"EB",X"01",
		X"E0",X"FF",X"09",X"EB",X"47",X"1A",X"FE",X"88",X"28",X"11",X"FE",X"89",X"28",X"09",X"FE",X"76",
		X"C0",X"B8",X"20",X"07",X"CD",X"33",X"1F",X"CD",X"15",X"1F",X"C9",X"CD",X"33",X"1F",X"C9",X"21",
		X"01",X"E0",X"CB",X"C6",X"CD",X"A3",X"1D",X"CD",X"15",X"1F",X"7E",X"E6",X"07",X"C0",X"44",X"4D",
		X"DD",X"56",X"01",X"DD",X"7E",X"03",X"D6",X"04",X"5F",X"CD",X"89",X"1D",X"EB",X"60",X"69",X"1A",
		X"FE",X"8A",X"28",X"0D",X"FE",X"76",X"28",X"09",X"FE",X"8B",X"20",X"08",X"CD",X"1E",X"1F",X"18",
		X"03",X"CD",X"27",X"1F",X"EB",X"01",X"E0",X"FF",X"09",X"EB",X"47",X"1A",X"FE",X"8A",X"28",X"11",
		X"FE",X"89",X"28",X"09",X"FE",X"76",X"C0",X"B8",X"20",X"07",X"CD",X"33",X"1F",X"CD",X"1E",X"1F",
		X"C9",X"CD",X"33",X"1F",X"C9",X"21",X"01",X"E0",X"CB",X"C6",X"CD",X"A3",X"1D",X"CD",X"33",X"1F",
		X"7E",X"E6",X"0E",X"C0",X"44",X"4D",X"DD",X"7E",X"01",X"C6",X"03",X"57",X"DD",X"5E",X"03",X"CD",
		X"89",X"1D",X"EB",X"60",X"69",X"1A",X"FE",X"8B",X"28",X"10",X"FE",X"88",X"28",X"07",X"FE",X"76",
		X"20",X"0B",X"CD",X"15",X"1F",X"CD",X"27",X"1F",X"18",X"03",X"CD",X"15",X"1F",X"1B",X"1A",X"FE",
		X"8B",X"28",X"0E",X"FE",X"8A",X"28",X"06",X"FE",X"76",X"C0",X"CD",X"1E",X"1F",X"CD",X"27",X"1F",
		X"C9",X"CD",X"1E",X"1F",X"C9",X"21",X"01",X"E0",X"CB",X"C6",X"CD",X"A3",X"1D",X"CD",X"27",X"1F",
		X"7E",X"E6",X"0B",X"C0",X"44",X"4D",X"DD",X"7E",X"01",X"D6",X"04",X"57",X"DD",X"5E",X"03",X"CD",
		X"89",X"1D",X"EB",X"60",X"69",X"1A",X"FE",X"89",X"28",X"10",X"FE",X"88",X"28",X"07",X"FE",X"76",
		X"20",X"0B",X"CD",X"15",X"1F",X"CD",X"33",X"1F",X"18",X"03",X"CD",X"15",X"1F",X"1B",X"1A",X"FE",
		X"89",X"28",X"0E",X"FE",X"8A",X"28",X"06",X"FE",X"76",X"C0",X"CD",X"1E",X"1F",X"CD",X"33",X"1F",
		X"C9",X"CD",X"1E",X"1F",X"C9",X"23",X"23",X"CB",X"CE",X"2B",X"2B",X"CB",X"DE",X"C9",X"2B",X"2B",
		X"CB",X"DE",X"23",X"23",X"CB",X"CE",X"C9",X"01",X"20",X"00",X"09",X"CB",X"C6",X"A7",X"ED",X"42",
		X"CB",X"D6",X"C9",X"01",X"E0",X"FF",X"09",X"CB",X"D6",X"A7",X"ED",X"42",X"CB",X"C6",X"C9",X"D9",
		X"21",X"80",X"E0",X"7E",X"A7",X"C8",X"47",X"23",X"FD",X"E5",X"11",X"31",X"00",X"FD",X"19",X"3E",
		X"0C",X"96",X"4F",X"87",X"87",X"87",X"91",X"5F",X"16",X"00",X"FD",X"E5",X"FD",X"19",X"D9",X"FD",
		X"70",X"00",X"FD",X"66",X"01",X"FD",X"6E",X"02",X"19",X"FD",X"74",X"01",X"FD",X"75",X"02",X"D9",
		X"FD",X"E1",X"23",X"10",X"DA",X"FD",X"E1",X"C9",X"FD",X"E5",X"11",X"31",X"00",X"FD",X"19",X"11",
		X"07",X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",X"80",X"20",X"20",X"FD",X"7E",X"01",X"DD",X"96",
		X"01",X"FE",X"09",X"38",X"04",X"FE",X"F8",X"38",X"12",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"FE",
		X"14",X"30",X"08",X"FE",X"10",X"38",X"04",X"FD",X"36",X"00",X"88",X"FD",X"19",X"10",X"D5",X"FD",
		X"E1",X"C9",X"DD",X"CB",X"00",X"76",X"20",X"51",X"FD",X"35",X"00",X"DD",X"36",X"00",X"E0",X"DD",
		X"36",X"02",X"00",X"DD",X"36",X"03",X"20",X"DD",X"36",X"04",X"00",X"DD",X"36",X"06",X"00",X"DD",
		X"36",X"07",X"80",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"10",X"00",X"DD",
		X"36",X"11",X"00",X"FD",X"36",X"0C",X"00",X"FD",X"36",X"10",X"00",X"21",X"01",X"E0",X"CB",X"C6",
		X"3E",X"19",X"06",X"00",X"CD",X"D9",X"02",X"3E",X"0F",X"06",X"00",X"CD",X"D9",X"02",X"DD",X"36",
		X"01",X"78",X"DD",X"36",X"05",X"3C",X"CD",X"EB",X"22",X"DD",X"CB",X"00",X"6E",X"28",X"10",X"DD",
		X"34",X"06",X"DD",X"7E",X"06",X"E6",X"0F",X"20",X"06",X"CD",X"09",X"23",X"CD",X"EB",X"22",X"DD",
		X"7E",X"05",X"A7",X"28",X"04",X"DD",X"35",X"05",X"C0",X"3A",X"00",X"E0",X"87",X"30",X"13",X"3A",
		X"02",X"A0",X"E6",X"04",X"20",X"0C",X"CD",X"6D",X"24",X"21",X"B6",X"E1",X"CB",X"FE",X"FD",X"36",
		X"30",X"00",X"CD",X"45",X"23",X"3A",X"00",X"E0",X"E6",X"40",X"20",X"08",X"DD",X"36",X"00",X"00",
		X"CD",X"6D",X"24",X"C9",X"3A",X"B6",X"E1",X"A7",X"C2",X"1A",X"22",X"CD",X"02",X"03",X"DD",X"CB",
		X"00",X"5E",X"C2",X"A5",X"22",X"DD",X"CB",X"00",X"66",X"C2",X"74",X"22",X"CD",X"5A",X"23",X"DD",
		X"CB",X"07",X"76",X"C2",X"8C",X"21",X"CD",X"32",X"23",X"2F",X"E6",X"0F",X"CA",X"6F",X"21",X"DD",
		X"34",X"08",X"1F",X"38",X"46",X"1F",X"38",X"2D",X"1F",X"38",X"16",X"DD",X"7E",X"01",X"D6",X"08",
		X"E6",X"0F",X"28",X"04",X"FE",X"0F",X"20",X"47",X"CD",X"63",X"23",X"D2",X"37",X"21",X"C3",X"3A",
		X"21",X"DD",X"7E",X"03",X"E6",X"0F",X"28",X"04",X"FE",X"0F",X"20",X"5F",X"CD",X"9A",X"23",X"D2",
		X"46",X"21",X"C3",X"49",X"21",X"DD",X"7E",X"01",X"D6",X"08",X"E6",X"0F",X"28",X"04",X"FE",X"0F",
		X"20",X"1D",X"CD",X"7F",X"23",X"D2",X"53",X"21",X"C3",X"56",X"21",X"DD",X"7E",X"03",X"E6",X"0F",
		X"28",X"04",X"FE",X"0F",X"20",X"35",X"CD",X"A5",X"23",X"D2",X"62",X"21",X"C3",X"65",X"21",X"47",
		X"DD",X"7E",X"00",X"E6",X"06",X"28",X"07",X"78",X"FE",X"0D",X"38",X"13",X"18",X"05",X"78",X"FE",
		X"04",X"38",X"0C",X"CD",X"9A",X"23",X"30",X"4E",X"CD",X"A5",X"23",X"30",X"65",X"18",X"66",X"CD",
		X"A5",X"23",X"30",X"5E",X"CD",X"9A",X"23",X"30",X"3D",X"18",X"3E",X"47",X"DD",X"7E",X"00",X"E6",
		X"06",X"FE",X"04",X"28",X"07",X"78",X"FE",X"0D",X"38",X"13",X"18",X"05",X"78",X"FE",X"04",X"38",
		X"0C",X"CD",X"63",X"23",X"30",X"11",X"CD",X"7F",X"23",X"30",X"28",X"18",X"29",X"CD",X"7F",X"23",
		X"30",X"21",X"CD",X"63",X"23",X"38",X"03",X"CD",X"95",X"24",X"DD",X"7E",X"00",X"E6",X"F9",X"F6",
		X"04",X"DD",X"77",X"00",X"18",X"29",X"CD",X"46",X"26",X"DD",X"7E",X"00",X"E6",X"F8",X"DD",X"77",
		X"00",X"18",X"1C",X"CD",X"6F",X"25",X"DD",X"7E",X"00",X"E6",X"F9",X"F6",X"06",X"DD",X"77",X"00",
		X"18",X"0D",X"CD",X"2C",X"27",X"DD",X"7E",X"00",X"E6",X"F8",X"F6",X"03",X"DD",X"77",X"00",X"DD",
		X"7E",X"07",X"E6",X"C0",X"FE",X"80",X"C2",X"1A",X"22",X"CD",X"32",X"23",X"E6",X"10",X"C2",X"1A",
		X"22",X"DD",X"CB",X"07",X"F6",X"DD",X"36",X"08",X"00",X"C3",X"1A",X"22",X"DD",X"34",X"08",X"DD",
		X"7E",X"08",X"FE",X"08",X"30",X"12",X"E6",X"04",X"0F",X"0F",X"C6",X"1E",X"DD",X"CB",X"00",X"56",
		X"28",X"02",X"C6",X"02",X"47",X"C3",X"52",X"22",X"DD",X"7E",X"07",X"E6",X"3C",X"DD",X"77",X"07",
		X"DD",X"36",X"08",X"00",X"FD",X"34",X"0C",X"21",X"D7",X"E1",X"06",X"09",X"DD",X"56",X"01",X"DD",
		X"5E",X"03",X"DD",X"7E",X"00",X"E6",X"07",X"FE",X"07",X"30",X"33",X"FE",X"06",X"30",X"28",X"FE",
		X"05",X"30",X"1D",X"FE",X"04",X"30",X"12",X"FE",X"02",X"30",X"07",X"7A",X"80",X"57",X"3E",X"81",
		X"18",X"21",X"7A",X"90",X"57",X"3E",X"83",X"18",X"1A",X"7B",X"80",X"5F",X"3E",X"80",X"18",X"13",
		X"7B",X"80",X"5F",X"3E",X"82",X"18",X"0C",X"7B",X"90",X"5F",X"3E",X"81",X"18",X"05",X"7B",X"90",
		X"5F",X"3E",X"83",X"77",X"23",X"72",X"23",X"36",X"00",X"23",X"73",X"23",X"36",X"00",X"23",X"36",
		X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"3E",X"00",X"DD",X"46",X"07",X"CB",
		X"68",X"20",X"16",X"CB",X"60",X"28",X"02",X"C6",X"0C",X"CB",X"78",X"28",X"02",X"C6",X"06",X"DD",
		X"CB",X"00",X"56",X"28",X"0C",X"C6",X"03",X"18",X"08",X"C6",X"18",X"CB",X"78",X"28",X"02",X"C6",
		X"03",X"47",X"DD",X"7E",X"08",X"E6",X"18",X"0F",X"0F",X"0F",X"FE",X"03",X"20",X"02",X"3E",X"01",
		X"80",X"47",X"DD",X"7E",X"00",X"E6",X"07",X"FE",X"04",X"30",X"04",X"E6",X"02",X"18",X"0A",X"E6",
		X"03",X"28",X"06",X"FE",X"03",X"28",X"02",X"EE",X"03",X"87",X"87",X"87",X"87",X"F6",X"02",X"4F",
		X"CD",X"97",X"02",X"C9",X"DD",X"CB",X"07",X"4E",X"20",X"24",X"DD",X"CB",X"07",X"CE",X"CD",X"6D",
		X"24",X"DD",X"7E",X"10",X"2F",X"E6",X"18",X"28",X"12",X"DD",X"7E",X"07",X"2F",X"E6",X"18",X"20",
		X"0D",X"DD",X"7E",X"00",X"E6",X"06",X"F6",X"18",X"DD",X"77",X"10",X"CD",X"03",X"1D",X"01",X"02",
		X"22",X"CD",X"97",X"02",X"C9",X"DD",X"CB",X"07",X"46",X"20",X"0F",X"DD",X"CB",X"07",X"C6",X"DD",
		X"36",X"08",X"FF",X"3E",X"24",X"06",X"00",X"CD",X"D9",X"02",X"DD",X"34",X"08",X"DD",X"7E",X"08",
		X"D6",X"1E",X"38",X"B0",X"FE",X"80",X"30",X"16",X"01",X"02",X"23",X"FE",X"10",X"38",X"0B",X"04",
		X"FE",X"20",X"38",X"06",X"04",X"FE",X"40",X"38",X"01",X"04",X"CD",X"97",X"02",X"C9",X"21",X"A9",
		X"E1",X"CB",X"FE",X"DD",X"36",X"00",X"00",X"CD",X"80",X"5A",X"C9",X"DD",X"7E",X"06",X"E6",X"F0",
		X"FE",X"60",X"30",X"10",X"0F",X"0F",X"0F",X"0F",X"F5",X"CD",X"20",X"23",X"CD",X"6C",X"04",X"F1",
		X"FD",X"BE",X"00",X"D8",X"DD",X"CB",X"00",X"AE",X"C9",X"DD",X"7E",X"06",X"E6",X"F0",X"0F",X"0F",
		X"0F",X"0F",X"3D",X"CD",X"20",X"23",X"3E",X"09",X"08",X"3E",X"2E",X"08",X"CD",X"42",X"04",X"C9",
		X"11",X"81",X"88",X"01",X"02",X"02",X"A7",X"C8",X"EB",X"11",X"40",X"00",X"19",X"3D",X"20",X"FC",
		X"EB",X"C9",X"3A",X"A5",X"E1",X"21",X"00",X"E0",X"CB",X"7E",X"C8",X"3A",X"00",X"A0",X"CB",X"46",
		X"C8",X"3A",X"01",X"A0",X"C9",X"DD",X"7E",X"0D",X"A7",X"C8",X"DD",X"35",X"0D",X"DD",X"56",X"0E",
		X"DD",X"5E",X"0F",X"01",X"0A",X"71",X"CD",X"9D",X"02",X"C9",X"FD",X"7E",X"10",X"A7",X"C8",X"FD",
		X"35",X"10",X"C9",X"DD",X"7E",X"03",X"FE",X"DF",X"3F",X"D8",X"DD",X"56",X"01",X"DD",X"7E",X"03",
		X"C6",X"07",X"5F",X"01",X"07",X"0B",X"CD",X"76",X"40",X"D8",X"CD",X"6D",X"24",X"A7",X"C9",X"DD",
		X"7E",X"03",X"FE",X"21",X"D8",X"DD",X"56",X"01",X"DD",X"7E",X"03",X"D6",X"07",X"5F",X"01",X"07",
		X"0B",X"CD",X"76",X"40",X"D8",X"CD",X"6D",X"24",X"A7",X"C9",X"DD",X"7E",X"01",X"FE",X"D7",X"3F",
		X"D8",X"0E",X"00",X"18",X"08",X"DD",X"7E",X"01",X"FE",X"29",X"D8",X"0E",X"03",X"DD",X"56",X"01",
		X"DD",X"5E",X"03",X"21",X"80",X"E0",X"36",X"00",X"23",X"D9",X"FD",X"E5",X"11",X"31",X"00",X"FD",
		X"19",X"11",X"07",X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",X"80",X"38",X"6D",X"FE",X"D0",X"28",
		X"04",X"FE",X"B8",X"30",X"65",X"D9",X"FD",X"7E",X"03",X"93",X"28",X"04",X"FE",X"01",X"20",X"3F",
		X"CB",X"49",X"20",X"06",X"FD",X"7E",X"01",X"92",X"18",X"04",X"7A",X"FD",X"96",X"01",X"28",X"49",
		X"FE",X"11",X"30",X"45",X"FE",X"0F",X"30",X"64",X"FD",X"7E",X"00",X"FE",X"A0",X"30",X"6A",X"3A",
		X"80",X"E0",X"3C",X"32",X"80",X"E0",X"D9",X"78",X"D9",X"77",X"23",X"FD",X"56",X"01",X"FD",X"5E",
		X"03",X"7A",X"FE",X"D8",X"30",X"53",X"FE",X"29",X"38",X"4F",X"D9",X"FD",X"E1",X"18",X"9B",X"FE",
		X"09",X"38",X"04",X"FE",X"F8",X"38",X"12",X"CB",X"41",X"20",X"06",X"FD",X"7E",X"01",X"92",X"18",
		X"04",X"7A",X"FD",X"96",X"01",X"FE",X"0F",X"38",X"30",X"D9",X"FD",X"19",X"10",X"88",X"3A",X"80",
		X"E0",X"A7",X"28",X"1E",X"D9",X"3E",X"07",X"CB",X"41",X"28",X"02",X"3E",X"F9",X"82",X"57",X"CD",
		X"AD",X"41",X"38",X"15",X"FD",X"E1",X"DD",X"CB",X"07",X"EE",X"A7",X"C9",X"3A",X"80",X"E0",X"A7",
		X"20",X"F2",X"FD",X"E1",X"CD",X"6D",X"24",X"A7",X"C9",X"FD",X"E1",X"37",X"C9",X"DD",X"7E",X"07",
		X"E6",X"20",X"C8",X"DD",X"CB",X"07",X"AE",X"FD",X"E5",X"11",X"31",X"00",X"FD",X"19",X"11",X"07",
		X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",X"98",X"20",X"04",X"FD",X"36",X"00",X"80",X"FD",X"19",
		X"10",X"F1",X"FD",X"E1",X"C9",X"DD",X"7E",X"00",X"E6",X"06",X"FE",X"04",X"28",X"35",X"DD",X"CB",
		X"11",X"BE",X"21",X"01",X"E0",X"CB",X"D6",X"DD",X"7E",X"10",X"47",X"E6",X"06",X"FE",X"04",X"20",
		X"11",X"DD",X"7E",X"07",X"E6",X"A0",X"B0",X"E6",X"B8",X"DD",X"77",X"07",X"DD",X"36",X"10",X"04",
		X"18",X"23",X"47",X"DD",X"7E",X"07",X"4F",X"E6",X"18",X"B0",X"DD",X"77",X"10",X"79",X"E6",X"A0",
		X"DD",X"77",X"07",X"DD",X"7E",X"10",X"2F",X"E6",X"18",X"20",X"0A",X"DD",X"7E",X"03",X"E6",X"07",
		X"FE",X"05",X"D4",X"03",X"1D",X"DD",X"7E",X"03",X"E6",X"0F",X"28",X"04",X"FE",X"0F",X"20",X"23",
		X"DD",X"CB",X"11",X"7E",X"20",X"21",X"DD",X"CB",X"11",X"FE",X"CD",X"A3",X"1D",X"CB",X"5E",X"28",
		X"09",X"CD",X"16",X"28",X"DD",X"36",X"10",X"04",X"18",X"48",X"CD",X"24",X"28",X"DD",X"36",X"10",
		X"14",X"18",X"3F",X"DD",X"CB",X"11",X"BE",X"DD",X"7E",X"07",X"47",X"E6",X"14",X"FE",X"10",X"20",
		X"2D",X"DD",X"7E",X"03",X"E6",X"07",X"CB",X"58",X"20",X"0A",X"FE",X"01",X"28",X"0E",X"FE",X"02",
		X"20",X"20",X"18",X"08",X"FE",X"05",X"28",X"04",X"FE",X"06",X"20",X"16",X"CD",X"9B",X"1A",X"CD",
		X"62",X"28",X"DD",X"7E",X"03",X"E6",X"0F",X"FE",X"0D",X"D4",X"C9",X"1D",X"18",X"04",X"DD",X"CB",
		X"07",X"96",X"CD",X"78",X"1F",X"CD",X"34",X"28",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"19",X"DD",
		X"74",X"03",X"DD",X"75",X"04",X"DD",X"7E",X"01",X"3C",X"E6",X"F8",X"DD",X"77",X"01",X"C9",X"DD",
		X"7E",X"00",X"E6",X"06",X"FE",X"06",X"28",X"35",X"DD",X"CB",X"11",X"BE",X"21",X"01",X"E0",X"CB",
		X"D6",X"DD",X"7E",X"10",X"47",X"E6",X"06",X"FE",X"06",X"20",X"11",X"DD",X"7E",X"07",X"E6",X"A0",
		X"B0",X"E6",X"B8",X"DD",X"77",X"07",X"DD",X"36",X"10",X"06",X"18",X"23",X"47",X"DD",X"7E",X"07",
		X"4F",X"E6",X"18",X"B0",X"DD",X"77",X"10",X"79",X"E6",X"A0",X"DD",X"77",X"07",X"DD",X"7E",X"10",
		X"2F",X"E6",X"18",X"20",X"0A",X"DD",X"7E",X"03",X"E6",X"07",X"FE",X"03",X"DC",X"03",X"1D",X"DD",
		X"7E",X"03",X"E6",X"0F",X"28",X"04",X"FE",X"0F",X"20",X"23",X"DD",X"CB",X"11",X"7E",X"20",X"21",
		X"DD",X"CB",X"11",X"FE",X"CD",X"A3",X"1D",X"CB",X"4E",X"28",X"09",X"CD",X"16",X"28",X"DD",X"36",
		X"10",X"06",X"18",X"48",X"CD",X"24",X"28",X"DD",X"36",X"10",X"16",X"18",X"3F",X"DD",X"CB",X"11",
		X"BE",X"DD",X"7E",X"07",X"47",X"E6",X"14",X"FE",X"10",X"20",X"2D",X"DD",X"7E",X"03",X"E6",X"07",
		X"CB",X"58",X"20",X"0A",X"FE",X"05",X"28",X"0E",X"FE",X"06",X"20",X"20",X"18",X"08",X"FE",X"01",
		X"28",X"04",X"FE",X"02",X"20",X"16",X"CD",X"D0",X"1A",X"CD",X"62",X"28",X"DD",X"7E",X"03",X"E6",
		X"0F",X"FE",X"03",X"DC",X"1F",X"1E",X"18",X"04",X"DD",X"CB",X"07",X"96",X"CD",X"4B",X"28",X"DD",
		X"66",X"03",X"DD",X"6E",X"04",X"19",X"DD",X"74",X"03",X"DD",X"75",X"04",X"DD",X"7E",X"01",X"3C",
		X"E6",X"F8",X"DD",X"77",X"01",X"C9",X"DD",X"7E",X"00",X"E6",X"06",X"28",X"33",X"DD",X"CB",X"11",
		X"BE",X"21",X"01",X"E0",X"CB",X"D6",X"DD",X"7E",X"10",X"47",X"E6",X"06",X"20",X"11",X"DD",X"7E",
		X"07",X"E6",X"A0",X"B0",X"E6",X"B8",X"DD",X"77",X"07",X"DD",X"36",X"10",X"00",X"18",X"23",X"47",
		X"DD",X"7E",X"07",X"4F",X"E6",X"18",X"B0",X"DD",X"77",X"10",X"79",X"E6",X"A0",X"DD",X"77",X"07",
		X"DD",X"7E",X"10",X"2F",X"E6",X"18",X"20",X"0A",X"DD",X"7E",X"01",X"E6",X"07",X"FE",X"05",X"D4",
		X"03",X"1D",X"DD",X"7E",X"01",X"E6",X"0F",X"FE",X"07",X"28",X"04",X"FE",X"08",X"20",X"23",X"DD",
		X"CB",X"11",X"7E",X"20",X"21",X"DD",X"CB",X"11",X"FE",X"CD",X"A3",X"1D",X"CB",X"56",X"28",X"09",
		X"CD",X"16",X"28",X"DD",X"36",X"10",X"00",X"18",X"4C",X"CD",X"24",X"28",X"DD",X"36",X"10",X"10",
		X"18",X"43",X"DD",X"CB",X"11",X"BE",X"DD",X"7E",X"07",X"47",X"E6",X"14",X"FE",X"10",X"20",X"31",
		X"DD",X"7E",X"01",X"E6",X"07",X"CB",X"58",X"20",X"0A",X"FE",X"01",X"28",X"0E",X"FE",X"02",X"20",
		X"24",X"18",X"08",X"FE",X"05",X"28",X"04",X"FE",X"06",X"20",X"1A",X"CD",X"05",X"1B",X"CD",X"62",
		X"28",X"DD",X"7E",X"01",X"E6",X"0F",X"FE",X"07",X"30",X"0B",X"FE",X"05",X"D4",X"75",X"1E",X"18",
		X"04",X"DD",X"CB",X"07",X"96",X"CD",X"78",X"1F",X"CD",X"34",X"28",X"DD",X"66",X"01",X"DD",X"6E",
		X"02",X"19",X"DD",X"74",X"01",X"DD",X"75",X"02",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"DD",X"77",
		X"03",X"DD",X"CB",X"07",X"6E",X"C8",X"06",X"98",X"CD",X"3F",X"1F",X"C9",X"DD",X"7E",X"00",X"E6",
		X"06",X"FE",X"02",X"28",X"35",X"DD",X"CB",X"11",X"BE",X"21",X"01",X"E0",X"CB",X"D6",X"DD",X"7E",
		X"10",X"47",X"E6",X"06",X"FE",X"02",X"20",X"11",X"DD",X"7E",X"07",X"E6",X"A0",X"B0",X"E6",X"B8",
		X"DD",X"77",X"07",X"DD",X"36",X"10",X"02",X"18",X"23",X"47",X"DD",X"7E",X"07",X"4F",X"E6",X"18",
		X"B0",X"DD",X"77",X"10",X"79",X"E6",X"A0",X"DD",X"77",X"07",X"DD",X"7E",X"10",X"2F",X"E6",X"18",
		X"20",X"0A",X"DD",X"7E",X"01",X"E6",X"07",X"FE",X"03",X"DC",X"03",X"1D",X"DD",X"7E",X"01",X"E6",
		X"0F",X"FE",X"07",X"28",X"04",X"FE",X"08",X"20",X"23",X"DD",X"CB",X"11",X"7E",X"20",X"21",X"DD",
		X"CB",X"11",X"FE",X"CD",X"A3",X"1D",X"CB",X"46",X"28",X"09",X"CD",X"16",X"28",X"DD",X"36",X"10",
		X"02",X"18",X"4C",X"CD",X"24",X"28",X"DD",X"36",X"10",X"12",X"18",X"43",X"DD",X"CB",X"11",X"BE",
		X"DD",X"7E",X"07",X"47",X"E6",X"14",X"FE",X"10",X"20",X"31",X"DD",X"7E",X"01",X"E6",X"07",X"CB",
		X"58",X"20",X"0A",X"FE",X"05",X"28",X"0E",X"FE",X"06",X"20",X"24",X"18",X"08",X"FE",X"01",X"28",
		X"04",X"FE",X"02",X"20",X"1A",X"CD",X"3B",X"1B",X"CD",X"62",X"28",X"DD",X"7E",X"01",X"E6",X"0F",
		X"FE",X"09",X"38",X"0B",X"FE",X"0B",X"DC",X"C5",X"1E",X"18",X"04",X"DD",X"CB",X"07",X"96",X"CD",
		X"78",X"1F",X"CD",X"4B",X"28",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"19",X"DD",X"74",X"01",X"DD",
		X"75",X"02",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"DD",X"77",X"03",X"DD",X"CB",X"07",X"6E",X"C8",
		X"06",X"98",X"CD",X"3F",X"1F",X"C9",X"21",X"01",X"E0",X"CB",X"C6",X"DD",X"7E",X"07",X"E6",X"E0",
		X"DD",X"77",X"07",X"C9",X"21",X"01",X"E0",X"CB",X"C6",X"DD",X"7E",X"07",X"E6",X"E0",X"F6",X"10",
		X"DD",X"77",X"07",X"C9",X"DD",X"7E",X"07",X"CB",X"6F",X"20",X"0C",X"E6",X"10",X"20",X"04",X"11",
		X"D5",X"00",X"C9",X"11",X"AB",X"00",X"C9",X"11",X"80",X"00",X"C9",X"DD",X"7E",X"07",X"CB",X"6F",
		X"20",X"0C",X"E6",X"10",X"20",X"04",X"11",X"2B",X"FF",X"C9",X"11",X"55",X"FF",X"C9",X"11",X"80",
		X"FF",X"C9",X"21",X"CE",X"E1",X"06",X"04",X"7E",X"FE",X"DC",X"38",X"17",X"FD",X"35",X"0B",X"FD",
		X"7E",X"0B",X"E6",X"03",X"20",X"0D",X"C5",X"E5",X"CD",X"94",X"28",X"E1",X"C1",X"FD",X"7E",X"0B",
		X"A7",X"28",X"04",X"23",X"10",X"E1",X"C9",X"21",X"B6",X"E1",X"CB",X"FE",X"FD",X"36",X"30",X"02",
		X"FD",X"34",X"09",X"C9",X"FD",X"7E",X"10",X"A7",X"20",X"10",X"FD",X"36",X"11",X"00",X"FD",X"36",
		X"10",X"1E",X"11",X"DB",X"28",X"CD",X"2A",X"03",X"18",X"24",X"FD",X"34",X"11",X"FD",X"7E",X"11",
		X"FE",X"08",X"30",X"E6",X"FE",X"07",X"38",X"E6",X"11",X"DE",X"28",X"CD",X"2A",X"03",X"DD",X"36",
		X"0D",X"1E",X"DD",X"7E",X"01",X"DD",X"77",X"0E",X"DD",X"7E",X"03",X"DD",X"77",X"0F",X"FD",X"7E",
		X"11",X"C6",X"01",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"00",X"00",X"50",X"00",X"05",X"00",X"DD",
		X"46",X"00",X"CB",X"58",X"C2",X"C4",X"2A",X"3A",X"00",X"E0",X"E6",X"40",X"20",X"05",X"DD",X"36",
		X"00",X"00",X"C9",X"3A",X"B6",X"E1",X"A7",X"C2",X"B2",X"2A",X"3A",X"C5",X"E1",X"E6",X"98",X"FE",
		X"80",X"C2",X"B2",X"2A",X"DD",X"34",X"08",X"FD",X"E5",X"FD",X"21",X"C5",X"E1",X"01",X"09",X"09",
		X"CD",X"D7",X"05",X"30",X"0B",X"FD",X"CB",X"07",X"FE",X"FD",X"E1",X"DD",X"36",X"00",X"00",X"C9",
		X"FD",X"21",X"1A",X"E2",X"11",X"15",X"00",X"06",X"08",X"FD",X"7E",X"00",X"E6",X"98",X"FE",X"80",
		X"20",X"15",X"C5",X"01",X"0A",X"0A",X"CD",X"D7",X"05",X"C1",X"30",X"0B",X"FD",X"CB",X"00",X"DE",
		X"DD",X"CB",X"00",X"DE",X"FD",X"E1",X"C9",X"FD",X"19",X"10",X"DE",X"FD",X"21",X"D3",X"E2",X"11",
		X"0F",X"00",X"06",X"03",X"FD",X"7E",X"00",X"E6",X"BC",X"FE",X"80",X"20",X"19",X"C5",X"01",X"0A",
		X"0A",X"CD",X"D7",X"05",X"C1",X"30",X"0F",X"FD",X"CB",X"00",X"DE",X"DD",X"CB",X"00",X"DE",X"FD",
		X"E1",X"FD",X"36",X"0C",X"01",X"C9",X"FD",X"19",X"10",X"DA",X"FD",X"21",X"C2",X"E2",X"FD",X"7E",
		X"00",X"E6",X"B8",X"FE",X"A0",X"20",X"17",X"01",X"0A",X"0A",X"CD",X"D7",X"05",X"30",X"0F",X"FD",
		X"CB",X"00",X"DE",X"DD",X"CB",X"00",X"DE",X"FD",X"E1",X"FD",X"36",X"0C",X"01",X"C9",X"FD",X"E1",
		X"11",X"31",X"00",X"FD",X"19",X"11",X"07",X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",X"80",X"38",
		X"12",X"FE",X"D0",X"28",X"04",X"FE",X"C8",X"30",X"0A",X"C5",X"01",X"08",X"08",X"CD",X"D7",X"05",
		X"38",X"07",X"C1",X"FD",X"19",X"10",X"E3",X"18",X"42",X"D1",X"FD",X"7E",X"00",X"FE",X"B8",X"38",
		X"09",X"FE",X"D0",X"28",X"05",X"DD",X"CB",X"00",X"DE",X"C9",X"DD",X"7E",X"00",X"EE",X"03",X"DD",
		X"77",X"00",X"CD",X"A1",X"2B",X"DD",X"6E",X"03",X"FD",X"56",X"01",X"FD",X"5E",X"03",X"CD",X"EF",
		X"05",X"30",X"04",X"DD",X"CB",X"00",X"E6",X"D5",X"CD",X"B5",X"2B",X"D1",X"6C",X"DD",X"66",X"01",
		X"CD",X"EF",X"05",X"30",X"04",X"DD",X"CB",X"00",X"EE",X"18",X"59",X"DD",X"7E",X"01",X"FE",X"24",
		X"38",X"04",X"FE",X"DB",X"38",X"04",X"DD",X"CB",X"00",X"EE",X"DD",X"7E",X"03",X"FE",X"1C",X"38",
		X"04",X"FE",X"E3",X"38",X"04",X"DD",X"CB",X"00",X"E6",X"DD",X"7E",X"00",X"E6",X"30",X"20",X"4F",
		X"DD",X"56",X"01",X"DD",X"5E",X"03",X"CD",X"C9",X"2B",X"DA",X"A0",X"2A",X"DD",X"7E",X"00",X"EE",
		X"03",X"DD",X"77",X"00",X"CD",X"A1",X"2B",X"EB",X"DD",X"5E",X"03",X"CD",X"C9",X"2B",X"38",X"04",
		X"DD",X"CB",X"00",X"E6",X"CD",X"B5",X"2B",X"DD",X"56",X"01",X"5C",X"CD",X"C9",X"2B",X"38",X"04",
		X"DD",X"CB",X"00",X"EE",X"DD",X"7E",X"00",X"EE",X"03",X"DD",X"77",X"00",X"E6",X"30",X"20",X"0F",
		X"CD",X"F4",X"02",X"E6",X"20",X"20",X"02",X"3E",X"10",X"DD",X"B6",X"00",X"DD",X"77",X"00",X"DD",
		X"34",X"07",X"20",X"05",X"DD",X"CB",X"00",X"DE",X"C9",X"3E",X"16",X"06",X"00",X"CD",X"D9",X"02",
		X"DD",X"7E",X"00",X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"03",X"A8",X"E6",X"83",X"DD",X"77",X"00",
		X"CD",X"A1",X"2B",X"DD",X"74",X"01",X"DD",X"75",X"02",X"CD",X"B5",X"2B",X"DD",X"74",X"03",X"DD",
		X"75",X"04",X"01",X"06",X"66",X"DD",X"7E",X"00",X"E6",X"03",X"87",X"87",X"87",X"87",X"B1",X"4F",
		X"CD",X"97",X"02",X"C9",X"DD",X"7E",X"06",X"E6",X"30",X"20",X"32",X"CD",X"B2",X"2C",X"DD",X"CB",
		X"06",X"E6",X"DD",X"36",X"05",X"01",X"DD",X"CB",X"01",X"3E",X"DD",X"CB",X"02",X"1E",X"DD",X"CB",
		X"01",X"3E",X"DD",X"CB",X"02",X"1E",X"DD",X"CB",X"03",X"3E",X"DD",X"CB",X"04",X"1E",X"DD",X"CB",
		X"03",X"3E",X"DD",X"CB",X"04",X"1E",X"3E",X"1B",X"06",X"00",X"CD",X"D9",X"02",X"DD",X"34",X"07",
		X"DD",X"35",X"05",X"C2",X"72",X"2B",X"DD",X"7E",X"06",X"E6",X"30",X"FE",X"20",X"CA",X"58",X"2B",
		X"DD",X"7E",X"06",X"E6",X"0F",X"FE",X"0A",X"D2",X"1F",X"2B",X"CD",X"5B",X"2C",X"18",X"53",X"DD",
		X"7E",X"06",X"C6",X"10",X"E6",X"30",X"DD",X"77",X"06",X"28",X"23",X"3A",X"01",X"E0",X"E6",X"40",
		X"28",X"04",X"3E",X"01",X"18",X"09",X"FD",X"7E",X"0C",X"FE",X"05",X"38",X"02",X"3E",X"04",X"5F",
		X"16",X"00",X"21",X"91",X"2E",X"19",X"7E",X"DD",X"77",X"05",X"CD",X"C8",X"2C",X"C9",X"DD",X"36",
		X"00",X"00",X"21",X"CC",X"E1",X"CB",X"FE",X"C9",X"CD",X"B2",X"2C",X"DD",X"36",X"06",X"30",X"DD",
		X"36",X"05",X"01",X"CD",X"38",X"2C",X"CD",X"C8",X"2C",X"C0",X"3E",X"1C",X"06",X"00",X"CD",X"D9",
		X"02",X"C9",X"DD",X"7E",X"06",X"E6",X"30",X"FE",X"30",X"CC",X"38",X"2C",X"06",X"05",X"11",X"0A",
		X"00",X"FD",X"21",X"E0",X"E1",X"DD",X"CB",X"07",X"46",X"28",X"04",X"FD",X"21",X"E5",X"E1",X"FD",
		X"CB",X"00",X"7E",X"28",X"07",X"C5",X"D5",X"CD",X"EB",X"2C",X"D1",X"C1",X"FD",X"19",X"10",X"EF",
		X"C9",X"DD",X"56",X"01",X"DD",X"5E",X"02",X"21",X"1F",X"02",X"DD",X"CB",X"00",X"4E",X"28",X"03",
		X"21",X"E1",X"FD",X"19",X"C9",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"21",X"1F",X"02",X"DD",X"CB",
		X"00",X"46",X"28",X"03",X"21",X"E1",X"FD",X"19",X"C9",X"D5",X"CD",X"89",X"1D",X"D1",X"7E",X"D6",
		X"72",X"D8",X"1F",X"F5",X"4F",X"06",X"00",X"21",X"F1",X"2B",X"09",X"F1",X"3E",X"10",X"30",X"02",
		X"3E",X"01",X"CB",X"52",X"20",X"02",X"87",X"87",X"CB",X"53",X"20",X"01",X"87",X"A6",X"C0",X"37",
		X"C9",X"00",X"00",X"0F",X"FF",X"FF",X"DE",X"B7",X"DE",X"B7",X"DE",X"B7",X"5C",X"A3",X"12",X"48",
		X"12",X"48",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"CC",X"AA",X"33",X"DB",X"7E",
		X"E7",X"BD",X"DB",X"7E",X"E7",X"BD",X"D7",X"ED",X"BE",X"7B",X"7D",X"DE",X"EB",X"B7",X"48",X"82",
		X"21",X"14",X"33",X"55",X"CC",X"AA",X"FF",X"FF",X"FF",X"FF",X"55",X"CC",X"AA",X"33",X"D7",X"ED",
		X"BE",X"7B",X"7D",X"DE",X"EB",X"B7",X"12",X"48",X"2A",X"C6",X"E1",X"CB",X"3D",X"CB",X"1C",X"CB",
		X"3D",X"CB",X"1C",X"DD",X"75",X"01",X"DD",X"74",X"02",X"2A",X"C8",X"E1",X"CB",X"3D",X"CB",X"1C",
		X"CB",X"3D",X"CB",X"1C",X"DD",X"75",X"03",X"DD",X"74",X"04",X"C9",X"DD",X"7E",X"06",X"E6",X"0F",
		X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"48",X"2E",X"19",X"7E",X"DD",X"77",X"05",X"44",X"4D",
		X"03",X"DD",X"CB",X"06",X"6E",X"28",X"01",X"03",X"0A",X"E6",X"F0",X"0F",X"0F",X"0F",X"21",X"66",
		X"2E",X"CD",X"C0",X"2C",X"D5",X"0A",X"E6",X"0F",X"87",X"21",X"66",X"2E",X"CD",X"C0",X"2C",X"DD",
		X"7E",X"06",X"E6",X"0F",X"47",X"87",X"87",X"80",X"4F",X"06",X"00",X"21",X"E0",X"E1",X"09",X"C1",
		X"DD",X"7E",X"06",X"F6",X"80",X"77",X"23",X"70",X"23",X"71",X"23",X"72",X"23",X"73",X"DD",X"34",
		X"06",X"C9",X"21",X"E0",X"E1",X"11",X"05",X"00",X"06",X"0A",X"36",X"00",X"19",X"10",X"FB",X"C9",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"C9",X"3A",X"00",X"E0",X"E6",X"40",X"28",X"0C",X"3A",
		X"B6",X"E1",X"A7",X"20",X"06",X"3A",X"C5",X"E1",X"E6",X"18",X"C8",X"DD",X"36",X"00",X"00",X"3E",
		X"FF",X"B7",X"C9",X"78",X"2F",X"47",X"79",X"2F",X"4F",X"03",X"C9",X"FD",X"CB",X"00",X"6E",X"20",
		X"48",X"FD",X"7E",X"01",X"FE",X"30",X"30",X"07",X"FD",X"7E",X"03",X"FE",X"36",X"38",X"05",X"FD",
		X"36",X"00",X"00",X"C9",X"CD",X"39",X"2E",X"0A",X"E6",X"F0",X"0F",X"0F",X"0F",X"21",X"80",X"2E",
		X"CD",X"C0",X"2C",X"FD",X"66",X"01",X"FD",X"6E",X"02",X"19",X"FD",X"74",X"01",X"FD",X"75",X"02",
		X"0A",X"E6",X"0F",X"87",X"21",X"80",X"2E",X"CD",X"C0",X"2C",X"FD",X"66",X"03",X"FD",X"6E",X"04",
		X"19",X"FD",X"74",X"03",X"FD",X"75",X"04",X"18",X"43",X"FD",X"CB",X"01",X"7E",X"20",X"C0",X"FD",
		X"CB",X"03",X"7E",X"20",X"BA",X"CD",X"39",X"2E",X"0A",X"E6",X"F0",X"0F",X"0F",X"0F",X"21",X"80",
		X"2E",X"CD",X"C0",X"2C",X"FD",X"66",X"01",X"FD",X"6E",X"02",X"A7",X"ED",X"52",X"FD",X"74",X"01",
		X"FD",X"75",X"02",X"0A",X"E6",X"0F",X"87",X"21",X"80",X"2E",X"CD",X"C0",X"2C",X"FD",X"66",X"03",
		X"FD",X"6E",X"04",X"A7",X"ED",X"52",X"FD",X"74",X"03",X"FD",X"75",X"04",X"01",X"0A",X"70",X"DD",
		X"CB",X"00",X"56",X"28",X"03",X"01",X"0A",X"79",X"C5",X"CD",X"A1",X"2D",X"C1",X"C5",X"CB",X"E1",
		X"CD",X"C0",X"2D",X"C1",X"CB",X"E9",X"C5",X"CD",X"E0",X"2D",X"C1",X"CB",X"E1",X"CD",X"00",X"2E",
		X"C9",X"FD",X"56",X"01",X"FD",X"5E",X"02",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"19",X"E5",X"FD",
		X"56",X"03",X"FD",X"5E",X"04",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"19",X"D1",X"C3",X"20",X"2E",
		X"FD",X"56",X"03",X"FD",X"5E",X"04",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"19",X"E5",X"FD",X"56",
		X"01",X"FD",X"5E",X"02",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"A7",X"ED",X"52",X"D1",X"18",X"40",
		X"FD",X"56",X"03",X"FD",X"5E",X"04",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"A7",X"ED",X"52",X"E5",
		X"FD",X"56",X"01",X"FD",X"5E",X"02",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"19",X"D1",X"18",X"20",
		X"FD",X"56",X"01",X"FD",X"5E",X"02",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"A7",X"ED",X"52",X"E5",
		X"FD",X"56",X"03",X"FD",X"5E",X"04",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"A7",X"ED",X"52",X"D1",
		X"7A",X"FE",X"06",X"D8",X"FE",X"3A",X"D0",X"7C",X"FE",X"01",X"D8",X"FE",X"3E",X"D0",X"EB",X"29",
		X"29",X"EB",X"29",X"29",X"5C",X"CD",X"9D",X"02",X"C9",X"FD",X"7E",X"00",X"E6",X"0F",X"5F",X"16",
		X"00",X"21",X"76",X"2E",X"19",X"44",X"4D",X"C9",X"02",X"00",X"01",X"04",X"00",X"22",X"03",X"00",
		X"34",X"01",X"56",X"43",X"02",X"00",X"01",X"08",X"77",X"22",X"03",X"00",X"34",X"03",X"56",X"43",
		X"04",X"00",X"22",X"1E",X"00",X"01",X"00",X"02",X"00",X"3E",X"6D",X"2C",X"B5",X"39",X"49",X"18",
		X"7B",X"05",X"65",X"03",X"D4",X"04",X"01",X"22",X"34",X"43",X"05",X"66",X"34",X"43",X"77",X"08",
		X"00",X"00",X"00",X"02",X"6A",X"01",X"52",X"02",X"EE",X"00",X"80",X"01",X"10",X"01",X"1F",X"02",
		X"80",X"03",X"01",X"78",X"B4",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"99",X"3A",X"00",X"E0",X"E6",X"40",X"20",X"05",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"CB",X"00",
		X"76",X"20",X"4A",X"11",X"CF",X"81",X"01",X"02",X"02",X"CD",X"6C",X"04",X"DD",X"CB",X"00",X"F6",
		X"DD",X"36",X"02",X"00",X"FD",X"7E",X"0A",X"DD",X"77",X"03",X"DD",X"36",X"04",X"00",X"DD",X"36",
		X"05",X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"FF",X"FD",X"36",X"12",X"00",X"FD",X"36",
		X"13",X"3C",X"CD",X"76",X"1A",X"FE",X"14",X"38",X"02",X"3E",X"13",X"5F",X"16",X"00",X"21",X"F9",
		X"31",X"19",X"7E",X"FD",X"77",X"0E",X"FD",X"36",X"0F",X"3C",X"C3",X"17",X"30",X"FD",X"7E",X"0E",
		X"A7",X"28",X"0C",X"FD",X"35",X"0F",X"20",X"07",X"FD",X"36",X"0F",X"3C",X"FD",X"35",X"0E",X"FD",
		X"35",X"13",X"20",X"12",X"FD",X"36",X"13",X"3C",X"FD",X"34",X"12",X"FD",X"7E",X"12",X"FE",X"40",
		X"38",X"04",X"FD",X"36",X"12",X"30",X"3A",X"B6",X"E1",X"A7",X"20",X"4E",X"3A",X"01",X"E0",X"E6",
		X"60",X"20",X"47",X"3A",X"00",X"E0",X"E6",X"08",X"20",X"40",X"3A",X"C5",X"E1",X"E6",X"98",X"FE",
		X"80",X"20",X"37",X"DD",X"7E",X"07",X"DD",X"36",X"07",X"FF",X"DD",X"CB",X"06",X"46",X"20",X"16",
		X"FE",X"51",X"30",X"26",X"DD",X"36",X"06",X"01",X"3E",X"0F",X"CD",X"EA",X"02",X"3E",X"10",X"06",
		X"00",X"CD",X"D9",X"02",X"18",X"14",X"FE",X"71",X"38",X"10",X"DD",X"36",X"06",X"00",X"3E",X"10",
		X"CD",X"EA",X"02",X"3E",X"0F",X"06",X"00",X"CD",X"D9",X"02",X"DD",X"CB",X"00",X"6E",X"C2",X"75",
		X"30",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"78",X"B1",X"28",X"09",X"0B",X"DD",X"70",X"01",X"DD",
		X"71",X"02",X"18",X"4B",X"DD",X"35",X"05",X"20",X"46",X"21",X"1A",X"E2",X"11",X"15",X"00",X"06",
		X"08",X"CB",X"7E",X"28",X"05",X"19",X"10",X"F9",X"18",X"4D",X"36",X"80",X"DD",X"34",X"04",X"DD",
		X"7E",X"04",X"DD",X"BE",X"03",X"30",X"40",X"CD",X"76",X"1A",X"FE",X"14",X"38",X"02",X"3E",X"13",
		X"87",X"5F",X"16",X"00",X"21",X"A1",X"31",X"19",X"5E",X"23",X"56",X"DD",X"6E",X"04",X"26",X"00",
		X"29",X"19",X"7E",X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"01",X"DD",X"36",X"05",X"30",X"06",
		X"2D",X"0E",X"02",X"DD",X"7E",X"05",X"FE",X"10",X"38",X"06",X"E6",X"08",X"20",X"02",X"06",X"6C",
		X"11",X"80",X"78",X"CD",X"9D",X"02",X"C9",X"DD",X"CB",X"00",X"EE",X"CD",X"58",X"31",X"5F",X"87",
		X"87",X"C6",X"00",X"08",X"16",X"00",X"21",X"0D",X"32",X"19",X"7E",X"01",X"02",X"02",X"11",X"CF",
		X"81",X"CD",X"42",X"04",X"C9",X"CD",X"80",X"31",X"DD",X"7E",X"00",X"CB",X"57",X"C0",X"E6",X"18",
		X"C2",X"13",X"31",X"CD",X"58",X"31",X"5F",X"C6",X"3D",X"47",X"16",X"00",X"21",X"19",X"32",X"19",
		X"4E",X"11",X"80",X"78",X"CD",X"9D",X"02",X"3A",X"C5",X"E1",X"E6",X"98",X"FE",X"80",X"C0",X"3A",
		X"C6",X"E1",X"67",X"3A",X"C8",X"E1",X"6F",X"11",X"80",X"78",X"01",X"05",X"05",X"CD",X"EF",X"05",
		X"D0",X"DD",X"CB",X"00",X"DE",X"21",X"00",X"E0",X"CB",X"DE",X"21",X"C5",X"E1",X"CB",X"BE",X"DD",
		X"36",X"02",X"1E",X"DD",X"36",X"01",X"01",X"11",X"CF",X"89",X"01",X"02",X"01",X"CD",X"6C",X"04",
		X"11",X"D0",X"81",X"01",X"02",X"01",X"CD",X"6C",X"04",X"CD",X"58",X"31",X"5F",X"16",X"00",X"21",
		X"25",X"32",X"19",X"7E",X"21",X"7D",X"E0",X"36",X"00",X"23",X"77",X"23",X"36",X"00",X"EB",X"CD",
		X"2A",X"03",X"FD",X"36",X"1B",X"03",X"3E",X"20",X"06",X"00",X"CD",X"D9",X"02",X"CD",X"58",X"31",
		X"C6",X"16",X"32",X"CF",X"85",X"3E",X"15",X"32",X"EF",X"85",X"3E",X"09",X"32",X"CF",X"81",X"32",
		X"EF",X"81",X"C9",X"DD",X"35",X"02",X"28",X"07",X"E6",X"18",X"FE",X"08",X"28",X"DF",X"C9",X"DD",
		X"36",X"02",X"1E",X"DD",X"35",X"01",X"C0",X"E6",X"18",X"FE",X"10",X"30",X"21",X"DD",X"7E",X"00",
		X"C6",X"08",X"DD",X"77",X"00",X"DD",X"36",X"01",X"09",X"21",X"C5",X"E1",X"CB",X"FE",X"21",X"17",
		X"0B",X"CD",X"D4",X"03",X"11",X"CF",X"81",X"01",X"02",X"01",X"CD",X"6C",X"04",X"C9",X"21",X"00",
		X"E0",X"CB",X"9E",X"DD",X"CB",X"00",X"D6",X"C9",X"FD",X"7E",X"08",X"FE",X"16",X"38",X"02",X"3E",
		X"15",X"5F",X"16",X"00",X"21",X"6A",X"31",X"19",X"7E",X"C9",X"00",X"01",X"02",X"03",X"04",X"04",
		X"05",X"05",X"06",X"06",X"07",X"07",X"08",X"08",X"08",X"09",X"09",X"09",X"0A",X"0A",X"0A",X"0B",
		X"DD",X"7E",X"00",X"E6",X"03",X"FE",X"02",X"D0",X"FE",X"01",X"30",X"0D",X"FD",X"7E",X"0A",X"3D",
		X"C0",X"DD",X"34",X"00",X"DD",X"36",X"05",X"FF",X"C9",X"DD",X"35",X"05",X"C0",X"DD",X"34",X"00",
		X"C9",X"C9",X"31",X"C9",X"31",X"C9",X"31",X"C9",X"31",X"C9",X"31",X"C9",X"31",X"C9",X"31",X"C9",
		X"31",X"C9",X"31",X"D9",X"31",X"D9",X"31",X"D9",X"31",X"D9",X"31",X"D9",X"31",X"D9",X"31",X"D9",
		X"31",X"D9",X"31",X"D9",X"31",X"D9",X"31",X"E9",X"31",X"C0",X"00",X"0C",X"00",X"C0",X"00",X"0C",
		X"00",X"C0",X"00",X"0C",X"00",X"C0",X"00",X"0C",X"00",X"84",X"00",X"0C",X"00",X"84",X"00",X"0C",
		X"00",X"84",X"00",X"0C",X"00",X"84",X"00",X"0C",X"00",X"48",X"00",X"0C",X"00",X"48",X"00",X"0C",
		X"00",X"48",X"00",X"0C",X"00",X"48",X"00",X"0C",X"00",X"1E",X"1C",X"1A",X"1A",X"18",X"18",X"16",
		X"16",X"14",X"14",X"12",X"12",X"10",X"10",X"0E",X"0E",X"0C",X"0C",X"0A",X"0A",X"95",X"B4",X"84",
		X"9D",X"BC",X"B0",X"B4",X"85",X"97",X"95",X"B4",X"82",X"03",X"03",X"09",X"03",X"0E",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"10",X"15",X"20",X"25",X"30",X"35",X"40",X"45",X"50",X"60",X"70",
		X"80",X"DD",X"CB",X"00",X"76",X"20",X"2C",X"DD",X"36",X"00",X"C3",X"DD",X"36",X"01",X"78",X"DD",
		X"36",X"02",X"00",X"DD",X"36",X"03",X"80",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"10",X"DD",
		X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"13",X"00",X"DD",
		X"36",X"14",X"00",X"DD",X"7E",X"00",X"1F",X"1F",X"1F",X"DA",X"A1",X"36",X"1F",X"DA",X"7A",X"36",
		X"1F",X"DA",X"59",X"36",X"47",X"3A",X"00",X"E0",X"E6",X"40",X"20",X"08",X"CD",X"69",X"1D",X"DD",
		X"36",X"00",X"00",X"C9",X"78",X"21",X"0E",X"33",X"E5",X"1F",X"DA",X"4D",X"36",X"3A",X"B6",X"E1",
		X"A7",X"C0",X"3A",X"C5",X"E1",X"E6",X"98",X"FE",X"80",X"C0",X"FD",X"E5",X"FD",X"21",X"C5",X"E1",
		X"01",X"07",X"07",X"CD",X"D7",X"05",X"30",X"0F",X"FD",X"CB",X"00",X"DE",X"DD",X"CB",X"00",X"EE",
		X"DD",X"36",X"06",X"1E",X"FD",X"E1",X"C9",X"FD",X"E1",X"3A",X"00",X"E0",X"E6",X"08",X"C2",X"D6",
		X"41",X"3A",X"01",X"E0",X"E6",X"60",X"C2",X"D6",X"41",X"CD",X"1F",X"43",X"DD",X"7E",X"05",X"E6",
		X"F0",X"FE",X"60",X"28",X"17",X"3A",X"12",X"E2",X"E6",X"02",X"28",X"10",X"DD",X"36",X"05",X"60",
		X"DD",X"CB",X"07",X"BE",X"DD",X"36",X"0D",X"FF",X"DD",X"36",X"0E",X"FF",X"DD",X"7E",X"05",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"00",X"33",X"19",X"5E",X"23",X"56",X"EB",X"E9",
		X"D2",X"35",X"9E",X"33",X"DF",X"35",X"81",X"35",X"A5",X"33",X"12",X"34",X"BE",X"34",X"DD",X"7E",
		X"13",X"FE",X"24",X"30",X"03",X"A7",X"20",X"4A",X"AF",X"DD",X"46",X"07",X"CB",X"68",X"20",X"08",
		X"CB",X"60",X"28",X"06",X"C6",X"06",X"18",X"02",X"C6",X"0C",X"47",X"DD",X"34",X"08",X"DD",X"7E",
		X"08",X"E6",X"18",X"0F",X"0F",X"FE",X"06",X"38",X"02",X"3E",X"02",X"80",X"5F",X"16",X"00",X"21",
		X"8C",X"33",X"19",X"46",X"23",X"4E",X"DD",X"7E",X"00",X"CB",X"4F",X"28",X"0B",X"04",X"04",X"04",
		X"E6",X"01",X"28",X"0A",X"CB",X"E1",X"18",X"06",X"E6",X"01",X"28",X"02",X"CB",X"E9",X"CD",X"97",
		X"02",X"C9",X"06",X"7A",X"0E",X"08",X"FE",X"18",X"30",X"06",X"04",X"FE",X"0C",X"30",X"01",X"04",
		X"DD",X"7E",X"00",X"CB",X"4F",X"20",X"08",X"E6",X"01",X"28",X"0D",X"CB",X"E9",X"18",X"09",X"04",
		X"04",X"04",X"E6",X"01",X"28",X"02",X"CB",X"E1",X"CD",X"97",X"02",X"C9",X"2D",X"02",X"2E",X"02",
		X"2F",X"02",X"33",X"02",X"34",X"08",X"35",X"0B",X"39",X"02",X"3A",X"02",X"3B",X"02",X"CD",X"5B",
		X"3B",X"A7",X"28",X"FA",X"C9",X"CD",X"B0",X"3D",X"28",X"40",X"CD",X"C1",X"3D",X"20",X"1D",X"DD",
		X"CB",X"07",X"7E",X"20",X"1B",X"CD",X"6C",X"42",X"A7",X"C2",X"35",X"36",X"CD",X"D6",X"3D",X"FE",
		X"04",X"30",X"2F",X"DD",X"36",X"14",X"00",X"CD",X"D7",X"3E",X"18",X"04",X"DD",X"CB",X"07",X"BE",
		X"CD",X"AA",X"40",X"38",X"04",X"CD",X"02",X"3A",X"C9",X"DD",X"7E",X"00",X"EE",X"01",X"DD",X"77",
		X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"07",X"00",X"C9",X"CD",X"5B",X"3B",X"DD",X"36",X"07",
		X"00",X"C9",X"DD",X"7E",X"14",X"A7",X"20",X"05",X"DD",X"36",X"14",X"1E",X"C9",X"DD",X"35",X"14",
		X"C0",X"DD",X"36",X"05",X"60",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"3C",X"DD",X"36",X"07",
		X"00",X"C9",X"DD",X"7E",X"05",X"E6",X"0F",X"20",X"03",X"DD",X"34",X"05",X"DD",X"7E",X"13",X"A7",
		X"20",X"12",X"CD",X"B0",X"3D",X"20",X"0D",X"CD",X"C1",X"3D",X"20",X"08",X"DD",X"36",X"07",X"00",
		X"CD",X"5B",X"3B",X"C9",X"DD",X"7E",X"05",X"E6",X"0F",X"FE",X"02",X"30",X"64",X"CD",X"C1",X"3D",
		X"20",X"1D",X"DD",X"CB",X"07",X"7E",X"20",X"1B",X"CD",X"6C",X"42",X"A7",X"C2",X"35",X"36",X"CD",
		X"D6",X"3D",X"FE",X"04",X"30",X"9C",X"DD",X"36",X"14",X"00",X"CD",X"D7",X"3E",X"18",X"04",X"DD",
		X"CB",X"07",X"BE",X"CD",X"AA",X"40",X"38",X"04",X"CD",X"02",X"3A",X"C9",X"DD",X"34",X"05",X"DD",
		X"7E",X"01",X"E6",X"F0",X"47",X"DD",X"7E",X"03",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"B0",X"DD",
		X"77",X"0F",X"DD",X"7E",X"00",X"CD",X"32",X"40",X"DD",X"77",X"12",X"DD",X"7E",X"00",X"EE",X"01",
		X"DD",X"77",X"00",X"CD",X"32",X"40",X"DD",X"77",X"10",X"DD",X"77",X"11",X"DD",X"36",X"07",X"00",
		X"C9",X"CD",X"BA",X"36",X"DD",X"CB",X"07",X"66",X"C0",X"DD",X"7E",X"05",X"E6",X"0F",X"FE",X"03",
		X"C0",X"DD",X"35",X"05",X"DD",X"7E",X"12",X"A7",X"C0",X"DD",X"36",X"05",X"51",X"C9",X"DD",X"7E",
		X"05",X"E6",X"0F",X"20",X"14",X"DD",X"34",X"05",X"DD",X"36",X"13",X"00",X"DD",X"36",X"14",X"00",
		X"DD",X"CB",X"07",X"66",X"28",X"03",X"DD",X"34",X"05",X"DD",X"7E",X"13",X"A7",X"20",X"2F",X"CD",
		X"B0",X"3D",X"20",X"0D",X"CD",X"C1",X"3D",X"20",X"25",X"DD",X"36",X"07",X"00",X"CD",X"5B",X"3B",
		X"C9",X"DD",X"7E",X"14",X"A7",X"20",X"13",X"DD",X"7E",X"0E",X"E6",X"3F",X"20",X"10",X"CD",X"F4",
		X"02",X"E6",X"03",X"20",X"09",X"DD",X"36",X"14",X"20",X"C9",X"DD",X"35",X"14",X"C9",X"DD",X"7E",
		X"05",X"E6",X"0F",X"FE",X"02",X"30",X"4D",X"CD",X"C1",X"3D",X"20",X"24",X"DD",X"CB",X"07",X"7E",
		X"20",X"22",X"CD",X"6C",X"42",X"A7",X"C2",X"35",X"36",X"CD",X"A2",X"37",X"DD",X"7E",X"05",X"E6",
		X"0F",X"FE",X"02",X"D0",X"CD",X"D6",X"3D",X"FE",X"04",X"30",X"16",X"CD",X"D7",X"3E",X"18",X"04",
		X"DD",X"CB",X"07",X"BE",X"CD",X"AA",X"40",X"38",X"04",X"CD",X"02",X"3A",X"C9",X"CD",X"6C",X"34",
		X"C9",X"DD",X"34",X"05",X"DD",X"36",X"0F",X"00",X"DD",X"7E",X"00",X"EE",X"01",X"CD",X"32",X"40",
		X"DD",X"77",X"10",X"C9",X"CD",X"BA",X"36",X"DD",X"CB",X"07",X"66",X"C0",X"DD",X"7E",X"05",X"E6",
		X"0F",X"FE",X"03",X"C0",X"DD",X"35",X"05",X"DD",X"7E",X"12",X"A7",X"C0",X"DD",X"36",X"05",X"60",
		X"C9",X"CD",X"B0",X"3D",X"28",X"44",X"CD",X"C1",X"3D",X"20",X"19",X"DD",X"CB",X"07",X"7E",X"20",
		X"17",X"CD",X"6C",X"42",X"A7",X"C2",X"35",X"36",X"CD",X"1A",X"3E",X"FE",X"04",X"30",X"12",X"CD",
		X"D7",X"3E",X"18",X"04",X"DD",X"CB",X"07",X"BE",X"CD",X"AA",X"40",X"38",X"15",X"CD",X"02",X"3A",
		X"C9",X"DD",X"36",X"05",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"B4",X"DD",X"36",X"07",
		X"00",X"C9",X"DD",X"7E",X"00",X"EE",X"01",X"DD",X"77",X"00",X"CD",X"5B",X"3B",X"DD",X"36",X"07",
		X"00",X"C9",X"CD",X"B0",X"3D",X"28",X"04",X"CD",X"D6",X"41",X"C9",X"CD",X"5B",X"3B",X"C9",X"CD",
		X"B0",X"3D",X"28",X"49",X"CD",X"C1",X"3D",X"20",X"2C",X"DD",X"CB",X"07",X"7E",X"20",X"2A",X"CD",
		X"6C",X"42",X"A7",X"20",X"40",X"CD",X"7C",X"3E",X"FE",X"04",X"30",X"31",X"DD",X"4E",X"00",X"CD",
		X"D7",X"3E",X"A9",X"E6",X"03",X"FE",X"01",X"20",X"10",X"DD",X"7E",X"05",X"DD",X"34",X"05",X"E6",
		X"0F",X"20",X"1A",X"18",X"1B",X"DD",X"CB",X"07",X"BE",X"CD",X"41",X"40",X"CD",X"76",X"40",X"38",
		X"04",X"CD",X"02",X"3A",X"C9",X"DD",X"7E",X"00",X"EE",X"01",X"DD",X"77",X"00",X"CD",X"5B",X"3B",
		X"DD",X"36",X"07",X"00",X"C9",X"CD",X"FF",X"42",X"C8",X"CD",X"D7",X"3E",X"CD",X"41",X"40",X"CD",
		X"76",X"40",X"38",X"04",X"CD",X"02",X"3A",X"C9",X"DD",X"CB",X"07",X"BE",X"C9",X"DD",X"35",X"06",
		X"C0",X"CD",X"69",X"1D",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"CB",X"07",X"4E",X"20",X"0E",X"DD",
		X"CB",X"07",X"CE",X"CD",X"69",X"1D",X"CD",X"A6",X"36",X"DD",X"36",X"06",X"00",X"DD",X"35",X"06",
		X"28",X"2F",X"06",X"3C",X"0E",X"02",X"CD",X"97",X"02",X"C9",X"DD",X"CB",X"07",X"46",X"20",X"14",
		X"DD",X"CB",X"07",X"C6",X"DD",X"36",X"06",X"1F",X"CD",X"69",X"1D",X"CD",X"A6",X"36",X"11",X"5A",
		X"3B",X"CD",X"2A",X"03",X"DD",X"35",X"06",X"28",X"08",X"06",X"71",X"0E",X"0A",X"CD",X"97",X"02",
		X"C9",X"DD",X"36",X"00",X"00",X"C9",X"FD",X"35",X"0A",X"C0",X"21",X"B6",X"E1",X"CB",X"FE",X"FD",
		X"36",X"30",X"01",X"FD",X"7E",X"08",X"FD",X"77",X"09",X"C9",X"CD",X"C1",X"3D",X"20",X"31",X"DD",
		X"CB",X"07",X"7E",X"20",X"2F",X"DD",X"7E",X"01",X"E6",X"F0",X"47",X"DD",X"7E",X"03",X"3C",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"B0",X"DD",X"BE",X"0F",X"28",X"06",X"DD",X"77",X"0F",X"CD",X"3C",
		X"37",X"CD",X"51",X"3F",X"FE",X"04",X"D0",X"CD",X"D7",X"3E",X"DD",X"CB",X"07",X"B6",X"18",X"04",
		X"DD",X"CB",X"07",X"BE",X"CD",X"AA",X"40",X"38",X"27",X"CD",X"80",X"38",X"DD",X"CB",X"07",X"F6",
		X"DD",X"CB",X"07",X"66",X"28",X"0C",X"DD",X"7E",X"05",X"E6",X"0F",X"FE",X"03",X"30",X"03",X"DD",
		X"34",X"05",X"DD",X"7E",X"13",X"A7",X"28",X"04",X"DD",X"35",X"13",X"C0",X"CD",X"02",X"3A",X"C9",
		X"DD",X"7E",X"00",X"CD",X"32",X"40",X"DD",X"B6",X"12",X"DD",X"77",X"12",X"CD",X"69",X"1D",X"DD",
		X"7E",X"00",X"EE",X"01",X"DD",X"77",X"00",X"DD",X"36",X"13",X"00",X"C9",X"DD",X"7E",X"00",X"EE",
		X"01",X"CD",X"32",X"40",X"DD",X"77",X"11",X"DD",X"36",X"12",X"00",X"DD",X"7E",X"10",X"CB",X"5F",
		X"20",X"36",X"CB",X"4F",X"20",X"22",X"CB",X"57",X"20",X"0F",X"DD",X"7E",X"01",X"E6",X"F0",X"47",
		X"3A",X"C6",X"E1",X"E6",X"F0",X"B8",X"38",X"2E",X"C9",X"3A",X"C6",X"E1",X"E6",X"F0",X"47",X"DD",
		X"7E",X"01",X"E6",X"F0",X"B8",X"38",X"1F",X"C9",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"47",X"3A",
		X"C8",X"E1",X"E6",X"F0",X"B8",X"38",X"0F",X"C9",X"3A",X"C8",X"E1",X"E6",X"F0",X"47",X"DD",X"7E",
		X"03",X"3C",X"E6",X"F0",X"B8",X"D0",X"DD",X"7E",X"00",X"EE",X"01",X"CD",X"32",X"40",X"DD",X"77",
		X"10",X"C9",X"DD",X"7E",X"01",X"E6",X"F0",X"0F",X"57",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"0F",
		X"5F",X"3A",X"C6",X"E1",X"E6",X"F0",X"0F",X"92",X"30",X"02",X"ED",X"44",X"57",X"3A",X"C8",X"E1",
		X"E6",X"F0",X"0F",X"93",X"30",X"02",X"ED",X"44",X"BA",X"38",X"0D",X"28",X"0B",X"CD",X"04",X"38",
		X"CD",X"23",X"38",X"CD",X"3A",X"38",X"18",X"09",X"CD",X"04",X"38",X"CD",X"3A",X"38",X"CD",X"23",
		X"38",X"CD",X"A3",X"1D",X"23",X"D9",X"7C",X"D9",X"BE",X"38",X"05",X"DD",X"36",X"05",X"61",X"C9",
		X"DD",X"36",X"05",X"62",X"AF",X"DD",X"77",X"0F",X"DD",X"7E",X"00",X"EE",X"01",X"CD",X"32",X"40",
		X"DD",X"77",X"10",X"C9",X"D9",X"21",X"00",X"00",X"D9",X"DD",X"7E",X"01",X"E6",X"F0",X"57",X"DD",
		X"7E",X"03",X"3C",X"E6",X"F0",X"5F",X"3A",X"C6",X"E1",X"E6",X"F0",X"47",X"3A",X"C8",X"E1",X"E6",
		X"F0",X"4F",X"C9",X"78",X"BA",X"C8",X"38",X"09",X"CD",X"51",X"38",X"7A",X"C6",X"10",X"57",X"18",
		X"F2",X"CD",X"51",X"38",X"7A",X"D6",X"10",X"57",X"18",X"E9",X"79",X"BB",X"C8",X"38",X"09",X"CD",
		X"51",X"38",X"7B",X"C6",X"10",X"5F",X"18",X"F2",X"CD",X"51",X"38",X"7B",X"D6",X"10",X"5F",X"18",
		X"E9",X"D5",X"CD",X"C0",X"1D",X"D1",X"7E",X"E6",X"0F",X"28",X"04",X"D9",X"24",X"D9",X"C9",X"D9",
		X"EB",X"CD",X"76",X"1A",X"EB",X"11",X"7F",X"38",X"FE",X"0F",X"30",X"0B",X"1B",X"FE",X"0A",X"30",
		X"06",X"1B",X"FE",X"05",X"30",X"01",X"1B",X"1A",X"84",X"67",X"D9",X"C9",X"05",X"04",X"03",X"02",
		X"DD",X"7E",X"00",X"E6",X"03",X"CA",X"7A",X"39",X"FE",X"01",X"CA",X"2A",X"39",X"FE",X"02",X"28",
		X"49",X"DD",X"CB",X"07",X"76",X"20",X"20",X"DD",X"7E",X"03",X"E6",X"0F",X"28",X"04",X"FE",X"0F",
		X"20",X"15",X"CD",X"A3",X"1D",X"CB",X"4E",X"28",X"08",X"CD",X"1B",X"28",X"DD",X"36",X"13",X"00",
		X"C9",X"CD",X"D2",X"39",X"CD",X"29",X"28",X"DD",X"7E",X"03",X"E6",X"03",X"FE",X"02",X"DA",X"CD",
		X"39",X"DD",X"7E",X"07",X"E6",X"14",X"FE",X"10",X"C0",X"CD",X"D0",X"1A",X"CD",X"E1",X"39",X"DD",
		X"7E",X"03",X"E6",X"0F",X"FE",X"04",X"DC",X"1F",X"1E",X"C9",X"CD",X"78",X"1F",X"DD",X"CB",X"07",
		X"76",X"20",X"21",X"DD",X"7E",X"03",X"E6",X"0F",X"28",X"04",X"FE",X"0F",X"20",X"16",X"CD",X"A3",
		X"1D",X"CB",X"5E",X"28",X"08",X"CD",X"1B",X"28",X"DD",X"36",X"13",X"00",X"C9",X"CD",X"D2",X"39",
		X"CD",X"29",X"28",X"C9",X"DD",X"7E",X"03",X"E6",X"03",X"CA",X"CD",X"39",X"FE",X"03",X"CA",X"CD",
		X"39",X"DD",X"7E",X"07",X"E6",X"14",X"FE",X"10",X"C0",X"CD",X"9B",X"1A",X"CD",X"E1",X"39",X"DD",
		X"7E",X"03",X"E6",X"0F",X"FE",X"0D",X"D4",X"C9",X"1D",X"C9",X"CD",X"78",X"1F",X"DD",X"CB",X"07",
		X"76",X"20",X"22",X"DD",X"7E",X"01",X"E6",X"0F",X"FE",X"07",X"28",X"04",X"FE",X"08",X"20",X"15",
		X"CD",X"A3",X"1D",X"CB",X"46",X"28",X"08",X"CD",X"1B",X"28",X"DD",X"36",X"13",X"00",X"C9",X"CD",
		X"D2",X"39",X"CD",X"29",X"28",X"DD",X"7E",X"01",X"E6",X"03",X"FE",X"02",X"38",X"6F",X"DD",X"7E",
		X"07",X"E6",X"14",X"FE",X"10",X"C0",X"CD",X"3B",X"1B",X"CD",X"E1",X"39",X"DD",X"7E",X"01",X"E6",
		X"0F",X"FE",X"0A",X"D8",X"FE",X"0D",X"DC",X"C5",X"1E",X"C9",X"CD",X"78",X"1F",X"DD",X"CB",X"07",
		X"76",X"20",X"23",X"DD",X"7E",X"01",X"E6",X"0F",X"FE",X"07",X"28",X"04",X"FE",X"08",X"20",X"16",
		X"CD",X"A3",X"1D",X"CB",X"56",X"28",X"08",X"CD",X"1B",X"28",X"DD",X"36",X"13",X"00",X"C9",X"CD",
		X"D2",X"39",X"CD",X"29",X"28",X"C9",X"DD",X"7E",X"01",X"E6",X"03",X"28",X"20",X"FE",X"03",X"28",
		X"1C",X"DD",X"7E",X"07",X"E6",X"14",X"FE",X"10",X"C0",X"CD",X"05",X"1B",X"CD",X"E1",X"39",X"DD",
		X"7E",X"01",X"E6",X"0F",X"FE",X"07",X"D0",X"FE",X"05",X"D4",X"75",X"1E",X"C9",X"DD",X"CB",X"07",
		X"96",X"C9",X"DD",X"CB",X"07",X"66",X"C0",X"DD",X"7E",X"13",X"A7",X"C0",X"DD",X"36",X"13",X"30",
		X"C9",X"DD",X"E5",X"E1",X"11",X"09",X"00",X"19",X"3E",X"DB",X"06",X"04",X"BE",X"30",X"05",X"FD",
		X"35",X"0B",X"28",X"04",X"23",X"10",X"F5",X"C9",X"21",X"B6",X"E1",X"CB",X"FE",X"FD",X"36",X"30",
		X"02",X"C9",X"DD",X"46",X"07",X"CB",X"68",X"20",X"32",X"CD",X"76",X"1A",X"FE",X"20",X"38",X"02",
		X"3E",X"1F",X"5F",X"16",X"00",X"21",X"88",X"3A",X"19",X"5E",X"FD",X"7E",X"0E",X"CB",X"60",X"20",
		X"0B",X"21",X"A8",X"3A",X"A7",X"20",X"0E",X"21",X"D4",X"3A",X"18",X"09",X"21",X"00",X"3B",X"A7",
		X"20",X"03",X"21",X"2C",X"3B",X"19",X"4E",X"23",X"46",X"18",X"03",X"01",X"55",X"00",X"DD",X"7E",
		X"00",X"CB",X"4F",X"28",X"1C",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"1F",X"DC",X"E3",X"2C",X"09",
		X"DD",X"74",X"03",X"DD",X"75",X"04",X"DD",X"7E",X"01",X"E6",X"F0",X"C6",X"08",X"DD",X"77",X"01",
		X"C9",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"1F",X"DC",X"E3",X"2C",X"09",X"DD",X"74",X"01",X"DD",
		X"75",X"02",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"DD",X"77",X"03",X"DD",X"CB",X"07",X"6E",X"C8",
		X"50",X"59",X"06",X"90",X"CD",X"3F",X"1F",X"C9",X"00",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0E",
		X"10",X"12",X"14",X"16",X"16",X"18",X"18",X"1A",X"1A",X"1C",X"1C",X"1E",X"1E",X"20",X"20",X"22",
		X"22",X"24",X"24",X"26",X"26",X"28",X"28",X"2A",X"D5",X"00",X"E2",X"00",X"EB",X"00",X"F3",X"00",
		X"FC",X"00",X"04",X"01",X"09",X"01",X"0D",X"01",X"11",X"01",X"13",X"01",X"15",X"01",X"17",X"01",
		X"1A",X"01",X"1C",X"01",X"1E",X"01",X"20",X"01",X"22",X"01",X"24",X"01",X"26",X"01",X"29",X"01",
		X"2B",X"01",X"33",X"01",X"00",X"01",X"0D",X"01",X"15",X"01",X"1A",X"01",X"1E",X"01",X"22",X"01",
		X"26",X"01",X"2B",X"01",X"2F",X"01",X"31",X"01",X"33",X"01",X"35",X"01",X"37",X"01",X"3A",X"01",
		X"3C",X"01",X"3E",X"01",X"40",X"01",X"42",X"01",X"44",X"01",X"49",X"01",X"4D",X"01",X"55",X"01",
		X"80",X"00",X"89",X"00",X"8D",X"00",X"91",X"00",X"95",X"00",X"9A",X"00",X"9E",X"00",X"A0",X"00",
		X"A2",X"00",X"A4",X"00",X"A6",X"00",X"A9",X"00",X"AB",X"00",X"AD",X"00",X"AF",X"00",X"B1",X"00",
		X"B3",X"00",X"B5",X"00",X"B7",X"00",X"BA",X"00",X"BC",X"00",X"C0",X"00",X"9A",X"00",X"A2",X"00",
		X"A6",X"00",X"AB",X"00",X"AF",X"00",X"B3",X"00",X"B7",X"00",X"BA",X"00",X"BC",X"00",X"BE",X"00",
		X"C0",X"00",X"C2",X"00",X"C4",X"00",X"C6",X"00",X"C9",X"00",X"CB",X"00",X"CD",X"00",X"CF",X"00",
		X"D1",X"00",X"D3",X"00",X"D5",X"00",X"DE",X"00",X"00",X"05",X"00",X"CD",X"F4",X"02",X"47",X"FD",
		X"7E",X"09",X"21",X"00",X"E0",X"CB",X"7E",X"28",X"0E",X"21",X"02",X"A0",X"CB",X"4E",X"20",X"07",
		X"FE",X"80",X"30",X"03",X"87",X"C6",X"01",X"FE",X"20",X"38",X"02",X"3E",X"1F",X"87",X"87",X"87",
		X"4F",X"FD",X"7E",X"12",X"E6",X"38",X"0F",X"0F",X"0F",X"81",X"5F",X"16",X"00",X"21",X"C0",X"3B",
		X"19",X"78",X"E6",X"07",X"86",X"5F",X"16",X"00",X"21",X"B8",X"3C",X"19",X"7E",X"CB",X"58",X"20",
		X"04",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"80",X"3D",
		X"19",X"7E",X"23",X"4E",X"23",X"46",X"DD",X"77",X"05",X"DD",X"70",X"0D",X"DD",X"71",X"0E",X"C9",
		X"08",X"10",X"20",X"30",X"40",X"50",X"80",X"80",X"08",X"18",X"30",X"40",X"48",X"70",X"80",X"80",
		X"08",X"20",X"38",X"48",X"58",X"78",X"88",X"88",X"08",X"28",X"40",X"50",X"68",X"80",X"88",X"88",
		X"08",X"30",X"48",X"58",X"70",X"88",X"90",X"90",X"10",X"38",X"50",X"60",X"78",X"88",X"90",X"90",
		X"10",X"40",X"58",X"68",X"80",X"90",X"98",X"98",X"10",X"48",X"60",X"70",X"88",X"90",X"98",X"98",
		X"10",X"50",X"68",X"78",X"88",X"98",X"A0",X"A0",X"10",X"58",X"70",X"80",X"90",X"98",X"A0",X"A0",
		X"18",X"60",X"78",X"88",X"90",X"A0",X"A8",X"A8",X"18",X"68",X"80",X"88",X"98",X"A0",X"A8",X"A8",
		X"18",X"70",X"80",X"90",X"98",X"A8",X"B0",X"B0",X"18",X"78",X"88",X"90",X"A0",X"A8",X"B0",X"B0",
		X"18",X"80",X"88",X"98",X"A0",X"B0",X"B8",X"B8",X"20",X"88",X"90",X"98",X"A8",X"B0",X"B8",X"B8",
		X"20",X"88",X"90",X"A0",X"A8",X"B8",X"C0",X"C0",X"20",X"90",X"98",X"A0",X"B0",X"B8",X"C0",X"C0",
		X"20",X"90",X"98",X"A8",X"B0",X"B8",X"C0",X"C0",X"20",X"98",X"A0",X"A8",X"B8",X"C0",X"C0",X"C0",
		X"28",X"98",X"A0",X"B0",X"B8",X"C0",X"C0",X"C0",X"28",X"A0",X"A8",X"B0",X"B8",X"C0",X"C0",X"C0",
		X"28",X"A0",X"A8",X"B8",X"C0",X"C0",X"C0",X"C0",X"28",X"A8",X"B0",X"B8",X"C0",X"C0",X"C0",X"C0",
		X"28",X"A8",X"B0",X"B8",X"C0",X"C0",X"C0",X"C0",X"30",X"B0",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"30",X"B0",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",X"30",X"B0",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"30",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"30",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"38",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"11",X"11",X"22",X"22",X"AB",X"EE",X"00",X"01",X"11",X"22",X"24",X"AB",X"BC",X"EF",
		X"00",X"00",X"11",X"12",X"23",X"4A",X"BE",X"EF",X"00",X"01",X"11",X"22",X"34",X"BE",X"FF",X"FF",
		X"00",X"01",X"11",X"22",X"24",X"7B",X"EF",X"FF",X"00",X"01",X"11",X"22",X"23",X"45",X"6B",X"EF",
		X"00",X"01",X"11",X"22",X"24",X"67",X"BE",X"EF",X"00",X"01",X"11",X"22",X"24",X"67",X"8B",X"EF",
		X"00",X"11",X"22",X"33",X"44",X"55",X"7B",X"EF",X"00",X"11",X"22",X"44",X"46",X"78",X"BE",X"EF",
		X"00",X"01",X"11",X"22",X"24",X"79",X"BE",X"FF",X"00",X"01",X"11",X"22",X"24",X"79",X"9B",X"EF",
		X"00",X"11",X"22",X"44",X"67",X"89",X"BE",X"EF",X"00",X"11",X"22",X"44",X"78",X"99",X"BE",X"EF",
		X"01",X"24",X"46",X"67",X"78",X"8A",X"BE",X"FF",X"00",X"11",X"22",X"44",X"79",X"99",X"BE",X"FF",
		X"01",X"24",X"46",X"67",X"79",X"9A",X"BE",X"FF",X"01",X"24",X"66",X"77",X"88",X"9B",X"EE",X"FF",
		X"01",X"24",X"47",X"78",X"89",X"99",X"BE",X"FF",X"01",X"24",X"67",X"78",X"89",X"99",X"9B",X"EF",
		X"01",X"24",X"67",X"89",X"99",X"99",X"9B",X"EF",X"01",X"46",X"79",X"99",X"99",X"99",X"9B",X"EF",
		X"01",X"79",X"99",X"99",X"99",X"99",X"9F",X"FF",X"17",X"99",X"99",X"99",X"99",X"99",X"9E",X"FF",
		X"40",X"3C",X"00",X"40",X"78",X"00",X"40",X"B4",X"00",X"50",X"3C",X"00",X"50",X"78",X"00",X"50",
		X"B4",X"00",X"60",X"3C",X"00",X"60",X"78",X"00",X"60",X"B4",X"00",X"60",X"FF",X"FF",X"20",X"3C",
		X"00",X"20",X"78",X"00",X"20",X"B4",X"00",X"20",X"2C",X"01",X"00",X"1E",X"00",X"30",X"58",X"02",
		X"DD",X"46",X"0D",X"DD",X"4E",X"0E",X"78",X"B1",X"C8",X"0B",X"DD",X"70",X"0D",X"DD",X"71",X"0E",
		X"C9",X"DD",X"7E",X"01",X"E6",X"0F",X"FE",X"07",X"28",X"03",X"FE",X"08",X"C0",X"DD",X"7E",X"03",
		X"E6",X"0F",X"C8",X"FE",X"0F",X"C9",X"CD",X"A3",X"1D",X"46",X"23",X"7E",X"CB",X"50",X"28",X"0B",
		X"EB",X"21",X"20",X"00",X"19",X"BE",X"EB",X"38",X"02",X"AF",X"C9",X"CB",X"40",X"28",X"0C",X"EB",
		X"21",X"E0",X"FF",X"19",X"BE",X"EB",X"38",X"03",X"3E",X"01",X"C9",X"CB",X"58",X"28",X"0A",X"23",
		X"23",X"BE",X"2B",X"2B",X"38",X"03",X"3E",X"02",X"C9",X"CB",X"48",X"28",X"0A",X"2B",X"2B",X"BE",
		X"23",X"23",X"38",X"03",X"3E",X"03",X"C9",X"3E",X"04",X"C9",X"CD",X"A3",X"1D",X"46",X"CB",X"70",
		X"28",X"B4",X"23",X"4E",X"CB",X"58",X"28",X"10",X"23",X"56",X"23",X"7E",X"2B",X"2B",X"CB",X"72",
		X"28",X"06",X"B9",X"38",X"03",X"3E",X"02",X"C9",X"CB",X"50",X"28",X"12",X"EB",X"21",X"20",X"00",
		X"19",X"7E",X"2B",X"CB",X"76",X"EB",X"28",X"06",X"B9",X"38",X"03",X"3E",X"00",X"C9",X"CB",X"48",
		X"28",X"11",X"2B",X"2B",X"7E",X"2B",X"CB",X"76",X"23",X"23",X"23",X"28",X"06",X"B9",X"38",X"03",
		X"3E",X"03",X"C9",X"CB",X"40",X"28",X"12",X"EB",X"21",X"E0",X"FF",X"19",X"7E",X"2B",X"CB",X"76",
		X"EB",X"28",X"06",X"B9",X"38",X"03",X"3E",X"01",X"C9",X"3E",X"04",X"C9",X"CD",X"A3",X"1D",X"46",
		X"23",X"0E",X"00",X"CB",X"58",X"28",X"0C",X"0C",X"23",X"23",X"7E",X"2B",X"2B",X"BE",X"38",X"03",
		X"3E",X"02",X"C9",X"CB",X"50",X"28",X"0E",X"0C",X"EB",X"21",X"20",X"00",X"19",X"EB",X"1A",X"BE",
		X"38",X"03",X"3E",X"00",X"C9",X"CB",X"48",X"28",X"0C",X"0C",X"2B",X"2B",X"7E",X"23",X"23",X"BE",
		X"38",X"03",X"3E",X"03",X"C9",X"CB",X"40",X"28",X"0E",X"0C",X"EB",X"21",X"E0",X"FF",X"19",X"EB",
		X"1A",X"BE",X"38",X"03",X"3E",X"01",X"C9",X"79",X"FE",X"02",X"30",X"08",X"DD",X"7E",X"00",X"EE",
		X"01",X"E6",X"03",X"C9",X"3E",X"04",X"C9",X"47",X"DD",X"7E",X"00",X"E6",X"FC",X"B0",X"DD",X"77",
		X"00",X"DD",X"CB",X"07",X"FE",X"C9",X"CD",X"A3",X"1D",X"46",X"23",X"4E",X"DD",X"7E",X"00",X"E6",
		X"03",X"FE",X"03",X"28",X"0F",X"CB",X"58",X"28",X"0B",X"23",X"23",X"7E",X"2B",X"2B",X"B9",X"38",
		X"03",X"3E",X"02",X"C9",X"DD",X"7E",X"00",X"E6",X"03",X"FE",X"01",X"28",X"11",X"CB",X"50",X"28",
		X"0D",X"EB",X"21",X"20",X"00",X"19",X"EB",X"1A",X"B9",X"38",X"03",X"3E",X"00",X"C9",X"DD",X"7E",
		X"00",X"E6",X"03",X"FE",X"02",X"28",X"0F",X"CB",X"48",X"28",X"0B",X"2B",X"2B",X"7E",X"23",X"23",
		X"B9",X"38",X"03",X"3E",X"03",X"C9",X"DD",X"7E",X"00",X"E6",X"03",X"28",X"11",X"CB",X"40",X"28",
		X"0D",X"EB",X"21",X"E0",X"FF",X"19",X"EB",X"1A",X"B9",X"38",X"03",X"3E",X"01",X"C9",X"3E",X"04",
		X"C9",X"DD",X"7E",X"01",X"3C",X"E6",X"FE",X"0F",X"57",X"DD",X"7E",X"03",X"3C",X"E6",X"FE",X"0F",
		X"5F",X"3A",X"C6",X"E1",X"E6",X"FE",X"0F",X"92",X"67",X"30",X"02",X"ED",X"44",X"57",X"3A",X"C8",
		X"E1",X"E6",X"FE",X"0F",X"93",X"6F",X"30",X"02",X"ED",X"44",X"5F",X"28",X"07",X"7A",X"A7",X"28",
		X"21",X"BB",X"30",X"1E",X"CB",X"7D",X"20",X"06",X"0E",X"08",X"16",X"02",X"18",X"04",X"0E",X"02",
		X"16",X"08",X"CB",X"7C",X"20",X"06",X"06",X"04",X"1E",X"01",X"18",X"22",X"06",X"01",X"1E",X"04",
		X"18",X"1C",X"CB",X"7C",X"20",X"06",X"0E",X"04",X"16",X"01",X"18",X"04",X"0E",X"01",X"16",X"04",
		X"CB",X"7D",X"20",X"06",X"06",X"08",X"1E",X"02",X"18",X"04",X"06",X"02",X"1E",X"08",X"21",X"8D",
		X"E0",X"70",X"23",X"71",X"23",X"72",X"23",X"73",X"21",X"8D",X"E0",X"06",X"04",X"DD",X"7E",X"10",
		X"DD",X"B6",X"11",X"DD",X"B6",X"12",X"2F",X"4F",X"79",X"A6",X"28",X"06",X"CD",X"FF",X"3F",X"FE",
		X"04",X"D8",X"23",X"10",X"F3",X"21",X"8D",X"E0",X"06",X"04",X"DD",X"7E",X"12",X"2F",X"4F",X"79",
		X"A6",X"28",X"06",X"CD",X"FF",X"3F",X"FE",X"04",X"D8",X"23",X"10",X"F3",X"3E",X"04",X"C9",X"CB",
		X"5F",X"20",X"25",X"CB",X"57",X"20",X"18",X"CB",X"4F",X"20",X"0A",X"DD",X"7E",X"01",X"FE",X"29",
		X"38",X"EA",X"3E",X"01",X"C9",X"DD",X"7E",X"03",X"FE",X"21",X"38",X"E0",X"3E",X"03",X"C9",X"DD",
		X"7E",X"01",X"FE",X"D7",X"30",X"D6",X"AF",X"C9",X"DD",X"7E",X"03",X"FE",X"DF",X"30",X"CD",X"3E",
		X"02",X"C9",X"E6",X"03",X"5F",X"16",X"00",X"21",X"3D",X"40",X"19",X"7E",X"C9",X"04",X"01",X"08",
		X"02",X"DD",X"56",X"01",X"DD",X"5E",X"03",X"DD",X"7E",X"00",X"E6",X"03",X"28",X"20",X"FE",X"01",
		X"28",X"14",X"FE",X"02",X"28",X"08",X"7B",X"D6",X"07",X"5F",X"01",X"07",X"0E",X"C9",X"7B",X"C6",
		X"07",X"5F",X"01",X"07",X"0E",X"C9",X"7A",X"D6",X"07",X"57",X"01",X"0E",X"07",X"C9",X"7A",X"C6",
		X"07",X"57",X"01",X"0E",X"07",X"C9",X"FD",X"E5",X"D9",X"11",X"31",X"00",X"FD",X"19",X"06",X"0C",
		X"11",X"07",X"00",X"D9",X"FD",X"7E",X"00",X"FE",X"80",X"38",X"16",X"FE",X"D0",X"28",X"04",X"FE",
		X"B8",X"30",X"0E",X"FD",X"66",X"01",X"FD",X"6E",X"03",X"CD",X"EF",X"05",X"30",X"03",X"FD",X"E1",
		X"C9",X"D9",X"FD",X"19",X"10",X"DD",X"FD",X"E1",X"A7",X"C9",X"DD",X"CB",X"00",X"4E",X"28",X"0B",
		X"CD",X"41",X"40",X"CD",X"76",X"40",X"DD",X"CB",X"07",X"AE",X"C9",X"DD",X"4E",X"00",X"DD",X"56",
		X"01",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"5F",X"21",X"80",X"E0",X"36",X"00",X"23",X"D9",X"FD",
		X"E5",X"11",X"31",X"00",X"FD",X"19",X"11",X"07",X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",X"80",
		X"38",X"6D",X"FE",X"D0",X"28",X"04",X"FE",X"B8",X"30",X"65",X"D9",X"FD",X"7E",X"03",X"93",X"20",
		X"43",X"CB",X"41",X"20",X"06",X"FD",X"7E",X"01",X"92",X"18",X"04",X"7A",X"FD",X"96",X"01",X"28",
		X"4D",X"FE",X"11",X"30",X"49",X"FE",X"0F",X"D2",X"9B",X"41",X"FD",X"7E",X"00",X"FE",X"90",X"D2",
		X"A9",X"41",X"3A",X"80",X"E0",X"3C",X"32",X"80",X"E0",X"D9",X"78",X"D9",X"77",X"23",X"FD",X"56",
		X"01",X"FD",X"5E",X"03",X"7A",X"FE",X"D8",X"D2",X"A9",X"41",X"FE",X"29",X"DA",X"A9",X"41",X"D9",
		X"FD",X"E1",X"18",X"9B",X"FE",X"09",X"38",X"04",X"FE",X"F8",X"38",X"12",X"CB",X"41",X"20",X"06",
		X"FD",X"7E",X"01",X"92",X"18",X"04",X"7A",X"FD",X"96",X"01",X"FE",X"0F",X"38",X"5B",X"D9",X"FD",
		X"19",X"10",X"88",X"3A",X"80",X"E0",X"A7",X"28",X"48",X"D9",X"3E",X"08",X"CB",X"41",X"28",X"02",
		X"3E",X"F8",X"D5",X"82",X"57",X"CD",X"0B",X"54",X"D1",X"38",X"3E",X"3E",X"07",X"CB",X"41",X"28",
		X"02",X"3E",X"F9",X"82",X"57",X"CD",X"AD",X"41",X"38",X"2F",X"3A",X"C5",X"E1",X"E6",X"98",X"FE",
		X"80",X"20",X"10",X"3A",X"C6",X"E1",X"67",X"3A",X"C8",X"E1",X"6F",X"01",X"0E",X"08",X"CD",X"EF",
		X"05",X"38",X"16",X"FD",X"E1",X"DD",X"CB",X"07",X"EE",X"A7",X"C9",X"3A",X"80",X"E0",X"A7",X"20",
		X"F2",X"FD",X"E1",X"DD",X"CB",X"07",X"AE",X"A7",X"C9",X"FD",X"E1",X"37",X"C9",X"01",X"02",X"06",
		X"D9",X"FD",X"21",X"1A",X"E2",X"11",X"15",X"00",X"06",X"08",X"D9",X"FD",X"7E",X"00",X"E6",X"98",
		X"FE",X"80",X"20",X"0A",X"FD",X"66",X"01",X"FD",X"6E",X"03",X"CD",X"EF",X"05",X"D8",X"D9",X"FD",
		X"19",X"10",X"E7",X"D9",X"A7",X"C9",X"DD",X"CB",X"07",X"66",X"C0",X"DD",X"7E",X"13",X"A7",X"C0",
		X"FD",X"E5",X"11",X"31",X"00",X"FD",X"19",X"11",X"07",X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",
		X"98",X"20",X"1A",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"28",X"04",X"FE",X"FF",X"38",X"0E",X"DD",
		X"7E",X"01",X"FD",X"96",X"01",X"FE",X"0E",X"38",X"0B",X"FE",X"F3",X"30",X"11",X"FD",X"19",X"10",
		X"DB",X"FD",X"E1",X"C9",X"DD",X"7E",X"00",X"E6",X"FC",X"DD",X"77",X"00",X"18",X"0A",X"DD",X"7E",
		X"00",X"E6",X"FC",X"F6",X"01",X"DD",X"77",X"00",X"FD",X"E1",X"CD",X"C1",X"3D",X"20",X"35",X"CD",
		X"A3",X"1D",X"DD",X"7E",X"00",X"E6",X"03",X"20",X"05",X"7E",X"E6",X"0E",X"18",X"03",X"7E",X"E6",
		X"0B",X"CB",X"57",X"20",X"17",X"CB",X"47",X"20",X"0F",X"CB",X"4F",X"20",X"07",X"CB",X"5F",X"C8",
		X"3E",X"02",X"18",X"09",X"3E",X"03",X"18",X"05",X"3E",X"01",X"18",X"01",X"AF",X"CD",X"D7",X"3E",
		X"DD",X"CB",X"07",X"BE",X"CD",X"AA",X"40",X"D8",X"CD",X"02",X"3A",X"C9",X"CD",X"A3",X"1D",X"FD",
		X"E5",X"11",X"31",X"00",X"FD",X"19",X"11",X"07",X"00",X"06",X"0C",X"FD",X"7E",X"00",X"FE",X"A0",
		X"38",X"32",X"FE",X"B8",X"30",X"2E",X"FD",X"7E",X"01",X"DD",X"96",X"01",X"30",X"02",X"ED",X"44",
		X"FE",X"0E",X"30",X"20",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"38",X"18",X"E6",X"F0",X"28",X"1C",
		X"0F",X"0F",X"0F",X"0F",X"4F",X"E5",X"7E",X"E6",X"0F",X"28",X"08",X"23",X"23",X"0D",X"20",X"F6",
		X"E1",X"18",X"09",X"E1",X"FD",X"19",X"10",X"C3",X"FD",X"E1",X"18",X"05",X"FD",X"E1",X"3E",X"07",
		X"C9",X"3A",X"D7",X"E1",X"E6",X"88",X"28",X"35",X"FE",X"80",X"28",X"07",X"3A",X"DD",X"E1",X"FE",
		X"20",X"30",X"2A",X"3A",X"D8",X"E1",X"DD",X"96",X"01",X"FE",X"20",X"38",X"08",X"FE",X"E0",X"38",
		X"1C",X"06",X"04",X"18",X"02",X"06",X"01",X"3A",X"DA",X"E1",X"DD",X"96",X"03",X"FE",X"20",X"38",
		X"08",X"FE",X"E0",X"38",X"08",X"78",X"F6",X"08",X"C9",X"78",X"F6",X"02",X"C9",X"AF",X"C9",X"F5",
		X"CD",X"A3",X"1D",X"F1",X"A6",X"C8",X"CB",X"57",X"20",X"0C",X"CB",X"47",X"20",X"0E",X"CB",X"4F",
		X"20",X"07",X"B7",X"3E",X"02",X"C9",X"3E",X"00",X"C9",X"3E",X"03",X"C9",X"3E",X"01",X"C9",X"DD",
		X"CB",X"07",X"66",X"20",X"0E",X"CD",X"A3",X"1D",X"23",X"7E",X"FE",X"08",X"D0",X"87",X"87",X"87",
		X"87",X"18",X"19",X"3A",X"C6",X"E1",X"DD",X"96",X"01",X"30",X"02",X"ED",X"44",X"47",X"3A",X"C8",
		X"E1",X"DD",X"96",X"03",X"30",X"02",X"ED",X"44",X"B8",X"30",X"01",X"78",X"21",X"19",X"E2",X"BE",
		X"D0",X"77",X"C9",X"DD",X"7E",X"00",X"CB",X"77",X"20",X"3E",X"DD",X"36",X"00",X"C0",X"DD",X"36",
		X"02",X"00",X"DD",X"36",X"03",X"F1",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",
		X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"DD",X"36",
		X"0A",X"00",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",
		X"0E",X"00",X"FD",X"CB",X"1B",X"8E",X"18",X"4B",X"DD",X"CB",X"00",X"6E",X"C2",X"4C",X"44",X"3A",
		X"00",X"E0",X"E6",X"40",X"20",X"05",X"DD",X"36",X"00",X"00",X"C9",X"3A",X"B6",X"E1",X"A7",X"C2",
		X"E0",X"44",X"FD",X"CB",X"1B",X"46",X"28",X"06",X"FD",X"CB",X"1B",X"86",X"18",X"52",X"CD",X"61",
		X"48",X"C2",X"E0",X"44",X"FD",X"CB",X"16",X"4E",X"20",X"10",X"FD",X"34",X"17",X"FD",X"7E",X"17",
		X"FE",X"04",X"38",X"0F",X"FD",X"CB",X"16",X"CE",X"18",X"09",X"FD",X"35",X"17",X"20",X"04",X"FD",
		X"CB",X"16",X"8E",X"21",X"AA",X"47",X"3A",X"00",X"E0",X"87",X"30",X"0A",X"3A",X"02",X"A0",X"E6",
		X"10",X"20",X"03",X"21",X"AE",X"47",X"CD",X"CD",X"47",X"17",X"30",X"02",X"23",X"23",X"7E",X"DD",
		X"77",X"10",X"23",X"7E",X"DD",X"77",X"0F",X"CD",X"C2",X"47",X"DD",X"77",X"01",X"C3",X"E0",X"44",
		X"DD",X"36",X"00",X"E3",X"DD",X"36",X"05",X"00",X"FD",X"7E",X"1A",X"FE",X"04",X"38",X"02",X"3E",
		X"03",X"87",X"5F",X"16",X"00",X"21",X"B2",X"47",X"3A",X"02",X"A0",X"E6",X"10",X"20",X"03",X"21",
		X"BA",X"47",X"19",X"7E",X"DD",X"77",X"10",X"23",X"7E",X"DD",X"77",X"0F",X"CD",X"DB",X"47",X"21",
		X"01",X"E0",X"CB",X"E6",X"3E",X"17",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"FD",X"46",X"14",X"FD",
		X"4E",X"15",X"78",X"B1",X"28",X"07",X"0B",X"FD",X"70",X"14",X"FD",X"71",X"15",X"FD",X"CB",X"1B",
		X"86",X"DD",X"7E",X"00",X"CB",X"57",X"C2",X"72",X"47",X"CB",X"5F",X"C2",X"20",X"47",X"E6",X"10",
		X"C2",X"FC",X"46",X"DD",X"CB",X"07",X"6E",X"C2",X"C1",X"46",X"CD",X"DB",X"47",X"3A",X"00",X"E0",
		X"E6",X"40",X"20",X"08",X"DD",X"36",X"00",X"00",X"CD",X"4F",X"05",X"C9",X"21",X"DD",X"44",X"E5",
		X"DD",X"CB",X"07",X"56",X"C2",X"B5",X"46",X"3A",X"B6",X"E1",X"A7",X"C0",X"3A",X"C5",X"E1",X"E6",
		X"98",X"FE",X"80",X"C0",X"FD",X"E5",X"FD",X"21",X"C5",X"E1",X"01",X"07",X"07",X"CD",X"D7",X"05",
		X"30",X"0F",X"FD",X"CB",X"00",X"DE",X"DD",X"CB",X"07",X"D6",X"DD",X"36",X"06",X"1E",X"FD",X"E1",
		X"C9",X"FD",X"E1",X"DD",X"7E",X"05",X"FE",X"40",X"D2",X"83",X"46",X"FE",X"30",X"D2",X"47",X"46",
		X"FE",X"20",X"D2",X"D2",X"45",X"FE",X"10",X"D2",X"46",X"45",X"C3",X"01",X"45",X"DD",X"34",X"08",
		X"DD",X"7E",X"08",X"FE",X"18",X"38",X"04",X"AF",X"DD",X"77",X"08",X"E6",X"18",X"0F",X"0F",X"0F",
		X"4F",X"FD",X"7E",X"17",X"47",X"87",X"80",X"81",X"C6",X"4D",X"47",X"0E",X"04",X"CD",X"97",X"02",
		X"C9",X"DD",X"7E",X"0D",X"A7",X"28",X"04",X"DD",X"35",X"0D",X"C9",X"DD",X"7E",X"05",X"E6",X"0F",
		X"20",X"06",X"CD",X"A5",X"49",X"DD",X"34",X"05",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"11",X"2B",
		X"FF",X"19",X"DD",X"74",X"03",X"DD",X"75",X"04",X"7C",X"FE",X"E1",X"D0",X"3A",X"01",X"E0",X"E6",
		X"40",X"20",X"06",X"DD",X"36",X"05",X"10",X"18",X"04",X"DD",X"36",X"05",X"20",X"DD",X"7E",X"0C",
		X"F6",X"E0",X"DD",X"77",X"00",X"C9",X"CD",X"61",X"48",X"20",X"0C",X"3A",X"01",X"E0",X"E6",X"40",
		X"20",X"05",X"DD",X"36",X"05",X"30",X"C9",X"CD",X"F2",X"48",X"D8",X"3A",X"CC",X"E1",X"87",X"30",
		X"4F",X"CD",X"C1",X"3D",X"20",X"42",X"DD",X"CB",X"07",X"7E",X"20",X"40",X"DD",X"CB",X"07",X"76",
		X"20",X"1C",X"CD",X"7C",X"3E",X"FE",X"04",X"D0",X"DD",X"4E",X"00",X"CD",X"D7",X"3E",X"A9",X"E6",
		X"03",X"FE",X"01",X"20",X"27",X"DD",X"CB",X"07",X"F6",X"DD",X"CB",X"07",X"BE",X"C9",X"CD",X"E6",
		X"3E",X"FE",X"04",X"30",X"08",X"CD",X"D7",X"3E",X"FD",X"CB",X"07",X"B6",X"C9",X"CD",X"D6",X"3D",
		X"FE",X"04",X"D0",X"CD",X"D7",X"3E",X"18",X"04",X"DD",X"CB",X"07",X"BE",X"CD",X"3F",X"49",X"C9",
		X"DD",X"CB",X"07",X"B6",X"CD",X"C1",X"3D",X"20",X"11",X"DD",X"CB",X"07",X"7E",X"20",X"0F",X"CD",
		X"D6",X"3D",X"FE",X"04",X"D0",X"CD",X"D7",X"3E",X"18",X"04",X"DD",X"CB",X"07",X"BE",X"CD",X"3F",
		X"49",X"C9",X"DD",X"7E",X"0E",X"FE",X"02",X"30",X"05",X"DD",X"36",X"05",X"10",X"C9",X"CD",X"61",
		X"48",X"CD",X"F2",X"48",X"D8",X"DD",X"7E",X"0D",X"A7",X"28",X"04",X"DD",X"35",X"0D",X"C9",X"FD",
		X"E5",X"FD",X"21",X"D3",X"E2",X"11",X"0F",X"00",X"06",X"03",X"D9",X"01",X"0E",X"0E",X"D9",X"FD",
		X"7E",X"00",X"E6",X"BC",X"FE",X"80",X"20",X"0E",X"D9",X"CD",X"D7",X"05",X"D9",X"30",X"07",X"FD",
		X"E1",X"DD",X"36",X"0D",X"1E",X"C9",X"FD",X"19",X"10",X"E5",X"FD",X"E1",X"CD",X"C1",X"3D",X"20",
		X"1E",X"DD",X"CB",X"07",X"7E",X"20",X"1C",X"CD",X"D6",X"3D",X"FE",X"04",X"D0",X"DD",X"4E",X"00",
		X"CD",X"D7",X"3E",X"A9",X"E6",X"03",X"FE",X"01",X"20",X"09",X"DD",X"36",X"0D",X"1E",X"C9",X"DD",
		X"CB",X"07",X"BE",X"CD",X"3F",X"49",X"C9",X"DD",X"7E",X"03",X"FE",X"DF",X"38",X"13",X"CD",X"C2",
		X"47",X"DD",X"BE",X"01",X"28",X"06",X"3D",X"DD",X"BE",X"01",X"20",X"05",X"DD",X"36",X"05",X"40",
		X"C9",X"CD",X"F2",X"48",X"D8",X"CD",X"C1",X"3D",X"20",X"11",X"DD",X"CB",X"07",X"7E",X"20",X"0F",
		X"CD",X"72",X"48",X"FE",X"04",X"D0",X"CD",X"D7",X"3E",X"18",X"04",X"DD",X"CB",X"07",X"BE",X"CD",
		X"3F",X"49",X"C9",X"DD",X"7E",X"05",X"E6",X"0F",X"20",X"07",X"DD",X"34",X"05",X"DD",X"36",X"00",
		X"E2",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"11",X"D5",X"00",X"19",X"DD",X"74",X"03",X"DD",X"75",
		X"04",X"7C",X"FE",X"F0",X"D8",X"CD",X"4F",X"05",X"CD",X"97",X"4D",X"3E",X"17",X"CD",X"EA",X"02",
		X"DD",X"36",X"00",X"80",X"C9",X"DD",X"35",X"06",X"C0",X"DD",X"36",X"00",X"00",X"CD",X"4F",X"05",
		X"C9",X"CD",X"D3",X"49",X"DD",X"7E",X"0A",X"FE",X"20",X"30",X"1C",X"06",X"2B",X"0E",X"04",X"DD",
		X"7E",X"00",X"CB",X"4F",X"20",X"08",X"E6",X"01",X"28",X"1E",X"CB",X"E9",X"18",X"1A",X"04",X"E6",
		X"01",X"28",X"15",X"CB",X"E1",X"18",X"11",X"06",X"49",X"0E",X"04",X"DD",X"7E",X"0B",X"D6",X"08",
		X"38",X"06",X"04",X"E6",X"08",X"28",X"01",X"04",X"CD",X"97",X"02",X"C9",X"DD",X"CB",X"07",X"4E",
		X"20",X"11",X"DD",X"CB",X"07",X"CE",X"CD",X"77",X"47",X"CD",X"97",X"4D",X"CD",X"AE",X"4D",X"DD",
		X"36",X"06",X"00",X"DD",X"35",X"06",X"28",X"5A",X"06",X"5C",X"0E",X"04",X"CD",X"97",X"02",X"C9",
		X"DD",X"CB",X"07",X"46",X"20",X"21",X"DD",X"CB",X"07",X"C6",X"DD",X"36",X"06",X"FF",X"CD",X"77",
		X"47",X"11",X"5A",X"3B",X"CD",X"2A",X"03",X"CD",X"97",X"4D",X"DD",X"CB",X"07",X"6E",X"28",X"07",
		X"DD",X"7E",X"0A",X"FE",X"10",X"28",X"28",X"DD",X"34",X"06",X"DD",X"7E",X"06",X"FE",X"26",X"30",
		X"21",X"FE",X"08",X"28",X"0F",X"30",X"10",X"06",X"67",X"0E",X"05",X"FE",X"04",X"30",X"01",X"04",
		X"CD",X"97",X"02",X"C9",X"CD",X"C6",X"4D",X"06",X"71",X"0E",X"0A",X"CD",X"97",X"02",X"C9",X"CD",
		X"AE",X"4D",X"DD",X"36",X"00",X"80",X"C9",X"FD",X"46",X"17",X"78",X"A7",X"3E",X"80",X"28",X"03",
		X"0F",X"10",X"FD",X"FD",X"B6",X"16",X"FD",X"77",X"16",X"CD",X"4F",X"05",X"3E",X"17",X"CD",X"EA",
		X"02",X"FD",X"7E",X"16",X"E6",X"F8",X"FE",X"F8",X"C0",X"3A",X"00",X"E0",X"87",X"D0",X"21",X"B6",
		X"E1",X"CB",X"FE",X"CB",X"DE",X"FD",X"36",X"30",X"04",X"C9",X"2C",X"01",X"3C",X"00",X"F0",X"00",
		X"78",X"00",X"B0",X"04",X"84",X"03",X"58",X"02",X"2C",X"01",X"C0",X"03",X"E0",X"01",X"F0",X"00",
		X"F0",X"00",X"FD",X"7E",X"17",X"87",X"87",X"47",X"87",X"80",X"C6",X"68",X"C9",X"FD",X"4E",X"16",
		X"FD",X"7E",X"17",X"47",X"A7",X"79",X"C8",X"87",X"10",X"FD",X"C9",X"FD",X"CB",X"1B",X"4E",X"C8",
		X"FD",X"CB",X"1B",X"8E",X"21",X"01",X"E0",X"CB",X"F6",X"3E",X"3C",X"CD",X"BE",X"06",X"DD",X"7E",
		X"05",X"A7",X"28",X"04",X"FE",X"40",X"38",X"0E",X"DD",X"36",X"05",X"00",X"CD",X"F4",X"02",X"E6",
		X"01",X"DD",X"77",X"0C",X"18",X"04",X"DD",X"36",X"05",X"20",X"DD",X"7E",X"00",X"E6",X"03",X"F6",
		X"80",X"47",X"DD",X"4E",X"01",X"DD",X"56",X"03",X"DD",X"5E",X"05",X"DD",X"66",X"0C",X"3E",X"1E",
		X"FD",X"E5",X"FD",X"21",X"D3",X"E2",X"D9",X"11",X"0F",X"00",X"D9",X"FD",X"70",X"00",X"FD",X"71",
		X"01",X"FD",X"36",X"02",X"00",X"FD",X"72",X"03",X"FD",X"36",X"04",X"00",X"FD",X"73",X"05",X"FD",
		X"74",X"0C",X"FD",X"77",X"0D",X"D9",X"FD",X"19",X"D9",X"C6",X"1E",X"FE",X"78",X"38",X"DC",X"FD",
		X"E1",X"DD",X"77",X"0D",X"DD",X"36",X"0E",X"03",X"FD",X"36",X"14",X"02",X"FD",X"36",X"15",X"D0",
		X"C9",X"DD",X"46",X"0F",X"DD",X"4E",X"10",X"78",X"B1",X"C8",X"0B",X"DD",X"70",X"0F",X"DD",X"71",
		X"10",X"C9",X"DD",X"7E",X"03",X"FE",X"DF",X"38",X"17",X"DD",X"7E",X"01",X"FE",X"67",X"38",X"10",
		X"FE",X"99",X"30",X"0C",X"4F",X"CD",X"C2",X"47",X"B9",X"38",X"02",X"AF",X"C9",X"3E",X"01",X"C9",
		X"CD",X"A3",X"1D",X"46",X"CB",X"68",X"CA",X"D6",X"3D",X"23",X"4E",X"CB",X"58",X"28",X"10",X"23",
		X"56",X"23",X"7E",X"2B",X"2B",X"CB",X"6A",X"28",X"06",X"B9",X"38",X"03",X"3E",X"02",X"C9",X"CB",
		X"50",X"28",X"11",X"EB",X"21",X"20",X"00",X"19",X"7E",X"2B",X"CB",X"6E",X"EB",X"28",X"05",X"B9",
		X"38",X"02",X"AF",X"C9",X"CB",X"48",X"28",X"11",X"2B",X"2B",X"7E",X"2B",X"CB",X"6E",X"23",X"23",
		X"23",X"28",X"06",X"B9",X"38",X"03",X"3E",X"03",X"C9",X"CB",X"40",X"28",X"12",X"EB",X"21",X"E0",
		X"FF",X"19",X"7E",X"2B",X"CB",X"6E",X"EB",X"28",X"06",X"B9",X"38",X"03",X"3E",X"01",X"C9",X"3E",
		X"04",X"C9",X"CD",X"41",X"40",X"FD",X"E5",X"D9",X"11",X"31",X"00",X"FD",X"19",X"06",X"0C",X"11",
		X"07",X"00",X"FD",X"7E",X"00",X"FE",X"80",X"38",X"17",X"FE",X"B8",X"30",X"13",X"E6",X"F8",X"FE",
		X"A8",X"28",X"0D",X"D9",X"FD",X"66",X"01",X"FD",X"6E",X"03",X"CD",X"EF",X"05",X"38",X"09",X"D9",
		X"FD",X"19",X"10",X"DE",X"FD",X"E1",X"A7",X"C9",X"DD",X"CB",X"07",X"EE",X"D9",X"DD",X"70",X"09",
		X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"0C",X"00",X"FD",X"E1",X"C9",X"01",
		X"D5",X"00",X"3A",X"01",X"E0",X"E6",X"40",X"28",X"20",X"01",X"B3",X"00",X"FD",X"7E",X"14",X"FD",
		X"B6",X"15",X"20",X"03",X"01",X"DE",X"00",X"FD",X"7E",X"08",X"FE",X"10",X"38",X"02",X"3E",X"0F",
		X"87",X"87",X"87",X"6F",X"26",X"00",X"09",X"44",X"4D",X"DD",X"CB",X"00",X"46",X"C4",X"E3",X"2C",
		X"DD",X"CB",X"00",X"4E",X"20",X"17",X"DD",X"66",X"01",X"DD",X"6E",X"02",X"09",X"DD",X"74",X"01",
		X"DD",X"75",X"02",X"DD",X"7E",X"03",X"3C",X"E6",X"F0",X"DD",X"77",X"03",X"C9",X"DD",X"66",X"03",
		X"DD",X"6E",X"04",X"09",X"DD",X"74",X"03",X"DD",X"75",X"04",X"DD",X"7E",X"01",X"E6",X"F0",X"C6",
		X"08",X"DD",X"77",X"01",X"C9",X"FD",X"7E",X"17",X"87",X"87",X"5F",X"16",X"00",X"21",X"BF",X"49",
		X"19",X"5E",X"23",X"56",X"23",X"46",X"23",X"4E",X"EB",X"3E",X"25",X"CD",X"5C",X"04",X"C9",X"9D",
		X"89",X"02",X"02",X"DD",X"89",X"02",X"01",X"FD",X"89",X"02",X"02",X"3D",X"8A",X"02",X"01",X"5D",
		X"8A",X"02",X"02",X"DD",X"7E",X"0A",X"FE",X"20",X"D2",X"DF",X"4A",X"FE",X"10",X"D2",X"8D",X"4A",
		X"FD",X"E5",X"CD",X"03",X"4B",X"FD",X"7E",X"00",X"FE",X"80",X"DA",X"82",X"4A",X"FE",X"B8",X"D2",
		X"82",X"4A",X"E6",X"F8",X"FE",X"A8",X"CA",X"82",X"4A",X"01",X"0E",X"0E",X"CD",X"D7",X"05",X"D2",
		X"82",X"4A",X"FD",X"7E",X"01",X"DD",X"96",X"01",X"38",X"04",X"FE",X"02",X"38",X"12",X"FD",X"7E",
		X"03",X"DD",X"96",X"03",X"38",X"04",X"FE",X"02",X"38",X"16",X"FD",X"E1",X"CD",X"3F",X"49",X"C9",
		X"FD",X"7E",X"03",X"DD",X"96",X"03",X"38",X"04",X"06",X"02",X"18",X"12",X"06",X"03",X"18",X"0E",
		X"FD",X"7E",X"01",X"DD",X"96",X"01",X"38",X"04",X"06",X"00",X"18",X"02",X"06",X"01",X"FD",X"7E",
		X"00",X"FD",X"36",X"00",X"D0",X"FD",X"36",X"06",X"00",X"FE",X"B0",X"28",X"04",X"FD",X"36",X"05",
		X"00",X"FD",X"E1",X"DD",X"36",X"0A",X"10",X"DD",X"7E",X"00",X"E6",X"03",X"B8",X"C8",X"DD",X"7E",
		X"00",X"E6",X"FC",X"B0",X"DD",X"77",X"00",X"78",X"EE",X"01",X"F6",X"80",X"DD",X"77",X"0C",X"C9",
		X"FD",X"36",X"00",X"00",X"FD",X"E1",X"DD",X"36",X"0A",X"20",X"3E",X"15",X"06",X"00",X"CD",X"D9",
		X"02",X"C9",X"FD",X"E1",X"DD",X"CB",X"07",X"AE",X"DD",X"CB",X"07",X"BE",X"C9",X"CD",X"C1",X"3D",
		X"20",X"13",X"CD",X"D6",X"3D",X"47",X"DD",X"7E",X"00",X"E6",X"03",X"B8",X"28",X"07",X"EE",X"01",
		X"F6",X"80",X"DD",X"77",X"0C",X"FD",X"E5",X"CD",X"03",X"4B",X"FD",X"7E",X"00",X"FE",X"D0",X"20",
		X"2A",X"FD",X"7E",X"01",X"DD",X"96",X"01",X"38",X"10",X"FE",X"02",X"30",X"0C",X"FD",X"7E",X"03",
		X"DD",X"96",X"03",X"38",X"04",X"FE",X"02",X"38",X"A7",X"01",X"0F",X"0F",X"CD",X"D7",X"05",X"30",
		X"06",X"FD",X"E1",X"CD",X"3F",X"49",X"C9",X"FD",X"36",X"00",X"88",X"FD",X"E1",X"18",X"09",X"DD",
		X"34",X"0B",X"DD",X"7E",X"0B",X"FE",X"40",X"D8",X"DD",X"CB",X"07",X"AE",X"DD",X"CB",X"07",X"BE",
		X"DD",X"7E",X"0C",X"CB",X"7F",X"C8",X"E6",X"03",X"47",X"DD",X"7E",X"00",X"E6",X"FC",X"B0",X"DD",
		X"77",X"00",X"C9",X"3E",X"0C",X"DD",X"96",X"09",X"4F",X"87",X"87",X"87",X"91",X"5F",X"16",X"00",
		X"21",X"31",X"00",X"19",X"EB",X"FD",X"19",X"C9",X"DD",X"CB",X"00",X"76",X"20",X"1C",X"DD",X"CB",
		X"00",X"F6",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",
		X"09",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"00",X"DD",X"7E",X"00",X"CB",X"57",X"C2",
		X"47",X"4D",X"CB",X"5F",X"C2",X"F8",X"4C",X"CB",X"6F",X"C2",X"4C",X"4D",X"E6",X"10",X"C2",X"D7",
		X"4C",X"DD",X"CB",X"07",X"6E",X"C2",X"92",X"4C",X"3A",X"00",X"E0",X"E6",X"40",X"20",X"05",X"DD",
		X"36",X"00",X"00",X"C9",X"21",X"CB",X"4B",X"E5",X"DD",X"CB",X"07",X"56",X"C2",X"89",X"4C",X"3A",
		X"01",X"E0",X"E6",X"40",X"20",X"05",X"DD",X"CB",X"00",X"EE",X"C9",X"3A",X"B6",X"E1",X"A7",X"C0",
		X"3A",X"C5",X"E1",X"E6",X"98",X"FE",X"80",X"C0",X"FD",X"E5",X"FD",X"21",X"C5",X"E1",X"01",X"07",
		X"07",X"CD",X"D7",X"05",X"30",X"0F",X"FD",X"CB",X"00",X"DE",X"DD",X"CB",X"07",X"D6",X"DD",X"36",
		X"06",X"1E",X"FD",X"E1",X"C9",X"FD",X"E1",X"DD",X"7E",X"0D",X"A7",X"28",X"14",X"DD",X"35",X"0D",
		X"C0",X"21",X"C9",X"E2",X"CB",X"66",X"C0",X"CB",X"E6",X"3E",X"11",X"06",X"00",X"CD",X"D9",X"02",
		X"C9",X"DD",X"7E",X"05",X"A7",X"C2",X"15",X"4C",X"C3",X"F4",X"4B",X"DD",X"34",X"08",X"06",X"27",
		X"0E",X"02",X"DD",X"7E",X"00",X"CB",X"4F",X"20",X"08",X"E6",X"01",X"28",X"0C",X"CB",X"E9",X"18",
		X"08",X"06",X"29",X"E6",X"01",X"28",X"02",X"CB",X"E1",X"DD",X"CB",X"08",X"5E",X"28",X"01",X"04",
		X"CD",X"97",X"02",X"C9",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"11",X"2B",X"FF",X"19",X"DD",X"74",
		X"03",X"DD",X"75",X"04",X"7C",X"FE",X"E1",X"D0",X"DD",X"36",X"05",X"10",X"DD",X"7E",X"0C",X"F6",
		X"C0",X"DD",X"77",X"00",X"C9",X"CD",X"F2",X"48",X"D8",X"CD",X"C1",X"3D",X"20",X"16",X"DD",X"CB",
		X"07",X"7E",X"20",X"14",X"CD",X"D6",X"3D",X"FE",X"04",X"30",X"11",X"DD",X"36",X"0E",X"00",X"CD",
		X"D7",X"3E",X"18",X"04",X"DD",X"CB",X"07",X"BE",X"CD",X"3F",X"49",X"C9",X"DD",X"7E",X"0E",X"A7",
		X"20",X"05",X"DD",X"36",X"0E",X"1E",X"C9",X"DD",X"35",X"0E",X"C0",X"3A",X"C6",X"E1",X"DD",X"96",
		X"01",X"FE",X"12",X"38",X"03",X"FE",X"EF",X"D8",X"47",X"3A",X"C8",X"E1",X"DD",X"96",X"03",X"FE",
		X"12",X"38",X"03",X"FE",X"EF",X"D8",X"B8",X"38",X"10",X"E6",X"80",X"20",X"06",X"3E",X"02",X"CD",
		X"D7",X"3E",X"C9",X"3E",X"03",X"CD",X"D7",X"3E",X"C9",X"CB",X"78",X"20",X"06",X"3E",X"00",X"CD",
		X"D7",X"3E",X"C9",X"3E",X"01",X"CD",X"D7",X"3E",X"C9",X"DD",X"35",X"06",X"C0",X"DD",X"36",X"00",
		X"00",X"C9",X"CD",X"D3",X"49",X"DD",X"7E",X"0A",X"FE",X"20",X"30",X"1C",X"06",X"2B",X"0E",X"04",
		X"DD",X"7E",X"00",X"CB",X"4F",X"20",X"08",X"E6",X"01",X"28",X"1E",X"CB",X"E9",X"18",X"1A",X"04",
		X"E6",X"01",X"28",X"15",X"CB",X"E1",X"18",X"11",X"06",X"49",X"0E",X"04",X"DD",X"7E",X"0B",X"D6",
		X"08",X"38",X"06",X"04",X"E6",X"08",X"28",X"01",X"04",X"CD",X"97",X"02",X"3A",X"01",X"E0",X"E6",
		X"40",X"C0",X"DD",X"CB",X"00",X"EE",X"C9",X"DD",X"CB",X"07",X"4E",X"20",X"0E",X"DD",X"CB",X"07",
		X"CE",X"CD",X"8D",X"4D",X"CD",X"AE",X"4D",X"DD",X"36",X"06",X"00",X"DD",X"35",X"06",X"28",X"57",
		X"06",X"4C",X"0E",X"02",X"CD",X"97",X"02",X"C9",X"DD",X"CB",X"07",X"46",X"20",X"1E",X"DD",X"CB",
		X"07",X"C6",X"DD",X"36",X"06",X"FF",X"CD",X"8D",X"4D",X"11",X"5A",X"3B",X"CD",X"2A",X"03",X"DD",
		X"CB",X"07",X"6E",X"28",X"07",X"DD",X"7E",X"0A",X"FE",X"10",X"28",X"28",X"DD",X"34",X"06",X"DD",
		X"7E",X"06",X"FE",X"26",X"30",X"21",X"FE",X"08",X"28",X"0F",X"30",X"10",X"06",X"67",X"0E",X"05",
		X"FE",X"04",X"38",X"01",X"04",X"CD",X"97",X"02",X"C9",X"CD",X"C6",X"4D",X"06",X"71",X"0E",X"0A",
		X"CD",X"97",X"02",X"C9",X"CD",X"AE",X"4D",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"CB",X"07",X"5E",
		X"20",X"0B",X"DD",X"CB",X"07",X"DE",X"DD",X"36",X"06",X"FF",X"CD",X"8D",X"4D",X"DD",X"34",X"06",
		X"DD",X"7E",X"06",X"D6",X"20",X"DA",X"CB",X"4B",X"FE",X"20",X"30",X"0D",X"06",X"67",X"0E",X"05",
		X"FE",X"10",X"38",X"01",X"04",X"CD",X"97",X"02",X"C9",X"DD",X"CB",X"07",X"6E",X"28",X"09",X"DD",
		X"7E",X"0A",X"FE",X"10",X"20",X"02",X"18",X"BC",X"CD",X"C6",X"4D",X"18",X"BA",X"21",X"D0",X"E2",
		X"35",X"C0",X"3E",X"11",X"CD",X"EA",X"02",X"21",X"00",X"E0",X"CB",X"76",X"C8",X"23",X"CB",X"76",
		X"C8",X"CB",X"B6",X"CB",X"EE",X"3E",X"40",X"32",X"05",X"E0",X"CD",X"A1",X"06",X"C9",X"DD",X"CB",
		X"07",X"6E",X"C8",X"FD",X"E5",X"CD",X"03",X"4B",X"FD",X"7E",X"00",X"FE",X"D0",X"20",X"04",X"FD",
		X"36",X"00",X"88",X"FD",X"E1",X"C9",X"FD",X"E5",X"11",X"31",X"00",X"FD",X"19",X"11",X"07",X"00",
		X"06",X"0C",X"FD",X"7E",X"00",X"A7",X"28",X"07",X"FD",X"19",X"10",X"F6",X"FD",X"E1",X"C9",X"FD",
		X"36",X"00",X"88",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"DD",X"7E",X"03",
		X"FD",X"77",X"03",X"FD",X"36",X"04",X"00",X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",X"00",X"FD",
		X"E1",X"C9",X"3A",X"00",X"E0",X"E6",X"40",X"20",X"04",X"DD",X"36",X"00",X"00",X"FD",X"E5",X"DD",
		X"E1",X"11",X"31",X"00",X"DD",X"19",X"11",X"07",X"00",X"06",X"0C",X"DD",X"CB",X"00",X"7E",X"28",
		X"07",X"C5",X"D5",X"CD",X"2D",X"4E",X"D1",X"C1",X"DD",X"19",X"10",X"EF",X"C9",X"21",X"44",X"4E",
		X"E5",X"DD",X"7E",X"00",X"E6",X"78",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"4C",X"4E",X"19",X"5E",
		X"23",X"56",X"EB",X"E9",X"06",X"5E",X"0E",X"05",X"CD",X"97",X"02",X"C9",X"62",X"4E",X"63",X"4E",
		X"98",X"4E",X"98",X"4E",X"B6",X"4E",X"08",X"4F",X"68",X"4F",X"10",X"50",X"3D",X"50",X"85",X"50",
		X"FA",X"50",X"C9",X"3A",X"C5",X"E1",X"87",X"30",X"1A",X"3A",X"C8",X"E1",X"DD",X"96",X"03",X"FE",
		X"ED",X"38",X"10",X"FE",X"F4",X"30",X"0C",X"3A",X"C6",X"E1",X"DD",X"96",X"01",X"FE",X"09",X"D8",
		X"FE",X"F8",X"D0",X"CD",X"A9",X"53",X"DD",X"7E",X"00",X"FE",X"88",X"D8",X"DD",X"77",X"05",X"DD",
		X"36",X"00",X"A0",X"DD",X"36",X"06",X"0A",X"C9",X"DD",X"46",X"00",X"C5",X"CD",X"A9",X"53",X"C1",
		X"DD",X"7E",X"00",X"FE",X"80",X"20",X"08",X"78",X"FE",X"98",X"C0",X"DD",X"77",X"00",X"C9",X"FE",
		X"B0",X"20",X"43",X"C3",X"52",X"4F",X"21",X"00",X"E3",X"CB",X"FE",X"DD",X"35",X"06",X"20",X"17",
		X"DD",X"34",X"00",X"DD",X"7E",X"00",X"E6",X"07",X"FE",X"04",X"28",X"20",X"DD",X"36",X"06",X"05",
		X"0F",X"38",X"04",X"DD",X"36",X"06",X"0A",X"DD",X"7E",X"00",X"E6",X"03",X"CB",X"47",X"28",X"02",
		X"E6",X"01",X"C6",X"5D",X"47",X"0E",X"05",X"CD",X"97",X"02",X"E1",X"C9",X"DD",X"7E",X"05",X"FE",
		X"B0",X"28",X"5F",X"DD",X"77",X"00",X"DD",X"36",X"05",X"00",X"1F",X"DD",X"7E",X"01",X"38",X"02",
		X"C6",X"08",X"E6",X"F8",X"DD",X"77",X"06",X"C9",X"21",X"00",X"E3",X"CB",X"FE",X"DD",X"7E",X"01",
		X"DD",X"BE",X"06",X"28",X"3A",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"21",X"95",X"FF",X"19",X"DD",
		X"74",X"03",X"DD",X"75",X"04",X"DD",X"56",X"01",X"DD",X"5E",X"02",X"21",X"B9",X"00",X"DD",X"CB",
		X"00",X"46",X"28",X"03",X"21",X"47",X"FF",X"19",X"DD",X"74",X"01",X"DD",X"75",X"02",X"06",X"5D",
		X"0E",X"05",X"DD",X"CB",X"00",X"46",X"28",X"02",X"06",X"5F",X"CD",X"97",X"02",X"E1",X"C9",X"CD",
		X"EF",X"51",X"DD",X"36",X"00",X"B0",X"DD",X"36",X"05",X"00",X"DD",X"7E",X"03",X"DD",X"77",X"06",
		X"3E",X"12",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"21",X"00",X"E3",X"CB",X"FE",X"FD",X"E5",X"11",
		X"31",X"00",X"FD",X"19",X"11",X"07",X"00",X"06",X"0C",X"D9",X"01",X"0E",X"0E",X"D9",X"FD",X"7E",
		X"00",X"FE",X"80",X"38",X"2B",X"FE",X"D0",X"28",X"04",X"FE",X"B0",X"30",X"23",X"D9",X"CD",X"D7",
		X"05",X"D9",X"30",X"1C",X"FD",X"36",X"00",X"C0",X"FD",X"E1",X"3E",X"12",X"CD",X"EA",X"02",X"DD",
		X"7E",X"05",X"E6",X"3F",X"20",X"05",X"DD",X"36",X"00",X"C0",X"C9",X"DD",X"36",X"00",X"B8",X"C9",
		X"FD",X"19",X"10",X"CA",X"FD",X"E1",X"CD",X"A9",X"53",X"DD",X"7E",X"00",X"FE",X"B0",X"20",X"1E",
		X"DD",X"7E",X"03",X"FE",X"21",X"38",X"17",X"CD",X"DF",X"51",X"CD",X"BE",X"52",X"DD",X"56",X"03",
		X"DD",X"5E",X"04",X"21",X"AB",X"FE",X"19",X"DD",X"74",X"03",X"DD",X"75",X"04",X"C9",X"DD",X"7E",
		X"03",X"3C",X"E6",X"F8",X"DD",X"77",X"03",X"DD",X"CB",X"05",X"BE",X"3E",X"12",X"CD",X"EA",X"02",
		X"DD",X"7E",X"05",X"E6",X"3F",X"20",X"B4",X"DD",X"7E",X"06",X"DD",X"46",X"03",X"90",X"FE",X"11",
		X"30",X"A4",X"78",X"FE",X"21",X"38",X"9F",X"DD",X"7E",X"00",X"FE",X"80",X"C2",X"F6",X"4E",X"C9",
		X"21",X"00",X"E3",X"CB",X"FE",X"DD",X"7E",X"00",X"E6",X"07",X"20",X"15",X"DD",X"34",X"00",X"DD",
		X"36",X"06",X"1E",X"DD",X"7E",X"05",X"E6",X"2F",X"28",X"07",X"3E",X"1A",X"06",X"00",X"CD",X"D9",
		X"02",X"DD",X"35",X"06",X"C0",X"DD",X"36",X"00",X"C8",X"CD",X"2A",X"51",X"C9",X"21",X"00",X"E3",
		X"CB",X"FE",X"DD",X"7E",X"00",X"E6",X"07",X"20",X"0E",X"DD",X"34",X"00",X"DD",X"36",X"06",X"00",
		X"3E",X"13",X"06",X"00",X"CD",X"D9",X"02",X"DD",X"34",X"06",X"DD",X"7E",X"06",X"E6",X"18",X"FE",
		X"18",X"CA",X"C4",X"50",X"0F",X"0F",X"C6",X"60",X"47",X"0E",X"05",X"DD",X"7E",X"01",X"D6",X"08",
		X"57",X"DD",X"5E",X"03",X"C5",X"D5",X"CD",X"9D",X"02",X"D1",X"C1",X"04",X"7A",X"C6",X"10",X"57",
		X"CD",X"9D",X"02",X"E1",X"C9",X"21",X"00",X"E3",X"CB",X"FE",X"DD",X"7E",X"00",X"E6",X"07",X"20",
		X"1C",X"DD",X"34",X"00",X"DD",X"36",X"06",X"1E",X"DD",X"7E",X"05",X"E6",X"0F",X"28",X"18",X"CD",
		X"91",X"51",X"DD",X"CB",X"05",X"66",X"28",X"05",X"21",X"C5",X"E1",X"CB",X"BE",X"DD",X"35",X"06",
		X"28",X"05",X"CD",X"B5",X"51",X"E1",X"C9",X"DD",X"CB",X"05",X"66",X"28",X"07",X"C3",X"C0",X"59",
		X"CB",X"FE",X"CB",X"DE",X"DD",X"36",X"00",X"00",X"E1",X"3A",X"00",X"E0",X"87",X"D0",X"3A",X"09",
		X"E3",X"A7",X"C0",X"CD",X"F4",X"02",X"3A",X"02",X"A0",X"E6",X"08",X"28",X"07",X"7D",X"E6",X"80",
		X"B4",X"C0",X"18",X"05",X"7D",X"E6",X"E0",X"B4",X"C0",X"21",X"09",X"E3",X"36",X"80",X"23",X"EB",
		X"DD",X"E5",X"E1",X"23",X"01",X"04",X"00",X"ED",X"B0",X"C9",X"21",X"00",X"E3",X"CB",X"FE",X"DD",
		X"7E",X"06",X"A7",X"20",X"1A",X"DD",X"34",X"06",X"CD",X"2A",X"51",X"DD",X"CB",X"05",X"66",X"28",
		X"05",X"21",X"C5",X"E1",X"CB",X"DE",X"CD",X"91",X"51",X"3E",X"12",X"CD",X"EA",X"02",X"C9",X"DD",
		X"7E",X"05",X"E6",X"0F",X"C8",X"CD",X"B5",X"51",X"E1",X"C9",X"DD",X"7E",X"05",X"E6",X"0F",X"C8",
		X"DD",X"CB",X"05",X"6E",X"28",X"07",X"21",X"C2",X"E2",X"CB",X"D6",X"3D",X"C8",X"4F",X"FD",X"E5",
		X"FD",X"21",X"1A",X"E2",X"11",X"15",X"00",X"06",X"08",X"FD",X"7E",X"00",X"E6",X"9C",X"FE",X"90",
		X"20",X"11",X"C5",X"01",X"FF",X"0E",X"CD",X"D7",X"05",X"C1",X"30",X"07",X"FD",X"CB",X"00",X"D6",
		X"0D",X"28",X"2B",X"FD",X"19",X"10",X"E2",X"FD",X"21",X"D3",X"E2",X"11",X"0F",X"00",X"06",X"03",
		X"FD",X"7E",X"00",X"E6",X"BC",X"FE",X"90",X"20",X"11",X"C5",X"01",X"FF",X"0E",X"CD",X"D7",X"05",
		X"C1",X"30",X"07",X"FD",X"CB",X"00",X"D6",X"0D",X"28",X"04",X"FD",X"19",X"10",X"E2",X"FD",X"E1",
		X"C9",X"DD",X"7E",X"05",X"E6",X"0F",X"C8",X"FE",X"06",X"38",X"02",X"3E",X"05",X"3D",X"5F",X"16",
		X"00",X"21",X"26",X"54",X"19",X"7E",X"21",X"7D",X"E0",X"36",X"00",X"23",X"77",X"23",X"36",X"00",
		X"EB",X"CD",X"2A",X"03",X"C9",X"DD",X"7E",X"05",X"E6",X"0F",X"FE",X"06",X"38",X"02",X"3E",X"05",
		X"C6",X"72",X"47",X"0E",X"0A",X"DD",X"7E",X"01",X"D6",X"08",X"57",X"DD",X"5E",X"03",X"D5",X"CD",
		X"9D",X"02",X"D1",X"7A",X"C6",X"10",X"57",X"06",X"72",X"0E",X"0A",X"CD",X"9D",X"02",X"C9",X"DD",
		X"7E",X"03",X"E6",X"07",X"28",X"09",X"FE",X"07",X"28",X"05",X"DD",X"CB",X"05",X"BE",X"C9",X"DD",
		X"CB",X"05",X"7E",X"C0",X"DD",X"CB",X"05",X"FE",X"DD",X"7E",X"01",X"C6",X"04",X"E6",X"F8",X"57",
		X"DD",X"7E",X"03",X"C6",X"07",X"5F",X"CD",X"0B",X"54",X"D8",X"2B",X"CD",X"0E",X"54",X"D8",X"11",
		X"E1",X"FF",X"19",X"CD",X"0E",X"54",X"D8",X"2B",X"CD",X"0E",X"54",X"D8",X"06",X"05",X"CD",X"87",
		X"1B",X"79",X"32",X"01",X"E3",X"CD",X"87",X"1B",X"79",X"32",X"02",X"E3",X"2B",X"CD",X"71",X"1B",
		X"79",X"32",X"03",X"E3",X"CD",X"71",X"1B",X"79",X"32",X"04",X"E3",X"11",X"20",X"00",X"19",X"05",
		X"CD",X"71",X"1B",X"79",X"32",X"05",X"E3",X"CD",X"71",X"1B",X"79",X"32",X"06",X"E3",X"23",X"CD",
		X"87",X"1B",X"79",X"32",X"07",X"E3",X"CD",X"87",X"1B",X"79",X"32",X"08",X"E3",X"21",X"01",X"E3",
		X"06",X"08",X"3E",X"DB",X"CD",X"EC",X"39",X"DD",X"7E",X"01",X"C6",X"04",X"E6",X"F8",X"57",X"E6",
		X"08",X"C8",X"DD",X"7E",X"03",X"3C",X"E6",X"F8",X"5F",X"E6",X"08",X"C0",X"DD",X"7E",X"05",X"DD",
		X"CB",X"05",X"F6",X"E6",X"40",X"C8",X"D5",X"21",X"01",X"E0",X"CB",X"C6",X"CD",X"C0",X"1D",X"CD",
		X"15",X"1F",X"D1",X"7E",X"E6",X"07",X"C0",X"44",X"4D",X"1D",X"CD",X"89",X"1D",X"EB",X"60",X"69",
		X"1A",X"FE",X"8A",X"28",X"04",X"FE",X"76",X"20",X"03",X"CD",X"27",X"1F",X"EB",X"01",X"E0",X"FF",
		X"09",X"EB",X"1A",X"FE",X"8A",X"28",X"03",X"FE",X"76",X"C0",X"CD",X"33",X"1F",X"C9",X"FD",X"E5",
		X"FD",X"21",X"1A",X"E2",X"11",X"15",X"00",X"06",X"08",X"D9",X"01",X"08",X"0E",X"D9",X"FD",X"7E",
		X"00",X"E6",X"9C",X"FE",X"90",X"28",X"04",X"FE",X"80",X"20",X"1E",X"D9",X"CD",X"D7",X"05",X"D9",
		X"30",X"17",X"FD",X"7E",X"00",X"E6",X"9C",X"FE",X"90",X"28",X"09",X"FD",X"CB",X"00",X"E6",X"DD",
		X"34",X"05",X"18",X"05",X"D9",X"CD",X"98",X"53",X"D9",X"FD",X"19",X"10",X"D1",X"FD",X"21",X"C2",
		X"E2",X"FD",X"7E",X"00",X"E6",X"B8",X"28",X"24",X"FE",X"B0",X"28",X"19",X"FE",X"A0",X"20",X"1C",
		X"01",X"08",X"0E",X"CD",X"D7",X"05",X"30",X"14",X"FD",X"CB",X"00",X"E6",X"DD",X"34",X"05",X"DD",
		X"CB",X"05",X"EE",X"18",X"07",X"DD",X"CB",X"05",X"6E",X"C4",X"98",X"53",X"FD",X"21",X"C5",X"E1",
		X"FD",X"7E",X"00",X"E6",X"98",X"28",X"21",X"FE",X"90",X"28",X"16",X"FE",X"80",X"20",X"19",X"01",
		X"09",X"09",X"CD",X"D7",X"05",X"30",X"11",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"05",X"E6",X"18",
		X"07",X"DD",X"CB",X"05",X"66",X"C4",X"98",X"53",X"FD",X"21",X"D3",X"E2",X"11",X"0F",X"00",X"06",
		X"03",X"D9",X"01",X"08",X"0E",X"D9",X"FD",X"7E",X"00",X"E6",X"BC",X"FE",X"90",X"28",X"04",X"FE",
		X"80",X"20",X"1E",X"D9",X"CD",X"D7",X"05",X"D9",X"30",X"17",X"FD",X"7E",X"00",X"E6",X"BC",X"FE",
		X"90",X"28",X"09",X"FD",X"CB",X"00",X"E6",X"DD",X"34",X"05",X"18",X"05",X"D9",X"CD",X"98",X"53",
		X"D9",X"FD",X"19",X"10",X"D1",X"FD",X"E1",X"C9",X"FD",X"56",X"03",X"FD",X"5E",X"04",X"21",X"AB",
		X"FE",X"19",X"FD",X"74",X"03",X"FD",X"75",X"04",X"C9",X"DD",X"56",X"01",X"DD",X"7E",X"03",X"D6",
		X"09",X"5F",X"D5",X"CD",X"0B",X"54",X"D1",X"38",X"4D",X"7A",X"C6",X"06",X"57",X"D5",X"CD",X"0B",
		X"54",X"D1",X"38",X"29",X"7A",X"D6",X"0D",X"57",X"D5",X"CD",X"0B",X"54",X"D1",X"38",X"05",X"DD",
		X"36",X"00",X"B0",X"C9",X"7A",X"C6",X"0F",X"57",X"D5",X"CD",X"0B",X"54",X"D1",X"38",X"27",X"7B",
		X"C6",X"08",X"5F",X"CD",X"0B",X"54",X"38",X"1E",X"DD",X"36",X"00",X"A8",X"C9",X"7A",X"D6",X"0E",
		X"57",X"D5",X"CD",X"0B",X"54",X"D1",X"38",X"0E",X"7B",X"C6",X"08",X"5F",X"CD",X"0B",X"54",X"38",
		X"05",X"DD",X"36",X"00",X"A9",X"C9",X"DD",X"36",X"00",X"80",X"C9",X"CD",X"89",X"1D",X"7E",X"FE",
		X"77",X"38",X"11",X"FE",X"7C",X"D8",X"FE",X"94",X"38",X"0A",X"FE",X"A4",X"D8",X"FE",X"DC",X"38",
		X"03",X"FE",X"E4",X"D8",X"A7",X"C9",X"10",X"20",X"40",X"60",X"80",X"3A",X"00",X"E0",X"E6",X"40",
		X"CA",X"BC",X"54",X"DD",X"CB",X"00",X"76",X"20",X"19",X"DD",X"CB",X"00",X"F6",X"DD",X"36",X"05",
		X"02",X"DD",X"36",X"06",X"58",X"DD",X"36",X"07",X"00",X"3E",X"23",X"06",X"00",X"CD",X"D9",X"02",
		X"18",X"1D",X"DD",X"CB",X"00",X"6E",X"20",X"6E",X"3A",X"B6",X"E1",X"A7",X"20",X"49",X"DD",X"46",
		X"05",X"DD",X"4E",X"06",X"0B",X"78",X"B1",X"28",X"53",X"DD",X"70",X"05",X"DD",X"71",X"06",X"3A",
		X"C5",X"E1",X"E6",X"98",X"FE",X"80",X"20",X"2F",X"FD",X"E5",X"FD",X"21",X"C5",X"E1",X"01",X"05",
		X"05",X"CD",X"D7",X"05",X"FD",X"E1",X"30",X"1F",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"07",X"1E",
		X"11",X"EB",X"54",X"CD",X"2A",X"03",X"3A",X"00",X"E0",X"87",X"D0",X"21",X"B6",X"E1",X"CB",X"FE",
		X"CB",X"EE",X"FD",X"36",X"30",X"03",X"C9",X"DD",X"34",X"07",X"DD",X"7E",X"07",X"E6",X"06",X"0F",
		X"FE",X"03",X"C8",X"C6",X"69",X"47",X"0E",X"07",X"CD",X"97",X"02",X"C9",X"DD",X"36",X"00",X"00",
		X"3E",X"23",X"CD",X"EA",X"02",X"C9",X"DD",X"35",X"07",X"28",X"F1",X"DD",X"7E",X"01",X"D6",X"08",
		X"57",X"DD",X"5E",X"03",X"06",X"77",X"0E",X"0A",X"C5",X"D5",X"CD",X"9D",X"02",X"D1",X"C1",X"7A",
		X"C6",X"10",X"57",X"06",X"72",X"CD",X"9D",X"02",X"C9",X"00",X"80",X"00",X"21",X"01",X"E0",X"CB",
		X"CE",X"CB",X"86",X"21",X"12",X"E4",X"11",X"06",X"00",X"0E",X"0C",X"06",X"0D",X"CB",X"BE",X"23",
		X"23",X"10",X"FA",X"19",X"0D",X"20",X"F4",X"21",X"00",X"00",X"22",X"D0",X"E5",X"22",X"10",X"E6",
		X"DD",X"21",X"C5",X"E1",X"CD",X"A3",X"1D",X"22",X"CE",X"E5",X"CB",X"FE",X"23",X"36",X"00",X"3E",
		X"01",X"32",X"31",X"E4",X"DD",X"21",X"CE",X"E5",X"FD",X"21",X"10",X"E6",X"EB",X"1B",X"1A",X"CB",
		X"5F",X"28",X"09",X"21",X"02",X"00",X"19",X"CB",X"7E",X"CC",X"9C",X"56",X"CB",X"57",X"28",X"09",
		X"21",X"20",X"00",X"19",X"CB",X"7E",X"CC",X"9C",X"56",X"CB",X"4F",X"28",X"09",X"21",X"FE",X"FF",
		X"19",X"CB",X"7E",X"CC",X"9C",X"56",X"CB",X"47",X"28",X"09",X"21",X"E0",X"FF",X"19",X"CB",X"7E",
		X"CC",X"9C",X"56",X"DD",X"23",X"DD",X"23",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"7A",X"B3",X"20",
		X"BD",X"21",X"31",X"E4",X"34",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"FD",X"E1",X"DD",X"5E",X"00",
		X"DD",X"56",X"01",X"7A",X"B3",X"20",X"A7",X"21",X"01",X"E0",X"CB",X"8E",X"CB",X"E6",X"21",X"01",
		X"E0",X"CB",X"DE",X"CB",X"96",X"21",X"12",X"E4",X"11",X"06",X"00",X"0E",X"0C",X"06",X"0D",X"CB",
		X"B6",X"23",X"23",X"10",X"FA",X"19",X"0D",X"20",X"F4",X"DD",X"21",X"C5",X"E1",X"CD",X"A3",X"1D",
		X"DD",X"7E",X"00",X"E6",X"06",X"28",X"32",X"FE",X"02",X"28",X"20",X"FE",X"04",X"28",X"0E",X"DD",
		X"7E",X"03",X"D6",X"18",X"E6",X"F0",X"28",X"42",X"11",X"FE",X"FF",X"18",X"28",X"3E",X"D8",X"DD",
		X"96",X"03",X"E6",X"F0",X"28",X"34",X"11",X"02",X"00",X"18",X"1A",X"DD",X"7E",X"01",X"D6",X"20",
		X"E6",X"F0",X"28",X"26",X"11",X"E0",X"FF",X"18",X"0C",X"3E",X"E0",X"DD",X"96",X"01",X"E6",X"F0",
		X"28",X"18",X"11",X"20",X"00",X"0F",X"0F",X"0F",X"0F",X"47",X"E5",X"19",X"7E",X"E6",X"0F",X"20",
		X"05",X"10",X"F8",X"E1",X"18",X"04",X"C1",X"18",X"01",X"2B",X"CB",X"F6",X"23",X"7E",X"A7",X"28",
		X"30",X"3D",X"2B",X"CB",X"5E",X"28",X"09",X"23",X"23",X"23",X"BE",X"28",X"EC",X"2B",X"2B",X"2B",
		X"CB",X"56",X"28",X"09",X"EB",X"21",X"21",X"00",X"19",X"BE",X"28",X"DD",X"EB",X"CB",X"4E",X"28",
		X"05",X"2B",X"BE",X"28",X"D4",X"23",X"CB",X"46",X"28",X"07",X"11",X"E1",X"FF",X"19",X"BE",X"28",
		X"C8",X"21",X"01",X"E0",X"CB",X"9E",X"C9",X"21",X"01",X"E0",X"CB",X"A6",X"21",X"12",X"E4",X"11",
		X"06",X"00",X"0E",X"0C",X"06",X"0D",X"CB",X"AE",X"23",X"23",X"10",X"FA",X"19",X"0D",X"20",X"F4",
		X"21",X"CA",X"E4",X"18",X"01",X"2B",X"CB",X"EE",X"23",X"7E",X"A7",X"C8",X"3D",X"2B",X"CB",X"5E",
		X"28",X"09",X"23",X"23",X"23",X"BE",X"28",X"ED",X"2B",X"2B",X"2B",X"CB",X"56",X"28",X"09",X"EB",
		X"21",X"21",X"00",X"19",X"BE",X"28",X"DE",X"EB",X"CB",X"4E",X"28",X"05",X"2B",X"BE",X"28",X"D5",
		X"23",X"CB",X"46",X"C8",X"11",X"E1",X"FF",X"19",X"BE",X"28",X"CA",X"C9",X"CB",X"FE",X"FD",X"2B",
		X"FD",X"2B",X"FD",X"75",X"00",X"FD",X"74",X"01",X"23",X"3A",X"31",X"E4",X"77",X"1A",X"C9",X"0E",
		X"22",X"AF",X"11",X"04",X"00",X"21",X"01",X"90",X"06",X"40",X"77",X"19",X"10",X"FC",X"0D",X"20",
		X"F4",X"AF",X"32",X"00",X"F0",X"32",X"00",X"F8",X"3E",X"29",X"08",X"3E",X"09",X"21",X"00",X"80",
		X"0E",X"04",X"06",X"04",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F9",X"08",X"0D",X"20",X"F3",X"3E",
		X"1B",X"32",X"90",X"8D",X"3E",X"18",X"32",X"B0",X"8D",X"3E",X"16",X"32",X"D0",X"8D",X"21",X"00",
		X"00",X"11",X"00",X"00",X"AF",X"06",X"20",X"86",X"2C",X"20",X"FC",X"24",X"10",X"F9",X"BB",X"28",
		X"24",X"16",X"FF",X"47",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"C6",X"00",X"32",X"50",X"8E",X"78",
		X"E6",X"0F",X"C6",X"00",X"32",X"70",X"8E",X"7B",X"C6",X"01",X"32",X"10",X"8E",X"01",X"00",X"00",
		X"0B",X"78",X"B1",X"20",X"FB",X"1C",X"7B",X"FE",X"04",X"38",X"C9",X"CB",X"7A",X"C2",X"00",X"00",
		X"3E",X"18",X"32",X"30",X"8E",X"3E",X"14",X"32",X"50",X"8E",X"01",X"00",X"00",X"0B",X"78",X"B1",
		X"20",X"FB",X"3E",X"1B",X"32",X"90",X"8D",X"3E",X"0A",X"32",X"B0",X"8D",X"3E",X"16",X"32",X"D0",
		X"8D",X"3E",X"29",X"32",X"30",X"8E",X"32",X"50",X"8E",X"06",X"00",X"78",X"D9",X"67",X"2E",X"00",
		X"11",X"00",X"E0",X"01",X"00",X"10",X"ED",X"B0",X"11",X"00",X"80",X"01",X"00",X"10",X"ED",X"B0",
		X"D9",X"78",X"D9",X"57",X"1E",X"00",X"21",X"00",X"E0",X"01",X"02",X"10",X"1A",X"BE",X"20",X"1C",
		X"13",X"2C",X"20",X"F8",X"24",X"10",X"F5",X"21",X"00",X"80",X"06",X"10",X"0D",X"20",X"ED",X"D9",
		X"78",X"C6",X"01",X"47",X"FE",X"61",X"38",X"C3",X"D9",X"21",X"00",X"00",X"D9",X"3E",X"29",X"08",
		X"3E",X"09",X"21",X"00",X"80",X"0E",X"04",X"06",X"04",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F9",
		X"08",X"0D",X"20",X"F3",X"3E",X"1B",X"32",X"90",X"8D",X"3E",X"0A",X"32",X"B0",X"8D",X"3E",X"16",
		X"32",X"D0",X"8D",X"D9",X"7C",X"B5",X"20",X"0C",X"3E",X"18",X"32",X"30",X"8E",X"3E",X"14",X"32",
		X"50",X"8E",X"18",X"1E",X"7C",X"FE",X"88",X"38",X"10",X"FE",X"90",X"38",X"10",X"FE",X"E8",X"30",
		X"04",X"3E",X"01",X"18",X"0A",X"3E",X"02",X"18",X"06",X"3E",X"03",X"18",X"02",X"3E",X"04",X"32",
		X"30",X"8E",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"7C",X"B5",X"D9",X"C2",X"00",X"00",
		X"31",X"80",X"EB",X"21",X"29",X"58",X"CD",X"03",X"04",X"21",X"01",X"98",X"36",X"9F",X"36",X"BF",
		X"36",X"DF",X"36",X"FF",X"21",X"02",X"98",X"36",X"9F",X"36",X"BF",X"36",X"DF",X"36",X"FF",X"01",
		X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"18",X"0D",X"70",X"89",X"09",X"09",X"1C",X"18",X"1E",
		X"17",X"0D",X"29",X"18",X"0F",X"0F",X"21",X"98",X"58",X"06",X"13",X"C5",X"CD",X"03",X"04",X"C1",
		X"10",X"F9",X"16",X"02",X"01",X"00",X"00",X"C5",X"D5",X"21",X"B9",X"8E",X"3A",X"00",X"A0",X"CD",
		X"77",X"58",X"3A",X"01",X"A0",X"CD",X"77",X"58",X"21",X"07",X"8E",X"3A",X"02",X"A0",X"CD",X"86",
		X"58",X"21",X"06",X"8E",X"3A",X"03",X"A0",X"CD",X"86",X"58",X"D1",X"C1",X"10",X"D9",X"0D",X"20",
		X"D6",X"15",X"20",X"D3",X"C3",X"46",X"59",X"06",X"08",X"87",X"38",X"04",X"36",X"00",X"18",X"02",
		X"36",X"01",X"2B",X"10",X"F4",X"C9",X"06",X"08",X"11",X"20",X"00",X"87",X"38",X"04",X"36",X"00",
		X"18",X"02",X"36",X"01",X"19",X"10",X"F4",X"C9",X"70",X"89",X"09",X"09",X"29",X"29",X"29",X"29",
		X"29",X"29",X"29",X"29",X"29",X"59",X"89",X"09",X"04",X"1D",X"12",X"15",X"1D",X"58",X"89",X"09",
		X"09",X"1C",X"0E",X"15",X"0E",X"0C",X"1D",X"29",X"02",X"19",X"37",X"8A",X"09",X"02",X"01",X"19",
		X"56",X"89",X"09",X"07",X"01",X"19",X"29",X"0F",X"12",X"1B",X"0E",X"B5",X"89",X"09",X"02",X"1E",
		X"19",X"B4",X"89",X"09",X"05",X"1B",X"12",X"10",X"11",X"1D",X"B3",X"89",X"09",X"04",X"0D",X"18",
		X"20",X"17",X"B2",X"89",X"09",X"04",X"15",X"0E",X"0F",X"1D",X"51",X"89",X"09",X"0A",X"0C",X"18",
		X"12",X"17",X"29",X"1B",X"12",X"10",X"11",X"1D",X"F0",X"89",X"09",X"04",X"15",X"0E",X"0F",X"1D",
		X"4F",X"89",X"09",X"08",X"17",X"18",X"1D",X"29",X"1E",X"1C",X"0E",X"0D",X"4E",X"89",X"09",X"07",
		X"02",X"19",X"29",X"0F",X"12",X"1B",X"0E",X"AD",X"89",X"09",X"02",X"1E",X"19",X"AC",X"89",X"09",
		X"05",X"1B",X"12",X"10",X"11",X"1D",X"AB",X"89",X"09",X"04",X"0D",X"18",X"20",X"17",X"AA",X"89",
		X"09",X"04",X"15",X"0E",X"0F",X"1D",X"07",X"89",X"09",X"07",X"0D",X"12",X"19",X"1C",X"20",X"29",
		X"0A",X"C6",X"89",X"09",X"01",X"0B",X"11",X"80",X"88",X"01",X"18",X"20",X"CD",X"6C",X"04",X"3E",
		X"F7",X"32",X"80",X"84",X"3E",X"F9",X"32",X"9F",X"84",X"3E",X"FD",X"32",X"60",X"87",X"3E",X"FF",
		X"32",X"7F",X"87",X"3E",X"F8",X"21",X"81",X"84",X"CD",X"AC",X"59",X"3E",X"FE",X"21",X"61",X"87",
		X"CD",X"AC",X"59",X"3E",X"FA",X"21",X"A0",X"84",X"CD",X"B3",X"59",X"3E",X"FC",X"21",X"BF",X"84",
		X"CD",X"B3",X"59",X"3E",X"FB",X"0E",X"16",X"21",X"A1",X"84",X"CD",X"AC",X"59",X"23",X"23",X"0D",
		X"20",X"F8",X"3E",X"89",X"0E",X"18",X"21",X"80",X"80",X"77",X"23",X"CD",X"AC",X"59",X"77",X"23",
		X"0D",X"20",X"F6",X"AF",X"32",X"00",X"F0",X"32",X"00",X"F8",X"18",X"FE",X"06",X"1E",X"77",X"23",
		X"10",X"FC",X"C9",X"06",X"16",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"C9",X"C4",X"FF",X"FF",
		X"21",X"C5",X"E1",X"CB",X"76",X"CA",X"C4",X"50",X"C3",X"C0",X"50",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"FF",X"32",X"26",X"EC",X"AF",X"21",X"00",X"EC",X"06",X"26",X"77",X"23",X"10",X"FC",X"C9",
		X"DD",X"21",X"00",X"EC",X"06",X"26",X"DD",X"CB",X"00",X"56",X"C4",X"F6",X"5A",X"DD",X"CB",X"00",
		X"46",X"C4",X"1D",X"5B",X"DD",X"CB",X"00",X"4E",X"C4",X"F6",X"5A",X"DD",X"23",X"10",X"E7",X"AF",
		X"32",X"74",X"EC",X"32",X"76",X"EC",X"21",X"26",X"EC",X"7E",X"FE",X"FF",X"28",X"1F",X"E5",X"47",
		X"87",X"87",X"80",X"4F",X"06",X"00",X"DD",X"21",X"00",X"60",X"DD",X"09",X"DD",X"5E",X"03",X"DD",
		X"56",X"04",X"D5",X"FD",X"E1",X"CD",X"98",X"5B",X"E1",X"23",X"23",X"18",X"DC",X"3A",X"74",X"EC",
		X"47",X"3E",X"9F",X"CB",X"00",X"38",X"03",X"32",X"01",X"98",X"CB",X"00",X"38",X"03",X"32",X"02",
		X"98",X"C6",X"20",X"30",X"EE",X"C9",X"DD",X"36",X"00",X"00",X"3E",X"26",X"90",X"4F",X"21",X"26",
		X"EC",X"7E",X"FE",X"FF",X"C8",X"B9",X"28",X"04",X"23",X"23",X"18",X"F5",X"54",X"5D",X"23",X"23",
		X"7E",X"12",X"FE",X"FF",X"C8",X"13",X"23",X"7E",X"12",X"13",X"23",X"18",X"F3",X"DD",X"7E",X"00",
		X"E6",X"F0",X"DD",X"77",X"00",X"C5",X"3E",X"26",X"90",X"4F",X"87",X"87",X"81",X"5F",X"16",X"00",
		X"FD",X"21",X"00",X"60",X"FD",X"19",X"06",X"01",X"21",X"26",X"EC",X"7E",X"23",X"FE",X"FF",X"28",
		X"1D",X"B9",X"28",X"2E",X"7E",X"23",X"FD",X"BE",X"00",X"38",X"F0",X"04",X"7E",X"23",X"FE",X"FF",
		X"28",X"0C",X"23",X"B9",X"20",X"F5",X"2B",X"54",X"5D",X"1B",X"1B",X"05",X"18",X"04",X"54",X"5D",
		X"23",X"23",X"1A",X"77",X"1B",X"2B",X"1A",X"77",X"1B",X"2B",X"10",X"F6",X"FD",X"7E",X"00",X"77",
		X"2B",X"71",X"FD",X"6E",X"01",X"FD",X"66",X"02",X"FD",X"5E",X"03",X"FD",X"56",X"04",X"79",X"12",
		X"13",X"7E",X"12",X"47",X"13",X"23",X"AF",X"C5",X"01",X"03",X"00",X"ED",X"B0",X"06",X"07",X"12",
		X"13",X"10",X"FC",X"C1",X"10",X"F1",X"C1",X"C9",X"FD",X"46",X"01",X"DD",X"E5",X"FD",X"E5",X"DD",
		X"E1",X"DD",X"23",X"DD",X"23",X"DD",X"7E",X"00",X"A7",X"20",X"07",X"11",X"0A",X"00",X"DD",X"19",
		X"18",X"F3",X"C5",X"CD",X"69",X"5C",X"C1",X"11",X"0A",X"00",X"DD",X"19",X"10",X"E7",X"DD",X"E1",
		X"FD",X"7E",X"01",X"A7",X"CA",X"5D",X"5C",X"3A",X"76",X"EC",X"FE",X"04",X"D0",X"A7",X"28",X"14",
		X"DD",X"4E",X"00",X"47",X"21",X"77",X"EC",X"7E",X"A9",X"57",X"E6",X"C0",X"C0",X"7A",X"E6",X"03",
		X"C8",X"23",X"10",X"F3",X"CD",X"10",X"5E",X"D0",X"21",X"76",X"EC",X"34",X"5E",X"16",X"00",X"19",
		X"DD",X"7E",X"00",X"77",X"3A",X"75",X"EC",X"32",X"74",X"EC",X"FD",X"46",X"01",X"FD",X"23",X"FD",
		X"23",X"FD",X"7E",X"00",X"A7",X"20",X"07",X"11",X"0A",X"00",X"FD",X"19",X"18",X"F3",X"C5",X"01",
		X"01",X"98",X"CB",X"47",X"28",X"03",X"01",X"02",X"98",X"E6",X"06",X"87",X"87",X"87",X"87",X"F6",
		X"80",X"57",X"FD",X"7E",X"00",X"E6",X"38",X"FE",X"20",X"38",X"04",X"FE",X"30",X"38",X"19",X"FD",
		X"5E",X"09",X"7B",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"B2",X"02",X"FD",X"7E",X"08",X"02",X"7B",
		X"E6",X"0F",X"B2",X"F6",X"10",X"02",X"18",X"0C",X"7A",X"FD",X"B6",X"08",X"02",X"7A",X"FD",X"B6",
		X"09",X"F6",X"10",X"02",X"C1",X"11",X"0A",X"00",X"FD",X"19",X"10",X"A5",X"C9",X"FD",X"4E",X"00",
		X"06",X"00",X"21",X"00",X"EC",X"09",X"CB",X"CE",X"C9",X"DD",X"7E",X"03",X"A7",X"28",X"23",X"DD",
		X"35",X"03",X"C0",X"DD",X"7E",X"00",X"E6",X"38",X"FE",X"30",X"30",X"16",X"DD",X"6E",X"01",X"DD",
		X"66",X"02",X"A7",X"28",X"05",X"FE",X"20",X"30",X"01",X"23",X"23",X"23",X"DD",X"75",X"01",X"DD",
		X"74",X"02",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"7E",X"FE",X"FF",X"CA",X"BB",X"5D",X"CB",X"7F",
		X"28",X"57",X"CB",X"77",X"28",X"1F",X"E6",X"07",X"87",X"87",X"87",X"47",X"DD",X"7E",X"00",X"E6",
		X"C7",X"B0",X"DD",X"77",X"00",X"23",X"DD",X"75",X"01",X"DD",X"74",X"02",X"AF",X"DD",X"77",X"08",
		X"DD",X"77",X"09",X"18",X"CD",X"EB",X"E6",X"30",X"0F",X"0F",X"0F",X"0F",X"C6",X"04",X"4F",X"06",
		X"00",X"DD",X"E5",X"E1",X"09",X"EB",X"1A",X"A7",X"20",X"10",X"7E",X"E6",X"0F",X"12",X"23",X"5E",
		X"23",X"56",X"DD",X"73",X"01",X"DD",X"72",X"02",X"18",X"A8",X"3D",X"12",X"20",X"F0",X"23",X"23",
		X"23",X"DD",X"75",X"01",X"DD",X"74",X"02",X"18",X"99",X"DD",X"7E",X"00",X"E6",X"38",X"28",X"14",
		X"FE",X"10",X"38",X"17",X"28",X"1D",X"FE",X"20",X"38",X"20",X"28",X"25",X"FE",X"30",X"38",X"28",
		X"28",X"2D",X"18",X"54",X"CD",X"C3",X"5D",X"CD",X"FA",X"5D",X"C9",X"CD",X"C3",X"5D",X"23",X"CD",
		X"08",X"5E",X"C9",X"CD",X"DD",X"5D",X"CD",X"FA",X"5D",X"C9",X"CD",X"DD",X"5D",X"CD",X"08",X"5E",
		X"C9",X"CD",X"E8",X"5D",X"CD",X"FA",X"5D",X"C9",X"CD",X"E8",X"5D",X"CD",X"08",X"5E",X"C9",X"DD",
		X"7E",X"08",X"DD",X"B6",X"09",X"28",X"29",X"23",X"23",X"E5",X"CD",X"08",X"5E",X"E1",X"23",X"56",
		X"23",X"5E",X"23",X"E5",X"DD",X"66",X"08",X"DD",X"6E",X"09",X"19",X"EB",X"E1",X"7E",X"23",X"6E",
		X"67",X"A7",X"ED",X"52",X"30",X"34",X"18",X"39",X"DD",X"7E",X"08",X"DD",X"B6",X"09",X"20",X"07",
		X"CD",X"DD",X"5D",X"CD",X"08",X"5E",X"C9",X"23",X"23",X"E5",X"CD",X"08",X"5E",X"E1",X"23",X"56",
		X"23",X"5E",X"23",X"E5",X"DD",X"66",X"08",X"DD",X"6E",X"09",X"A7",X"ED",X"52",X"EB",X"E1",X"7E",
		X"23",X"6E",X"67",X"A7",X"ED",X"52",X"28",X"02",X"30",X"07",X"DD",X"72",X"08",X"DD",X"73",X"09",
		X"C9",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"11",X"07",X"00",X"19",X"DD",X"75",X"01",X"DD",X"74",
		X"02",X"AF",X"DD",X"77",X"08",X"DD",X"77",X"09",X"C3",X"92",X"5C",X"DD",X"36",X"00",X"00",X"FD",
		X"35",X"01",X"C9",X"7E",X"87",X"5F",X"16",X"00",X"E5",X"21",X"14",X"5F",X"19",X"5E",X"23",X"56",
		X"E1",X"23",X"7E",X"E6",X"0F",X"B3",X"DD",X"72",X"08",X"DD",X"77",X"09",X"C9",X"7E",X"DD",X"77",
		X"08",X"23",X"7E",X"DD",X"77",X"09",X"23",X"C9",X"7E",X"E6",X"70",X"0F",X"0F",X"0F",X"0F",X"DD",
		X"77",X"08",X"7E",X"E6",X"0F",X"DD",X"77",X"09",X"23",X"C9",X"7E",X"E6",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"5F",X"16",X"00",X"21",X"04",X"5F",X"19",X"56",X"CD",X"D4",X"5E",X"DD",X"72",X"03",X"C9",
		X"3A",X"74",X"EC",X"32",X"75",X"EC",X"FD",X"E5",X"FD",X"46",X"01",X"FD",X"23",X"FD",X"23",X"FD",
		X"7E",X"00",X"E6",X"F8",X"20",X"07",X"11",X"0A",X"00",X"FD",X"19",X"18",X"F2",X"4F",X"E6",X"C0",
		X"FE",X"C0",X"28",X"68",X"FE",X"80",X"28",X"22",X"3A",X"75",X"EC",X"67",X"11",X"00",X"80",X"7C",
		X"A2",X"28",X"0B",X"CB",X"3A",X"1C",X"7B",X"FE",X"06",X"38",X"F4",X"C3",X"D0",X"5E",X"7C",X"B2",
		X"32",X"75",X"EC",X"7B",X"B1",X"FD",X"77",X"00",X"18",X"69",X"E1",X"E5",X"23",X"7E",X"90",X"28",
		X"16",X"FD",X"E5",X"E1",X"11",X"F6",X"FF",X"19",X"7E",X"FE",X"C0",X"38",X"0A",X"E6",X"07",X"C6",
		X"02",X"B1",X"FD",X"77",X"00",X"18",X"4C",X"3A",X"75",X"EC",X"CB",X"4F",X"20",X"0D",X"CB",X"CF",
		X"32",X"75",X"EC",X"79",X"F6",X"06",X"FD",X"77",X"00",X"18",X"38",X"CB",X"47",X"20",X"41",X"CB",
		X"C7",X"32",X"75",X"EC",X"79",X"F6",X"07",X"FD",X"77",X"00",X"18",X"27",X"3A",X"75",X"EC",X"57",
		X"E6",X"0A",X"20",X"0E",X"7A",X"F6",X"0A",X"32",X"75",X"EC",X"79",X"F6",X"04",X"FD",X"77",X"00",
		X"18",X"11",X"7A",X"E6",X"05",X"20",X"19",X"7A",X"F6",X"05",X"32",X"75",X"EC",X"79",X"F6",X"05",
		X"FD",X"77",X"00",X"11",X"0A",X"00",X"FD",X"19",X"05",X"C2",X"1F",X"5E",X"FD",X"E1",X"37",X"C9",
		X"FD",X"E1",X"A7",X"C9",X"FD",X"4E",X"00",X"06",X"00",X"21",X"00",X"EC",X"09",X"7E",X"E6",X"F0",
		X"C8",X"6F",X"26",X"00",X"29",X"7A",X"EB",X"CD",X"F5",X"5E",X"EB",X"CB",X"7B",X"28",X"01",X"14",
		X"7A",X"A7",X"C0",X"14",X"C9",X"21",X"00",X"00",X"06",X"08",X"0F",X"30",X"01",X"19",X"EB",X"29",
		X"EB",X"10",X"F7",X"C9",X"48",X"24",X"18",X"12",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",
		X"04",X"03",X"02",X"01",X"40",X"3F",X"C0",X"3B",X"60",X"38",X"30",X"35",X"40",X"32",X"60",X"2F",
		X"C0",X"2C",X"40",X"2A",X"E0",X"27",X"A0",X"25",X"80",X"23",X"80",X"21",X"A0",X"1F",X"E0",X"1D",
		X"30",X"1C",X"A0",X"1A",X"20",X"19",X"B0",X"17",X"60",X"16",X"20",X"15",X"F0",X"13",X"D0",X"12",
		X"C0",X"11",X"C0",X"10",X"D0",X"0F",X"F0",X"0E",X"10",X"0E",X"50",X"0D",X"90",X"0C",X"E0",X"0B",
		X"30",X"0B",X"90",X"0A",X"F0",X"09",X"60",X"09",X"E0",X"08",X"60",X"08",X"F0",X"07",X"70",X"07",
		X"10",X"07",X"A0",X"06",X"40",X"06",X"F0",X"05",X"90",X"05",X"40",X"05",X"00",X"05",X"B0",X"04",
		X"70",X"04",X"30",X"04",X"F0",X"03",X"C0",X"03",X"80",X"03",X"50",X"03",X"20",X"03",X"F0",X"02",
		X"D0",X"02",X"A0",X"02",X"80",X"02",X"60",X"02",X"40",X"02",X"20",X"02",X"00",X"02",X"E0",X"01",
		X"C0",X"01",X"B0",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"BE",X"60",X"7B",X"EC",X"C0",X"C2",X"60",X"87",X"EC",X"C0",X"C6",X"60",X"93",X"EC",X"C0",
		X"CA",X"60",X"9F",X"EC",X"C0",X"CE",X"60",X"AB",X"EC",X"C0",X"D2",X"60",X"B7",X"EC",X"C0",X"D6",
		X"60",X"C3",X"EC",X"C0",X"DA",X"60",X"CF",X"EC",X"C0",X"DE",X"60",X"DB",X"EC",X"FF",X"E2",X"60",
		X"E7",X"EC",X"FF",X"E6",X"60",X"F3",X"EC",X"FF",X"EA",X"60",X"FF",X"EC",X"FF",X"EE",X"60",X"0B",
		X"ED",X"FF",X"F2",X"60",X"17",X"ED",X"FF",X"F6",X"60",X"23",X"ED",X"FF",X"FA",X"60",X"2F",X"ED",
		X"FF",X"01",X"61",X"45",X"ED",X"F7",X"08",X"61",X"5B",X"ED",X"CA",X"0F",X"61",X"71",X"ED",X"C6",
		X"16",X"61",X"87",X"ED",X"00",X"1D",X"61",X"9D",X"ED",X"C2",X"24",X"61",X"B3",X"ED",X"C1",X"2B",
		X"61",X"C9",X"ED",X"FB",X"32",X"61",X"DF",X"ED",X"C3",X"39",X"61",X"F5",X"ED",X"01",X"40",X"61",
		X"0B",X"EE",X"C2",X"4A",X"61",X"2B",X"EE",X"C1",X"54",X"61",X"4B",X"EE",X"C1",X"5E",X"61",X"6B",
		X"EE",X"02",X"68",X"61",X"8B",X"EE",X"42",X"72",X"61",X"AB",X"EE",X"41",X"7C",X"61",X"CB",X"EE",
		X"80",X"86",X"61",X"EB",X"EE",X"01",X"90",X"61",X"0B",X"EF",X"01",X"9A",X"61",X"2B",X"EF",X"40",
		X"A4",X"61",X"4B",X"EF",X"03",X"B1",X"61",X"75",X"EF",X"FF",X"BE",X"61",X"9F",X"EF",X"01",X"40",
		X"FF",X"6F",X"01",X"40",X"D0",X"61",X"01",X"40",X"E0",X"61",X"01",X"40",X"F0",X"61",X"01",X"40",
		X"00",X"62",X"01",X"40",X"10",X"62",X"01",X"40",X"20",X"62",X"01",X"40",X"30",X"62",X"01",X"40",
		X"40",X"62",X"01",X"40",X"FF",X"6F",X"01",X"40",X"FF",X"6F",X"01",X"40",X"FF",X"6F",X"01",X"40",
		X"FF",X"6F",X"01",X"40",X"FF",X"6F",X"01",X"40",X"FF",X"6F",X"02",X"40",X"D0",X"7C",X"40",X"40",
		X"7D",X"02",X"40",X"D0",X"69",X"40",X"40",X"6A",X"02",X"40",X"70",X"62",X"40",X"A0",X"62",X"02",
		X"40",X"D0",X"63",X"40",X"10",X"64",X"02",X"40",X"E0",X"67",X"40",X"F0",X"67",X"02",X"40",X"70",
		X"63",X"40",X"A0",X"63",X"02",X"40",X"50",X"62",X"40",X"60",X"62",X"02",X"40",X"50",X"64",X"40",
		X"70",X"64",X"02",X"40",X"A0",X"66",X"40",X"00",X"67",X"02",X"40",X"FF",X"6F",X"40",X"FF",X"6F",
		X"03",X"40",X"C0",X"68",X"40",X"00",X"69",X"40",X"40",X"69",X"03",X"40",X"00",X"6B",X"40",X"10",
		X"6B",X"40",X"20",X"6B",X"03",X"40",X"90",X"64",X"40",X"B0",X"64",X"40",X"D0",X"64",X"03",X"40",
		X"F0",X"64",X"40",X"10",X"65",X"40",X"30",X"65",X"03",X"40",X"30",X"6B",X"40",X"B0",X"6B",X"40",
		X"70",X"6C",X"03",X"40",X"30",X"6D",X"40",X"B0",X"6D",X"40",X"30",X"6E",X"03",X"40",X"B0",X"6E",
		X"40",X"30",X"6F",X"40",X"A0",X"6F",X"03",X"40",X"D0",X"62",X"40",X"E0",X"62",X"40",X"F0",X"62",
		X"03",X"40",X"10",X"68",X"40",X"50",X"68",X"40",X"90",X"68",X"03",X"40",X"70",X"69",X"40",X"90",
		X"69",X"40",X"B0",X"69",X"04",X"40",X"60",X"67",X"40",X"80",X"67",X"40",X"A0",X"67",X"40",X"C0",
		X"67",X"04",X"40",X"40",X"66",X"40",X"70",X"66",X"40",X"00",X"63",X"40",X"20",X"63",X"04",X"40",
		X"50",X"65",X"40",X"A0",X"65",X"40",X"F0",X"65",X"40",X"FF",X"6F",X"FF",X"FF",X"70",X"13",X"FA",
		X"C0",X"19",X"D0",X"25",X"D0",X"82",X"D0",X"61",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"1B",X"D0",X"27",X"D0",X"82",X"E0",X"61",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"1D",X"D0",X"29",X"D0",X"82",X"F0",X"61",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"1E",X"D0",X"2A",X"D0",X"82",X"00",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"20",X"D0",X"2C",X"D0",X"82",X"10",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"22",X"D0",X"2E",X"D0",X"82",X"20",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"24",X"D0",X"30",X"D0",X"82",X"30",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"25",X"D0",X"31",X"D0",X"84",X"40",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0D",X"A0",X"00",X"DF",X"25",X"C0",X"26",X"C0",X"82",X"50",X"62",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"14",X"A0",X"00",X"DF",X"23",X"C0",X"24",X"C0",X"82",X"60",X"62",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"12",X"80",X"00",X"8F",X"17",X"C0",X"00",X"CF",X"17",X"C0",X"00",X"CF",X"14",X"C0",X"00",
		X"CF",X"17",X"C0",X"00",X"CF",X"17",X"C0",X"00",X"CF",X"14",X"C0",X"00",X"CF",X"80",X"70",X"62",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0F",X"C0",X"00",X"CF",X"0F",X"C0",X"00",X"CF",X"0B",X"C0",X"00",X"CF",X"0F",X"C0",X"00",
		X"CF",X"10",X"C0",X"00",X"CF",X"10",X"C0",X"00",X"CF",X"0B",X"C0",X"00",X"CF",X"10",X"C0",X"00",
		X"CF",X"80",X"A0",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"2F",X"91",X"2B",X"91",X"32",X"91",X"26",X"91",X"2B",X"91",X"00",X"2F",X"00",X"FF",X"FF",
		X"C0",X"2E",X"91",X"2A",X"91",X"31",X"91",X"25",X"91",X"2A",X"91",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"3D",X"91",X"3B",X"91",X"3A",X"91",X"38",X"91",X"36",X"91",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"31",X"80",X"35",X"80",X"00",X"6F",X"1E",X"80",X"20",X"80",X"00",X"6F",X"2D",X"80",X"23",
		X"80",X"00",X"6F",X"1C",X"80",X"19",X"A0",X"19",X"A2",X"19",X"A4",X"19",X"A8",X"FF",X"FF",X"FF",
		X"C0",X"00",X"0F",X"80",X"20",X"63",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"B2",X"02",X"B4",X"02",X"68",X"00",X"0F",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"26",X"E3",X"2B",X"E2",X"28",X"E1",X"2D",X"E0",X"2B",X"E0",X"2F",X"E0",X"2D",X"E1",X"32",
		X"E2",X"2F",X"E3",X"34",X"E4",X"32",X"E5",X"37",X"E6",X"34",X"E7",X"39",X"E8",X"37",X"E9",X"3B",
		X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"28",X"E3",X"2D",X"E2",X"2B",X"E1",X"2F",X"E0",X"2D",X"E0",X"32",X"E0",X"2F",X"E1",X"34",
		X"E2",X"32",X"E3",X"37",X"E4",X"34",X"E5",X"39",X"E6",X"37",X"E7",X"3B",X"E8",X"39",X"E9",X"3E",
		X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"30",X"C0",X"2F",X"C0",X"2E",X"C0",X"2D",X"C0",X"2C",X"C0",X"2B",X"C0",X"2A",X"C0",X"29",
		X"C0",X"28",X"C1",X"27",X"C1",X"26",X"C2",X"25",X"C2",X"24",X"C3",X"23",X"C3",X"22",X"C4",X"21",
		X"C4",X"20",X"C5",X"1F",X"C5",X"1E",X"C6",X"1D",X"C6",X"1C",X"C7",X"1B",X"C7",X"1A",X"C8",X"19",
		X"C8",X"18",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"30",X"C0",X"2F",X"C0",X"2E",X"C0",X"2D",X"C0",X"2C",X"C0",X"2B",X"C0",X"2A",X"C0",X"29",
		X"C0",X"28",X"C1",X"27",X"C1",X"26",X"C2",X"25",X"C2",X"24",X"C3",X"23",X"C3",X"22",X"C4",X"21",
		X"C4",X"20",X"C5",X"1F",X"C5",X"1E",X"C6",X"1D",X"C6",X"1C",X"C7",X"1B",X"C7",X"1A",X"C8",X"19",
		X"C8",X"18",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"11",X"F1",X"11",X"F0",X"11",X"F1",X"11",X"F2",X"11",X"F3",X"11",X"F4",X"11",X"F5",X"11",
		X"F6",X"11",X"F7",X"11",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0D",X"F1",X"0D",X"F0",X"0D",X"F1",X"0D",X"F2",X"0D",X"F3",X"0D",X"F4",X"0D",X"F5",X"0D",
		X"F6",X"0D",X"F7",X"0D",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0D",X"D2",X"16",X"D1",X"12",X"D0",X"19",X"D0",X"16",X"D0",X"1E",X"D0",X"19",X"D0",X"22",
		X"D1",X"1E",X"D2",X"25",X"D3",X"22",X"D4",X"2A",X"D5",X"25",X"D6",X"2E",X"D7",X"FF",X"FF",X"FF",
		X"C0",X"00",X"AF",X"16",X"D2",X"1E",X"D1",X"19",X"D0",X"22",X"D0",X"1E",X"D0",X"25",X"D0",X"22",
		X"D0",X"2A",X"D1",X"25",X"D2",X"2E",X"D3",X"2A",X"D4",X"31",X"D5",X"2E",X"D6",X"36",X"D7",X"FF",
		X"C0",X"00",X"4F",X"1E",X"D2",X"25",X"D1",X"22",X"D0",X"2A",X"D0",X"25",X"D0",X"2E",X"D0",X"2A",
		X"D0",X"31",X"D1",X"2E",X"D2",X"36",X"D3",X"31",X"D4",X"3A",X"D5",X"36",X"D6",X"3D",X"D7",X"FF",
		X"C0",X"3D",X"D7",X"36",X"D6",X"3A",X"D5",X"31",X"D4",X"36",X"D3",X"2E",X"D2",X"31",X"D1",X"2A",
		X"D0",X"2E",X"D0",X"25",X"D0",X"2A",X"D0",X"22",X"D0",X"25",X"D1",X"1E",X"D2",X"FF",X"FF",X"FF",
		X"C0",X"00",X"AF",X"36",X"D7",X"2E",X"D6",X"31",X"D5",X"2A",X"D4",X"2E",X"D3",X"25",X"D2",X"2A",
		X"D1",X"22",X"D0",X"25",X"D0",X"1E",X"D0",X"22",X"D0",X"19",X"D0",X"1E",X"D1",X"16",X"D2",X"FF",
		X"C0",X"00",X"4F",X"2E",X"D7",X"25",X"D6",X"2A",X"D5",X"22",X"D4",X"25",X"D3",X"1E",X"D2",X"22",
		X"D1",X"19",X"D0",X"1E",X"D0",X"16",X"D0",X"19",X"D0",X"12",X"D0",X"16",X"D1",X"0D",X"D2",X"FF",
		X"C0",X"19",X"C4",X"00",X"CF",X"1D",X"C6",X"00",X"CF",X"1D",X"C6",X"00",X"CF",X"1D",X"C6",X"00",
		X"CF",X"1B",X"C3",X"00",X"CF",X"1E",X"C5",X"00",X"CF",X"1E",X"C5",X"00",X"CF",X"1E",X"C5",X"00",
		X"CF",X"1D",X"C2",X"00",X"CF",X"20",X"C4",X"00",X"CF",X"20",X"C3",X"00",X"CF",X"20",X"C2",X"00",
		X"CF",X"20",X"C2",X"00",X"CF",X"1E",X"C4",X"00",X"CF",X"1D",X"C6",X"00",X"CF",X"1B",X"C8",X"00",
		X"CF",X"80",X"50",X"65",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"19",X"C4",X"00",X"CF",X"20",X"C6",X"00",X"CF",X"20",X"C6",X"00",X"CF",X"20",X"C6",X"00",
		X"CF",X"1B",X"C5",X"00",X"CF",X"22",X"C5",X"00",X"CF",X"22",X"C5",X"00",X"CF",X"22",X"C5",X"00",
		X"CF",X"1D",X"C2",X"00",X"CF",X"24",X"C4",X"00",X"CF",X"24",X"C3",X"00",X"CF",X"24",X"C2",X"00",
		X"CF",X"24",X"C2",X"00",X"CF",X"22",X"C4",X"00",X"CF",X"20",X"C6",X"00",X"CF",X"1E",X"C8",X"00",
		X"CF",X"80",X"A0",X"65",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"8F",X"25",X"C0",X"00",X"CF",X"29",X"C0",X"00",X"CF",X"2A",X"C0",X"00",X"CF",X"2C",
		X"80",X"00",X"8F",X"31",X"80",X"00",X"8F",X"30",X"80",X"00",X"8F",X"2E",X"80",X"00",X"8F",X"29",
		X"20",X"00",X"8F",X"00",X"8F",X"29",X"C0",X"00",X"CF",X"2A",X"C0",X"00",X"CF",X"29",X"C0",X"00",
		X"CF",X"27",X"20",X"00",X"8F",X"00",X"8F",X"27",X"C0",X"00",X"CF",X"29",X"C0",X"00",X"CF",X"2A",
		X"C0",X"00",X"CF",X"2C",X"20",X"00",X"8F",X"80",X"F0",X"65",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"38",X"80",X"3C",X"80",X"00",X"6F",X"15",X"80",X"1B",X"80",X"00",X"6F",X"27",X"80",X"2D",
		X"80",X"00",X"6F",X"04",X"80",X"01",X"A0",X"01",X"A2",X"01",X"A4",X"01",X"A8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"35",X"80",X"38",X"80",X"00",X"6F",X"1A",X"80",X"18",X"80",X"00",X"6F",X"2A",X"80",X"28",
		X"80",X"00",X"6F",X"10",X"80",X"0D",X"A0",X"0D",X"A2",X"0D",X"A4",X"0D",X"A8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"25",X"A2",X"00",X"CF",X"20",X"A3",X"00",X"CF",X"20",X"A3",X"00",X"CF",X"20",X"A3",X"00",
		X"CF",X"81",X"A1",X"66",X"22",X"A2",X"00",X"CF",X"1E",X"A3",X"00",X"CF",X"1E",X"A3",X"00",X"CF",
		X"1E",X"A3",X"00",X"CF",X"81",X"B4",X"66",X"20",X"A2",X"00",X"CF",X"24",X"A3",X"00",X"CF",X"24",
		X"A3",X"00",X"CF",X"24",X"A3",X"00",X"CF",X"81",X"C7",X"66",X"24",X"A2",X"00",X"CF",X"27",X"A3",
		X"00",X"CF",X"27",X"A3",X"00",X"CF",X"27",X"A3",X"00",X"CF",X"27",X"A2",X"00",X"CF",X"25",X"A3",
		X"00",X"CF",X"25",X"A3",X"00",X"3F",X"90",X"A0",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"19",X"D2",X"00",X"EF",X"14",X"D2",X"00",X"EF",X"87",X"00",X"67",X"16",X"D2",X"00",X"EF",
		X"12",X"D2",X"00",X"EF",X"87",X"0C",X"67",X"14",X"D2",X"00",X"EF",X"18",X"D2",X"00",X"EF",X"87",
		X"17",X"67",X"18",X"D2",X"00",X"EF",X"1B",X"D2",X"00",X"EF",X"83",X"22",X"67",X"27",X"A2",X"00",
		X"CF",X"22",X"A3",X"00",X"CF",X"22",X"A3",X"00",X"3F",X"90",X"00",X"67",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"38",X"A0",X"38",X"A2",X"38",X"A4",X"00",X"AF",X"3B",X"A0",X"3B",X"A2",X"3B",X"A4",X"00",
		X"AF",X"3D",X"A0",X"3D",X"A2",X"00",X"FF",X"80",X"60",X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"AF",X"39",X"A0",X"39",X"A2",X"39",X"A4",X"00",X"AF",X"39",X"A0",X"39",X"A2",X"39",
		X"A4",X"00",X"AF",X"3B",X"A0",X"00",X"FF",X"80",X"80",X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"AF",X"00",X"AF",X"00",X"AF",X"3D",X"A0",X"3D",X"A2",X"3D",X"A4",X"00",X"AF",X"39",
		X"A0",X"39",X"A2",X"39",X"A4",X"00",X"FF",X"80",X"A0",X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"AF",X"00",X"AF",X"3A",X"A0",X"3A",X"A2",X"3A",X"A4",X"00",X"AF",X"38",X"A0",X"38",
		X"A2",X"38",X"A4",X"00",X"AF",X"00",X"FF",X"80",X"C0",X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0D",X"A0",X"00",X"DF",X"25",X"C0",X"26",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"14",X"A0",X"00",X"DF",X"23",X"C0",X"24",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"1E",X"70",X"00",X"7F",X"25",X"90",X"00",X"EF",X"25",X"90",X"00",X"EF",X"22",X"30",X"1E",
		X"70",X"00",X"7F",X"1E",X"70",X"00",X"7F",X"25",X"90",X"00",X"EF",X"25",X"90",X"00",X"EF",X"22",
		X"30",X"1E",X"70",X"00",X"7F",X"20",X"70",X"00",X"7F",X"25",X"90",X"00",X"EF",X"25",X"90",X"00",
		X"EF",X"25",X"10",X"00",X"3F",X"19",X"70",X"00",X"7F",X"1E",X"70",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"12",X"76",X"00",X"7F",X"0D",X"96",X"00",X"EF",X"0D",X"96",X"00",X"EF",X"0F",X"36",X"12",
		X"76",X"00",X"7F",X"12",X"76",X"00",X"7F",X"0D",X"96",X"00",X"EF",X"0D",X"96",X"00",X"EF",X"0F",
		X"36",X"12",X"76",X"00",X"7F",X"14",X"76",X"00",X"7F",X"0D",X"96",X"00",X"EF",X"0D",X"96",X"00",
		X"EF",X"0D",X"16",X"00",X"3F",X"0D",X"76",X"00",X"7F",X"12",X"76",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"16",X"33",X"19",X"33",X"16",X"33",X"19",X"33",X"16",X"33",X"19",X"33",X"16",X"33",X"19",
		X"33",X"14",X"33",X"19",X"33",X"14",X"33",X"19",X"33",X"00",X"3F",X"01",X"74",X"00",X"7F",X"06",
		X"74",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"2C",X"A3",X"00",X"CF",X"25",X"A3",X"00",X"CF",X"82",X"C5",X"68",X"2A",X"A3",X"00",X"CF",
		X"24",X"A3",X"00",X"CF",X"82",X"D0",X"68",X"2C",X"A3",X"00",X"CF",X"2A",X"A3",X"00",X"CF",X"29",
		X"A3",X"00",X"CF",X"27",X"A3",X"00",X"CF",X"25",X"43",X"00",X"3F",X"00",X"4F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"11",X"A3",X"00",X"CF",X"83",X"01",X"69",X"0F",X"A3",X"00",X"CF",X"83",X"08",X"69",X"11",
		X"A3",X"00",X"CF",X"0F",X"A3",X"00",X"CF",X"0D",X"A3",X"00",X"CF",X"0C",X"A3",X"00",X"CF",X"0A",
		X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"20",X"A3",X"00",X"CF",X"1D",X"A3",X"00",X"CF",X"82",X"45",X"69",X"1E",X"A3",X"00",X"CF",
		X"1B",X"A3",X"00",X"CF",X"82",X"50",X"69",X"20",X"A3",X"00",X"CF",X"1E",X"A3",X"00",X"CF",X"1D",
		X"A3",X"00",X"CF",X"1B",X"A3",X"00",X"CF",X"19",X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"19",X"C2",X"00",X"CF",X"1E",X"C2",X"00",X"CF",X"22",X"C2",X"00",X"CF",X"25",X"72",X"00",
		X"7F",X"22",X"D2",X"00",X"DF",X"25",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0A",X"C2",X"00",X"CF",X"0D",X"C2",X"00",X"CF",X"12",X"C2",X"00",X"CF",X"16",X"72",X"00",
		X"7F",X"12",X"D2",X"00",X"DF",X"16",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"25",X"C2",X"00",X"CF",X"2A",X"C2",X"00",X"CF",X"2E",X"C2",X"00",X"CF",X"31",X"72",X"00",
		X"7F",X"2E",X"D2",X"00",X"DF",X"31",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0D",X"30",X"00",X"AF",X"0F",X"C0",X"00",X"EF",X"12",X"C0",X"00",X"EF",X"11",X"C0",X"00",
		X"EF",X"0F",X"C0",X"00",X"EF",X"14",X"A0",X"00",X"AF",X"14",X"A0",X"00",X"AF",X"14",X"C0",X"00",
		X"EF",X"16",X"C0",X"00",X"EF",X"11",X"C0",X"00",X"EF",X"12",X"C0",X"00",X"EF",X"0F",X"A0",X"00",
		X"AF",X"0F",X"A0",X"00",X"AF",X"0F",X"C0",X"00",X"EF",X"12",X"C0",X"00",X"EF",X"11",X"C0",X"00",
		X"EF",X"0F",X"C0",X"00",X"EF",X"0D",X"C0",X"00",X"EF",X"19",X"C0",X"00",X"EF",X"18",X"C0",X"00",
		X"EF",X"16",X"C0",X"00",X"EF",X"14",X"C0",X"00",X"EF",X"12",X"C0",X"00",X"EF",X"11",X"C0",X"00",
		X"EF",X"0F",X"C0",X"00",X"EF",X"80",X"D0",X"69",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"1D",X"C2",X"00",X"EF",X"20",X"C2",X"00",X"EF",X"1D",X"C2",X"00",X"EF",X"20",X"C2",X"00",
		X"EF",X"1E",X"C2",X"00",X"EF",X"1B",X"C2",X"00",X"EF",X"20",X"C2",X"00",X"EF",X"1E",X"C2",X"00",
		X"EF",X"1D",X"C2",X"00",X"EF",X"19",X"C2",X"00",X"EF",X"1D",X"C2",X"00",X"EF",X"19",X"C2",X"00",
		X"EF",X"1D",X"C2",X"00",X"EF",X"1E",X"C2",X"00",X"EF",X"19",X"C2",X"00",X"EF",X"1B",X"C2",X"00",
		X"EF",X"1E",X"C2",X"00",X"EF",X"20",X"C2",X"00",X"EF",X"1E",X"C2",X"00",X"EF",X"20",X"C2",X"00",
		X"EF",X"1E",X"C2",X"00",X"EF",X"1B",X"C2",X"00",X"EF",X"20",X"C2",X"00",X"EF",X"1E",X"C2",X"00",
		X"EF",X"1D",X"C2",X"00",X"EF",X"14",X"C2",X"00",X"EF",X"1B",X"C2",X"00",X"EF",X"1E",X"C2",X"00",
		X"EF",X"1D",X"C2",X"00",X"EF",X"1B",X"C2",X"00",X"EF",X"19",X"C2",X"00",X"EF",X"1E",X"C2",X"00",
		X"EF",X"80",X"40",X"6A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1B",X"A2",X"1E",X"A2",X"20",X"A2",X"1E",X"A2",X"20",X"A2",X"1E",X"A2",X"1B",X"A2",X"20",X"A2",
		X"1E",X"A2",X"1D",X"A2",X"14",X"A2",X"1B",X"A2",X"1E",X"A2",X"1D",X"C0",X"00",X"EF",X"1B",X"C0",
		X"00",X"EF",X"19",X"C0",X"00",X"EF",X"1E",X"C0",X"00",X"EF",X"80",X"B1",X"6A",X"FF",X"FF",X"FF",
		X"C0",X"29",X"B0",X"00",X"DF",X"35",X"C0",X"00",X"DF",X"33",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"31",X"90",X"00",X"DF",X"3D",X"C0",X"00",X"DF",X"3C",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"2C",X"70",X"00",X"DF",X"38",X"C0",X"00",X"DF",X"36",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"2C",X"41",X"00",X"FF",X"2C",X"41",X"00",X"FF",X"2A",X"41",X"00",X"FF",X"2A",X"41",X"00",
		X"FF",X"29",X"41",X"00",X"FF",X"29",X"41",X"00",X"FF",X"27",X"21",X"00",X"EF",X"2C",X"41",X"00",
		X"FF",X"2C",X"41",X"00",X"FF",X"2A",X"41",X"00",X"FF",X"2A",X"41",X"00",X"FF",X"29",X"41",X"00",
		X"FF",X"29",X"41",X"00",X"FF",X"27",X"21",X"00",X"EF",X"19",X"41",X"00",X"FF",X"19",X"41",X"00",
		X"FF",X"20",X"41",X"00",X"FF",X"20",X"41",X"00",X"FF",X"22",X"41",X"00",X"FF",X"22",X"41",X"00",
		X"FF",X"20",X"21",X"00",X"EF",X"1E",X"41",X"00",X"FF",X"1E",X"41",X"00",X"FF",X"1D",X"41",X"00",
		X"FF",X"1D",X"41",X"00",X"FF",X"1B",X"41",X"00",X"FF",X"1B",X"41",X"00",X"FF",X"19",X"21",X"00",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"31",X"A2",X"38",X"A2",X"00",X"FF",X"35",X"A2",X"38",X"A2",X"00",X"FF",X"30",X"A2",X"38",
		X"A2",X"00",X"FF",X"33",X"A2",X"38",X"A2",X"00",X"FF",X"31",X"A2",X"38",X"A2",X"00",X"FF",X"35",
		X"A2",X"38",X"A2",X"00",X"FF",X"30",X"A2",X"38",X"A2",X"33",X"A2",X"38",X"A2",X"00",X"EF",X"31",
		X"A2",X"38",X"A2",X"00",X"FF",X"35",X"A2",X"38",X"A2",X"00",X"FF",X"30",X"A2",X"38",X"A2",X"00",
		X"FF",X"33",X"A2",X"38",X"A2",X"00",X"FF",X"31",X"A2",X"38",X"A2",X"00",X"FF",X"35",X"A2",X"38",
		X"A2",X"00",X"FF",X"30",X"A2",X"38",X"A2",X"33",X"A2",X"38",X"A2",X"00",X"EF",X"0D",X"A2",X"14",
		X"A2",X"00",X"FF",X"11",X"A2",X"14",X"A2",X"00",X"FF",X"0D",X"A2",X"14",X"A2",X"00",X"FF",X"11",
		X"A2",X"14",X"A2",X"00",X"FF",X"0D",X"A2",X"16",X"A2",X"00",X"FF",X"13",X"A2",X"16",X"A2",X"00",
		X"FF",X"0D",X"A2",X"14",X"A2",X"11",X"A2",X"14",X"A2",X"00",X"EF",X"0C",X"A2",X"14",X"A2",X"00",
		X"FF",X"0F",X"A2",X"14",X"A2",X"00",X"FF",X"0D",X"A2",X"14",X"A2",X"00",X"FF",X"11",X"A2",X"14",
		X"A2",X"00",X"FF",X"0C",X"A2",X"14",X"A2",X"00",X"FF",X"12",X"A2",X"14",X"A2",X"00",X"FF",X"11",
		X"A2",X"14",X"A2",X"0D",X"42",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"38",X"A0",X"35",X"A0",X"00",X"FF",X"38",X"A0",X"35",X"A0",X"00",X"FF",X"36",X"A0",X"33",
		X"A0",X"00",X"FF",X"36",X"A0",X"33",X"A0",X"00",X"FF",X"35",X"A0",X"36",X"A0",X"00",X"FF",X"38",
		X"A0",X"35",X"A0",X"00",X"FF",X"33",X"A0",X"35",X"A0",X"33",X"40",X"00",X"EF",X"38",X"A0",X"35",
		X"A0",X"00",X"FF",X"38",X"A0",X"35",X"A0",X"00",X"FF",X"36",X"A0",X"33",X"A0",X"00",X"FF",X"36",
		X"A0",X"33",X"A0",X"00",X"FF",X"35",X"A0",X"36",X"A0",X"00",X"FF",X"38",X"A0",X"35",X"A0",X"00",
		X"FF",X"33",X"A0",X"35",X"A0",X"33",X"40",X"00",X"EF",X"31",X"A0",X"35",X"A0",X"00",X"FF",X"31",
		X"A0",X"35",X"A0",X"00",X"FF",X"38",X"A0",X"35",X"A0",X"00",X"FF",X"38",X"A0",X"35",X"A0",X"00",
		X"FF",X"3A",X"A0",X"3C",X"A0",X"00",X"FF",X"3D",X"A0",X"3A",X"A0",X"00",X"FF",X"38",X"A0",X"35",
		X"A0",X"31",X"40",X"00",X"EF",X"36",X"A0",X"38",X"A0",X"00",X"FF",X"3A",X"A0",X"36",X"A0",X"00",
		X"FF",X"35",X"A0",X"36",X"A0",X"00",X"FF",X"38",X"A0",X"35",X"A0",X"00",X"FF",X"33",X"A0",X"35",
		X"A0",X"00",X"FF",X"36",X"A0",X"33",X"A0",X"00",X"FF",X"31",X"A0",X"35",X"A0",X"31",X"40",X"00",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"1D",X"30",X"00",X"FF",X"1D",X"30",X"00",X"FF",X"1D",X"70",X"1E",X"30",X"00",X"FF",
		X"1F",X"70",X"20",X"10",X"20",X"70",X"00",X"FF",X"20",X"70",X"00",X"FF",X"1F",X"70",X"00",X"FF",
		X"20",X"70",X"22",X"30",X"00",X"FF",X"22",X"30",X"00",X"FF",X"22",X"70",X"24",X"30",X"00",X"FF",
		X"25",X"70",X"29",X"10",X"00",X"FF",X"00",X"3F",X"2A",X"70",X"00",X"FF",X"29",X"70",X"00",X"FF",
		X"27",X"10",X"22",X"30",X"00",X"FF",X"29",X"70",X"00",X"FF",X"27",X"70",X"00",X"FF",X"25",X"10",
		X"20",X"30",X"00",X"FF",X"1F",X"70",X"00",X"FF",X"20",X"70",X"00",X"FF",X"22",X"30",X"00",X"FF",
		X"22",X"30",X"00",X"FF",X"24",X"70",X"22",X"30",X"00",X"FF",X"20",X"70",X"25",X"10",X"25",X"70",
		X"00",X"FF",X"00",X"7F",X"00",X"FF",X"25",X"60",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"0D",X"72",X"14",X"72",X"00",X"FF",X"11",X"72",X"14",X"72",X"00",X"FF",X"0D",X"72",X"14",
		X"72",X"11",X"72",X"00",X"FF",X"14",X"72",X"0D",X"72",X"14",X"72",X"11",X"72",X"14",X"72",X"0D",
		X"72",X"00",X"FF",X"14",X"72",X"00",X"FF",X"11",X"72",X"00",X"FF",X"14",X"72",X"0D",X"72",X"16",
		X"72",X"00",X"FF",X"12",X"72",X"16",X"72",X"00",X"FF",X"0D",X"72",X"16",X"72",X"12",X"72",X"00",
		X"FF",X"16",X"72",X"0D",X"72",X"19",X"72",X"14",X"72",X"19",X"72",X"00",X"FF",X"11",X"72",X"19",
		X"72",X"16",X"72",X"00",X"FF",X"19",X"72",X"00",X"FF",X"12",X"32",X"12",X"32",X"12",X"32",X"12",
		X"F2",X"00",X"3F",X"00",X"EF",X"11",X"32",X"11",X"32",X"11",X"32",X"11",X"F2",X"00",X"3F",X"00",
		X"EF",X"11",X"72",X"16",X"72",X"00",X"FF",X"13",X"72",X"16",X"72",X"00",X"FF",X"11",X"72",X"14",
		X"72",X"12",X"72",X"00",X"FF",X"14",X"72",X"0D",X"72",X"11",X"72",X"14",X"72",X"11",X"72",X"0D",
		X"72",X"00",X"FF",X"00",X"7F",X"00",X"FF",X"0D",X"62",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"1F",X"00",X"1F",X"00",X"DF",X"00",X"1F",X"00",X"1F",X"00",X"DF",X"00",X"1F",X"00",
		X"1F",X"00",X"DF",X"00",X"1F",X"00",X"1F",X"00",X"DF",X"00",X"7F",X"1B",X"82",X"00",X"FF",X"1B",
		X"82",X"00",X"FF",X"1B",X"82",X"00",X"FF",X"1B",X"32",X"00",X"FF",X"00",X"3F",X"00",X"EF",X"00",
		X"7F",X"19",X"82",X"00",X"FF",X"19",X"82",X"00",X"FF",X"19",X"82",X"00",X"FF",X"19",X"32",X"00",
		X"FF",X"00",X"3F",X"00",X"EF",X"00",X"1F",X"00",X"1F",X"00",X"DF",X"00",X"1F",X"00",X"3F",X"00",
		X"EF",X"11",X"62",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"2B",X"A0",X"2C",X"A0",X"00",X"FF",X"29",X"80",X"00",X"BF",X"82",X"B7",X"6E",X"2B",X"A0",
		X"2C",X"A0",X"00",X"FF",X"29",X"80",X"00",X"BF",X"29",X"80",X"00",X"BF",X"35",X"80",X"00",X"BF",
		X"33",X"A0",X"00",X"FF",X"31",X"A0",X"00",X"FF",X"30",X"A0",X"00",X"FF",X"2E",X"A0",X"00",X"FF",
		X"2C",X"40",X"2A",X"40",X"29",X"80",X"00",X"BF",X"2A",X"80",X"00",X"BF",X"2C",X"40",X"00",X"9F",
		X"00",X"9F",X"2B",X"A0",X"2C",X"A0",X"00",X"FF",X"29",X"80",X"00",X"BF",X"82",X"F8",X"6E",X"2B",
		X"A0",X"2C",X"A0",X"00",X"FF",X"29",X"80",X"00",X"BF",X"29",X"80",X"00",X"BF",X"35",X"80",X"00",
		X"BF",X"33",X"A0",X"00",X"FF",X"31",X"A0",X"00",X"FF",X"30",X"A0",X"00",X"FF",X"2E",X"A0",X"00",
		X"FF",X"2C",X"40",X"30",X"40",X"31",X"80",X"00",X"BF",X"35",X"80",X"00",X"BF",X"31",X"40",X"FF",
		X"C0",X"13",X"A2",X"14",X"A2",X"00",X"FF",X"11",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",X"0D",
		X"82",X"00",X"BF",X"81",X"31",X"6F",X"0C",X"A2",X"00",X"FF",X"0A",X"A2",X"00",X"FF",X"08",X"A2",
		X"00",X"FF",X"06",X"A2",X"00",X"FF",X"05",X"42",X"03",X"42",X"01",X"82",X"00",X"BF",X"03",X"82",
		X"00",X"BF",X"05",X"82",X"00",X"BF",X"05",X"82",X"00",X"BF",X"13",X"A2",X"14",X"A2",X"00",X"FF",
		X"11",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",X"0D",X"82",X"00",X"BF",X"81",X"6A",X"6F",X"0C",
		X"A2",X"00",X"FF",X"0A",X"A2",X"00",X"FF",X"08",X"A2",X"00",X"FF",X"06",X"A2",X"00",X"FF",X"05",
		X"42",X"03",X"42",X"05",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",X"05",X"40",X"00",X"3F",X"FF",
		X"C0",X"01",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",X"05",X"82",X"00",X"BF",X"01",X"82",X"00",
		X"BF",X"82",X"A1",X"6F",X"01",X"82",X"00",X"BF",X"05",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",
		X"01",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",X"01",X"82",X"00",X"BF",X"05",X"82",X"00",X"BF",
		X"01",X"82",X"00",X"BF",X"82",X"C4",X"6F",X"01",X"82",X"00",X"BF",X"05",X"82",X"00",X"BF",X"01",
		X"40",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C2",X"DD",X"7E",X"03",X"FE",X"03",X"30",X"26",X"FE",X"02",X"30",X"0F",X"DD",X"7E",X"04",X"A7",
		X"20",X"09",X"11",X"B4",X"80",X"01",X"16",X"07",X"CD",X"6C",X"04",X"DD",X"7E",X"04",X"32",X"00",
		X"F8",X"E6",X"07",X"CC",X"36",X"70",X"DD",X"35",X"04",X"C0",X"DD",X"34",X"03",X"C9",X"DD",X"34",
		X"02",X"DD",X"36",X"03",X"00",X"C9",X"DD",X"7E",X"04",X"E6",X"F8",X"D6",X"E8",X"6F",X"26",X"00",
		X"29",X"29",X"11",X"14",X"80",X"19",X"EB",X"E6",X"08",X"0F",X"0F",X"4F",X"06",X"00",X"21",X"6A",
		X"70",X"09",X"7E",X"EB",X"01",X"01",X"07",X"C5",X"D5",X"E5",X"CD",X"5C",X"04",X"E1",X"D1",X"C1",
		X"13",X"1A",X"11",X"00",X"04",X"19",X"CD",X"5C",X"04",X"C9",X"5B",X"26",X"66",X"27",X"11",X"94",
		X"88",X"01",X"18",X"07",X"3E",X"40",X"CD",X"6D",X"04",X"08",X"3E",X"10",X"08",X"3E",X"8E",X"01",
		X"06",X"04",X"11",X"D7",X"88",X"CD",X"42",X"04",X"01",X"07",X"07",X"11",X"94",X"89",X"CD",X"42",
		X"04",X"01",X"04",X"05",X"CD",X"42",X"04",X"01",X"03",X"07",X"CD",X"42",X"04",X"21",X"94",X"80",
		X"01",X"18",X"07",X"3E",X"40",X"CD",X"5C",X"04",X"C9",X"DD",X"7E",X"03",X"A7",X"20",X"68",X"DD",
		X"34",X"03",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"FD",X"36",X"00",X"00",X"FD",X"36",
		X"04",X"01",X"FD",X"36",X"08",X"00",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"02",X"FD",X"36",
		X"16",X"00",X"FD",X"36",X"17",X"00",X"FD",X"36",X"1A",X"00",X"CD",X"85",X"04",X"CD",X"86",X"10",
		X"3A",X"E6",X"06",X"01",X"12",X"0E",X"21",X"C3",X"80",X"CD",X"5C",X"04",X"3A",X"E7",X"06",X"01",
		X"12",X"0E",X"21",X"C3",X"84",X"CD",X"5C",X"04",X"11",X"1E",X"71",X"CD",X"34",X"07",X"CD",X"6C",
		X"71",X"CD",X"6E",X"70",X"21",X"A0",X"71",X"CD",X"03",X"04",X"DD",X"36",X"01",X"1E",X"21",X"00",
		X"E0",X"CB",X"F6",X"23",X"CB",X"B6",X"C9",X"CD",X"AF",X"71",X"CD",X"58",X"72",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"45",X"55",X"55",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"E5",X"E1",X"11",
		X"31",X"00",X"19",X"E5",X"11",X"07",X"00",X"06",X"0C",X"36",X"00",X"19",X"10",X"FB",X"D1",X"21",
		X"92",X"71",X"01",X"07",X"00",X"ED",X"B0",X"01",X"07",X"00",X"ED",X"B0",X"3E",X"80",X"32",X"00",
		X"E3",X"C9",X"80",X"88",X"00",X"60",X"00",X"00",X"00",X"80",X"A8",X"00",X"60",X"00",X"00",X"00",
		X"52",X"89",X"3E",X"0B",X"12",X"17",X"1C",X"1D",X"1B",X"1E",X"0C",X"1D",X"12",X"18",X"17",X"DD",
		X"7E",X"03",X"FE",X"02",X"30",X"4D",X"DD",X"34",X"03",X"DD",X"36",X"04",X"FF",X"DD",X"36",X"05",
		X"1E",X"DD",X"E5",X"DD",X"21",X"C5",X"E1",X"DD",X"36",X"00",X"C0",X"DD",X"36",X"01",X"48",X"DD",
		X"36",X"02",X"00",X"DD",X"36",X"03",X"70",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"DD",
		X"36",X"07",X"80",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"10",X"00",X"DD",
		X"36",X"11",X"00",X"DD",X"E1",X"FD",X"36",X"0C",X"00",X"FD",X"36",X"0D",X"FF",X"21",X"01",X"E0",
		X"CB",X"C6",X"C9",X"DD",X"35",X"05",X"C0",X"DD",X"7E",X"03",X"FE",X"16",X"30",X"15",X"87",X"5F",
		X"16",X"00",X"21",X"2C",X"72",X"19",X"7E",X"DD",X"77",X"04",X"23",X"7E",X"DD",X"77",X"05",X"DD",
		X"34",X"03",X"C9",X"DD",X"34",X"02",X"DD",X"36",X"03",X"00",X"21",X"00",X"E0",X"CB",X"B6",X"C9",
		X"EF",X"01",X"FF",X"B3",X"EF",X"01",X"FF",X"EF",X"EF",X"01",X"FF",X"B3",X"EF",X"01",X"FF",X"B3",
		X"EF",X"01",X"FF",X"B3",X"FD",X"30",X"FB",X"60",X"FF",X"04",X"FB",X"18",X"FF",X"50",X"FB",X"30",
		X"FF",X"5C",X"FE",X"14",X"FD",X"28",X"FF",X"50",X"DD",X"7E",X"07",X"A7",X"28",X"04",X"DD",X"35",
		X"07",X"C9",X"DD",X"7E",X"06",X"FE",X"12",X"D0",X"FE",X"11",X"D2",X"93",X"73",X"FE",X"10",X"D2",
		X"6F",X"73",X"FE",X"07",X"D2",X"31",X"73",X"FE",X"06",X"D2",X"29",X"73",X"FE",X"01",X"30",X"44",
		X"DD",X"E5",X"DD",X"21",X"1A",X"E2",X"DD",X"36",X"00",X"C1",X"DD",X"36",X"01",X"A8",X"DD",X"36",
		X"02",X"00",X"DD",X"36",X"03",X"70",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"40",X"DD",X"36",
		X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0D",X"FF",X"DD",X"36",
		X"0E",X"FF",X"DD",X"36",X"13",X"00",X"DD",X"36",X"14",X"00",X"DD",X"E1",X"DD",X"34",X"06",X"DD",
		X"36",X"07",X"B4",X"C9",X"DD",X"7E",X"06",X"3D",X"FD",X"77",X"17",X"DD",X"E5",X"DD",X"21",X"C2",
		X"E2",X"DD",X"36",X"00",X"E1",X"DD",X"36",X"01",X"A8",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",
		X"70",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"20",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",
		X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",
		X"00",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"03",X"DD",X"36",X"0F",
		X"FF",X"DD",X"36",X"10",X"FF",X"DD",X"E1",X"DD",X"36",X"07",X"B4",X"DD",X"34",X"06",X"DD",X"7E",
		X"06",X"FE",X"06",X"D8",X"DD",X"36",X"07",X"E6",X"C9",X"DD",X"36",X"07",X"50",X"DD",X"34",X"06",
		X"C9",X"3E",X"2E",X"08",X"3E",X"09",X"01",X"02",X"02",X"11",X"29",X"8B",X"CD",X"42",X"04",X"DD",
		X"CB",X"06",X"46",X"28",X"15",X"CD",X"4F",X"05",X"DD",X"34",X"06",X"DD",X"36",X"07",X"14",X"DD",
		X"7E",X"06",X"FE",X"0F",X"D8",X"DD",X"36",X"07",X"2A",X"C9",X"01",X"0A",X"02",X"11",X"7D",X"89",
		X"CD",X"6C",X"04",X"DD",X"34",X"06",X"DD",X"36",X"07",X"08",X"AF",X"32",X"C2",X"E2",X"C9",X"DD",
		X"E5",X"DD",X"21",X"09",X"E3",X"DD",X"36",X"00",X"80",X"DD",X"36",X"01",X"A8",X"DD",X"36",X"02",
		X"00",X"DD",X"36",X"03",X"30",X"DD",X"36",X"04",X"00",X"DD",X"E1",X"DD",X"34",X"06",X"DD",X"36",
		X"07",X"46",X"C9",X"3E",X"32",X"08",X"3E",X"4D",X"01",X"02",X"02",X"11",X"25",X"8B",X"CD",X"42",
		X"04",X"DD",X"34",X"06",X"C9",X"DD",X"7E",X"02",X"FE",X"04",X"D2",X"EF",X"74",X"FE",X"03",X"30",
		X"6E",X"FE",X"02",X"30",X"3C",X"FE",X"01",X"30",X"16",X"CD",X"85",X"04",X"DD",X"36",X"01",X"04",
		X"DD",X"34",X"02",X"DD",X"36",X"03",X"00",X"3E",X"1D",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"DD",
		X"7E",X"03",X"21",X"FB",X"74",X"CD",X"25",X"04",X"DD",X"36",X"01",X"04",X"DD",X"34",X"03",X"DD",
		X"7E",X"03",X"FE",X"0F",X"D8",X"DD",X"36",X"01",X"08",X"DD",X"34",X"02",X"DD",X"36",X"03",X"00",
		X"C9",X"DD",X"7E",X"03",X"87",X"5F",X"16",X"00",X"21",X"0E",X"75",X"19",X"5E",X"23",X"56",X"EB",
		X"CD",X"03",X"04",X"DD",X"36",X"01",X"08",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"06",X"D8",
		X"DD",X"34",X"02",X"DD",X"36",X"01",X"0C",X"DD",X"36",X"03",X"48",X"DD",X"36",X"04",X"00",X"DD",
		X"7E",X"03",X"FE",X"48",X"20",X"5C",X"CD",X"B4",X"7C",X"3E",X"B6",X"08",X"3E",X"BE",X"01",X"12",
		X"04",X"11",X"E7",X"88",X"CD",X"42",X"04",X"21",X"4A",X"75",X"CD",X"03",X"04",X"3A",X"06",X"E0",
		X"FE",X"0A",X"38",X"02",X"3E",X"09",X"32",X"65",X"8E",X"3E",X"5E",X"08",X"3E",X"9B",X"01",X"04",
		X"03",X"11",X"AC",X"80",X"CD",X"42",X"04",X"3E",X"72",X"08",X"3E",X"91",X"01",X"03",X"0A",X"11",
		X"CF",X"80",X"CD",X"42",X"04",X"3E",X"91",X"01",X"04",X"06",X"11",X"31",X"81",X"CD",X"42",X"04",
		X"06",X"6D",X"0E",X"0C",X"11",X"90",X"D0",X"CD",X"9D",X"02",X"DD",X"36",X"05",X"D0",X"DD",X"36",
		X"06",X"90",X"CD",X"56",X"75",X"DD",X"7E",X"03",X"CD",X"B4",X"7C",X"A7",X"28",X"03",X"DD",X"34",
		X"03",X"DD",X"7E",X"03",X"A7",X"28",X"0C",X"FE",X"C8",X"30",X"08",X"FE",X"94",X"D8",X"DD",X"35",
		X"05",X"18",X"0A",X"DD",X"7E",X"06",X"FE",X"2C",X"38",X"11",X"DD",X"35",X"06",X"06",X"6D",X"0E",
		X"0C",X"DD",X"56",X"05",X"DD",X"5E",X"06",X"CD",X"9D",X"02",X"C9",X"21",X"0B",X"77",X"06",X"42",
		X"AF",X"86",X"23",X"10",X"FC",X"FE",X"DF",X"20",X"03",X"3A",X"06",X"E0",X"C6",X"01",X"27",X"32",
		X"06",X"E0",X"FE",X"0A",X"38",X"02",X"3E",X"09",X"32",X"65",X"8E",X"21",X"01",X"E0",X"CB",X"FE",
		X"3E",X"14",X"06",X"00",X"CD",X"D9",X"02",X"DD",X"34",X"02",X"DD",X"36",X"05",X"E0",X"C9",X"CD",
		X"56",X"75",X"DD",X"35",X"05",X"C0",X"DD",X"CB",X"00",X"AE",X"C9",X"1A",X"89",X"3E",X"0F",X"0C",
		X"18",X"17",X"10",X"1B",X"0A",X"1D",X"1E",X"15",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"1A",X"75",
		X"21",X"75",X"28",X"75",X"33",X"75",X"3A",X"75",X"42",X"75",X"D5",X"89",X"0B",X"03",X"22",X"18",
		X"1E",X"55",X"8A",X"0B",X"03",X"20",X"12",X"17",X"94",X"8A",X"2C",X"07",X"1C",X"19",X"0E",X"0C",
		X"12",X"0A",X"15",X"D2",X"89",X"0B",X"03",X"18",X"17",X"0E",X"52",X"8A",X"0B",X"04",X"16",X"18",
		X"1B",X"0E",X"91",X"8A",X"22",X"04",X"10",X"0A",X"16",X"0E",X"85",X"89",X"0B",X"08",X"0C",X"1B",
		X"0E",X"0D",X"12",X"1D",X"29",X"29",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"03",X"38",X"04",
		X"AF",X"DD",X"77",X"04",X"21",X"78",X"75",X"A7",X"28",X"0A",X"21",X"80",X"75",X"FE",X"01",X"28",
		X"03",X"21",X"88",X"75",X"CD",X"03",X"04",X"C9",X"AE",X"80",X"9B",X"04",X"60",X"63",X"66",X"69",
		X"AE",X"80",X"9B",X"04",X"6A",X"6B",X"6C",X"6D",X"AE",X"80",X"9B",X"04",X"6E",X"6F",X"70",X"71",
		X"DD",X"7E",X"02",X"FE",X"04",X"D2",X"0B",X"77",X"FE",X"03",X"D2",X"FD",X"76",X"FE",X"02",X"D2",
		X"D6",X"76",X"FE",X"01",X"D2",X"99",X"76",X"DD",X"34",X"02",X"CD",X"85",X"04",X"DD",X"36",X"03",
		X"00",X"DD",X"36",X"04",X"C0",X"DD",X"36",X"05",X"00",X"DD",X"36",X"06",X"00",X"DD",X"7E",X"04",
		X"CB",X"2F",X"CD",X"B4",X"7C",X"3E",X"51",X"01",X"20",X"0A",X"21",X"03",X"80",X"CD",X"5C",X"04",
		X"3E",X"64",X"01",X"20",X"0A",X"21",X"03",X"84",X"CD",X"5C",X"04",X"3E",X"09",X"01",X"16",X"05",
		X"21",X"0D",X"80",X"CD",X"5C",X"04",X"3E",X"A5",X"01",X"16",X"05",X"21",X"0D",X"84",X"CD",X"5C",
		X"04",X"3E",X"0B",X"01",X"20",X"0B",X"21",X"12",X"80",X"CD",X"5C",X"04",X"3E",X"2F",X"01",X"20",
		X"0B",X"21",X"12",X"84",X"CD",X"5C",X"04",X"3E",X"2E",X"08",X"3E",X"0B",X"01",X"11",X"02",X"11",
		X"10",X"80",X"CD",X"42",X"04",X"3E",X"6C",X"01",X"04",X"03",X"11",X"2D",X"82",X"CD",X"42",X"04",
		X"3E",X"2C",X"01",X"04",X"02",X"11",X"30",X"82",X"CD",X"42",X"04",X"3E",X"51",X"01",X"0A",X"05",
		X"11",X"A8",X"82",X"CD",X"42",X"04",X"3E",X"09",X"01",X"06",X"03",X"11",X"CD",X"82",X"CD",X"42",
		X"04",X"3E",X"0B",X"01",X"04",X"04",X"11",X"B0",X"82",X"CD",X"42",X"04",X"3E",X"6C",X"01",X"03",
		X"02",X"11",X"30",X"83",X"CD",X"42",X"04",X"3E",X"0B",X"01",X"03",X"02",X"11",X"32",X"83",X"CD",
		X"42",X"04",X"3E",X"6C",X"01",X"04",X"05",X"11",X"8D",X"83",X"CD",X"42",X"04",X"3E",X"2C",X"01",
		X"04",X"02",X"11",X"92",X"83",X"CD",X"42",X"04",X"3E",X"82",X"08",X"3E",X"89",X"01",X"04",X"06",
		X"11",X"08",X"89",X"CD",X"42",X"04",X"3E",X"89",X"01",X"02",X"01",X"21",X"2C",X"89",X"CD",X"5C",
		X"04",X"3E",X"1E",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",
		X"A4",X"30",X"0D",X"CD",X"4D",X"77",X"CD",X"85",X"77",X"CD",X"91",X"78",X"CD",X"52",X"79",X"C9",
		X"DD",X"34",X"02",X"DD",X"36",X"03",X"00",X"DD",X"36",X"06",X"DC",X"3E",X"E0",X"08",X"3E",X"51",
		X"01",X"04",X"01",X"11",X"AC",X"82",X"CD",X"42",X"04",X"3E",X"09",X"01",X"04",X"02",X"11",X"AD",
		X"82",X"CD",X"42",X"04",X"18",X"0A",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"90",X"30",X"0A",
		X"CD",X"EA",X"77",X"CD",X"07",X"79",X"CD",X"52",X"79",X"C9",X"FD",X"34",X"00",X"CD",X"AA",X"05",
		X"21",X"01",X"E0",X"CB",X"FE",X"DD",X"34",X"02",X"DD",X"36",X"03",X"00",X"C9",X"CD",X"07",X"79",
		X"CD",X"52",X"79",X"DD",X"34",X"03",X"C0",X"DD",X"34",X"02",X"C9",X"CD",X"07",X"79",X"CD",X"52",
		X"79",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"24",X"D8",X"11",X"70",X"8C",X"3E",X"A5",X"12",
		X"13",X"21",X"45",X"77",X"06",X"04",X"7E",X"12",X"23",X"3A",X"03",X"98",X"E6",X"7E",X"BE",X"20",
		X"0C",X"13",X"23",X"10",X"F1",X"FD",X"34",X"1A",X"FD",X"7E",X"16",X"E6",X"02",X"FD",X"77",X"16",
		X"DD",X"CB",X"00",X"9E",X"C9",X"A5",X"40",X"C2",X"4C",X"36",X"2A",X"6F",X"66",X"DD",X"7E",X"03",
		X"FE",X"10",X"D8",X"FE",X"91",X"D0",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"CB",X"2F",X"CD",X"B4",
		X"7C",X"DD",X"7E",X"04",X"3D",X"47",X"E6",X"0F",X"C0",X"21",X"77",X"77",X"CB",X"60",X"28",X"03",
		X"21",X"7E",X"77",X"CD",X"03",X"04",X"C9",X"08",X"89",X"89",X"03",X"82",X"88",X"8E",X"08",X"89",
		X"89",X"03",X"9A",X"9B",X"9C",X"DD",X"7E",X"03",X"FE",X"88",X"D8",X"20",X"2A",X"3E",X"9D",X"08",
		X"3E",X"89",X"01",X"02",X"03",X"11",X"49",X"89",X"CD",X"42",X"04",X"DD",X"36",X"07",X"05",X"DD",
		X"36",X"08",X"58",X"DD",X"36",X"09",X"00",X"DD",X"36",X"0A",X"60",X"DD",X"36",X"0B",X"00",X"DD",
		X"36",X"0C",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"34",X"08",X"DD",X"34",X"08",X"DD",X"CB",X"07",
		X"46",X"28",X"13",X"DD",X"35",X"0A",X"DD",X"35",X"0A",X"DD",X"7E",X"0A",X"FE",X"41",X"30",X"0C",
		X"DD",X"CB",X"07",X"86",X"18",X"06",X"DD",X"34",X"0A",X"DD",X"34",X"0A",X"06",X"78",X"0E",X"06",
		X"DD",X"56",X"08",X"DD",X"5E",X"0A",X"CD",X"9D",X"02",X"C9",X"DD",X"7E",X"03",X"FE",X"78",X"30",
		X"60",X"FE",X"3C",X"28",X"19",X"A7",X"20",X"35",X"DD",X"36",X"07",X"04",X"DD",X"36",X"08",X"26",
		X"DD",X"36",X"0A",X"18",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0D",X"10",X"18",X"1C",X"FD",X"7E",
		X"00",X"FE",X"06",X"38",X"02",X"3E",X"05",X"87",X"87",X"C6",X"0A",X"DD",X"77",X"08",X"DD",X"36",
		X"0A",X"0A",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0D",X"30",X"CD",X"B2",X"2C",X"DD",X"E5",X"DD",
		X"21",X"BD",X"E1",X"DD",X"34",X"07",X"DD",X"35",X"05",X"20",X"0C",X"DD",X"7E",X"06",X"E6",X"0F",
		X"FE",X"0A",X"30",X"03",X"CD",X"5B",X"2C",X"FD",X"E5",X"CD",X"7C",X"2B",X"FD",X"E1",X"DD",X"E1",
		X"C9",X"DD",X"7E",X"03",X"FE",X"78",X"20",X"16",X"DD",X"CB",X"08",X"26",X"DD",X"CB",X"08",X"26",
		X"DD",X"CB",X"0A",X"26",X"DD",X"CB",X"0A",X"26",X"DD",X"36",X"0C",X"00",X"18",X"06",X"DD",X"35",
		X"0A",X"DD",X"34",X"0C",X"DD",X"7E",X"0C",X"E6",X"18",X"0F",X"0F",X"0F",X"FE",X"03",X"20",X"02",
		X"3E",X"01",X"C6",X"06",X"47",X"0E",X"02",X"DD",X"56",X"08",X"DD",X"5E",X"0A",X"CD",X"9D",X"02",
		X"C9",X"DD",X"7E",X"03",X"FE",X"04",X"D8",X"DD",X"7E",X"05",X"DD",X"34",X"05",X"FE",X"3C",X"30",
		X"10",X"47",X"E6",X"03",X"C0",X"78",X"E6",X"3C",X"0F",X"0F",X"21",X"CB",X"78",X"CD",X"25",X"04",
		X"C9",X"47",X"E6",X"07",X"C0",X"78",X"D6",X"40",X"E6",X"18",X"0F",X"0F",X"5F",X"16",X"00",X"21",
		X"DE",X"78",X"19",X"5E",X"23",X"56",X"EB",X"CD",X"03",X"04",X"C9",X"1A",X"89",X"3E",X"0F",X"0C",
		X"18",X"17",X"10",X"1B",X"0A",X"1D",X"1E",X"15",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"E6",X"78",
		X"ED",X"78",X"F4",X"78",X"FD",X"78",X"18",X"89",X"00",X"03",X"22",X"18",X"1E",X"98",X"89",X"00",
		X"03",X"20",X"12",X"17",X"77",X"89",X"00",X"05",X"0E",X"21",X"1D",X"1B",X"0A",X"37",X"8A",X"2E",
		X"06",X"60",X"61",X"62",X"63",X"64",X"65",X"DD",X"34",X"06",X"DD",X"7E",X"02",X"FE",X"03",X"30",
		X"05",X"DD",X"CB",X"06",X"7E",X"C0",X"DD",X"7E",X"06",X"E6",X"0F",X"C0",X"DD",X"CB",X"06",X"66",
		X"20",X"18",X"3E",X"A3",X"08",X"3E",X"D1",X"01",X"03",X"03",X"11",X"EA",X"89",X"CD",X"42",X"04",
		X"01",X"03",X"02",X"11",X"E8",X"89",X"CD",X"6C",X"04",X"C9",X"3E",X"AC",X"08",X"3E",X"D1",X"01",
		X"03",X"03",X"11",X"E8",X"89",X"CD",X"42",X"04",X"01",X"03",X"02",X"11",X"EB",X"89",X"CD",X"6C",
		X"04",X"C9",X"DD",X"7E",X"03",X"E6",X"1F",X"28",X"0D",X"FE",X"14",X"C0",X"01",X"0A",X"02",X"11",
		X"7D",X"89",X"CD",X"6C",X"04",X"C9",X"CD",X"4F",X"05",X"C9",X"DD",X"7E",X"02",X"FE",X"05",X"D2",
		X"51",X"7A",X"FE",X"04",X"D2",X"04",X"7A",X"FE",X"03",X"D2",X"F9",X"79",X"FE",X"02",X"30",X"5F",
		X"DD",X"34",X"02",X"DD",X"36",X"01",X"1E",X"DD",X"36",X"03",X"00",X"DD",X"36",X"05",X"00",X"CD",
		X"85",X"04",X"FD",X"35",X"04",X"FD",X"35",X"04",X"FD",X"E5",X"E1",X"11",X"1C",X"00",X"19",X"11",
		X"BA",X"88",X"CD",X"38",X"7C",X"FD",X"34",X"04",X"01",X"07",X"00",X"09",X"1B",X"1B",X"CD",X"38",
		X"7C",X"FD",X"34",X"04",X"01",X"07",X"00",X"09",X"1B",X"1B",X"CD",X"38",X"7C",X"21",X"5D",X"7A",
		X"CD",X"03",X"04",X"DD",X"7E",X"03",X"CD",X"B4",X"7C",X"3E",X"A8",X"08",X"3E",X"95",X"01",X"04",
		X"04",X"11",X"08",X"80",X"CD",X"42",X"04",X"3E",X"1F",X"06",X"00",X"CD",X"D9",X"02",X"C9",X"DD",
		X"35",X"03",X"DD",X"7E",X"03",X"CD",X"B4",X"7C",X"CD",X"6C",X"7A",X"DD",X"7E",X"03",X"FE",X"98",
		X"C0",X"DD",X"34",X"02",X"DD",X"36",X"04",X"3C",X"C9",X"CD",X"6C",X"7A",X"DD",X"35",X"04",X"C0",
		X"DD",X"34",X"02",X"C9",X"DD",X"7E",X"03",X"FE",X"68",X"28",X"14",X"FE",X"98",X"20",X"29",X"3E",
		X"B8",X"08",X"3E",X"89",X"01",X"04",X"04",X"11",X"68",X"82",X"CD",X"42",X"04",X"18",X"19",X"3E",
		X"C8",X"08",X"3E",X"91",X"01",X"04",X"04",X"11",X"A8",X"81",X"CD",X"42",X"04",X"3E",X"89",X"01",
		X"04",X"05",X"11",X"28",X"81",X"CD",X"42",X"04",X"DD",X"35",X"03",X"DD",X"7E",X"03",X"CD",X"B4",
		X"7C",X"CD",X"6C",X"7A",X"DD",X"7E",X"03",X"A7",X"C0",X"DD",X"34",X"02",X"DD",X"36",X"04",X"4A",
		X"C9",X"CD",X"6C",X"7A",X"DD",X"35",X"04",X"C0",X"DD",X"36",X"02",X"00",X"C9",X"51",X"89",X"2C",
		X"0B",X"1F",X"0E",X"1B",X"22",X"29",X"10",X"18",X"18",X"0D",X"29",X"25",X"DD",X"34",X"05",X"DD",
		X"7E",X"05",X"E6",X"0F",X"C0",X"DD",X"CB",X"05",X"66",X"20",X"19",X"21",X"AD",X"7A",X"CD",X"03",
		X"04",X"DD",X"7E",X"03",X"FE",X"98",X"D0",X"CD",X"D4",X"03",X"DD",X"7E",X"03",X"FE",X"48",X"D0",
		X"CD",X"D4",X"03",X"C9",X"21",X"C7",X"7A",X"CD",X"03",X"04",X"DD",X"7E",X"03",X"FE",X"98",X"D0",
		X"CD",X"D4",X"03",X"DD",X"7E",X"03",X"FE",X"48",X"D0",X"CD",X"D4",X"03",X"C9",X"08",X"80",X"95",
		X"04",X"A8",X"AC",X"B0",X"B4",X"88",X"82",X"89",X"03",X"02",X"BC",X"BD",X"C0",X"C1",X"C4",X"C5",
		X"28",X"81",X"89",X"01",X"02",X"D8",X"D9",X"08",X"80",X"15",X"04",X"F9",X"FA",X"FB",X"FC",X"88",
		X"82",X"89",X"03",X"02",X"EC",X"ED",X"EE",X"EF",X"F0",X"F1",X"28",X"81",X"89",X"01",X"02",X"F2",
		X"F3",X"DD",X"7E",X"02",X"FE",X"07",X"D2",X"A7",X"7B",X"CD",X"85",X"04",X"CD",X"A1",X"06",X"3A",
		X"83",X"80",X"01",X"02",X"02",X"21",X"CF",X"81",X"CD",X"5C",X"04",X"3A",X"83",X"84",X"01",X"02",
		X"02",X"21",X"CF",X"85",X"CD",X"5C",X"04",X"11",X"2A",X"81",X"01",X"0D",X"03",X"CD",X"6C",X"04",
		X"11",X"93",X"80",X"01",X"18",X"0A",X"CD",X"6C",X"04",X"FD",X"E5",X"E1",X"11",X"2A",X"00",X"19",
		X"11",X"BA",X"88",X"CD",X"38",X"7C",X"21",X"B0",X"7B",X"CD",X"03",X"04",X"CD",X"03",X"04",X"CD",
		X"03",X"04",X"FD",X"E5",X"E1",X"23",X"11",X"B7",X"89",X"0E",X"2C",X"CD",X"A1",X"03",X"23",X"0E",
		X"2C",X"CD",X"90",X"7C",X"FD",X"E5",X"E1",X"23",X"11",X"91",X"E0",X"01",X"03",X"00",X"ED",X"B0",
		X"FD",X"46",X"04",X"CD",X"D3",X"7B",X"21",X"94",X"E0",X"11",X"B5",X"89",X"0E",X"22",X"CD",X"A1",
		X"03",X"FD",X"56",X"05",X"FD",X"5E",X"06",X"CD",X"1E",X"7C",X"21",X"91",X"E0",X"36",X"00",X"23",
		X"72",X"23",X"73",X"FD",X"46",X"04",X"CD",X"D3",X"7B",X"21",X"94",X"E0",X"11",X"91",X"E0",X"01",
		X"03",X"00",X"ED",X"B0",X"06",X"60",X"CD",X"D3",X"7B",X"21",X"92",X"E0",X"3A",X"96",X"E0",X"77",
		X"11",X"75",X"8A",X"0E",X"22",X"CD",X"90",X"7C",X"3E",X"1F",X"06",X"00",X"CD",X"D9",X"02",X"DD",
		X"34",X"02",X"DD",X"36",X"01",X"F0",X"C9",X"DD",X"36",X"02",X"00",X"DD",X"36",X"01",X"B4",X"C9",
		X"B7",X"88",X"2C",X"05",X"1D",X"18",X"1D",X"0A",X"15",X"B5",X"88",X"22",X"07",X"0A",X"1F",X"0E",
		X"1B",X"0A",X"10",X"0E",X"4B",X"89",X"3E",X"0B",X"20",X"18",X"17",X"0D",X"0E",X"1B",X"0F",X"1E",
		X"15",X"29",X"25",X"21",X"93",X"E0",X"11",X"94",X"E0",X"AF",X"12",X"13",X"12",X"13",X"12",X"B8",
		X"20",X"02",X"06",X"99",X"7E",X"90",X"27",X"77",X"2B",X"7E",X"DE",X"00",X"27",X"77",X"2B",X"7E",
		X"DE",X"00",X"27",X"77",X"23",X"23",X"38",X"15",X"1A",X"C6",X"01",X"27",X"12",X"1B",X"1A",X"CE",
		X"00",X"27",X"12",X"1B",X"1A",X"CE",X"00",X"27",X"12",X"13",X"13",X"18",X"D7",X"7E",X"80",X"27",
		X"77",X"2B",X"7E",X"CE",X"00",X"27",X"77",X"2B",X"7E",X"CE",X"00",X"27",X"77",X"C9",X"06",X"3C",
		X"21",X"00",X"00",X"7A",X"CD",X"2F",X"7C",X"10",X"FA",X"7B",X"CD",X"2F",X"7C",X"EB",X"C9",X"85",
		X"27",X"6F",X"7C",X"CE",X"00",X"27",X"67",X"C9",X"D5",X"E5",X"21",X"89",X"7C",X"CD",X"07",X"04",
		X"21",X"C0",X"00",X"19",X"EB",X"FD",X"E5",X"E1",X"01",X"04",X"00",X"09",X"AF",X"06",X"02",X"0E",
		X"09",X"CD",X"A4",X"03",X"E1",X"E5",X"0E",X"09",X"CD",X"A1",X"03",X"0E",X"09",X"CD",X"90",X"7C",
		X"23",X"7B",X"E6",X"1F",X"87",X"87",X"87",X"C6",X"04",X"5F",X"16",X"D0",X"7E",X"A7",X"28",X"0E",
		X"87",X"4F",X"06",X"00",X"21",X"7F",X"7C",X"09",X"46",X"23",X"4E",X"CD",X"9D",X"02",X"E1",X"D1",
		X"C9",X"2D",X"02",X"6E",X"0D",X"69",X"07",X"51",X"04",X"09",X"05",X"1C",X"0C",X"0E",X"17",X"0E",
		X"E5",X"21",X"20",X"00",X"19",X"EB",X"E1",X"AF",X"06",X"02",X"CD",X"A4",X"03",X"79",X"12",X"E5",
		X"21",X"00",X"04",X"19",X"36",X"2D",X"21",X"20",X"00",X"19",X"EB",X"E1",X"3E",X"80",X"06",X"02",
		X"CD",X"A4",X"03",X"C9",X"21",X"00",X"E0",X"CB",X"46",X"28",X"02",X"ED",X"44",X"32",X"00",X"F8",
		X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"3F",X"0D",X"21",X"00",X"4F",X"0F",X"B1",X"00",X"CF",X"12",X"B1",X"00",X"CF",X"11",
		X"B1",X"00",X"CF",X"0F",X"B1",X"00",X"CF",X"14",X"71",X"00",X"7F",X"14",X"71",X"00",X"7F",X"14",
		X"B1",X"00",X"CF",X"16",X"B1",X"00",X"CF",X"11",X"B1",X"00",X"CF",X"12",X"B1",X"00",X"CF",X"0F",
		X"71",X"00",X"7F",X"0F",X"71",X"00",X"7F",X"0F",X"B1",X"00",X"CF",X"12",X"B1",X"00",X"CF",X"11",
		X"B1",X"00",X"CF",X"0F",X"B1",X"00",X"CF",X"0D",X"B1",X"00",X"CF",X"19",X"B1",X"00",X"CF",X"18",
		X"B1",X"00",X"CF",X"16",X"B1",X"00",X"CF",X"14",X"B1",X"00",X"CF",X"12",X"B1",X"00",X"CF",X"11",
		X"B1",X"00",X"CF",X"0F",X"B1",X"00",X"CF",X"80",X"D3",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"3F",X"1D",X"B3",X"00",X"CF",X"20",X"B3",X"00",X"CF",X"1D",X"B3",X"00",X"CF",X"20",
		X"B3",X"00",X"CF",X"1E",X"B3",X"00",X"CF",X"1B",X"B3",X"00",X"CF",X"20",X"B3",X"00",X"CF",X"1E",
		X"B3",X"00",X"CF",X"1D",X"B3",X"00",X"CF",X"19",X"B3",X"00",X"CF",X"1D",X"B3",X"00",X"CF",X"19",
		X"B3",X"00",X"CF",X"1D",X"B3",X"00",X"CF",X"1E",X"B3",X"00",X"CF",X"19",X"B3",X"00",X"CF",X"1B",
		X"B3",X"00",X"CF",X"1E",X"B3",X"00",X"CF",X"20",X"B3",X"00",X"CF",X"1E",X"B3",X"00",X"CF",X"20",
		X"B3",X"00",X"CF",X"1E",X"B3",X"00",X"CF",X"1B",X"B3",X"00",X"CF",X"20",X"B3",X"00",X"CF",X"1E",
		X"B3",X"00",X"CF",X"1D",X"B3",X"00",X"CF",X"14",X"B3",X"00",X"CF",X"1B",X"B3",X"00",X"CF",X"1E",
		X"B3",X"00",X"CF",X"1D",X"B3",X"00",X"CF",X"1B",X"B3",X"00",X"CF",X"19",X"B3",X"00",X"CF",X"1E",
		X"B3",X"00",X"CF",X"80",X"43",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
