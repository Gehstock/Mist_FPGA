library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bios is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bios is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"13",X"E0",X"C3",X"55",X"E8",X"C3",X"CB",X"F1",X"C3",X"72",X"E2",X"C3",X"CC",X"E2",X"C3",
		X"F5",X"F1",X"32",X"F3",X"3E",X"AA",X"D3",X"10",X"D3",X"11",X"D3",X"12",X"D3",X"13",X"3E",X"80",
		X"D3",X"6B",X"3E",X"30",X"D3",X"63",X"3E",X"76",X"D3",X"63",X"3E",X"94",X"D3",X"63",X"3E",X"0D",
		X"D3",X"62",X"3E",X"90",X"D3",X"47",X"3E",X"F0",X"D3",X"46",X"3E",X"15",X"D3",X"79",X"3E",X"40",
		X"D3",X"79",X"3E",X"FE",X"D3",X"79",X"3E",X"16",X"D3",X"74",X"3E",X"DF",X"D3",X"75",X"3E",X"FF",
		X"D3",X"75",X"AF",X"D3",X"6A",X"32",X"FE",X"DF",X"32",X"FF",X"DF",X"3E",X"C3",X"32",X"04",X"DF",
		X"21",X"13",X"E0",X"22",X"05",X"DF",X"FB",X"01",X"00",X"60",X"3E",X"E9",X"D3",X"61",X"3E",X"07",
		X"D3",X"61",X"3E",X"15",X"D3",X"79",X"0B",X"79",X"B0",X"C2",X"76",X"E0",X"3E",X"25",X"D3",X"79",
		X"01",X"FF",X"FF",X"0B",X"79",X"B0",X"C2",X"83",X"E0",X"31",X"00",X"DF",X"CD",X"66",X"EE",X"01",
		X"20",X"DF",X"21",X"26",X"DF",X"CD",X"55",X"F0",X"7A",X"FE",X"DC",X"CC",X"3C",X"F8",X"3A",X"FF",
		X"DF",X"B7",X"C2",X"9E",X"E0",X"31",X"00",X"DF",X"CD",X"10",X"FF",X"3E",X"25",X"D3",X"79",X"3E",
		X"FF",X"D3",X"75",X"3E",X"20",X"D3",X"74",X"CD",X"04",X"E9",X"21",X"19",X"E1",X"CD",X"C2",X"E3",
		X"21",X"25",X"E1",X"CD",X"C2",X"E3",X"31",X"00",X"DF",X"21",X"8C",X"E1",X"CD",X"C2",X"E3",X"CD",
		X"72",X"E2",X"21",X"C6",X"E0",X"E5",X"FE",X"3F",X"CA",X"AB",X"E0",X"FE",X"0D",X"C8",X"FE",X"53",
		X"CA",X"05",X"E2",X"FE",X"52",X"CA",X"53",X"E2",X"FE",X"57",X"CA",X"5A",X"E2",X"FE",X"4C",X"CA",
		X"6A",X"E3",X"FE",X"47",X"CA",X"41",X"E2",X"FE",X"59",X"CA",X"53",X"E3",X"FE",X"55",X"CA",X"60",
		X"E3",X"CD",X"07",X"E1",X"C3",X"C6",X"E0",X"21",X"0D",X"E1",X"C3",X"C2",X"E3",X"0D",X"0A",X"2D",
		X"DE",X"E8",X"D8",X"D1",X"DA",X"D0",X"2D",X"0D",X"00",X"1B",X"42",X"B7",X"B0",X"B3",X"C0",X"C3",
		X"B7",X"C7",X"B8",X"BA",X"00",X"C4",X"E3",X"DD",X"DA",X"E6",X"D8",X"D8",X"3A",X"0D",X"0A",X"53",
		X"2D",X"E3",X"E1",X"E2",X"D0",X"DD",X"DE",X"D2",X"DA",X"D0",X"20",X"EF",X"E7",X"D5",X"D9",X"DA",
		X"D8",X"0D",X"0A",X"4C",X"2D",X"D7",X"D0",X"D3",X"E0",X"E3",X"D7",X"DA",X"D0",X"20",X"D8",X"D7",
		X"20",X"BF",X"B7",X"C3",X"0D",X"0A",X"52",X"2D",X"E7",X"E2",X"D5",X"DD",X"D8",X"D5",X"20",X"E1",
		X"20",X"BC",X"BB",X"0D",X"0A",X"57",X"2D",X"D7",X"D0",X"DF",X"D8",X"E1",X"EC",X"20",X"DD",X"D0",
		X"20",X"BC",X"BB",X"0D",X"0A",X"47",X"2D",X"D2",X"EB",X"DF",X"DE",X"DB",X"DD",X"D8",X"E2",X"EC",
		X"20",X"DF",X"E0",X"DE",X"D3",X"E0",X"D0",X"DC",X"DC",X"E3",X"0D",X"00",X"0A",X"3E",X"00",X"0D",
		X"0A",X"BF",X"DE",X"D4",X"D3",X"DE",X"E2",X"DE",X"D2",X"EC",X"E2",X"D5",X"20",X"DC",X"D0",X"D3",
		X"DD",X"D8",X"E2",X"DE",X"E4",X"DE",X"DD",X"20",X"D4",X"DB",X"EF",X"20",X"00",X"B7",X"B0",X"BF",
		X"B8",X"C1",X"B8",X"00",X"C7",X"C2",X"B5",X"BD",X"B8",X"CF",X"00",X"0D",X"0A",X"D8",X"20",X"DD",
		X"D0",X"D6",X"DC",X"D8",X"E2",X"D5",X"20",X"3C",X"B2",X"BA",X"3E",X"00",X"0A",X"2A",X"B7",X"B0",
		X"BF",X"B8",X"C1",X"CC",X"2A",X"0D",X"00",X"0A",X"2A",X"C7",X"C2",X"B5",X"BD",X"B8",X"B5",X"2A",
		X"0D",X"00",X"0A",X"2A",X"DE",X"E8",X"D8",X"D1",X"DA",X"D0",X"20",X"BA",X"C1",X"2A",X"0D",X"00",
		X"0A",X"D2",X"EB",X"DA",X"DB",X"EE",X"E7",X"D8",X"20",X"DC",X"D0",X"D3",X"DD",X"D8",X"E2",X"DE",
		X"E4",X"DE",X"DD",X"0D",X"00",X"CD",X"CC",X"E2",X"3D",X"C2",X"01",X"E1",X"2A",X"1A",X"DF",X"CD",
		X"41",X"E3",X"E5",X"CD",X"46",X"E3",X"CD",X"4E",X"E3",X"E1",X"7E",X"E5",X"CD",X"D5",X"E3",X"CD",
		X"4E",X"E3",X"CD",X"72",X"E2",X"E1",X"FE",X"0D",X"CA",X"3D",X"E2",X"FE",X"2E",X"C8",X"E5",X"CD",
		X"CF",X"E2",X"2A",X"1A",X"DF",X"7C",X"B7",X"C2",X"01",X"E1",X"7D",X"E1",X"77",X"23",X"C3",X"0F",
		X"E2",X"CD",X"CC",X"E2",X"3D",X"C2",X"01",X"E1",X"31",X"00",X"DF",X"21",X"C6",X"E0",X"E5",X"2A",
		X"1A",X"DF",X"E9",X"CD",X"61",X"E2",X"CD",X"E2",X"EF",X"C9",X"CD",X"61",X"E2",X"CD",X"A8",X"EF",
		X"C9",X"CD",X"CC",X"E2",X"FE",X"02",X"C2",X"01",X"E1",X"2A",X"1A",X"DF",X"44",X"4D",X"2A",X"1C",
		X"DF",X"C9",X"11",X"DA",X"DF",X"06",X"00",X"CD",X"6F",X"E4",X"FE",X"0D",X"CA",X"89",X"E2",X"FE",
		X"7F",X"CA",X"9D",X"E2",X"FE",X"20",X"DA",X"77",X"E2",X"CD",X"CE",X"E3",X"12",X"13",X"FE",X"0D",
		X"CA",X"AC",X"E2",X"04",X"78",X"FE",X"20",X"CA",X"AC",X"E2",X"C3",X"77",X"E2",X"AF",X"B0",X"CA",
		X"77",X"E2",X"05",X"1B",X"3E",X"7F",X"CD",X"CE",X"E3",X"C3",X"77",X"E2",X"21",X"DA",X"DF",X"22",
		X"17",X"DF",X"78",X"32",X"16",X"DF",X"E5",X"21",X"16",X"DF",X"7E",X"B7",X"3E",X"0D",X"CA",X"CA",
		X"E2",X"35",X"2A",X"17",X"DF",X"7E",X"23",X"22",X"17",X"DF",X"E1",X"C9",X"CD",X"B6",X"E2",X"21",
		X"19",X"DF",X"36",X"00",X"23",X"FE",X"0D",X"CA",X"01",X"E3",X"CD",X"08",X"E3",X"CD",X"20",X"E3",
		X"FE",X"0D",X"CA",X"01",X"E3",X"CD",X"B6",X"E2",X"CD",X"08",X"E3",X"CD",X"20",X"E3",X"FE",X"0D",
		X"CA",X"01",X"E3",X"CD",X"B6",X"E2",X"CD",X"08",X"E3",X"CD",X"20",X"E3",X"FE",X"0D",X"C2",X"01",
		X"E1",X"11",X"19",X"DF",X"1A",X"13",X"B7",X"C9",X"EB",X"21",X"00",X"00",X"CD",X"2B",X"E3",X"29",
		X"29",X"29",X"29",X"B5",X"6F",X"CD",X"B6",X"E2",X"CD",X"38",X"E3",X"C2",X"0C",X"E3",X"EB",X"C9",
		X"73",X"23",X"72",X"23",X"E5",X"21",X"19",X"DF",X"34",X"E1",X"C9",X"D6",X"30",X"FE",X"0A",X"D8",
		X"C6",X"F9",X"FE",X"10",X"D8",X"C3",X"01",X"E1",X"FE",X"0D",X"C8",X"FE",X"2C",X"C8",X"FE",X"20",
		X"C9",X"3E",X"0A",X"C3",X"CE",X"E3",X"7C",X"CD",X"D5",X"E3",X"7D",X"C3",X"D5",X"E3",X"3E",X"20",
		X"C3",X"CE",X"E3",X"CD",X"61",X"E2",X"CD",X"44",X"E4",X"CD",X"F1",X"E3",X"C2",X"07",X"E1",X"C9",
		X"CD",X"61",X"E2",X"CD",X"44",X"E4",X"CD",X"1C",X"E4",X"C9",X"CD",X"CC",X"E2",X"FE",X"03",X"C2",
		X"01",X"E1",X"2A",X"1A",X"DF",X"44",X"4D",X"2A",X"1C",X"DF",X"E5",X"2A",X"1E",X"DF",X"54",X"5D",
		X"E1",X"3E",X"90",X"D3",X"47",X"7B",X"D3",X"45",X"7A",X"F6",X"C0",X"D3",X"46",X"7A",X"E6",X"C0",
		X"C2",X"A1",X"E3",X"3E",X"0C",X"D3",X"47",X"DB",X"44",X"F5",X"3E",X"0D",X"D3",X"47",X"C3",X"AC",
		X"E3",X"3E",X"0E",X"D3",X"47",X"DB",X"44",X"F5",X"3E",X"0F",X"D3",X"47",X"F1",X"02",X"13",X"CD",
		X"B6",X"E3",X"DA",X"85",X"E3",X"C9",X"78",X"94",X"DA",X"BF",X"E3",X"C0",X"79",X"95",X"D0",X"03",
		X"37",X"C9",X"F5",X"7E",X"CD",X"CE",X"E3",X"23",X"B7",X"C2",X"C3",X"E3",X"F1",X"C9",X"C5",X"4F",
		X"CD",X"D7",X"E7",X"C1",X"C9",X"F5",X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",X"CD",X"E2",X"E3",X"F1",
		X"E6",X"0F",X"FE",X"0A",X"D2",X"EC",X"E3",X"C6",X"30",X"C3",X"CE",X"E3",X"C6",X"37",X"C3",X"CE",
		X"E3",X"C5",X"CD",X"65",X"E4",X"C0",X"DB",X"78",X"B7",X"C0",X"CD",X"65",X"E4",X"C0",X"DB",X"78",
		X"FE",X"FF",X"C0",X"CD",X"65",X"E4",X"C0",X"DB",X"78",X"02",X"CD",X"B6",X"E3",X"DA",X"03",X"E4",
		X"CD",X"65",X"E4",X"C0",X"DB",X"78",X"C1",X"CD",X"55",X"F0",X"BA",X"C9",X"C5",X"CD",X"55",X"F0",
		X"C1",X"D5",X"CD",X"5D",X"E4",X"AF",X"D3",X"78",X"CD",X"5D",X"E4",X"3E",X"FF",X"D3",X"78",X"CD",
		X"5D",X"E4",X"0A",X"D3",X"78",X"CD",X"B6",X"E3",X"DA",X"2F",X"E4",X"CD",X"5D",X"E4",X"DB",X"78",
		X"F1",X"D3",X"78",X"C9",X"3E",X"96",X"D3",X"63",X"3E",X"07",X"D3",X"62",X"3E",X"15",X"D3",X"79",
		X"3E",X"40",X"D3",X"79",X"3E",X"FE",X"D3",X"79",X"3E",X"27",X"D3",X"79",X"C9",X"DB",X"79",X"E6",
		X"05",X"CA",X"5D",X"E4",X"C9",X"DB",X"79",X"E6",X"3A",X"CA",X"65",X"E4",X"FE",X"02",X"C9",X"C5",
		X"D5",X"3E",X"FF",X"32",X"D7",X"DF",X"CD",X"AF",X"E4",X"FE",X"FF",X"CA",X"76",X"E4",X"4F",X"3A",
		X"45",X"DF",X"B7",X"CA",X"9D",X"E4",X"11",X"00",X"08",X"CD",X"FC",X"E6",X"CA",X"96",X"E4",X"1B",
		X"7B",X"B2",X"C2",X"89",X"E4",X"2F",X"32",X"45",X"DF",X"79",X"D1",X"C1",X"C9",X"11",X"00",X"20",
		X"C3",X"89",X"E4",X"AF",X"32",X"D7",X"DF",X"CD",X"AF",X"E4",X"FE",X"FF",X"C0",X"2F",X"C9",X"C5",
		X"D5",X"E5",X"3A",X"25",X"DF",X"B7",X"CA",X"CB",X"E4",X"2A",X"6E",X"DF",X"7E",X"32",X"25",X"DF",
		X"B7",X"CA",X"AC",X"E6",X"23",X"22",X"6E",X"DF",X"C3",X"B4",X"E6",X"3E",X"04",X"F5",X"06",X"58",
		X"16",X"00",X"1E",X"7F",X"21",X"01",X"28",X"F3",X"3E",X"02",X"D3",X"6A",X"4E",X"3A",X"FE",X"DF",
		X"D3",X"6A",X"FB",X"3E",X"01",X"F5",X"A1",X"C2",X"09",X"E5",X"14",X"7A",X"B8",X"FA",X"F5",X"E4",
		X"16",X"00",X"C3",X"13",X"E5",X"F1",X"07",X"D2",X"E5",X"E4",X"7D",X"07",X"D2",X"05",X"E5",X"21",
		X"01",X"29",X"C3",X"D7",X"E4",X"6F",X"C3",X"D7",X"E4",X"7B",X"FE",X"7F",X"C2",X"13",X"E5",X"5A",
		X"C3",X"EA",X"E4",X"F1",X"3A",X"D6",X"DF",X"BA",X"7A",X"32",X"D6",X"DF",X"CA",X"23",X"E5",X"F1",
		X"C3",X"CB",X"E4",X"F1",X"3D",X"C2",X"CD",X"E4",X"7B",X"FE",X"7F",X"CA",X"B2",X"E6",X"7A",X"B7",
		X"CA",X"63",X"E5",X"FE",X"38",X"FA",X"B2",X"E6",X"FE",X"40",X"7B",X"FA",X"4F",X"E5",X"FE",X"38",
		X"FA",X"B2",X"E6",X"FE",X"40",X"F2",X"B2",X"E6",X"CD",X"C7",X"E6",X"5A",X"C3",X"30",X"E6",X"FE",
		X"38",X"FA",X"5C",X"E5",X"FE",X"40",X"F2",X"B2",X"E6",X"C3",X"8B",X"E6",X"7A",X"CD",X"C7",X"E6",
		X"C3",X"7A",X"E5",X"06",X"00",X"7B",X"FE",X"38",X"FA",X"7A",X"E5",X"FE",X"40",X"F2",X"30",X"E6",
		X"FE",X"3C",X"C2",X"B2",X"E6",X"3E",X"1B",X"C3",X"B4",X"E6",X"16",X"00",X"3A",X"26",X"DF",X"4F",
		X"A8",X"E6",X"04",X"CA",X"8C",X"E5",X"2A",X"27",X"DF",X"C3",X"DF",X"E5",X"21",X"87",X"E7",X"78",
		X"00",X"E6",X"10",X"C2",X"DF",X"E5",X"7B",X"FE",X"20",X"D2",X"EA",X"E5",X"21",X"1F",X"E7",X"79",
		X"A8",X"06",X"00",X"E6",X"03",X"CA",X"D9",X"E5",X"FE",X"01",X"C2",X"CF",X"E5",X"7B",X"FE",X"05",
		X"CA",X"D9",X"E5",X"FE",X"07",X"CA",X"D9",X"E5",X"FE",X"0F",X"CA",X"D9",X"E5",X"FE",X"11",X"CA",
		X"D9",X"E5",X"FE",X"18",X"CA",X"D9",X"E5",X"FE",X"1B",X"CA",X"D9",X"E5",X"C3",X"D7",X"E5",X"21",
		X"67",X"E7",X"FE",X"02",X"CA",X"D9",X"E5",X"06",X"20",X"19",X"7E",X"80",X"C3",X"B4",X"E6",X"7B",
		X"06",X"00",X"FE",X"30",X"D2",X"B2",X"E6",X"C3",X"D9",X"E5",X"D6",X"20",X"FE",X"10",X"D2",X"20",
		X"E6",X"5F",X"FE",X"0B",X"C2",X"0B",X"E6",X"79",X"A8",X"E6",X"02",X"CA",X"0B",X"E6",X"79",X"A8",
		X"E6",X"01",X"3E",X"F1",X"C2",X"B4",X"E6",X"3D",X"C3",X"B4",X"E6",X"79",X"A8",X"06",X"00",X"E6",
		X"01",X"C2",X"1A",X"E6",X"21",X"3F",X"E7",X"C3",X"D9",X"E5",X"21",X"57",X"E7",X"C3",X"D9",X"E5",
		X"D6",X"10",X"FE",X"08",X"D2",X"B2",X"E6",X"5F",X"21",X"4F",X"E7",X"06",X"00",X"C3",X"D9",X"E5",
		X"3A",X"26",X"DF",X"4F",X"7B",X"16",X"00",X"D6",X"40",X"FE",X"10",X"DA",X"5C",X"E6",X"D6",X"18",
		X"2F",X"3C",X"5F",X"79",X"A8",X"E6",X"01",X"C2",X"4C",X"E6",X"16",X"05",X"7B",X"82",X"11",X"0A",
		X"00",X"21",X"68",X"DF",X"19",X"3D",X"C2",X"54",X"E6",X"C3",X"BC",X"E4",X"5F",X"FE",X"08",X"CA",
		X"6C",X"E6",X"FE",X"0A",X"CA",X"6C",X"E6",X"FE",X"0B",X"C2",X"76",X"E6",X"79",X"A8",X"E6",X"01",
		X"C2",X"83",X"E6",X"C3",X"7D",X"E6",X"79",X"A8",X"E6",X"08",X"C2",X"83",X"E6",X"21",X"B7",X"E7",
		X"C3",X"86",X"E6",X"21",X"C7",X"E7",X"06",X"00",X"C3",X"D9",X"E5",X"3A",X"D7",X"DF",X"B7",X"CA",
		X"B2",X"E6",X"7A",X"FE",X"39",X"7B",X"CA",X"9F",X"E6",X"FE",X"39",X"7A",X"C2",X"B2",X"E6",X"CD",
		X"C7",X"E6",X"3A",X"26",X"DF",X"A8",X"32",X"26",X"DF",X"CD",X"7F",X"EB",X"CD",X"FC",X"E6",X"C2",
		X"AC",X"E6",X"3E",X"FF",X"4F",X"FE",X"FF",X"CA",X"C3",X"E6",X"3A",X"26",X"DF",X"E6",X"10",X"C4",
		X"39",X"F8",X"79",X"E1",X"D1",X"C1",X"C9",X"06",X"00",X"FE",X"38",X"CA",X"D3",X"E6",X"FE",X"3F",
		X"C2",X"D6",X"E6",X"06",X"01",X"C9",X"FE",X"3E",X"C2",X"DE",X"E6",X"06",X"02",X"C9",X"FE",X"3D",
		X"C2",X"E6",X"E6",X"06",X"04",X"C9",X"FE",X"3B",X"C2",X"EE",X"E6",X"06",X"08",X"C9",X"FE",X"3A",
		X"C2",X"F6",X"E6",X"06",X"10",X"C9",X"FE",X"3C",X"C0",X"06",X"20",X"C9",X"F3",X"3E",X"02",X"D3",
		X"6A",X"3A",X"7F",X"28",X"B7",X"C2",X"14",X"E7",X"3A",X"80",X"28",X"E6",X"12",X"C2",X"14",X"E7",
		X"3A",X"FF",X"29",X"B7",X"3A",X"FE",X"DF",X"D3",X"6A",X"FB",X"3E",X"00",X"C8",X"2F",X"C9",X"55",
		X"41",X"54",X"4C",X"57",X"60",X"46",X"7E",X"4A",X"59",X"56",X"4B",X"52",X"51",X"42",X"7B",X"44",
		X"5B",X"45",X"4E",X"43",X"48",X"5A",X"47",X"7D",X"58",X"4F",X"5D",X"49",X"50",X"53",X"4D",X"2A",
		X"26",X"5E",X"25",X"24",X"23",X"40",X"5F",X"3C",X"27",X"2B",X"FF",X"21",X"7C",X"29",X"28",X"20",
		X"09",X"7F",X"1C",X"1D",X"03",X"1F",X"0D",X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"2D",X"2C",
		X"3B",X"3D",X"FF",X"31",X"5C",X"30",X"39",X"B3",X"C4",X"B5",X"B4",X"C6",X"B1",X"B0",X"CE",X"BE",
		X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"C5",X"B2",X"B6",X"C3",X"C2",X"C1",X"C0",X"CF",X"BF",X"CA",
		X"C7",X"C9",X"CD",X"C8",X"B7",X"CB",X"CC",X"15",X"01",X"14",X"0C",X"17",X"FF",X"06",X"FF",X"0A",
		X"19",X"16",X"0B",X"12",X"11",X"02",X"FF",X"04",X"1B",X"05",X"0E",X"03",X"08",X"1A",X"07",X"FF",
		X"18",X"0F",X"1D",X"09",X"10",X"13",X"0D",X"FF",X"FF",X"1E",X"FF",X"FF",X"FF",X"00",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"1C",X"FF",X"FF",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"30",X"3F",
		X"2E",X"22",X"3E",X"FF",X"FF",X"39",X"38",X"0C",X"18",X"11",X"08",X"15",X"1A",X"16",X"17",X"2F",
		X"10",X"3A",X"2E",X"FF",X"FF",X"14",X"19",X"F3",X"F5",X"C5",X"D5",X"E5",X"CD",X"55",X"E8",X"21",
		X"4C",X"E8",X"E5",X"C3",X"35",X"DF",X"79",X"FE",X"1B",X"C2",X"F8",X"E7",X"3E",X"C3",X"32",X"35",
		X"DF",X"21",X"64",X"EC",X"22",X"36",X"DF",X"C9",X"FE",X"08",X"C2",X"02",X"E8",X"3E",X"12",X"C3",
		X"1B",X"E8",X"FE",X"0C",X"C2",X"0C",X"E8",X"3E",X"13",X"C3",X"1B",X"E8",X"FE",X"1B",X"D2",X"24",
		X"E8",X"FE",X"11",X"CA",X"24",X"E8",X"FE",X"10",X"DA",X"24",X"E8",X"C6",X"31",X"4F",X"CD",X"EC",
		X"E7",X"C3",X"35",X"DF",X"FE",X"7F",X"CA",X"7C",X"E8",X"FE",X"09",X"CA",X"85",X"E8",X"FE",X"0A",
		X"CA",X"C2",X"E8",X"FE",X"0D",X"CA",X"EA",X"E8",X"FE",X"1F",X"CA",X"04",X"E9",X"FE",X"07",X"CA",
		X"BE",X"E8",X"FE",X"20",X"D8",X"E1",X"CD",X"C9",X"E9",X"CD",X"9D",X"E9",X"CD",X"55",X"E8",X"E1",
		X"D1",X"C1",X"F1",X"FB",X"C9",X"F5",X"2A",X"38",X"DF",X"CD",X"48",X"EA",X"E5",X"3E",X"02",X"CD",
		X"6A",X"E8",X"E1",X"3E",X"03",X"CD",X"6A",X"E8",X"F1",X"C9",X"D3",X"6A",X"06",X"0A",X"7E",X"2F",
		X"77",X"2C",X"05",X"C2",X"6E",X"E8",X"3A",X"FE",X"DF",X"D3",X"6A",X"C9",X"CD",X"B4",X"E9",X"3E",
		X"20",X"CD",X"C9",X"E9",X"C9",X"3A",X"43",X"DF",X"47",X"3A",X"3E",X"DF",X"B8",X"CA",X"B7",X"E8",
		X"47",X"AF",X"B8",X"CA",X"99",X"E8",X"D2",X"9E",X"E8",X"C6",X"08",X"C3",X"92",X"E8",X"47",X"00",
		X"3A",X"43",X"DF",X"B8",X"DA",X"A8",X"E8",X"78",X"32",X"3E",X"DF",X"47",X"3A",X"3F",X"DF",X"4F",
		X"CD",X"C3",X"ED",X"22",X"38",X"DF",X"C9",X"CD",X"EA",X"E8",X"CD",X"C2",X"E8",X"C9",X"CD",X"39",
		X"F8",X"C9",X"3A",X"41",X"DF",X"47",X"3A",X"3F",X"DF",X"FE",X"17",X"CA",X"DF",X"E8",X"B8",X"C8",
		X"3C",X"32",X"3F",X"DF",X"2A",X"38",X"DF",X"7D",X"C6",X"0A",X"6F",X"22",X"38",X"DF",X"C9",X"3A",
		X"26",X"DF",X"E6",X"20",X"CA",X"EC",X"EA",X"C2",X"88",X"E9",X"3A",X"42",X"DF",X"47",X"3A",X"3E",
		X"DF",X"B8",X"C8",X"2A",X"38",X"DF",X"90",X"25",X"3D",X"C2",X"F7",X"E8",X"78",X"32",X"3E",X"DF",
		X"22",X"38",X"DF",X"C9",X"F5",X"C5",X"D5",X"E5",X"21",X"06",X"44",X"22",X"3A",X"DF",X"21",X"EC",
		X"44",X"22",X"3C",X"DF",X"CD",X"6E",X"E9",X"CD",X"25",X"E9",X"CD",X"88",X"E9",X"CD",X"7F",X"EB",
		X"E1",X"D1",X"C1",X"F1",X"C9",X"E5",X"F5",X"3E",X"FF",X"D3",X"10",X"D3",X"11",X"D3",X"12",X"D3",
		X"13",X"21",X"00",X"40",X"E5",X"3E",X"02",X"CD",X"5D",X"E9",X"E1",X"3E",X"03",X"CD",X"5D",X"E9",
		X"3A",X"21",X"DF",X"D3",X"10",X"3A",X"22",X"DF",X"D3",X"11",X"3A",X"23",X"DF",X"D3",X"12",X"3A",
		X"24",X"DF",X"D3",X"13",X"AF",X"32",X"44",X"DF",X"D3",X"69",X"F1",X"E1",X"C9",X"D3",X"6A",X"36",
		X"00",X"23",X"7C",X"FE",X"70",X"C2",X"5F",X"E9",X"3A",X"FE",X"DF",X"D3",X"6A",X"C9",X"AF",X"32",
		X"42",X"DF",X"32",X"40",X"DF",X"3E",X"27",X"32",X"43",X"DF",X"3E",X"17",X"32",X"41",X"DF",X"3A",
		X"26",X"DF",X"E6",X"1F",X"32",X"26",X"DF",X"C9",X"3A",X"42",X"DF",X"32",X"3E",X"DF",X"47",X"3A",
		X"40",X"DF",X"32",X"3F",X"DF",X"4F",X"CD",X"C3",X"ED",X"22",X"38",X"DF",X"C9",X"3A",X"43",X"DF",
		X"47",X"3A",X"3E",X"DF",X"B8",X"CA",X"B7",X"E8",X"3C",X"32",X"3E",X"DF",X"2A",X"38",X"DF",X"24",
		X"22",X"38",X"DF",X"C9",X"3A",X"42",X"DF",X"47",X"3A",X"3E",X"DF",X"B8",X"C8",X"3D",X"32",X"3E",
		X"DF",X"2A",X"38",X"DF",X"25",X"22",X"38",X"DF",X"C9",X"F5",X"AF",X"32",X"D9",X"DF",X"CD",X"48",
		X"EA",X"11",X"D9",X"DF",X"06",X"01",X"CD",X"5A",X"EA",X"F1",X"CD",X"EB",X"E9",X"06",X"08",X"CD",
		X"5A",X"EA",X"06",X"01",X"11",X"D9",X"DF",X"CD",X"5A",X"EA",X"C9",X"E5",X"21",X"32",X"EA",X"E5",
		X"01",X"29",X"DF",X"FE",X"40",X"D2",X"FB",X"E9",X"D6",X"20",X"C9",X"03",X"03",X"FE",X"60",X"D2",
		X"05",X"EA",X"D6",X"40",X"C9",X"03",X"03",X"FE",X"80",X"D2",X"0F",X"EA",X"D6",X"60",X"C9",X"03",
		X"03",X"FE",X"B0",X"D2",X"19",X"EA",X"D6",X"80",X"C9",X"03",X"03",X"FE",X"D0",X"D2",X"23",X"EA",
		X"D6",X"B0",X"C9",X"03",X"03",X"FE",X"F3",X"D2",X"2D",X"EA",X"D6",X"D0",X"C9",X"01",X"29",X"DF",
		X"AF",X"E1",X"F5",X"0A",X"6F",X"03",X"0A",X"67",X"F1",X"11",X"08",X"00",X"B7",X"CA",X"45",X"EA",
		X"19",X"3D",X"C3",X"3C",X"EA",X"EB",X"E1",X"C9",X"D5",X"F5",X"2A",X"38",X"DF",X"EB",X"2A",X"3A",
		X"DF",X"7D",X"83",X"6F",X"7C",X"82",X"67",X"F1",X"D1",X"C9",X"1A",X"4F",X"D5",X"11",X"D5",X"EA",
		X"D5",X"3A",X"20",X"DF",X"FE",X"01",X"C2",X"6D",X"EA",X"16",X"00",X"59",X"C9",X"FE",X"02",X"C2",
		X"76",X"EA",X"51",X"1E",X"00",X"C9",X"FE",X"03",X"C2",X"7E",X"EA",X"51",X"59",X"C9",X"FE",X"04",
		X"C2",X"89",X"EA",X"16",X"00",X"79",X"2F",X"5F",X"C9",X"FE",X"06",X"C2",X"93",X"EA",X"51",X"79",
		X"2F",X"5F",X"C9",X"FE",X"07",X"C2",X"9C",X"EA",X"51",X"1E",X"FF",X"C9",X"FE",X"08",X"C2",X"A7",
		X"EA",X"79",X"2F",X"57",X"1E",X"00",X"C9",X"FE",X"09",X"C2",X"B1",X"EA",X"79",X"2F",X"57",X"59",
		X"C9",X"FE",X"0B",X"C2",X"BA",X"EA",X"16",X"FF",X"59",X"C9",X"FE",X"0C",X"C2",X"C4",X"EA",X"79",
		X"2F",X"57",X"5F",X"C9",X"FE",X"0D",X"C2",X"CF",X"EA",X"79",X"2F",X"57",X"1E",X"FF",X"C9",X"D1",
		X"16",X"FF",X"79",X"2F",X"5F",X"3E",X"02",X"D3",X"6A",X"72",X"3E",X"03",X"D3",X"6A",X"73",X"3A",
		X"FE",X"DF",X"D3",X"6A",X"D1",X"13",X"2C",X"05",X"C2",X"5A",X"EA",X"C9",X"21",X"00",X"00",X"39",
		X"22",X"EC",X"DF",X"21",X"EC",X"DF",X"F9",X"2A",X"3C",X"DF",X"7D",X"C6",X"0A",X"6F",X"22",X"3C",
		X"DF",X"3E",X"02",X"F5",X"D3",X"6A",X"06",X"1A",X"E5",X"0E",X"28",X"36",X"00",X"24",X"0D",X"C2",
		X"0B",X"EB",X"E1",X"2C",X"05",X"C2",X"08",X"EB",X"F1",X"3D",X"CA",X"2F",X"EB",X"F5",X"3E",X"06",
		X"32",X"07",X"EB",X"2A",X"3A",X"DF",X"7D",X"C6",X"04",X"6F",X"3E",X"03",X"C3",X"04",X"EB",X"3E",
		X"1A",X"32",X"07",X"EB",X"2A",X"3C",X"DF",X"E5",X"D1",X"7D",X"C6",X"0A",X"6F",X"DB",X"74",X"E6",
		X"01",X"C2",X"3D",X"EB",X"3A",X"44",X"DF",X"C6",X"0A",X"D3",X"69",X"32",X"44",X"DF",X"3E",X"03",
		X"D3",X"6A",X"06",X"0A",X"E5",X"D5",X"0E",X"28",X"1A",X"77",X"AF",X"12",X"14",X"24",X"0D",X"C2",
		X"58",X"EB",X"D1",X"E1",X"2C",X"1C",X"05",X"C2",X"54",X"EB",X"2A",X"3A",X"DF",X"7D",X"C6",X"0A",
		X"6F",X"22",X"3A",X"DF",X"2A",X"EC",X"DF",X"F9",X"3A",X"FE",X"DF",X"D3",X"6A",X"C9",X"0D",X"F5",
		X"C5",X"D5",X"E5",X"3A",X"20",X"DF",X"F5",X"3E",X"04",X"32",X"20",X"DF",X"21",X"46",X"DF",X"3A",
		X"26",X"DF",X"E6",X"04",X"C2",X"B1",X"EB",X"3A",X"26",X"DF",X"E6",X"02",X"C2",X"A8",X"EB",X"01",
		X"52",X"EC",X"CD",X"44",X"EC",X"C3",X"B7",X"EB",X"01",X"55",X"EC",X"CD",X"44",X"EC",X"C3",X"B7",
		X"EB",X"01",X"58",X"EC",X"CD",X"44",X"EC",X"36",X"2F",X"23",X"3A",X"26",X"DF",X"E6",X"01",X"CA",
		X"C7",X"EB",X"36",X"48",X"C3",X"C9",X"EB",X"36",X"42",X"23",X"36",X"50",X"23",X"36",X"2F",X"23",
		X"3A",X"26",X"DF",X"E6",X"08",X"C2",X"DE",X"EB",X"01",X"5B",X"EC",X"C3",X"E1",X"EB",X"01",X"5E",
		X"EC",X"CD",X"44",X"EC",X"3A",X"26",X"DF",X"E6",X"20",X"C2",X"F8",X"EB",X"36",X"2F",X"23",X"01",
		X"61",X"EC",X"CD",X"44",X"EC",X"C3",X"01",X"EC",X"36",X"20",X"23",X"01",X"4F",X"EC",X"CD",X"44",
		X"EC",X"06",X"28",X"11",X"46",X"DF",X"AF",X"32",X"D9",X"DF",X"2A",X"38",X"DF",X"E5",X"2A",X"3C",
		X"DF",X"3E",X"0B",X"85",X"6F",X"22",X"38",X"DF",X"C5",X"E5",X"D5",X"11",X"D9",X"DF",X"06",X"01",
		X"CD",X"5A",X"EA",X"D1",X"1A",X"D5",X"CD",X"EB",X"E9",X"06",X"08",X"CD",X"5A",X"EA",X"D1",X"E1",
		X"24",X"C1",X"13",X"05",X"C2",X"15",X"EC",X"E1",X"22",X"38",X"DF",X"F1",X"32",X"20",X"DF",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"16",X"03",X"0A",X"77",X"23",X"03",X"15",X"C2",X"46",X"EC",X"C9",X"20",
		X"20",X"20",X"BB",X"D0",X"E2",X"C0",X"E3",X"E1",X"B3",X"E0",X"E4",X"C6",X"E4",X"E0",X"C3",X"DF",
		X"BA",X"C0",X"E3",X"DB",X"79",X"D6",X"41",X"FE",X"1A",X"D2",X"AD",X"EC",X"5F",X"16",X"00",X"21",
		X"79",X"EC",X"19",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"5E",X"EF",X"2E",X"ED",X"73",X"ED",X"79",
		X"ED",X"82",X"EF",X"8C",X"EF",X"7C",X"EF",X"6F",X"EF",X"6D",X"ED",X"52",X"ED",X"67",X"ED",X"7F",
		X"ED",X"AD",X"EC",X"66",X"EE",X"85",X"ED",X"E5",X"EE",X"AD",X"EC",X"AD",X"EC",X"AD",X"EC",X"B9",
		X"EC",X"1D",X"EE",X"AD",X"EC",X"EF",X"EC",X"0A",X"EF",X"9B",X"EE",X"AD",X"EC",X"3E",X"C3",X"32",
		X"35",X"DF",X"21",X"E6",X"E7",X"22",X"36",X"DF",X"C9",X"AF",X"32",X"D8",X"DF",X"21",X"C4",X"EC",
		X"22",X"36",X"DF",X"C9",X"3A",X"D8",X"DF",X"B7",X"C2",X"DE",X"EC",X"21",X"68",X"DF",X"79",X"32",
		X"D8",X"DF",X"11",X"0A",X"00",X"19",X"3D",X"C2",X"D5",X"EC",X"22",X"17",X"DF",X"C9",X"79",X"2A",
		X"17",X"DF",X"77",X"23",X"22",X"17",X"DF",X"B7",X"C0",X"32",X"D8",X"DF",X"C3",X"AD",X"EC",X"3E",
		X"03",X"32",X"D8",X"DF",X"21",X"01",X"ED",X"22",X"36",X"DF",X"21",X"29",X"DF",X"22",X"EC",X"DF",
		X"C9",X"3A",X"D8",X"DF",X"2A",X"EC",X"DF",X"FE",X"03",X"C2",X"1B",X"ED",X"F5",X"79",X"3D",X"07",
		X"5F",X"16",X"00",X"19",X"22",X"EC",X"DF",X"F1",X"C3",X"26",X"ED",X"FE",X"02",X"C2",X"24",X"ED",
		X"71",X"C3",X"26",X"ED",X"23",X"71",X"3D",X"32",X"D8",X"DF",X"C0",X"C3",X"AD",X"EC",X"CD",X"8E",
		X"EE",X"21",X"3E",X"ED",X"22",X"36",X"DF",X"21",X"55",X"DF",X"22",X"17",X"DF",X"C9",X"79",X"B7",
		X"CA",X"4C",X"ED",X"2A",X"17",X"DF",X"77",X"23",X"22",X"17",X"DF",X"C9",X"CD",X"7F",X"EB",X"C3",
		X"AD",X"EC",X"3A",X"40",X"DF",X"47",X"3A",X"3F",X"DF",X"B8",X"CA",X"AD",X"EC",X"3D",X"F5",X"3A",
		X"3E",X"DF",X"47",X"F1",X"C3",X"68",X"EF",X"CD",X"C2",X"E8",X"C3",X"AD",X"EC",X"CD",X"9D",X"E9",
		X"C3",X"AD",X"EC",X"CD",X"B4",X"E9",X"C3",X"AD",X"EC",X"CD",X"88",X"E9",X"C3",X"AD",X"EC",X"CD",
		X"6E",X"E9",X"C3",X"AD",X"EC",X"3A",X"20",X"DF",X"F5",X"0F",X"0F",X"E6",X"03",X"F5",X"3A",X"42",
		X"DF",X"47",X"3A",X"40",X"DF",X"4F",X"CD",X"C3",X"ED",X"11",X"06",X"44",X"19",X"F1",X"F5",X"E6",
		X"01",X"32",X"20",X"DF",X"E5",X"3E",X"02",X"32",X"D9",X"DF",X"CD",X"DC",X"ED",X"E1",X"F1",X"E6",
		X"02",X"32",X"20",X"DF",X"3E",X"03",X"32",X"D9",X"DF",X"CD",X"DC",X"ED",X"F1",X"32",X"20",X"DF",
		X"C3",X"AD",X"EC",X"21",X"00",X"00",X"78",X"B7",X"CA",X"D0",X"ED",X"24",X"3D",X"C2",X"CB",X"ED",
		X"79",X"B7",X"C8",X"7D",X"C6",X"0A",X"0D",X"C2",X"D4",X"ED",X"6F",X"C9",X"3A",X"42",X"DF",X"47",
		X"3A",X"43",X"DF",X"90",X"3C",X"4F",X"3A",X"40",X"DF",X"47",X"3A",X"41",X"DF",X"90",X"3C",X"47",
		X"C5",X"E5",X"3A",X"D9",X"DF",X"D3",X"6A",X"3A",X"20",X"DF",X"B7",X"C2",X"02",X"EE",X"57",X"C3",
		X"04",X"EE",X"16",X"FF",X"3E",X"0A",X"72",X"2C",X"3D",X"C2",X"06",X"EE",X"05",X"C2",X"04",X"EE",
		X"3A",X"FE",X"DF",X"D3",X"6A",X"E1",X"24",X"C1",X"0D",X"C2",X"F0",X"ED",X"C9",X"3E",X"04",X"32",
		X"D8",X"DF",X"21",X"31",X"EE",X"22",X"36",X"DF",X"3A",X"26",X"DF",X"F6",X"20",X"32",X"26",X"DF",
		X"C9",X"3A",X"D8",X"DF",X"F5",X"0D",X"21",X"5D",X"EE",X"E5",X"FE",X"04",X"C2",X"44",X"EE",X"79",
		X"32",X"42",X"DF",X"C9",X"FE",X"03",X"C2",X"4E",X"EE",X"79",X"32",X"40",X"DF",X"C9",X"FE",X"02",
		X"C2",X"58",X"EE",X"79",X"32",X"43",X"DF",X"C9",X"79",X"32",X"41",X"DF",X"E1",X"F1",X"3D",X"32",
		X"D8",X"DF",X"CA",X"79",X"ED",X"C9",X"3E",X"0A",X"01",X"F6",X"FF",X"21",X"D6",X"DF",X"09",X"77",
		X"23",X"36",X"00",X"2B",X"3D",X"C2",X"6E",X"EE",X"0E",X"15",X"11",X"93",X"EF",X"21",X"20",X"DF",
		X"1A",X"77",X"13",X"23",X"0D",X"C2",X"80",X"EE",X"CD",X"8E",X"EE",X"C3",X"AD",X"EC",X"21",X"54",
		X"DF",X"3E",X"1A",X"36",X"20",X"23",X"3D",X"C2",X"93",X"EE",X"C9",X"3E",X"02",X"32",X"D8",X"DF",
		X"21",X"A7",X"EE",X"22",X"36",X"DF",X"C9",X"3A",X"D8",X"DF",X"0D",X"F5",X"FE",X"02",X"C2",X"C1",
		X"EE",X"79",X"D6",X"20",X"FE",X"18",X"DA",X"BB",X"EE",X"3E",X"17",X"32",X"3F",X"DF",X"C3",X"CE",
		X"EE",X"79",X"D6",X"20",X"FE",X"28",X"DA",X"CB",X"EE",X"3E",X"27",X"32",X"3E",X"DF",X"F1",X"3D",
		X"32",X"D8",X"DF",X"C0",X"3A",X"3E",X"DF",X"47",X"3A",X"3F",X"DF",X"4F",X"CD",X"C3",X"ED",X"22",
		X"38",X"DF",X"C3",X"AD",X"EC",X"21",X"EC",X"EE",X"22",X"36",X"DF",X"C9",X"79",X"E6",X"0F",X"F5",
		X"F5",X"0F",X"0F",X"E6",X"03",X"47",X"F1",X"E6",X"03",X"B8",X"C2",X"03",X"EF",X"F1",X"3E",X"02",
		X"C3",X"04",X"EF",X"F1",X"32",X"20",X"DF",X"C3",X"AD",X"EC",X"3E",X"04",X"32",X"D8",X"DF",X"21",
		X"16",X"EF",X"22",X"36",X"DF",X"C9",X"3A",X"D8",X"DF",X"F5",X"21",X"55",X"EF",X"E5",X"FE",X"04",
		X"C2",X"2D",X"EF",X"79",X"FE",X"80",X"C8",X"32",X"22",X"DF",X"D3",X"11",X"C9",X"FE",X"03",X"C2",
		X"3C",X"EF",X"79",X"FE",X"80",X"C8",X"32",X"23",X"DF",X"D3",X"12",X"C9",X"FE",X"02",X"C2",X"4B",
		X"EF",X"79",X"FE",X"80",X"C8",X"32",X"24",X"DF",X"D3",X"13",X"C9",X"79",X"FE",X"80",X"C8",X"32",
		X"21",X"DF",X"D3",X"10",X"E1",X"F1",X"3D",X"32",X"D8",X"DF",X"CA",X"AD",X"EC",X"C9",X"3A",X"43",
		X"DF",X"32",X"3E",X"DF",X"47",X"3A",X"41",X"DF",X"32",X"3F",X"DF",X"4F",X"C3",X"DC",X"EE",X"3A",
		X"42",X"DF",X"32",X"3E",X"DF",X"47",X"3A",X"3F",X"DF",X"C3",X"6B",X"EF",X"3A",X"43",X"DF",X"C3",
		X"72",X"EF",X"3A",X"3E",X"DF",X"47",X"3A",X"40",X"DF",X"C3",X"68",X"EF",X"3A",X"3E",X"DF",X"47",
		X"C3",X"65",X"EF",X"02",X"FF",X"CD",X"1E",X"F0",X"00",X"00",X"1F",X"E7",X"EF",X"F2",X"EF",X"F3",
		X"EF",X"F4",X"EF",X"F2",X"EF",X"F5",X"EF",X"F6",X"F5",X"D5",X"E5",X"C5",X"CD",X"55",X"F0",X"21",
		X"8F",X"E1",X"CD",X"C2",X"E3",X"21",X"AD",X"E1",X"CD",X"C2",X"E3",X"21",X"BB",X"E1",X"CD",X"C2",
		X"E3",X"CD",X"6F",X"E4",X"FE",X"0D",X"CA",X"CE",X"EF",X"C1",X"E1",X"C3",X"2B",X"F0",X"21",X"CC",
		X"E1",X"CD",X"C2",X"E3",X"C1",X"E1",X"1E",X"B0",X"CD",X"63",X"F0",X"3E",X"0D",X"D3",X"62",X"C3",
		X"2B",X"F0",X"22",X"1E",X"DF",X"21",X"00",X"00",X"39",X"22",X"17",X"DF",X"2A",X"1E",X"DF",X"F5",
		X"D5",X"E5",X"C5",X"21",X"8F",X"E1",X"CD",X"C2",X"E3",X"21",X"B4",X"E1",X"CD",X"C2",X"E3",X"21",
		X"BB",X"E1",X"CD",X"C2",X"E3",X"CD",X"6F",X"E4",X"FE",X"0D",X"C2",X"C9",X"EF",X"21",X"D7",X"E1",
		X"CD",X"C2",X"E3",X"AF",X"C1",X"E1",X"CD",X"86",X"F0",X"F3",X"C2",X"47",X"F0",X"7A",X"CD",X"55",
		X"F0",X"BA",X"CA",X"2B",X"F0",X"21",X"E2",X"E1",X"CD",X"C2",X"E3",X"21",X"13",X"E0",X"22",X"05",
		X"DF",X"CD",X"38",X"F0",X"D1",X"F1",X"FB",X"C9",X"3E",X"FF",X"D3",X"75",X"3E",X"20",X"D3",X"74",
		X"21",X"F0",X"E1",X"CD",X"C2",X"E3",X"C9",X"21",X"B7",X"F1",X"CD",X"C2",X"E3",X"CD",X"38",X"F0",
		X"2A",X"17",X"DF",X"F9",X"C9",X"F5",X"16",X"00",X"0A",X"82",X"57",X"CD",X"B6",X"E3",X"DA",X"58",
		X"F0",X"F1",X"C9",X"F5",X"C5",X"E5",X"D5",X"C5",X"CD",X"AC",X"F0",X"7D",X"91",X"4F",X"7C",X"98",
		X"47",X"03",X"E1",X"56",X"CD",X"DB",X"F0",X"23",X"0B",X"78",X"B1",X"C2",X"73",X"F0",X"D1",X"CD",
		X"DB",X"F0",X"E1",X"C1",X"F1",X"C9",X"F5",X"C5",X"E5",X"E5",X"C5",X"CD",X"2D",X"F1",X"C1",X"E1",
		X"0B",X"03",X"C5",X"CD",X"5C",X"F1",X"C1",X"7A",X"02",X"79",X"AD",X"C2",X"91",X"F0",X"78",X"AC",
		X"C2",X"91",X"F0",X"C5",X"CD",X"5C",X"F1",X"C1",X"E1",X"C1",X"F1",X"C9",X"F3",X"E5",X"21",X"22",
		X"F1",X"22",X"05",X"DF",X"21",X"40",X"1F",X"3E",X"9E",X"D3",X"63",X"3E",X"02",X"D3",X"62",X"3E",
		X"10",X"D3",X"63",X"3E",X"FD",X"D3",X"75",X"3E",X"0D",X"CD",X"22",X"F1",X"3E",X"0C",X"76",X"3E",
		X"0D",X"76",X"2B",X"7C",X"B5",X"C2",X"CC",X"F0",X"E1",X"F3",X"C9",X"3E",X"0C",X"FB",X"76",X"3E",
		X"0C",X"76",X"3E",X"0D",X"76",X"3E",X"0D",X"76",X"3E",X"08",X"F5",X"3E",X"0C",X"76",X"7A",X"0F",
		X"57",X"3E",X"06",X"17",X"76",X"7A",X"07",X"57",X"3E",X"06",X"3F",X"17",X"76",X"7A",X"0F",X"57",
		X"3E",X"0D",X"76",X"F1",X"3D",X"C2",X"EA",X"F0",X"3E",X"0C",X"76",X"3E",X"0D",X"76",X"3E",X"0C",
		X"76",X"3E",X"0D",X"76",X"3E",X"0C",X"76",X"3E",X"0D",X"76",X"3E",X"0C",X"76",X"3E",X"0D",X"76",
		X"F3",X"C9",X"D3",X"6B",X"7B",X"D3",X"60",X"3E",X"61",X"D3",X"74",X"FB",X"C9",X"21",X"47",X"F0",
		X"22",X"05",X"DF",X"F3",X"3E",X"10",X"D3",X"63",X"3E",X"FD",X"D3",X"75",X"21",X"E8",X"03",X"CD",
		X"85",X"F1",X"2B",X"7C",X"B5",X"C2",X"3F",X"F1",X"44",X"5C",X"FB",X"CD",X"85",X"F1",X"09",X"1D",
		X"C2",X"4B",X"F1",X"24",X"24",X"24",X"7C",X"A7",X"1F",X"84",X"5F",X"C9",X"CD",X"85",X"F1",X"CD",
		X"85",X"F1",X"79",X"93",X"DA",X"5F",X"F1",X"06",X"08",X"16",X"00",X"CD",X"85",X"F1",X"79",X"93",
		X"D2",X"78",X"F1",X"F5",X"CD",X"85",X"F1",X"F1",X"7A",X"1F",X"57",X"05",X"C2",X"6B",X"F1",X"CD",
		X"85",X"F1",X"CD",X"85",X"F1",X"DB",X"74",X"E6",X"10",X"CA",X"85",X"F1",X"DB",X"74",X"E6",X"10",
		X"C2",X"8C",X"F1",X"AF",X"D3",X"63",X"DB",X"60",X"2F",X"4F",X"3E",X"10",X"D3",X"63",X"3E",X"FF",
		X"D3",X"60",X"C9",X"C5",X"D5",X"CD",X"5C",X"F1",X"7A",X"D1",X"C1",X"C9",X"F5",X"D5",X"1E",X"B0",
		X"51",X"CD",X"DB",X"F0",X"D1",X"F1",X"C9",X"0A",X"2A",X"20",X"DE",X"E8",X"D8",X"D1",X"DA",X"D0",
		X"20",X"E7",X"E2",X"D5",X"DD",X"D8",X"EF",X"20",X"2A",X"0D",X"00",X"11",X"00",X"00",X"01",X"00",
		X"C0",X"21",X"01",X"C0",X"CD",X"81",X"E3",X"2A",X"00",X"C0",X"7C",X"BD",X"C8",X"03",X"21",X"FF",
		X"C3",X"CD",X"81",X"E3",X"CD",X"59",X"E2",X"2A",X"00",X"C0",X"2B",X"7E",X"23",X"CD",X"C2",X"E3",
		X"B7",X"CA",X"2D",X"F2",X"57",X"06",X"00",X"CD",X"6F",X"E4",X"FE",X"0D",X"CA",X"20",X"F2",X"FE",
		X"19",X"C2",X"0E",X"F2",X"4F",X"78",X"B7",X"CA",X"F7",X"F1",X"05",X"C3",X"1A",X"F2",X"FE",X"1A",
		X"C2",X"F7",X"F1",X"4F",X"78",X"BA",X"CA",X"F7",X"F1",X"04",X"CD",X"D7",X"E7",X"C3",X"F7",X"F1",
		X"78",X"01",X"08",X"00",X"B7",X"CA",X"2D",X"F2",X"09",X"3D",X"C3",X"24",X"F2",X"5E",X"23",X"56",
		X"D5",X"23",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"D5",X"23",X"5E",X"23",X"56",X"EB",X"D1",
		X"CD",X"81",X"E3",X"CD",X"66",X"EE",X"E1",X"E9",X"DB",X"74",X"E6",X"04",X"C8",X"3E",X"FF",X"C9",
		X"F5",X"C5",X"CD",X"48",X"F2",X"CA",X"52",X"F2",X"79",X"FE",X"80",X"D4",X"6B",X"F2",X"2F",X"D3",
		X"68",X"3E",X"09",X"D3",X"6B",X"3D",X"D3",X"6B",X"C1",X"F1",X"C9",X"FE",X"F0",X"C2",X"75",X"F2",
		X"3E",X"B5",X"C3",X"7C",X"F2",X"FE",X"F1",X"C2",X"7C",X"F2",X"3E",X"D5",X"FE",X"D0",X"D2",X"88",
		X"F2",X"D6",X"B0",X"0E",X"00",X"C3",X"8C",X"F2",X"D6",X"D0",X"0E",X"01",X"E5",X"D5",X"21",X"A1",
		X"F2",X"16",X"00",X"5F",X"19",X"5E",X"79",X"B7",X"7B",X"C2",X"9E",X"F2",X"C6",X"20",X"D1",X"E1",
		X"C9",X"C1",X"C2",X"D7",X"C7",X"C4",X"C5",X"D6",X"DA",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",
		X"D0",X"D2",X"D3",X"D4",X"D5",X"C6",X"C8",X"C3",X"DE",X"DB",X"DD",X"DF",X"D9",X"D8",X"DC",X"C0",
		X"D1",X"C5",X"0E",X"40",X"C3",X"CA",X"F2",X"C5",X"0E",X"80",X"F3",X"06",X"F6",X"3E",X"0B",X"D3",
		X"6B",X"3D",X"D3",X"6B",X"DB",X"74",X"04",X"A1",X"CA",X"D4",X"F2",X"78",X"A7",X"F2",X"EB",X"F2",
		X"2F",X"3C",X"FE",X"0A",X"06",X"00",X"FA",X"EB",X"F2",X"06",X"7F",X"78",X"C1",X"FB",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"1E",X"0C",X"0C",X"00",X"0C",X"00",X"36",
		X"36",X"36",X"00",X"00",X"00",X"00",X"00",X"36",X"36",X"7F",X"36",X"7F",X"36",X"36",X"00",X"00",
		X"18",X"7C",X"06",X"3C",X"60",X"37",X"18",X"00",X"63",X"33",X"18",X"0C",X"66",X"63",X"00",X"1C",
		X"36",X"1C",X"6E",X"3B",X"33",X"6E",X"00",X"06",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"18",
		X"0C",X"06",X"06",X"06",X"0C",X"18",X"00",X"06",X"0C",X"18",X"18",X"18",X"0C",X"06",X"00",X"00",
		X"66",X"3C",X"FF",X"3C",X"66",X"00",X"00",X"00",X"0C",X"0C",X"3F",X"0C",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"06",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"3E",
		X"63",X"73",X"7B",X"6F",X"67",X"3E",X"00",X"0C",X"0E",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"1E",
		X"33",X"30",X"1C",X"06",X"33",X"3F",X"00",X"3F",X"33",X"18",X"1C",X"30",X"33",X"1E",X"00",X"38",
		X"3C",X"36",X"33",X"7F",X"30",X"78",X"00",X"3F",X"03",X"1F",X"30",X"30",X"33",X"1E",X"00",X"1C",
		X"06",X"03",X"1F",X"33",X"33",X"1E",X"00",X"3F",X"33",X"30",X"18",X"0C",X"0C",X"0C",X"00",X"1E",
		X"33",X"33",X"1E",X"33",X"33",X"1E",X"00",X"1E",X"33",X"33",X"3E",X"30",X"18",X"0E",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"0C",X"0C",X"00",X"00",X"0C",X"0C",X"00",X"00",X"0C",X"0C",X"06",X"18",
		X"0C",X"06",X"03",X"06",X"0C",X"18",X"00",X"00",X"00",X"3F",X"00",X"3F",X"00",X"00",X"00",X"06",
		X"0C",X"18",X"30",X"18",X"0C",X"06",X"00",X"1E",X"33",X"30",X"18",X"0C",X"00",X"0C",X"00",X"3E",
		X"63",X"7B",X"7B",X"03",X"1E",X"00",X"00",X"0C",X"1E",X"33",X"33",X"3F",X"33",X"33",X"00",X"3F",
		X"66",X"66",X"3E",X"66",X"66",X"3F",X"00",X"3C",X"66",X"03",X"03",X"03",X"66",X"3C",X"00",X"1F",
		X"36",X"66",X"66",X"66",X"36",X"1F",X"00",X"7F",X"46",X"16",X"1E",X"16",X"46",X"7F",X"00",X"7F",
		X"46",X"16",X"1E",X"16",X"06",X"0F",X"00",X"3C",X"66",X"03",X"03",X"73",X"66",X"7C",X"00",X"33",
		X"33",X"33",X"3F",X"33",X"33",X"33",X"00",X"1E",X"0C",X"0C",X"0C",X"0C",X"0C",X"1E",X"00",X"78",
		X"30",X"30",X"30",X"33",X"33",X"1E",X"00",X"67",X"66",X"36",X"1E",X"36",X"66",X"67",X"00",X"0F",
		X"06",X"06",X"06",X"46",X"66",X"7F",X"00",X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"63",
		X"67",X"6F",X"7B",X"73",X"63",X"63",X"00",X"1C",X"36",X"63",X"63",X"63",X"36",X"1C",X"00",X"3F",
		X"66",X"66",X"3E",X"06",X"06",X"0F",X"00",X"1E",X"33",X"33",X"33",X"3B",X"1E",X"38",X"00",X"7F",
		X"66",X"66",X"3E",X"36",X"66",X"67",X"00",X"1E",X"33",X"06",X"0C",X"18",X"33",X"1E",X"00",X"3F",
		X"2D",X"0C",X"0C",X"0C",X"0C",X"1E",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"1E",X"00",X"33",
		X"33",X"33",X"33",X"33",X"1E",X"0C",X"00",X"63",X"63",X"63",X"6B",X"7F",X"77",X"63",X"00",X"63",
		X"63",X"36",X"1C",X"1C",X"36",X"63",X"00",X"33",X"33",X"33",X"1E",X"0C",X"0C",X"1E",X"00",X"7F",
		X"63",X"31",X"18",X"4C",X"66",X"7F",X"00",X"1E",X"06",X"06",X"06",X"06",X"06",X"1E",X"00",X"03",
		X"06",X"0C",X"18",X"30",X"60",X"40",X"00",X"1E",X"18",X"18",X"18",X"18",X"18",X"1E",X"00",X"08",
		X"1C",X"36",X"63",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"0C",
		X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"30",X"3E",X"33",X"6E",X"00",X"07",
		X"06",X"06",X"3E",X"66",X"66",X"3B",X"00",X"00",X"00",X"1E",X"33",X"03",X"33",X"1E",X"00",X"38",
		X"30",X"30",X"3E",X"33",X"33",X"6E",X"00",X"00",X"00",X"1E",X"33",X"3F",X"03",X"1E",X"00",X"1C",
		X"36",X"06",X"0F",X"06",X"06",X"0F",X"00",X"00",X"00",X"6E",X"33",X"33",X"3E",X"30",X"1F",X"07",
		X"06",X"36",X"6E",X"66",X"66",X"67",X"00",X"0C",X"00",X"0E",X"0C",X"0C",X"0C",X"1E",X"00",X"30",
		X"00",X"30",X"30",X"30",X"33",X"33",X"1E",X"07",X"06",X"66",X"36",X"1E",X"36",X"67",X"00",X"0E",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"1E",X"00",X"00",X"00",X"33",X"7F",X"7F",X"6B",X"63",X"00",X"00",
		X"00",X"1F",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"1E",X"33",X"33",X"33",X"1E",X"00",X"00",
		X"00",X"3B",X"66",X"66",X"3E",X"06",X"0F",X"00",X"00",X"6E",X"33",X"33",X"3E",X"30",X"78",X"00",
		X"00",X"3B",X"6E",X"66",X"06",X"0F",X"00",X"00",X"00",X"3E",X"03",X"1E",X"30",X"1F",X"00",X"08",
		X"0C",X"3E",X"0C",X"0C",X"2C",X"18",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"6E",X"00",X"00",
		X"00",X"33",X"33",X"33",X"1E",X"0C",X"00",X"00",X"00",X"63",X"6B",X"7F",X"7F",X"36",X"00",X"00",
		X"00",X"63",X"36",X"1C",X"36",X"63",X"00",X"00",X"00",X"33",X"33",X"33",X"3E",X"30",X"1F",X"00",
		X"00",X"3F",X"19",X"0C",X"26",X"3F",X"00",X"38",X"0C",X"0C",X"07",X"0C",X"0C",X"38",X"00",X"08",
		X"08",X"08",X"00",X"00",X"08",X"08",X"08",X"07",X"0C",X"0C",X"38",X"0C",X"0C",X"07",X"00",X"6E",
		X"3B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"36",X"63",X"63",X"7F",X"00",X"0C",
		X"1E",X"33",X"33",X"3F",X"33",X"33",X"00",X"7F",X"06",X"06",X"3E",X"66",X"66",X"3F",X"00",X"3F",
		X"66",X"66",X"3E",X"66",X"66",X"3F",X"00",X"7F",X"66",X"06",X"06",X"06",X"06",X"0F",X"00",X"3C",
		X"36",X"36",X"36",X"36",X"36",X"7F",X"63",X"7F",X"46",X"16",X"1E",X"16",X"46",X"7F",X"00",X"6B",
		X"6B",X"3E",X"1C",X"3E",X"69",X"6B",X"00",X"3E",X"63",X"60",X"38",X"60",X"63",X"3E",X"00",X"63",
		X"63",X"73",X"7B",X"6F",X"67",X"63",X"00",X"1C",X"63",X"73",X"7B",X"6F",X"67",X"63",X"00",X"63",
		X"33",X"1B",X"0F",X"1B",X"33",X"63",X"00",X"78",X"6C",X"66",X"66",X"66",X"66",X"63",X"00",X"63",
		X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"33",X"33",X"33",X"3F",X"33",X"33",X"33",X"00",X"3E",
		X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"7F",X"63",X"63",X"63",X"63",X"63",X"63",X"00",X"3F",
		X"66",X"66",X"3E",X"06",X"06",X"0F",X"00",X"3C",X"66",X"03",X"03",X"03",X"66",X"3C",X"00",X"3F",
		X"2D",X"0C",X"0C",X"0C",X"0C",X"1E",X"00",X"63",X"63",X"63",X"7E",X"60",X"20",X"1E",X"00",X"18",
		X"7E",X"DB",X"DB",X"7E",X"18",X"3C",X"00",X"63",X"36",X"1C",X"1C",X"36",X"63",X"63",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"7F",X"60",X"63",X"63",X"63",X"7E",X"60",X"60",X"60",X"00",X"63",
		X"6B",X"6B",X"6B",X"6B",X"6B",X"7F",X"00",X"63",X"6B",X"6B",X"6B",X"6B",X"6B",X"7F",X"60",X"07",
		X"06",X"06",X"36",X"66",X"66",X"36",X"00",X"63",X"63",X"63",X"6F",X"5B",X"5B",X"6F",X"00",X"03",
		X"03",X"03",X"3F",X"63",X"63",X"3F",X"00",X"3E",X"63",X"60",X"7C",X"60",X"63",X"3E",X"00",X"33",
		X"6B",X"6B",X"6F",X"6B",X"6B",X"33",X"00",X"7E",X"63",X"63",X"7E",X"6C",X"66",X"63",X"00",X"00",
		X"00",X"1E",X"30",X"3E",X"33",X"7E",X"00",X"00",X"00",X"3F",X"03",X"3F",X"63",X"3F",X"00",X"00",
		X"00",X"1F",X"33",X"1F",X"33",X"1F",X"00",X"00",X"00",X"3F",X"03",X"03",X"03",X"03",X"00",X"00",
		X"00",X"3C",X"36",X"36",X"36",X"7F",X"63",X"00",X"00",X"1E",X"33",X"3F",X"03",X"1E",X"00",X"00",
		X"00",X"6B",X"6B",X"3E",X"6B",X"6B",X"00",X"00",X"00",X"1E",X"33",X"18",X"33",X"1E",X"00",X"00",
		X"00",X"63",X"63",X"73",X"7F",X"66",X"00",X"00",X"18",X"63",X"63",X"73",X"7F",X"66",X"00",X"00",
		X"00",X"33",X"1B",X"0F",X"1B",X"73",X"00",X"00",X"00",X"78",X"6C",X"66",X"66",X"67",X"00",X"00",
		X"00",X"63",X"77",X"7F",X"6B",X"63",X"00",X"00",X"00",X"63",X"63",X"7F",X"63",X"63",X"00",X"00",
		X"00",X"3E",X"63",X"63",X"63",X"3E",X"00",X"00",X"00",X"7F",X"63",X"63",X"63",X"63",X"00",X"00",
		X"00",X"3F",X"63",X"63",X"3F",X"03",X"03",X"00",X"00",X"3E",X"63",X"03",X"63",X"3E",X"00",X"00",
		X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"63",X"66",X"7C",X"60",X"3E",X"00",X"00",
		X"00",X"18",X"7E",X"DB",X"7E",X"18",X"18",X"00",X"00",X"63",X"36",X"1C",X"36",X"63",X"00",X"00",
		X"00",X"33",X"33",X"33",X"33",X"7F",X"60",X"00",X"00",X"33",X"33",X"3E",X"30",X"30",X"00",X"00",
		X"00",X"6B",X"6B",X"6B",X"6B",X"7F",X"00",X"00",X"00",X"6B",X"6B",X"6B",X"6B",X"7F",X"60",X"00",
		X"00",X"07",X"06",X"3E",X"66",X"3E",X"00",X"00",X"00",X"63",X"63",X"6F",X"5B",X"6F",X"00",X"00",
		X"00",X"03",X"03",X"3F",X"63",X"3F",X"00",X"00",X"00",X"3F",X"60",X"78",X"60",X"3F",X"00",X"00",
		X"00",X"33",X"6B",X"6F",X"6B",X"33",X"00",X"00",X"00",X"7E",X"63",X"7E",X"66",X"63",X"00",X"14",
		X"7F",X"46",X"16",X"1E",X"16",X"46",X"7F",X"00",X"12",X"1E",X"33",X"3F",X"03",X"1E",X"00",X"64",
		X"C3",X"A3",X"E4",X"C3",X"6F",X"E4",X"C3",X"A3",X"F1",X"C3",X"D7",X"E7",X"C3",X"AC",X"F1",X"C3",
		X"50",X"F2",X"C3",X"FC",X"E6",X"C3",X"48",X"F2",X"C3",X"C2",X"E3",X"C3",X"F1",X"E3",X"C3",X"2D",
		X"F1",X"C3",X"AC",X"F0",X"C3",X"E2",X"EF",X"C3",X"A8",X"EF",X"C3",X"55",X"F0",X"C3",X"1C",X"E4",
		X"C3",X"A5",X"E0",X"C3",X"1C",X"FD",X"C3",X"40",X"FD",X"C3",X"2E",X"FD",X"C3",X"35",X"FD",X"C3",
		X"80",X"F8",X"C3",X"F0",X"F8",X"C3",X"AB",X"F9",X"C3",X"80",X"FA",X"C3",X"16",X"FB",X"C3",X"72",
		X"FB",X"C3",X"BE",X"FB",X"C3",X"05",X"FC",X"C3",X"39",X"FC",X"C3",X"A0",X"FC",X"C3",X"25",X"E9",
		X"C3",X"04",X"E9",X"C3",X"81",X"E3",X"C3",X"FF",X"FF",X"C3",X"B6",X"E3",X"C3",X"7E",X"F8",X"C3",
		X"7E",X"F8",X"C3",X"44",X"E4",X"C3",X"D5",X"E3",X"C3",X"C1",X"F2",X"C3",X"C7",X"F2",X"C9",X"FF",
		X"CD",X"BA",X"F8",X"D8",X"E5",X"D5",X"C5",X"7A",X"1F",X"7B",X"1F",X"1F",X"1F",X"E6",X"3F",X"C6",
		X"40",X"57",X"4B",X"58",X"79",X"E6",X"07",X"4F",X"06",X"00",X"21",X"E8",X"F8",X"09",X"46",X"EB",
		X"3A",X"DC",X"DF",X"4F",X"CD",X"C5",X"F8",X"78",X"32",X"DF",X"DF",X"22",X"DD",X"DF",X"C1",X"E1",
		X"D1",X"22",X"EF",X"DF",X"78",X"32",X"F1",X"DF",X"EB",X"C9",X"78",X"C6",X"0A",X"D8",X"3E",X"7F",
		X"93",X"3E",X"01",X"9A",X"C9",X"16",X"02",X"F3",X"3E",X"02",X"D3",X"6A",X"79",X"A2",X"78",X"CA",
		X"D6",X"F8",X"B6",X"C3",X"D8",X"F8",X"2F",X"A6",X"77",X"3E",X"03",X"D3",X"6A",X"15",X"C2",X"CC",
		X"F8",X"3A",X"FE",X"DF",X"D3",X"6A",X"FB",X"C9",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",
		X"CD",X"BA",X"F8",X"D8",X"E5",X"D5",X"C5",X"2A",X"EF",X"DF",X"7B",X"95",X"6F",X"7A",X"9C",X"67",
		X"DC",X"A3",X"F9",X"0E",X"02",X"DA",X"0A",X"F9",X"0E",X"00",X"3A",X"F1",X"DF",X"EB",X"90",X"6F",
		X"DC",X"A3",X"F9",X"3E",X"00",X"67",X"DA",X"1B",X"F9",X"3E",X"40",X"B1",X"4F",X"7B",X"95",X"7A",
		X"9C",X"3E",X"01",X"D2",X"29",X"F9",X"EB",X"3E",X"80",X"B1",X"32",X"E0",X"DF",X"29",X"CD",X"A3",
		X"F9",X"2B",X"22",X"E3",X"DF",X"EB",X"22",X"E5",X"DF",X"54",X"5D",X"29",X"22",X"E1",X"DF",X"3A",
		X"DC",X"DF",X"4F",X"3A",X"DF",X"DF",X"47",X"2A",X"DD",X"DF",X"7C",X"D6",X"40",X"DA",X"37",X"FA",
		X"3E",X"70",X"94",X"DA",X"37",X"FA",X"7A",X"B3",X"CA",X"A7",X"F8",X"1B",X"D5",X"E5",X"2A",X"E3",
		X"DF",X"EB",X"2A",X"E5",X"DF",X"23",X"19",X"3A",X"E0",X"DF",X"DA",X"74",X"F9",X"F6",X"81",X"EB",
		X"2A",X"E1",X"DF",X"19",X"22",X"E5",X"DF",X"E1",X"57",X"0F",X"D2",X"90",X"F9",X"0F",X"78",X"D2",
		X"8A",X"F9",X"0F",X"D2",X"8F",X"F9",X"25",X"C3",X"8F",X"F9",X"07",X"D2",X"8F",X"F9",X"24",X"47",
		X"7A",X"07",X"D2",X"9C",X"F9",X"07",X"2D",X"DA",X"9C",X"F9",X"2C",X"2C",X"CD",X"C5",X"F8",X"D1",
		X"C3",X"56",X"F9",X"7C",X"2F",X"67",X"7D",X"2F",X"6F",X"23",X"C9",X"CD",X"BA",X"F8",X"D8",X"E5",
		X"D5",X"C5",X"EB",X"22",X"E9",X"DF",X"68",X"26",X"00",X"22",X"EB",X"DF",X"3A",X"F7",X"DF",X"47",
		X"2A",X"F8",X"DF",X"EB",X"CD",X"91",X"FA",X"DA",X"37",X"FA",X"59",X"16",X"00",X"3A",X"EE",X"DF",
		X"6F",X"62",X"EB",X"A7",X"C4",X"A8",X"FA",X"22",X"D7",X"DF",X"59",X"3A",X"ED",X"DF",X"6F",X"62",
		X"EB",X"A7",X"C4",X"A8",X"FA",X"22",X"F5",X"DF",X"48",X"CD",X"C5",X"FA",X"E5",X"2A",X"F5",X"DF",
		X"CD",X"A8",X"FA",X"24",X"22",X"F3",X"DF",X"2A",X"D7",X"DF",X"EB",X"CD",X"A8",X"FA",X"22",X"D9",
		X"DF",X"EB",X"D1",X"CD",X"A8",X"FA",X"22",X"D7",X"DF",X"2A",X"F5",X"DF",X"CD",X"A8",X"FA",X"22",
		X"F5",X"DF",X"3A",X"F9",X"DF",X"4F",X"CD",X"3B",X"FA",X"CD",X"80",X"F8",X"DA",X"37",X"FA",X"0C",
		X"3E",X"48",X"A9",X"C2",X"27",X"FA",X"4F",X"CD",X"3B",X"FA",X"CD",X"F0",X"F8",X"DA",X"37",X"FA",
		X"3A",X"F8",X"DF",X"A9",X"C2",X"1F",X"FA",X"C1",X"D1",X"E1",X"C9",X"CD",X"C5",X"FA",X"22",X"E1",
		X"DF",X"EB",X"22",X"E5",X"DF",X"2A",X"D9",X"DF",X"CD",X"9D",X"FA",X"E5",X"2A",X"E5",X"DF",X"EB",
		X"2A",X"F5",X"DF",X"CD",X"9D",X"FA",X"D1",X"19",X"EB",X"2A",X"EB",X"DF",X"19",X"7C",X"C6",X"FF",
		X"D8",X"45",X"2A",X"E5",X"DF",X"EB",X"2A",X"F3",X"DF",X"CD",X"9D",X"FA",X"E5",X"2A",X"E1",X"DF",
		X"EB",X"2A",X"D7",X"DF",X"CD",X"9D",X"FA",X"D1",X"19",X"EB",X"2A",X"E9",X"DF",X"19",X"EB",X"C9",
		X"CD",X"91",X"FA",X"D8",X"22",X"ED",X"DF",X"EB",X"22",X"F8",X"DF",X"EB",X"78",X"32",X"F7",X"DF",
		X"C9",X"7A",X"C6",X"B9",X"D8",X"7B",X"C6",X"B9",X"D8",X"78",X"C6",X"B9",X"C9",X"CD",X"A8",X"FA",
		X"7C",X"26",X"00",X"0F",X"DC",X"A3",X"F9",X"C9",X"D5",X"C5",X"7C",X"AA",X"47",X"7D",X"21",X"FF",
		X"00",X"54",X"0E",X"08",X"0F",X"D2",X"B9",X"FA",X"19",X"EB",X"29",X"EB",X"0D",X"C2",X"B4",X"FA",
		X"6C",X"60",X"C1",X"D1",X"C9",X"C5",X"79",X"01",X"00",X"00",X"16",X"12",X"92",X"FA",X"DC",X"FA",
		X"0C",X"92",X"FA",X"DC",X"FA",X"04",X"92",X"FA",X"DC",X"FA",X"0D",X"92",X"82",X"07",X"6F",X"26",
		X"00",X"11",X"F0",X"FA",X"19",X"5E",X"23",X"6E",X"60",X"51",X"7C",X"AA",X"C1",X"C8",X"EB",X"C9",
		X"00",X"FF",X"16",X"FF",X"2C",X"FC",X"42",X"F7",X"58",X"F1",X"6C",X"E8",X"80",X"DE",X"93",X"D2",
		X"A5",X"C4",X"B5",X"B5",X"C4",X"A5",X"D2",X"93",X"DE",X"80",X"E8",X"6C",X"F1",X"58",X"F7",X"42",
		X"FC",X"2C",X"FF",X"16",X"FF",X"00",X"78",X"C6",X"F0",X"D8",X"C5",X"D5",X"E5",X"CD",X"61",X"FB",
		X"0E",X"20",X"F3",X"1A",X"CD",X"53",X"FB",X"47",X"3E",X"02",X"D3",X"6A",X"70",X"3A",X"FE",X"DF",
		X"D3",X"6A",X"13",X"1A",X"CD",X"53",X"FB",X"47",X"3E",X"03",X"D3",X"6A",X"70",X"3A",X"FE",X"DF",
		X"D3",X"6A",X"13",X"23",X"0D",X"C2",X"23",X"FB",X"FB",X"3A",X"FE",X"DF",X"D3",X"6A",X"AF",X"E1",
		X"D1",X"C1",X"C9",X"E5",X"C5",X"67",X"06",X"08",X"29",X"1F",X"05",X"C2",X"58",X"FB",X"C1",X"E1",
		X"C9",X"78",X"0F",X"0F",X"0F",X"47",X"E6",X"F0",X"4F",X"78",X"E6",X"03",X"47",X"21",X"00",X"3C",
		X"09",X"C9",X"78",X"C6",X"F0",X"D8",X"7A",X"C6",X"D1",X"D8",X"7B",X"C6",X"8C",X"D8",X"C5",X"D5",
		X"E5",X"CD",X"61",X"FB",X"7B",X"07",X"5F",X"3E",X"40",X"82",X"57",X"06",X"02",X"D5",X"0E",X"10",
		X"F3",X"3E",X"02",X"D3",X"6A",X"1A",X"24",X"24",X"77",X"25",X"25",X"B6",X"12",X"3E",X"03",X"D3",
		X"6A",X"1A",X"24",X"24",X"77",X"25",X"25",X"B6",X"12",X"23",X"13",X"0D",X"C2",X"91",X"FB",X"3A",
		X"FE",X"DF",X"D3",X"6A",X"FB",X"D1",X"14",X"05",X"C2",X"8D",X"FB",X"C3",X"4E",X"FB",X"78",X"C6",
		X"F0",X"D8",X"7A",X"C6",X"D1",X"D8",X"7B",X"C6",X"8C",X"D8",X"C5",X"D5",X"E5",X"7B",X"07",X"6F",
		X"3E",X"40",X"82",X"67",X"E5",X"CD",X"61",X"FB",X"11",X"00",X"02",X"19",X"EB",X"E1",X"06",X"02",
		X"E5",X"0E",X"10",X"F3",X"3E",X"02",X"D3",X"6A",X"1A",X"77",X"3E",X"03",X"D3",X"6A",X"1A",X"77",
		X"13",X"23",X"0D",X"C2",X"E4",X"FB",X"3A",X"FE",X"DF",X"D3",X"6A",X"FB",X"E1",X"24",X"05",X"C2",
		X"E0",X"FB",X"C3",X"4E",X"FB",X"CD",X"BA",X"F8",X"D8",X"C5",X"D5",X"E5",X"CD",X"34",X"FC",X"CD",
		X"BA",X"F8",X"DA",X"30",X"FC",X"78",X"91",X"D4",X"34",X"FC",X"05",X"04",X"CD",X"84",X"F8",X"CD",
		X"34",X"FC",X"C5",X"41",X"CD",X"F0",X"F8",X"C1",X"CD",X"34",X"FC",X"4F",X"B8",X"C2",X"1B",X"FC",
		X"E1",X"D1",X"C1",X"C9",X"EB",X"78",X"41",X"4F",X"C9",X"CD",X"8A",X"FC",X"D8",X"C5",X"E5",X"E5",
		X"7C",X"C6",X"40",X"67",X"47",X"4D",X"CD",X"7A",X"FC",X"DA",X"6C",X"FC",X"F3",X"3E",X"02",X"D3",
		X"6A",X"0A",X"77",X"2B",X"77",X"3E",X"03",X"D3",X"6A",X"0A",X"77",X"23",X"77",X"7C",X"25",X"05",
		X"D6",X"40",X"92",X"C2",X"4D",X"FC",X"3A",X"FE",X"DF",X"D3",X"6A",X"FB",X"E1",X"7D",X"2D",X"93",
		X"C2",X"3F",X"FC",X"E1",X"CD",X"7A",X"FC",X"A7",X"C1",X"C9",X"7D",X"2E",X"F5",X"93",X"07",X"D8",
		X"3C",X"83",X"D8",X"C6",X"0A",X"D8",X"D6",X"0A",X"6F",X"C9",X"7A",X"C6",X"D1",X"D8",X"7B",X"C6",
		X"0B",X"D8",X"7C",X"C6",X"D0",X"D8",X"7D",X"C6",X"0A",X"D8",X"7C",X"92",X"D8",X"7D",X"93",X"C9",
		X"CD",X"8A",X"FC",X"D8",X"C5",X"E5",X"E5",X"7C",X"C6",X"40",X"47",X"4D",X"CD",X"DD",X"FC",X"DA",
		X"CF",X"FC",X"7C",X"C6",X"40",X"67",X"D5",X"3E",X"02",X"32",X"D6",X"DF",X"CD",X"EA",X"FC",X"3E",
		X"03",X"32",X"D6",X"DF",X"CD",X"EA",X"FC",X"D1",X"7D",X"2D",X"0D",X"93",X"C2",X"B6",X"FC",X"E1",
		X"7C",X"25",X"92",X"C2",X"A6",X"FC",X"E1",X"CD",X"DD",X"FC",X"A7",X"C1",X"C9",X"7C",X"92",X"07",
		X"3C",X"82",X"67",X"3E",X"2F",X"94",X"D0",X"26",X"2F",X"C9",X"F3",X"E5",X"3A",X"D6",X"DF",X"D3",
		X"6A",X"0A",X"21",X"00",X"00",X"16",X"08",X"29",X"29",X"07",X"D2",X"00",X"FD",X"2C",X"2C",X"2C",
		X"15",X"C2",X"F7",X"FC",X"55",X"5C",X"3A",X"FE",X"DF",X"D3",X"6A",X"E1",X"3A",X"D6",X"DF",X"D3",
		X"6A",X"73",X"25",X"72",X"3A",X"FE",X"DF",X"D3",X"6A",X"24",X"FB",X"C9",X"F5",X"E6",X"04",X"CA",
		X"29",X"FD",X"F1",X"3A",X"20",X"DF",X"C3",X"2A",X"FD",X"F1",X"32",X"DC",X"DF",X"C9",X"E5",X"21",
		X"39",X"FE",X"C3",X"39",X"FD",X"E5",X"21",X"32",X"FE",X"C5",X"01",X"00",X"20",X"C3",X"42",X"FD",
		X"E5",X"C5",X"3E",X"88",X"32",X"FF",X"DF",X"32",X"FA",X"DF",X"79",X"32",X"FD",X"DF",X"3E",X"25",
		X"D3",X"79",X"3E",X"A6",X"D3",X"63",X"78",X"D3",X"62",X"3E",X"10",X"D3",X"63",X"3E",X"76",X"D3",
		X"63",X"3E",X"C3",X"32",X"04",X"DF",X"22",X"FB",X"DF",X"21",X"71",X"FD",X"22",X"05",X"DF",X"C1",
		X"E1",X"F5",X"C5",X"D5",X"E5",X"3A",X"FA",X"DF",X"A7",X"C2",X"94",X"FD",X"3C",X"32",X"FA",X"DF",
		X"D3",X"60",X"3E",X"25",X"D3",X"79",X"3E",X"FD",X"D3",X"75",X"3E",X"61",X"D3",X"74",X"FB",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"AF",X"32",X"FA",X"DF",X"2A",X"FB",X"DF",X"7E",X"A7",X"C2",X"C6",X"FD",
		X"3E",X"FF",X"D3",X"75",X"AF",X"32",X"FF",X"DF",X"3E",X"76",X"D3",X"63",X"3E",X"96",X"D3",X"63",
		X"3E",X"0D",X"D3",X"62",X"3E",X"FF",X"D3",X"75",X"3E",X"20",X"D3",X"74",X"21",X"00",X"E0",X"22",
		X"05",X"DF",X"FB",X"C3",X"8F",X"FD",X"F2",X"D0",X"FD",X"32",X"FF",X"DF",X"23",X"C3",X"9B",X"FD",
		X"E6",X"70",X"0F",X"0F",X"0F",X"0F",X"4F",X"3A",X"FD",X"DF",X"81",X"E6",X"07",X"4F",X"7E",X"23",
		X"22",X"FB",X"DF",X"E6",X"0F",X"FE",X"0D",X"F2",X"0E",X"FE",X"3D",X"07",X"5F",X"16",X"00",X"21",
		X"1A",X"FE",X"19",X"56",X"23",X"5E",X"0D",X"CA",X"04",X"FE",X"A7",X"7A",X"1F",X"57",X"7B",X"1F",
		X"5F",X"C3",X"F6",X"FD",X"7B",X"D3",X"61",X"7A",X"D3",X"61",X"3E",X"05",X"D3",X"79",X"3A",X"FF",
		X"DF",X"E6",X"7F",X"07",X"3D",X"D3",X"60",X"C3",X"86",X"FD",X"EE",X"EA",X"E1",X"78",X"D4",X"E0",
		X"C8",X"D6",X"BD",X"A0",X"B2",X"FB",X"A8",X"EB",X"9F",X"70",X"96",X"88",X"8E",X"0C",X"86",X"01",
		X"7D",X"E1",X"90",X"5B",X"90",X"51",X"A0",X"65",X"00",X"88",X"5B",X"00",X"3E",X"AF",X"D3",X"1A",
		X"3E",X"FF",X"D3",X"1B",X"07",X"D3",X"1B",X"07",X"D3",X"1B",X"07",X"D3",X"1B",X"07",X"D3",X"1B",
		X"07",X"D3",X"1B",X"07",X"D3",X"1B",X"07",X"D3",X"1B",X"C9",X"3E",X"FF",X"D3",X"1B",X"D3",X"1B",
		X"D3",X"1B",X"D3",X"1B",X"D3",X"1B",X"D3",X"1B",X"D3",X"1B",X"D3",X"1B",X"DB",X"1B",X"C9",X"21",
		X"00",X"00",X"11",X"00",X"00",X"4F",X"CD",X"40",X"FE",X"79",X"CD",X"42",X"FE",X"7A",X"CD",X"42",
		X"FE",X"7B",X"CD",X"42",X"FE",X"7C",X"CD",X"42",X"FE",X"7D",X"CD",X"42",X"FE",X"3E",X"95",X"CD",
		X"42",X"FE",X"11",X"80",X"80",X"21",X"20",X"4E",X"CD",X"5A",X"FE",X"4F",X"92",X"BB",X"79",X"D0",
		X"2B",X"7C",X"B5",X"C2",X"98",X"FE",X"D6",X"01",X"C9",X"C5",X"D5",X"E5",X"11",X"FF",X"00",X"CD",
		X"95",X"FE",X"E1",X"D1",X"C1",X"C9",X"CD",X"3D",X"FE",X"06",X"10",X"CD",X"40",X"FE",X"05",X"C2",
		X"BB",X"FE",X"CD",X"3C",X"FE",X"3E",X"40",X"CD",X"6F",X"FE",X"FE",X"01",X"C0",X"3E",X"77",X"CD",
		X"6F",X"FE",X"E6",X"FE",X"C0",X"3E",X"69",X"CD",X"6F",X"FE",X"FE",X"01",X"CA",X"CD",X"FE",X"B7",
		X"C9",X"CD",X"A9",X"FE",X"D8",X"E5",X"EB",X"29",X"5C",X"65",X"AF",X"57",X"6F",X"3E",X"51",X"CD",
		X"75",X"FE",X"E1",X"D8",X"06",X"00",X"E5",X"11",X"01",X"FF",X"CD",X"95",X"FE",X"E1",X"FE",X"FE",
		X"C0",X"CD",X"5A",X"FE",X"77",X"23",X"CD",X"5A",X"FE",X"77",X"23",X"05",X"C2",X"01",X"FF",X"C9",
		X"3E",X"02",X"D3",X"6A",X"3A",X"80",X"28",X"E6",X"04",X"C0",X"AF",X"D3",X"6A",X"CD",X"24",X"FF",
		X"DA",X"3D",X"FE",X"E9",X"CD",X"B6",X"FE",X"37",X"C0",X"11",X"00",X"00",X"21",X"00",X"C0",X"CD",
		X"E1",X"FE",X"D8",X"CD",X"42",X"FF",X"D0",X"2A",X"C6",X"C1",X"EB",X"21",X"00",X"C0",X"CD",X"E1",
		X"FE",X"D8",X"CD",X"BA",X"FF",X"37",X"C0",X"2A",X"16",X"C0",X"EB",X"2A",X"0E",X"C0",X"3A",X"10",
		X"C0",X"19",X"3D",X"C2",X"51",X"FF",X"EB",X"2A",X"1C",X"C0",X"19",X"22",X"F0",X"C1",X"EB",X"2A",
		X"11",X"C0",X"4D",X"44",X"29",X"29",X"29",X"29",X"E5",X"79",X"E6",X"0F",X"C5",X"CC",X"9E",X"FF",
		X"D5",X"E5",X"06",X"0B",X"11",X"CB",X"FF",X"1A",X"BE",X"C2",X"AA",X"FF",X"13",X"23",X"05",X"C2",
		X"77",X"FF",X"C1",X"C1",X"C1",X"11",X"0F",X"00",X"19",X"5E",X"23",X"56",X"1B",X"1B",X"2A",X"F0",
		X"C1",X"3A",X"0D",X"C0",X"19",X"3D",X"C2",X"94",X"FF",X"D1",X"5A",X"57",X"19",X"EB",X"D5",X"21",
		X"00",X"C2",X"E5",X"CD",X"E1",X"FE",X"E1",X"D1",X"13",X"C9",X"E1",X"11",X"20",X"00",X"19",X"D1",
		X"C1",X"0B",X"78",X"B1",X"C2",X"69",X"FF",X"C1",X"37",X"C9",X"21",X"36",X"C0",X"7E",X"23",X"FE",
		X"46",X"C0",X"7E",X"23",X"FE",X"41",X"C0",X"7E",X"FE",X"54",X"C9",X"42",X"4F",X"4F",X"54",X"20",
		X"20",X"20",X"20",X"52",X"4F",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"59",X"2C",X"2C",X"2D",X"DE",X"E8",X"D8",
		X"D1",X"DA",X"D0",X"20",X"D7",X"D0",X"D3",X"E0",X"E3",X"D7",X"DA",X"D8",X"2D",X"00",X"FF",X"F6");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
