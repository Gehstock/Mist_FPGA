library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_1N is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_1N is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"02",X"61",X"C3",X"37",X"61",X"C3",X"74",X"61",X"C3",X"A6",X"61",X"C3",X"09",X"62",X"C3",
		X"81",X"62",X"C3",X"BE",X"62",X"C3",X"E5",X"62",X"C3",X"26",X"63",X"C3",X"9A",X"63",X"C3",X"BF",
		X"63",X"C3",X"79",X"64",X"C3",X"D8",X"64",X"C3",X"24",X"65",X"C3",X"69",X"65",X"C3",X"90",X"65",
		X"C3",X"FB",X"66",X"C3",X"18",X"67",X"C3",X"81",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C9",X"21",X"7A",X"82",X"11",X"18",X"85",X"06",X"09",X"C5",X"01",X"04",X"00",X"2B",X"2B",
		X"7E",X"FE",X"20",X"23",X"23",X"C2",X"29",X"61",X"2B",X"7E",X"FE",X"0C",X"23",X"D2",X"29",X"61",
		X"13",X"13",X"13",X"13",X"ED",X"B0",X"C3",X"2F",X"61",X"ED",X"B0",X"13",X"13",X"13",X"13",X"01",
		X"15",X"00",X"09",X"C1",X"10",X"D4",X"C9",X"3A",X"8D",X"80",X"B7",X"C2",X"73",X"61",X"DD",X"5E",
		X"0E",X"DD",X"56",X"0F",X"D5",X"01",X"80",X"01",X"21",X"10",X"00",X"EB",X"B7",X"ED",X"42",X"7D",
		X"B4",X"E1",X"C2",X"58",X"61",X"11",X"08",X"00",X"19",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"DD",
		X"5E",X"0A",X"DD",X"56",X"0B",X"19",X"DD",X"5E",X"07",X"DD",X"56",X"05",X"19",X"DD",X"75",X"07",
		X"DD",X"74",X"05",X"C9",X"78",X"92",X"57",X"79",X"93",X"5F",X"AF",X"B2",X"F2",X"8C",X"61",X"23",
		X"ED",X"44",X"57",X"7E",X"23",X"92",X"DA",X"A4",X"61",X"C3",X"91",X"61",X"7E",X"23",X"C3",X"84",
		X"61",X"AF",X"B3",X"F2",X"9A",X"61",X"23",X"ED",X"44",X"5F",X"7E",X"93",X"DA",X"A4",X"61",X"3E",
		X"01",X"C3",X"A5",X"61",X"AF",X"C9",X"3A",X"8D",X"80",X"B7",X"C2",X"08",X"62",X"DD",X"7E",X"11",
		X"FE",X"02",X"D2",X"C3",X"61",X"DD",X"5E",X"08",X"DD",X"56",X"09",X"DD",X"66",X"04",X"DD",X"6E",
		X"06",X"18",X"0F",X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"DD",X"66",X"05",X"DD",X"6E",X"07",X"3D",
		X"E6",X"01",X"B7",X"C2",X"D9",X"61",X"19",X"18",X"03",X"B7",X"ED",X"52",X"3E",X"01",X"DD",X"BE",
		X"11",X"DA",X"F7",X"61",X"7C",X"DD",X"BE",X"04",X"CA",X"EF",X"61",X"DD",X"36",X"18",X"00",X"DD",
		X"74",X"04",X"DD",X"75",X"06",X"18",X"11",X"7C",X"DD",X"BE",X"05",X"CA",X"02",X"62",X"DD",X"36",
		X"18",X"00",X"DD",X"74",X"05",X"DD",X"75",X"07",X"C9",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"DD",X"21",X"28",X"C8",X"3A",X"A0",X"81",X"3D",X"01",X"06",X"00",X"21",X"3B",X"DE",X"CD",X"F6",
		X"00",X"7E",X"87",X"16",X"00",X"5F",X"DD",X"19",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"E5",X"DD",
		X"E1",X"FD",X"21",X"80",X"84",X"0E",X"00",X"79",X"FE",X"18",X"CA",X"75",X"62",X"FD",X"71",X"00",
		X"21",X"C8",X"C9",X"16",X"00",X"DD",X"7E",X"00",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"5F",X"19",X"7E",X"FD",X"77",X"01",X"21",X"C8",X"C9",X"16",X"00",X"DD",X"7E",X"00",X"E6",X"0F",
		X"5F",X"19",X"7E",X"FD",X"77",X"02",X"0C",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"FD",X"23",X"18",X"C2",X"FD",X"36",X"00",X"FF",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",
		X"C9",X"C5",X"D5",X"E5",X"F5",X"3A",X"70",X"80",X"B7",X"20",X"16",X"3A",X"17",X"80",X"B7",X"C2",
		X"A1",X"62",X"3A",X"13",X"80",X"CB",X"7F",X"28",X"20",X"F1",X"F5",X"E6",X"7F",X"FE",X"20",X"20",
		X"18",X"21",X"01",X"87",X"01",X"01",X"00",X"3A",X"00",X"87",X"CD",X"F6",X"00",X"F1",X"77",X"3A",
		X"00",X"87",X"3C",X"32",X"00",X"87",X"C3",X"BA",X"62",X"F1",X"E1",X"D1",X"C1",X"C9",X"3A",X"00",
		X"87",X"B7",X"C8",X"21",X"01",X"87",X"7E",X"32",X"00",X"B8",X"3A",X"00",X"87",X"3D",X"32",X"00",
		X"87",X"C8",X"47",X"21",X"01",X"87",X"E5",X"DD",X"E1",X"DD",X"23",X"DD",X"7E",X"00",X"77",X"23",
		X"DD",X"23",X"10",X"F7",X"C9",X"3A",X"70",X"80",X"FE",X"00",X"28",X"08",X"3A",X"14",X"80",X"E6",
		X"18",X"0F",X"0F",X"0F",X"21",X"01",X"63",X"16",X"00",X"5F",X"19",X"7E",X"32",X"A8",X"81",X"18",
		X"04",X"00",X"01",X"03",X"07",X"3A",X"70",X"80",X"FE",X"00",X"28",X"08",X"3A",X"14",X"80",X"E6",
		X"60",X"07",X"07",X"07",X"21",X"21",X"63",X"16",X"00",X"5F",X"19",X"7E",X"32",X"A9",X"81",X"18",
		X"04",X"00",X"00",X"01",X"03",X"C9",X"C5",X"D5",X"E5",X"FE",X"11",X"D2",X"96",X"63",X"32",X"86",
		X"89",X"FE",X"10",X"CA",X"91",X"63",X"FE",X"08",X"D2",X"69",X"63",X"21",X"3A",X"DE",X"01",X"06",
		X"00",X"3A",X"A0",X"81",X"3D",X"CD",X"F6",X"00",X"7E",X"F5",X"21",X"00",X"D7",X"01",X"10",X"00",
		X"CD",X"F6",X"00",X"11",X"A0",X"8C",X"ED",X"B0",X"F1",X"21",X"80",X"D7",X"01",X"10",X"00",X"CD",
		X"F6",X"00",X"11",X"80",X"8C",X"ED",X"B0",X"18",X"28",X"D6",X"08",X"87",X"21",X"81",X"63",X"16",
		X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",X"11",X"70",X"8C",X"01",X"10",X"00",X"ED",X"B0",X"18",
		X"10",X"00",X"D8",X"10",X"D8",X"20",X"D8",X"30",X"D8",X"40",X"D8",X"50",X"D8",X"60",X"D8",X"70",
		X"D8",X"3E",X"01",X"32",X"85",X"89",X"E1",X"D1",X"C1",X"C9",X"3A",X"85",X"89",X"B7",X"C8",X"3A",
		X"86",X"89",X"FE",X"10",X"CA",X"B4",X"63",X"F5",X"21",X"70",X"8C",X"11",X"70",X"9C",X"01",X"40",
		X"00",X"ED",X"B0",X"F1",X"CB",X"E7",X"32",X"00",X"9E",X"3E",X"00",X"32",X"85",X"89",X"C9",X"F5",
		X"E5",X"DD",X"E5",X"D5",X"3A",X"9E",X"81",X"E6",X"0F",X"5F",X"F5",X"3A",X"AC",X"81",X"57",X"C5",
		X"B7",X"CB",X"38",X"CB",X"19",X"B7",X"CB",X"38",X"CB",X"19",X"B7",X"CB",X"38",X"CB",X"19",X"B7",
		X"CB",X"38",X"CB",X"19",X"B7",X"2A",X"B1",X"81",X"7D",X"81",X"27",X"6F",X"7C",X"88",X"27",X"67",
		X"22",X"B1",X"81",X"C1",X"21",X"9C",X"81",X"7E",X"81",X"27",X"77",X"23",X"7E",X"88",X"27",X"77",
		X"23",X"7E",X"CE",X"00",X"27",X"77",X"23",X"7E",X"CE",X"00",X"27",X"77",X"3A",X"AE",X"81",X"FE",
		X"FF",X"28",X"10",X"3A",X"9E",X"81",X"E6",X"0F",X"BB",X"28",X"08",X"5F",X"3A",X"AD",X"81",X"3C",
		X"32",X"AD",X"81",X"7A",X"FE",X"00",X"28",X"04",X"15",X"C3",X"CF",X"63",X"3A",X"27",X"80",X"B7",
		X"CA",X"3A",X"64",X"DD",X"21",X"61",X"CA",X"C3",X"3E",X"64",X"DD",X"21",X"4F",X"CA",X"3A",X"70",
		X"80",X"B7",X"CA",X"48",X"64",X"CD",X"D5",X"00",X"F1",X"3A",X"B2",X"81",X"FE",X"05",X"38",X"20",
		X"D6",X"05",X"27",X"FE",X"05",X"30",X"F9",X"32",X"B2",X"81",X"3A",X"88",X"80",X"FE",X"00",X"20",
		X"0F",X"3A",X"AC",X"81",X"FE",X"04",X"30",X"08",X"3A",X"00",X"89",X"CB",X"C7",X"32",X"00",X"89",
		X"CD",X"DD",X"5F",X"D1",X"DD",X"E1",X"E1",X"F1",X"C9",X"CD",X"24",X"65",X"CD",X"D8",X"64",X"3A",
		X"13",X"80",X"E6",X"03",X"FE",X"00",X"20",X"06",X"DD",X"21",X"2B",X"66",X"18",X"18",X"FE",X"01",
		X"20",X"06",X"DD",X"21",X"4B",X"66",X"18",X"0E",X"FE",X"02",X"20",X"06",X"DD",X"21",X"6B",X"66",
		X"18",X"04",X"DD",X"21",X"8B",X"66",X"CD",X"D2",X"00",X"DD",X"21",X"AB",X"66",X"CD",X"D2",X"00",
		X"3E",X"20",X"CD",X"FC",X"00",X"01",X"00",X"00",X"3E",X"01",X"32",X"6E",X"80",X"3E",X"02",X"32",
		X"8C",X"80",X"3A",X"6E",X"80",X"FE",X"00",X"20",X"F9",X"03",X"78",X"FE",X"02",X"20",X"E9",X"79",
		X"FE",X"58",X"20",X"E4",X"CD",X"69",X"65",X"C9",X"C3",X"00",X"6A",X"DD",X"E5",X"DD",X"21",X"00",
		X"85",X"06",X"A8",X"0E",X"06",X"26",X"21",X"79",X"FE",X"00",X"28",X"32",X"FE",X"04",X"20",X"02",
		X"06",X"B4",X"DD",X"70",X"00",X"DD",X"36",X"01",X"24",X"DD",X"74",X"02",X"DD",X"36",X"03",X"20",
		X"04",X"11",X"08",X"00",X"DD",X"19",X"DD",X"70",X"00",X"DD",X"36",X"01",X"24",X"DD",X"74",X"02",
		X"DD",X"36",X"03",X"40",X"DD",X"19",X"04",X"0D",X"3E",X"20",X"84",X"67",X"18",X"C9",X"DD",X"E1",
		X"E1",X"D1",X"C1",X"C9",X"C5",X"D5",X"E5",X"3A",X"64",X"88",X"F6",X"80",X"32",X"64",X"88",X"21",
		X"1A",X"0F",X"11",X"00",X"88",X"01",X"0A",X"00",X"ED",X"B0",X"21",X"FF",X"0F",X"22",X"42",X"8C",
		X"21",X"0F",X"00",X"22",X"44",X"8C",X"21",X"AF",X"00",X"22",X"46",X"8C",X"21",X"0F",X"08",X"22",
		X"48",X"8C",X"21",X"AD",X"0F",X"11",X"4A",X"8C",X"01",X"06",X"00",X"ED",X"B0",X"3A",X"00",X"88",
		X"E6",X"7F",X"32",X"00",X"88",X"E1",X"D1",X"C1",X"C9",X"C5",X"D5",X"E5",X"3A",X"00",X"88",X"F6",
		X"80",X"32",X"00",X"88",X"11",X"42",X"8C",X"21",X"42",X"D5",X"01",X"0E",X"00",X"ED",X"B0",X"3A",
		X"64",X"88",X"E6",X"7F",X"32",X"64",X"88",X"3E",X"00",X"CD",X"F6",X"4F",X"E1",X"D1",X"C1",X"C9",
		X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"CB",X"00",X"76",X"CA",X"22",X"66",X"DD",
		X"7E",X"03",X"FE",X"00",X"C2",X"22",X"66",X"DD",X"7E",X"04",X"FE",X"00",X"CA",X"22",X"66",X"FE",
		X"01",X"20",X"45",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"CD",X"DE",X"00",X"E5",X"FD",X"E1",X"3A",
		X"AC",X"81",X"26",X"00",X"6F",X"29",X"29",X"29",X"11",X"D3",X"66",X"19",X"7E",X"FD",X"77",X"E0",
		X"23",X"7E",X"FD",X"77",X"E1",X"23",X"7E",X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"01",X"11",
		X"00",X"04",X"FD",X"19",X"23",X"7E",X"FD",X"77",X"E0",X"23",X"7E",X"FD",X"77",X"E1",X"23",X"7E",
		X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"01",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"1F",
		X"38",X"20",X"DD",X"36",X"04",X"00",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"CD",X"DE",X"00",X"E5",
		X"FD",X"E1",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"E1",X"00",X"FD",X"36",
		X"E0",X"00",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"13",X"09",X"31",X"05",X"43",
		X"00",X"4F",X"00",X"49",X"00",X"4E",X"00",X"02",X"FF",X"00",X"00",X"31",X"05",X"43",X"00",X"52",
		X"00",X"45",X"00",X"44",X"00",X"49",X"00",X"54",X"00",X"FF",X"FF",X"13",X"09",X"31",X"05",X"43",
		X"00",X"4F",X"00",X"49",X"00",X"4E",X"00",X"02",X"FF",X"00",X"00",X"32",X"05",X"43",X"00",X"52",
		X"00",X"45",X"00",X"44",X"00",X"49",X"00",X"54",X"00",X"FF",X"FF",X"13",X"09",X"31",X"05",X"43",
		X"00",X"4F",X"00",X"49",X"00",X"4E",X"00",X"02",X"FF",X"00",X"00",X"33",X"05",X"43",X"00",X"52",
		X"00",X"45",X"00",X"44",X"00",X"49",X"00",X"54",X"00",X"FF",X"FF",X"13",X"09",X"31",X"05",X"43",
		X"00",X"4F",X"00",X"49",X"00",X"4E",X"00",X"02",X"FF",X"00",X"00",X"36",X"05",X"43",X"00",X"52",
		X"00",X"45",X"00",X"44",X"00",X"49",X"00",X"54",X"00",X"FF",X"FF",X"1C",X"07",X"3A",X"05",X"3B",
		X"05",X"31",X"05",X"39",X"05",X"38",X"05",X"34",X"05",X"00",X"00",X"54",X"0F",X"45",X"0F",X"48",
		X"0F",X"4B",X"0F",X"41",X"0F",X"4E",X"0F",X"00",X"00",X"4C",X"05",X"54",X"05",X"44",X"05",X"2E",
		X"05",X"FF",X"FF",X"80",X"81",X"82",X"83",X"15",X"15",X"15",X"15",X"90",X"91",X"92",X"93",X"15",
		X"15",X"15",X"15",X"94",X"95",X"96",X"97",X"15",X"15",X"15",X"15",X"98",X"99",X"9A",X"9B",X"15",
		X"15",X"15",X"15",X"9C",X"9D",X"9E",X"9F",X"15",X"15",X"15",X"15",X"F5",X"E5",X"21",X"00",X"00",
		X"22",X"9F",X"80",X"22",X"A1",X"80",X"22",X"A3",X"80",X"3A",X"6D",X"67",X"32",X"00",X"85",X"3A",
		X"6E",X"67",X"32",X"01",X"85",X"E1",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"DD",X"21",X"9F",X"80",X"DD",X"7E",X"00",X"FE",X"0E",X"38",X"36",X"FD",X"21",X"6D",X"67",X"ED",
		X"5B",X"A0",X"80",X"B7",X"FD",X"19",X"FD",X"7E",X"00",X"FE",X"FF",X"20",X"0C",X"FD",X"21",X"6D",
		X"67",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"FD",X"7E",X"00",X"32",X"00",X"85",X"FD",
		X"7E",X"01",X"32",X"01",X"85",X"DD",X"36",X"00",X"00",X"2A",X"A0",X"80",X"23",X"23",X"22",X"A0",
		X"80",X"DD",X"34",X"00",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"31",X"00",X"32",
		X"00",X"31",X"00",X"32",X"80",X"31",X"00",X"33",X"00",X"31",X"00",X"33",X"00",X"FF",X"FF",X"FF",
		X"FF",X"DD",X"21",X"10",X"85",X"3A",X"02",X"89",X"FE",X"FF",X"28",X"3E",X"3E",X"FF",X"32",X"02",
		X"89",X"DD",X"36",X"00",X"18",X"DD",X"36",X"01",X"0B",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",
		X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"3A",X"9B",X"81",X"3C",X"32",X"9B",X"81",
		X"FE",X"08",X"38",X"02",X"3E",X"07",X"4F",X"0D",X"06",X"10",X"79",X"FE",X"00",X"28",X"07",X"78",
		X"C6",X"10",X"47",X"0D",X"18",X"F4",X"78",X"32",X"03",X"89",X"3A",X"13",X"85",X"FE",X"F0",X"CA",
		X"FE",X"67",X"3A",X"12",X"85",X"FE",X"78",X"28",X"16",X"30",X"08",X"3C",X"FE",X"78",X"28",X"09",
		X"3C",X"18",X"06",X"3D",X"FE",X"78",X"28",X"01",X"3D",X"32",X"12",X"85",X"C3",X"7A",X"68",X"3A",
		X"13",X"85",X"3C",X"FE",X"F0",X"28",X"01",X"3C",X"32",X"13",X"85",X"C3",X"7A",X"68",X"3A",X"04",
		X"89",X"FE",X"01",X"28",X"24",X"3A",X"03",X"89",X"47",X"3A",X"12",X"85",X"B8",X"28",X"08",X"3D",
		X"B8",X"28",X"04",X"3D",X"B8",X"20",X"0C",X"47",X"3E",X"01",X"32",X"04",X"89",X"3E",X"30",X"32",
		X"05",X"89",X"78",X"32",X"12",X"85",X"C3",X"7A",X"68",X"3A",X"05",X"89",X"3D",X"32",X"05",X"89",
		X"FE",X"00",X"C2",X"7A",X"68",X"3E",X"1F",X"CD",X"FC",X"00",X"21",X"00",X"00",X"22",X"10",X"85",
		X"DD",X"46",X"02",X"DD",X"4E",X"03",X"CD",X"DE",X"00",X"E5",X"FD",X"E1",X"FD",X"36",X"00",X"0E",
		X"FD",X"36",X"01",X"0F",X"FD",X"36",X"E0",X"0C",X"FD",X"36",X"E1",X"0D",X"11",X"00",X"04",X"B7",
		X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"E0",X"00",X"FD",X"36",
		X"E1",X"00",X"3E",X"00",X"32",X"02",X"89",X"32",X"88",X"80",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C5",X"D5",X"E5",X"CD",X"CF",X"00",X"10",X"6A",X"02",X"C3",X"DB",X"64",X"00",X"00",X"00",X"00",
		X"20",X"6A",X"60",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"04",X"22",X"14",X"20",X"14",X"26",X"14",X"24",X"14",X"2A",X"14",X"28",X"14",X"2E",X"14",
		X"2C",X"14",X"32",X"14",X"30",X"14",X"36",X"14",X"34",X"14",X"3A",X"14",X"38",X"14",X"3E",X"14",
		X"3C",X"14",X"42",X"14",X"40",X"14",X"46",X"14",X"44",X"14",X"4A",X"14",X"48",X"14",X"4E",X"14",
		X"4C",X"14",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"04",X"23",X"14",X"21",X"14",X"27",X"14",X"25",X"14",X"2B",X"14",X"29",X"14",X"2F",X"14",
		X"2D",X"14",X"33",X"14",X"31",X"14",X"37",X"14",X"35",X"14",X"3B",X"14",X"39",X"14",X"3F",X"14",
		X"3D",X"14",X"43",X"14",X"41",X"14",X"47",X"14",X"45",X"14",X"4B",X"14",X"49",X"14",X"4F",X"14",
		X"4D",X"14",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"08",X"06",X"10",X"1E",X"00",X"02",X"05",X"05",X"15",X"02",X"11",X"03",X"01",X"04",X"11",
		X"05",X"01",X"05",X"11",X"04",X"05",X"03",X"15",X"0A",X"05",X"04",X"15",X"04",X"05",X"05",X"15",
		X"06",X"05",X"03",X"01",X"42",X"09",X"01",X"08",X"01",X"00",X"45",X"06",X"02",X"16",X"3A",X"02",
		X"02",X"16",X"28",X"02",X"02",X"15",X"27",X"05",X"15",X"00",X"02",X"15",X"70",X"05",X"02",X"16",
		X"33",X"06",X"02",X"10",X"0E",X"0A",X"30",X"00",X"02",X"10",X"05",X"00",X"02",X"10",X"10",X"00",
		X"02",X"10",X"05",X"00",X"02",X"10",X"60",X"00",X"0A",X"01",X"0A",X"02",X"02",X"16",X"21",X"06",
		X"02",X"10",X"10",X"01",X"2D",X"0A",X"40",X"09",X"02",X"16",X"10",X"06",X"02",X"16",X"02",X"06",
		X"02",X"16",X"35",X"06",X"70",X"00",X"02",X"14",X"42",X"04",X"30",X"05",X"25",X"00",X"53",X"09",
		X"53",X"0A",X"0A",X"00",X"98",X"00",X"30",X"02",X"02",X"16",X"20",X"06",X"05",X"05",X"10",X"06",
		X"1C",X"05",X"02",X"15",X"24",X"08",X"02",X"10",X"05",X"00",X"02",X"10",X"10",X"00",X"02",X"10",
		X"05",X"00",X"02",X"10",X"10",X"00",X"02",X"10",X"05",X"00",X"02",X"10",X"10",X"00",X"05",X"01",
		X"02",X"11",X"20",X"01",X"02",X"11",X"40",X"01",X"42",X"08",X"27",X"02",X"02",X"16",X"35",X"06",
		X"30",X"08",X"60",X"01",X"02",X"10",X"20",X"04",X"10",X"06",X"10",X"05",X"18",X"04",X"02",X"16",
		X"30",X"06",X"02",X"15",X"30",X"05",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"06",X"05",
		X"1E",X"05",X"0E",X"02",X"02",X"10",X"1E",X"00",X"03",X"05",X"03",X"15",X"03",X"05",X"10",X"05",
		X"01",X"00",X"10",X"16",X"10",X"06",X"10",X"16",X"05",X"06",X"05",X"16",X"05",X"06",X"05",X"16",
		X"30",X"05",X"10",X"00",X"03",X"10",X"28",X"00",X"08",X"02",X"05",X"16",X"05",X"06",X"05",X"16",
		X"05",X"02",X"05",X"16",X"02",X"06",X"02",X"16",X"02",X"06",X"02",X"16",X"02",X"06",X"02",X"16",
		X"05",X"06",X"05",X"16",X"05",X"06",X"02",X"16",X"02",X"06",X"02",X"16",X"02",X"06",X"02",X"16",
		X"02",X"06",X"02",X"16",X"02",X"06",X"02",X"16",X"05",X"06",X"05",X"16",X"08",X"00",X"02",X"15",
		X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"15",X"02",X"05",
		X"80",X"05",X"50",X"00",X"45",X"02",X"40",X"00",X"02",X"10",X"53",X"00",X"05",X"15",X"05",X"05",
		X"02",X"15",X"05",X"06",X"02",X"16",X"02",X"06",X"03",X"16",X"03",X"06",X"03",X"16",X"03",X"06",
		X"03",X"16",X"03",X"06",X"03",X"16",X"03",X"06",X"03",X"16",X"18",X"06",X"32",X"08",X"01",X"00",
		X"02",X"10",X"2A",X"04",X"02",X"15",X"35",X"05",X"1C",X"00",X"05",X"16",X"05",X"06",X"05",X"16",
		X"05",X"02",X"03",X"12",X"10",X"00",X"03",X"02",X"02",X"05",X"02",X"05",X"02",X"05",X"18",X"01",
		X"50",X"00",X"02",X"10",X"13",X"00",X"02",X"15",X"05",X"00",X"3D",X"09",X"60",X"00",X"30",X"01",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"06",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",
		X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",X"02",X"05",X"02",X"15",
		X"02",X"05",X"02",X"15",X"02",X"05",X"40",X"01",X"30",X"00",X"40",X"02",X"02",X"10",X"10",X"04",
		X"18",X"05",X"02",X"15",X"20",X"01",X"10",X"02",X"02",X"10",X"20",X"04",X"02",X"10",X"05",X"05",
		X"05",X"15",X"05",X"05",X"05",X"15",X"10",X"05",X"20",X"02",X"20",X"08",X"02",X"10",X"20",X"04",
		X"02",X"10",X"10",X"01",X"20",X"00",X"02",X"10",X"02",X"00",X"02",X"10",X"05",X"00",X"02",X"10",
		X"02",X"00",X"02",X"10",X"05",X"00",X"02",X"10",X"02",X"00",X"02",X"10",X"05",X"00",X"02",X"10",
		X"02",X"00",X"02",X"10",X"05",X"00",X"15",X"0A",X"15",X"08",X"18",X"01",X"44",X"00",X"0C",X"01",
		X"28",X"02",X"22",X"0A",X"10",X"08",X"02",X"14",X"16",X"04",X"13",X"06",X"02",X"12",X"10",X"02",
		X"10",X"01",X"02",X"00",X"10",X"01",X"0E",X"00",X"02",X"14",X"02",X"06",X"02",X"16",X"02",X"06",
		X"02",X"16",X"02",X"06",X"02",X"16",X"12",X"06",X"40",X"00",X"44",X"01",X"10",X"00",X"02",X"10",
		X"40",X"04",X"02",X"16",X"0A",X"06",X"33",X"08",X"02",X"10",X"20",X"04",X"1E",X"05",X"02",X"10",
		X"05",X"06",X"05",X"16",X"05",X"06",X"05",X"16",X"05",X"06",X"05",X"16",X"05",X"06",X"05",X"16",
		X"05",X"06",X"05",X"16",X"05",X"06",X"05",X"16",X"10",X"06",X"08",X"00",X"05",X"15",X"05",X"05",
		X"05",X"15",X"05",X"05",X"05",X"15",X"05",X"05",X"10",X"08",X"10",X"0A",X"10",X"00",X"10",X"01",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"2C",X"70",
		X"58",X"70",X"84",X"70",X"94",X"70",X"C0",X"70",X"D0",X"70",X"C0",X"70",X"F8",X"70",X"08",X"71",
		X"18",X"71",X"44",X"71",X"54",X"71",X"6C",X"71",X"7C",X"71",X"A8",X"71",X"09",X"06",X"12",X"0B",
		X"10",X"0B",X"12",X"1B",X"10",X"1B",X"12",X"1B",X"10",X"1B",X"12",X"1B",X"10",X"1B",X"12",X"1B",
		X"10",X"1B",X"12",X"1B",X"10",X"1B",X"12",X"1B",X"10",X"1B",X"12",X"1B",X"10",X"1B",X"12",X"1B",
		X"10",X"1B",X"1E",X"0B",X"1C",X"0B",X"FF",X"FF",X"0A",X"06",X"13",X"0B",X"11",X"0B",X"13",X"1B",
		X"11",X"1B",X"13",X"1B",X"11",X"1B",X"13",X"1B",X"11",X"1B",X"13",X"1B",X"11",X"1B",X"13",X"1B",
		X"11",X"1B",X"13",X"1B",X"11",X"1B",X"13",X"1B",X"11",X"1B",X"13",X"1B",X"11",X"1B",X"1F",X"0B",
		X"1D",X"0B",X"FF",X"FF",X"0B",X"06",X"16",X"1B",X"14",X"1B",X"10",X"FF",X"00",X"00",X"1E",X"1B",
		X"1C",X"1B",X"FF",X"FF",X"0C",X"06",X"17",X"1B",X"15",X"1B",X"00",X"00",X"59",X"00",X"4F",X"00",
		X"55",X"00",X"3D",X"00",X"56",X"00",X"45",X"00",X"00",X"00",X"47",X"00",X"4F",X"00",X"54",X"00",
		X"54",X"00",X"45",X"00",X"4E",X"00",X"00",X"00",X"00",X"00",X"1F",X"1B",X"1D",X"1B",X"FF",X"FF",
		X"0D",X"06",X"16",X"1B",X"14",X"1B",X"10",X"FF",X"00",X"00",X"1E",X"1B",X"1C",X"1B",X"FF",X"FF",
		X"0E",X"06",X"17",X"1B",X"15",X"1B",X"04",X"FF",X"00",X"00",X"46",X"00",X"49",X"00",X"52",X"00",
		X"45",X"00",X"00",X"00",X"42",X"00",X"4F",X"00",X"4D",X"00",X"42",X"00",X"53",X"00",X"2E",X"00",
		X"00",X"00",X"1F",X"1B",X"1D",X"1B",X"FF",X"FF",X"0F",X"06",X"16",X"1B",X"14",X"1B",X"10",X"FF",
		X"00",X"00",X"1E",X"1B",X"1C",X"1B",X"FF",X"FF",X"10",X"06",X"17",X"1B",X"15",X"1B",X"10",X"FF",
		X"00",X"00",X"1F",X"1B",X"1D",X"1B",X"FF",X"FF",X"11",X"06",X"16",X"1B",X"14",X"1B",X"00",X"00",
		X"53",X"05",X"50",X"05",X"45",X"05",X"43",X"05",X"49",X"05",X"41",X"05",X"4C",X"05",X"00",X"00",
		X"42",X"05",X"4F",X"05",X"4E",X"05",X"55",X"05",X"53",X"05",X"00",X"00",X"00",X"00",X"1E",X"1B",
		X"1C",X"1B",X"FF",X"FF",X"12",X"06",X"17",X"1B",X"15",X"1B",X"10",X"FF",X"00",X"00",X"1F",X"1B",
		X"1D",X"1B",X"FF",X"FF",X"13",X"06",X"16",X"1B",X"14",X"1B",X"0A",X"FF",X"00",X"00",X"3E",X"05",
		X"3C",X"05",X"04",X"FF",X"00",X"00",X"1E",X"1B",X"1C",X"1B",X"FF",X"FF",X"14",X"06",X"17",X"1B",
		X"15",X"1B",X"10",X"FF",X"00",X"00",X"1F",X"1B",X"1D",X"1B",X"FF",X"FF",X"15",X"06",X"16",X"0B",
		X"14",X"0B",X"1A",X"1B",X"18",X"1B",X"1A",X"1B",X"18",X"1B",X"1A",X"1B",X"18",X"1B",X"1A",X"1B",
		X"18",X"1B",X"1A",X"1B",X"18",X"1B",X"1A",X"1B",X"18",X"1B",X"1A",X"1B",X"18",X"1B",X"1A",X"1B",
		X"18",X"1B",X"1A",X"0B",X"18",X"0B",X"FF",X"FF",X"16",X"06",X"17",X"0B",X"15",X"0B",X"1B",X"1B",
		X"19",X"1B",X"1B",X"1B",X"19",X"1B",X"1B",X"1B",X"19",X"1B",X"1B",X"1B",X"19",X"1B",X"1B",X"1B",
		X"19",X"1B",X"1B",X"1B",X"19",X"1B",X"1B",X"1B",X"19",X"1B",X"1B",X"1B",X"19",X"1B",X"1B",X"0B",
		X"19",X"0B",X"FF",X"FF",X"E4",X"71",X"EC",X"71",X"FC",X"71",X"04",X"72",X"14",X"72",X"1C",X"72",
		X"2C",X"72",X"34",X"72",X"0E",X"09",X"32",X"0F",X"30",X"0F",X"FF",X"FF",X"13",X"0B",X"00",X"00",
		X"31",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",X"FF",X"FF",X"0E",X"09",X"32",X"0F",
		X"31",X"0F",X"FF",X"FF",X"13",X"0B",X"00",X"00",X"32",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",
		X"30",X"0F",X"FF",X"FF",X"0E",X"09",X"32",X"0F",X"32",X"0F",X"FF",X"FF",X"13",X"0B",X"00",X"00",
		X"33",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",X"FF",X"FF",X"0E",X"09",X"32",X"0F",
		X"33",X"0F",X"FF",X"FF",X"13",X"0B",X"00",X"00",X"35",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",
		X"30",X"0F",X"FF",X"FF",X"13",X"0B",X"82",X"89",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"73",X"1C",X"73",X"28",X"73",X"38",X"73",X"44",X"73",X"08",X"11",X"60",X"09",X"62",X"09",
		X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"0B",X"08",X"60",X"09",
		X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"14",X"0E",X"60",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"17",X"05",X"60",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"1A",X"12",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"6E",X"73",X"82",X"73",X"8E",X"73",
		X"9A",X"73",X"A6",X"73",X"B2",X"73",X"BE",X"73",X"CA",X"73",X"D6",X"73",X"E2",X"73",X"08",X"0C",
		X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",
		X"FF",X"FF",X"0C",X"08",X"64",X"09",X"0E",X"FF",X"00",X"00",X"64",X"09",X"FF",X"FF",X"0D",X"08",
		X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"0E",X"08",X"67",X"09",X"0E",X"FF",
		X"00",X"00",X"67",X"09",X"FF",X"FF",X"0F",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",
		X"FF",X"FF",X"10",X"08",X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"11",X"08",
		X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"12",X"08",X"67",X"09",X"0E",X"FF",
		X"00",X"00",X"67",X"09",X"FF",X"FF",X"13",X"08",X"65",X"09",X"0E",X"FF",X"00",X"00",X"65",X"09",
		X"FF",X"FF",X"17",X"0C",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",
		X"63",X"09",X"61",X"09",X"FF",X"FF",X"08",X"74",X"16",X"74",X"2C",X"74",X"3C",X"74",X"42",X"74",
		X"48",X"74",X"4E",X"74",X"54",X"74",X"5A",X"74",X"08",X"0F",X"60",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"61",X"09",X"FF",X"FF",X"0B",X"02",X"6C",X"09",X"62",X"09",X"63",X"09",X"62",X"09",
		X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"0E",X"14",X"68",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"0F",X"14",X"66",X"09",
		X"FF",X"FF",X"10",X"14",X"67",X"09",X"FF",X"FF",X"11",X"14",X"66",X"09",X"FF",X"FF",X"12",X"14",
		X"67",X"09",X"FF",X"FF",X"13",X"14",X"66",X"09",X"FF",X"FF",X"14",X"08",X"60",X"09",X"62",X"09",
		X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",
		X"63",X"09",X"62",X"09",X"6B",X"09",X"FF",X"FF",X"90",X"74",X"9C",X"74",X"A8",X"74",X"B4",X"74",
		X"C0",X"74",X"CC",X"74",X"EC",X"74",X"0C",X"75",X"18",X"75",X"24",X"75",X"30",X"75",X"3C",X"75",
		X"06",X"0B",X"64",X"09",X"08",X"FF",X"00",X"00",X"64",X"09",X"FF",X"FF",X"07",X"0B",X"66",X"09",
		X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"08",X"0B",X"67",X"09",X"08",X"FF",X"00",X"00",
		X"67",X"09",X"FF",X"FF",X"09",X"0B",X"66",X"09",X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",
		X"0A",X"0B",X"67",X"09",X"08",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"0B",X"06",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"6B",X"09",X"08",X"FF",X"00",X"00",X"6A",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"14",X"06",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"69",X"09",X"08",X"FF",X"00",X"00",X"68",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"15",X"0B",X"66",X"09",
		X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"16",X"0B",X"67",X"09",X"08",X"FF",X"00",X"00",
		X"67",X"09",X"FF",X"FF",X"17",X"0B",X"66",X"09",X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",
		X"18",X"0B",X"67",X"09",X"08",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"19",X"0B",X"65",X"09",
		X"08",X"FF",X"00",X"00",X"65",X"09",X"FF",X"FF",X"50",X"75",X"74",X"75",X"90",X"75",X"B4",X"75",
		X"08",X"05",X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"05",X"FF",X"00",X"00",X"60",X"09",
		X"62",X"09",X"63",X"09",X"61",X"09",X"05",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"0E",X"09",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",
		X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",
		X"14",X"05",X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"05",X"FF",X"00",X"00",X"60",X"09",
		X"62",X"09",X"63",X"09",X"61",X"09",X"05",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"1A",X"09",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",
		X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",
		X"D8",X"75",X"E4",X"75",X"04",X"76",X"24",X"76",X"08",X"0E",X"60",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"0E",X"08",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"11",X"08",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"17",X"0E",X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",
		X"34",X"76",X"50",X"76",X"08",X"06",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",
		X"0A",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",
		X"17",X"06",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"0A",X"FF",X"00",X"00",
		X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"72",X"76",X"8E",X"76",
		X"9A",X"76",X"08",X"09",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"04",X"FF",
		X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"14",X"0E",
		X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"17",X"05",X"60",X"09",X"62",X"09",
		X"63",X"09",X"61",X"09",X"0E",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",
		X"FF",X"FF",X"CC",X"76",X"F0",X"76",X"FC",X"76",X"08",X"77",X"14",X"77",X"20",X"77",X"2C",X"77",
		X"38",X"77",X"44",X"77",X"50",X"77",X"5C",X"77",X"68",X"77",X"74",X"77",X"08",X"08",X"68",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"69",X"09",X"FF",X"FF",
		X"09",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"0A",X"08",X"67",X"09",
		X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"0B",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",
		X"66",X"09",X"FF",X"FF",X"0C",X"08",X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",
		X"0D",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"0E",X"08",X"67",X"09",
		X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"0F",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",
		X"66",X"09",X"FF",X"FF",X"10",X"08",X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",
		X"11",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"12",X"08",X"67",X"09",
		X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"13",X"08",X"65",X"09",X"0E",X"FF",X"00",X"00",
		X"65",X"09",X"FF",X"FF",X"14",X"0E",X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",
		X"A0",X"77",X"AA",X"77",X"B0",X"77",X"B6",X"77",X"C2",X"77",X"D4",X"77",X"DA",X"77",X"E0",X"77",
		X"EC",X"77",X"04",X"78",X"10",X"78",X"16",X"78",X"1C",X"78",X"3A",X"78",X"40",X"78",X"46",X"78",
		X"05",X"0E",X"68",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"06",X"0E",X"66",X"09",X"FF",X"FF",
		X"07",X"0E",X"67",X"09",X"FF",X"FF",X"08",X"0E",X"6A",X"09",X"62",X"09",X"63",X"09",X"61",X"09",
		X"FF",X"FF",X"0B",X"0B",X"60",X"09",X"62",X"09",X"63",X"09",X"6E",X"09",X"63",X"09",X"62",X"09",
		X"61",X"09",X"FF",X"FF",X"0C",X"0E",X"66",X"09",X"FF",X"FF",X"0D",X"0E",X"67",X"09",X"FF",X"FF",
		X"0E",X"0E",X"6A",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"11",X"0E",X"68",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"61",X"09",X"FF",X"FF",X"14",X"0E",X"6A",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",
		X"12",X"0E",X"66",X"09",X"FF",X"FF",X"13",X"0E",X"67",X"09",X"FF",X"FF",X"17",X"05",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"6E",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"18",X"0E",X"66",X"09",X"FF",X"FF",
		X"19",X"0E",X"67",X"09",X"FF",X"FF",X"1A",X"0E",X"6A",X"09",X"62",X"09",X"63",X"09",X"61",X"09",
		X"FF",X"FF",X"58",X"78",X"78",X"78",X"94",X"78",X"0B",X"02",X"6C",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"61",X"09",X"10",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"6D",X"09",X"FF",X"FF",X"11",X"06",X"60",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"61",X"09",X"0A",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",
		X"61",X"09",X"FF",X"FF",X"17",X"09",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",
		X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",
		X"D0",X"78",X"F2",X"78",X"FE",X"78",X"0A",X"79",X"16",X"79",X"22",X"79",X"2E",X"79",X"3A",X"79",
		X"46",X"79",X"52",X"79",X"5E",X"79",X"6A",X"79",X"76",X"79",X"82",X"79",X"8E",X"79",X"9A",X"79",
		X"08",X"08",X"68",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"61",X"09",X"03",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"69",X"09",
		X"FF",X"FF",X"09",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"0A",X"08",
		X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"0B",X"08",X"66",X"09",X"0E",X"FF",
		X"00",X"00",X"66",X"09",X"FF",X"FF",X"0C",X"08",X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",
		X"FF",X"FF",X"0D",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"0E",X"08",
		X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"0F",X"08",X"66",X"09",X"0E",X"FF",
		X"00",X"00",X"66",X"09",X"FF",X"FF",X"10",X"08",X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",
		X"FF",X"FF",X"11",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"12",X"08",
		X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"13",X"08",X"66",X"09",X"0E",X"FF",
		X"00",X"00",X"66",X"09",X"FF",X"FF",X"14",X"08",X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",
		X"FF",X"FF",X"15",X"08",X"66",X"09",X"0E",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"16",X"08",
		X"67",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"17",X"08",X"6A",X"09",X"62",X"09",
		X"63",X"09",X"61",X"09",X"03",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",
		X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"6B",X"09",X"FF",X"FF",X"E8",X"79",X"00",X"7A",
		X"06",X"7A",X"0C",X"7A",X"18",X"7A",X"24",X"7A",X"30",X"7A",X"3C",X"7A",X"42",X"7A",X"48",X"7A",
		X"60",X"7A",X"6C",X"7A",X"78",X"7A",X"90",X"7A",X"96",X"7A",X"9C",X"7A",X"A8",X"7A",X"B4",X"7A",
		X"C0",X"7A",X"CC",X"7A",X"D2",X"7A",X"D8",X"7A",X"05",X"08",X"60",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"69",X"09",X"FF",X"FF",
		X"06",X"11",X"66",X"09",X"FF",X"FF",X"07",X"11",X"67",X"09",X"FF",X"FF",X"08",X"11",X"66",X"09",
		X"08",X"FF",X"00",X"00",X"64",X"09",X"FF",X"FF",X"09",X"11",X"67",X"09",X"08",X"FF",X"00",X"00",
		X"66",X"09",X"FF",X"FF",X"0A",X"11",X"66",X"09",X"08",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",
		X"0B",X"11",X"65",X"09",X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"0C",X"1A",X"67",X"09",
		X"FF",X"FF",X"0D",X"1A",X"66",X"09",X"FF",X"FF",X"0E",X"05",X"68",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"0E",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",
		X"0F",X"05",X"66",X"09",X"14",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"10",X"05",X"67",X"09",
		X"14",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"11",X"05",X"66",X"09",X"0E",X"FF",X"00",X"00",
		X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"6B",X"09",X"FF",X"FF",
		X"12",X"05",X"67",X"09",X"FF",X"FF",X"13",X"05",X"66",X"09",X"FF",X"FF",X"14",X"05",X"67",X"09",
		X"08",X"FF",X"00",X"00",X"64",X"09",X"FF",X"FF",X"15",X"05",X"66",X"09",X"08",X"FF",X"00",X"00",
		X"66",X"09",X"FF",X"FF",X"16",X"05",X"67",X"09",X"08",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",
		X"17",X"05",X"65",X"09",X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"18",X"0E",X"67",X"09",
		X"FF",X"FF",X"19",X"0E",X"66",X"09",X"FF",X"FF",X"1A",X"0E",X"6A",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",
		X"FC",X"7A",X"0C",X"7B",X"1C",X"7B",X"2C",X"7B",X"3C",X"7B",X"4C",X"7B",X"08",X"18",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"6D",X"09",X"FF",X"FF",X"0B",X"02",X"6C",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"0E",X"18",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"6D",X"09",X"FF",X"FF",X"11",X"02",X"6C",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"14",X"18",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"6D",X"09",X"FF",X"FF",X"17",X"02",X"6C",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"FF",X"FF",X"7C",X"7B",X"98",X"7B",
		X"A4",X"7B",X"B0",X"7B",X"C8",X"7B",X"D4",X"7B",X"E0",X"7B",X"EC",X"7B",X"F8",X"7B",X"04",X"7C",
		X"10",X"7C",X"1C",X"7C",X"28",X"7C",X"40",X"7C",X"4C",X"7C",X"58",X"7C",X"05",X"09",X"60",X"09",
		X"62",X"09",X"63",X"09",X"62",X"09",X"61",X"09",X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",
		X"63",X"09",X"62",X"09",X"61",X"09",X"FF",X"FF",X"09",X"05",X"64",X"09",X"14",X"FF",X"00",X"00",
		X"64",X"09",X"FF",X"FF",X"0A",X"05",X"66",X"09",X"14",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",
		X"0B",X"05",X"67",X"09",X"08",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",
		X"08",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",X"0C",X"05",X"66",X"09",X"14",X"FF",X"00",X"00",
		X"66",X"09",X"FF",X"FF",X"0D",X"05",X"65",X"09",X"14",X"FF",X"00",X"00",X"65",X"09",X"FF",X"FF",
		X"0E",X"0B",X"64",X"09",X"08",X"FF",X"00",X"00",X"64",X"09",X"FF",X"FF",X"0F",X"0B",X"66",X"09",
		X"08",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"10",X"0B",X"67",X"09",X"08",X"FF",X"00",X"00",
		X"67",X"09",X"FF",X"FF",X"11",X"0B",X"65",X"09",X"08",X"FF",X"00",X"00",X"65",X"09",X"FF",X"FF",
		X"12",X"05",X"64",X"09",X"14",X"FF",X"00",X"00",X"64",X"09",X"FF",X"FF",X"13",X"05",X"66",X"09",
		X"14",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"14",X"05",X"67",X"09",X"08",X"FF",X"00",X"00",
		X"60",X"09",X"62",X"09",X"63",X"09",X"61",X"09",X"08",X"FF",X"00",X"00",X"67",X"09",X"FF",X"FF",
		X"15",X"05",X"66",X"09",X"14",X"FF",X"00",X"00",X"66",X"09",X"FF",X"FF",X"16",X"05",X"65",X"09",
		X"14",X"FF",X"00",X"00",X"65",X"09",X"FF",X"FF",X"1A",X"09",X"60",X"09",X"62",X"09",X"63",X"09",
		X"62",X"09",X"61",X"09",X"04",X"FF",X"00",X"00",X"60",X"09",X"62",X"09",X"63",X"09",X"62",X"09",
		X"61",X"09",X"FF",X"FF",X"94",X"7C",X"9E",X"7C",X"A8",X"7C",X"B2",X"7C",X"BC",X"7C",X"C0",X"7C",
		X"CB",X"7C",X"D5",X"7C",X"DF",X"7C",X"EA",X"7C",X"F4",X"7C",X"FE",X"7C",X"09",X"7D",X"13",X"7D",
		X"1D",X"7D",X"28",X"7D",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"00",X"73",X"05",X"C9",X"CD",X"32",
		X"7D",X"CD",X"CF",X"00",X"5A",X"73",X"0A",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"F6",X"73",
		X"09",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"78",X"74",X"0C",X"C9",X"CD",X"32",X"7D",X"C9",
		X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"48",X"75",X"04",X"00",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",
		X"00",X"D0",X"75",X"04",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"30",X"76",X"02",X"C9",X"CD",
		X"32",X"7D",X"CD",X"CF",X"00",X"6C",X"76",X"03",X"00",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",
		X"B2",X"76",X"0D",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"80",X"77",X"10",X"C9",X"CD",X"32",
		X"7D",X"CD",X"CF",X"00",X"52",X"78",X"03",X"00",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"B0",
		X"78",X"10",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"BC",X"79",X"16",X"C9",X"CD",X"32",X"7D",
		X"CD",X"CF",X"00",X"F0",X"7A",X"06",X"00",X"C9",X"CD",X"32",X"7D",X"CD",X"CF",X"00",X"5C",X"7B",
		X"10",X"C9",X"3E",X"09",X"CD",X"F0",X"4F",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
