library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity popeye_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of popeye_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"FF",X"00",X"1F",X"00",X"0F",X"00",X"1F",X"00",X"1F",X"00",X"3F",X"00",X"3F",X"00",
		X"3F",X"00",X"3F",X"00",X"1F",X"00",X"0F",X"00",X"0F",X"00",X"1F",X"00",X"3F",X"00",X"3F",X"00",
		X"3F",X"00",X"3F",X"00",X"7E",X"01",X"7E",X"03",X"38",X"07",X"08",X"0F",X"00",X"07",X"00",X"03",
		X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"80",X"C0",X"F0",X"F8",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"01",X"03",X"0F",X"1F",X"1F",X"3F",X"7F",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"C3",X"C7",X"CF",X"DF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"27",X"73",X"F3",X"33",X"13",X"63",X"97",X"D7",X"67",
		X"3F",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"60",
		X"60",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"80",X"C0",X"C0",X"40",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"1F",X"0F",X"03",X"01",X"01",X"01",X"01",X"07",X"07",X"07",X"01",X"01",X"04",
		X"02",X"04",X"02",X"00",X"91",X"48",X"28",X"00",X"20",X"43",X"03",X"04",X"02",X"00",X"61",X"7E",
		X"3B",X"3B",X"18",X"03",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"18",X"38",X"3C",X"1C",X"00",X"00",X"60",X"30",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"80",X"00",X"04",X"36",X"7E",X"FE",X"FC",X"7C",X"3E",X"1E",X"05",X"C0",
		X"F0",X"E0",X"F8",X"00",X"00",X"00",X"00",X"08",X"90",X"60",X"C0",X"A0",X"E0",X"E0",X"C0",X"00",
		X"04",X"86",X"00",X"00",X"00",X"00",X"1C",X"3F",X"7F",X"BF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",
		X"00",X"08",X"00",X"F0",X"E0",X"80",X"00",X"00",X"01",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"07",X"03",X"00",X"00",X"B8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"26",X"2F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"BE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"00",
		X"00",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"06",X"8F",X"DF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",X"17",X"1F",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",
		X"C0",X"E0",X"F0",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"7C",X"7C",X"7C",X"7C",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"60",X"C0",X"C0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"3E",X"FF",X"FF",X"BF",X"8F",X"6F",X"0F",X"1F",X"1F",
		X"1F",X"1F",X"3F",X"3F",X"FF",X"C3",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"1C",X"1E",X"9E",X"9E",X"CE",X"C7",X"E7",X"E3",X"F3",X"F9",X"38",X"0D",X"0E",X"03",X"00",
		X"12",X"0A",X"81",X"D0",X"C0",X"C0",X"80",X"02",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"80",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"9E",X"9E",X"DE",X"CE",X"6F",X"E7",X"E3",X"F1",X"F8",X"FD",X"FE",X"8F",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"3F",X"3F",X"1F",X"1F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"70",X"70",X"78",X"38",X"38",X"38",X"38",X"38",X"78",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"03",X"06",X"04",X"01",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"60",X"38",X"0E",X"07",X"0F",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"07",X"03",X"00",X"00",X"00",
		X"00",X"0E",X"3C",X"78",X"F0",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"38",
		X"00",X"00",X"80",X"40",X"C0",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"EF",X"EE",X"C7",X"87",X"83",X"01",X"83",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"87",X"C7",X"8F",X"0D",X"09",X"08",X"98",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"FE",X"FE",X"06",X"06",X"FE",X"FE",
		X"00",X"00",X"06",X"06",X"00",X"00",X"0C",X"18",X"38",X"30",X"70",X"70",X"60",X"60",X"00",X"00",
		X"00",X"00",X"CF",X"CF",X"C3",X"C3",X"C3",X"CF",X"CF",X"C3",X"C3",X"C3",X"CF",X"CF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FC",X"FA",X"FA",X"FA",X"F6",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"1C",
		X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",
		X"00",X"00",X"FE",X"FE",X"FE",X"1E",X"1E",X"FE",X"FE",X"FE",X"1E",X"1E",X"FE",X"FE",X"FE",X"00",
		X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"1E",X"FE",X"FE",X"FE",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",
		X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"1E",X"FE",X"FE",X"1E",X"1E",X"1E",X"1E",X"FE",X"FE",X"00",
		X"00",X"00",X"33",X"33",X"30",X"30",X"30",X"F0",X"F0",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"33",X"33",X"33",X"33",X"3F",X"3F",X"3F",X"33",X"33",X"33",X"33",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"F8",X"F0",X"C0",X"C0",X"B8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"3C",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"8C",X"CC",X"E4",X"F6",X"F7",X"F7",X"FE",X"7C",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"DE",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"98",X"00",X"00",X"98",X"98",X"98",X"98",X"98",X"98",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"FE",X"FD",X"FD",X"FD",X"FB",
		X"FE",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"20",X"F0",X"90",X"B0",X"D0",X"90",X"F0",X"F4",X"F8",X"00",X"08",X"50",X"20",X"00",
		X"F0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FB",X"F3",X"E3",X"66",X"BC",X"C8",X"60",X"E0",X"F0",X"C0",
		X"0C",X"FE",X"FF",X"FD",X"FF",X"FC",X"E4",X"E4",X"BC",X"1C",X"38",X"70",X"E0",X"C0",X"80",X"00",
		X"F0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FB",X"F3",X"E3",X"C6",X"CC",X"58",X"70",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"F0",X"FE",X"FF",X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"3E",X"3E",X"1F",X"1F",X"3F",X"1F",X"1F",X"1F",X"1F",X"2F",X"7F",X"EF",X"F7",X"FF",X"F7",
		X"F7",X"EF",X"EF",X"FF",X"EE",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"60",X"60",X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"FE",X"FF",X"F0",X"FE",
		X"FF",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"F3",
		X"E1",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"FF",X"F0",X"FC",
		X"FE",X"FF",X"0F",X"03",X"00",X"00",X"00",X"80",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",
		X"DF",X"EF",X"8F",X"87",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"20",X"40",X"80",X"C0",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"01",
		X"03",X"AF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"0F",X"1F",X"1F",X"1F",X"17",X"03",
		X"03",X"03",X"07",X"07",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"C0",X"E0",X"F8",
		X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"73",X"03",X"07",X"07",X"0F",X"1F",X"1F",X"0F",X"03",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"07",X"1F",X"3F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"4F",X"67",X"F3",X"33",X"13",X"03",X"63",X"B7",X"D7",X"67",
		X"04",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B8",X"5C",X"4C",X"24",X"20",X"40",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"07",X"FE",X"FE",X"FC",
		X"00",X"00",X"F8",X"80",X"04",X"2C",X"EC",X"EC",X"E8",X"E4",X"8C",X"6C",X"EC",X"EC",X"E8",X"E4",
		X"8C",X"6C",X"EC",X"EC",X"E8",X"E0",X"00",X"00",X"10",X"10",X"10",X"30",X"60",X"C0",X"80",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"00",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7E",
		X"FC",X"7C",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"78",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"03",X"03",X"03",X"07",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"7E",X"4F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DE",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"E0",X"DF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"48",X"48",X"88",X"88",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"20",X"00",X"40",X"83",X"0F",X"1E",X"3C",X"BC",X"F8",X"FF",X"E7",X"CB",X"F5",X"7A",X"3C",X"76",
		X"03",X"43",X"A3",X"EA",X"CD",X"09",X"19",X"FB",X"FF",X"FF",X"FF",X"FF",X"7F",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"7E",
		X"F3",X"FB",X"FF",X"FE",X"FE",X"FC",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"80",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"90",
		X"F8",X"BD",X"BF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"F3",X"F2",X"FD",X"FD",X"FD",X"3B",X"27",X"DF",X"EF",X"DF",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FB",X"FB",X"FB",X"FB",X"7B",X"8F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",
		X"07",X"07",X"07",X"07",X"07",X"4F",X"8F",X"8F",X"CF",X"5F",X"7F",X"7F",X"7F",X"FF",X"DF",X"C7",
		X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"01",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"FF",X"FF",X"FB",X"F7",X"7F",X"EF",X"DF",X"BF",X"7F",X"7F",
		X"78",X"70",X"E0",X"E9",X"FE",X"C6",X"B3",X"B9",X"9C",X"EE",X"F7",X"FB",X"9C",X"0C",X"8F",X"5F",
		X"82",X"A4",X"C8",X"10",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"C0",X"00",X"00",X"40",X"80",X"00",X"01",X"11",X"39",
		X"F9",X"3F",X"03",X"00",X"00",X"24",X"1F",X"9F",X"F1",X"75",X"65",X"69",X"CB",X"13",X"66",X"0C",
		X"34",X"00",X"03",X"02",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"FF",X"FF",X"FF",X"DF",X"BF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"EF",X"CD",X"8D",X"07",X"07",X"03",X"07",X"06",X"03",X"03",X"03",X"01",X"00",X"03",X"06",
		X"0F",X"0F",X"0F",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"07",X"01",X"03",X"03",X"0F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0E",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"3E",X"3F",X"3F",X"3F",X"3F",X"1F",X"1E",X"1E",X"1F",X"0F",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"FC",X"7C",X"BA",X"B1",X"B2",X"30",X"71",X"70",X"D2",X"85",X"02",X"01",X"01",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",
		X"40",X"80",X"C0",X"C0",X"C0",X"C0",X"40",X"80",X"C0",X"C0",X"C0",X"40",X"00",X"80",X"00",X"00",
		X"62",X"7F",X"FF",X"FF",X"E7",X"E7",X"FF",X"E0",X"80",X"0F",X"5F",X"DF",X"DF",X"DF",X"C0",X"1F",
		X"DF",X"DF",X"DF",X"DF",X"C0",X"1F",X"DF",X"DF",X"DF",X"DF",X"C0",X"00",X"1F",X"3F",X"00",X"00",
		X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",
		X"C0",X"C0",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"DF",
		X"6F",X"70",X"FD",X"FE",X"BE",X"BF",X"9F",X"9F",X"8F",X"87",X"83",X"81",X"82",X"81",X"C3",X"CF",
		X"C7",X"EF",X"E7",X"77",X"16",X"1C",X"01",X"02",X"0E",X"0C",X"0C",X"06",X"07",X"03",X"01",X"00",
		X"1F",X"3F",X"37",X"33",X"1E",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"98",X"88",X"41",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"23",X"40",X"E4",X"F8",
		X"07",X"07",X"0B",X"0B",X"1B",X"1D",X"1E",X"1F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"80",X"80",X"40",X"30",X"40",X"80",X"00",
		X"F8",X"7C",X"3E",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"C0",X"88",
		X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"80",X"80",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"FB",X"FB",X"FD",X"0E",
		X"03",X"03",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",
		X"2F",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"78",X"B8",X"B0",X"F0",X"E0",
		X"C0",X"C0",X"D2",X"FC",X"FF",X"80",X"85",X"F1",X"3D",X"1E",X"3B",X"81",X"A1",X"51",X"75",X"66",
		X"04",X"8C",X"FE",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"07",X"07",X"07",X"05",X"24",X"2C",X"28",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"FE",X"F8",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FE",X"FE",X"FF",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",
		X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"F7",X"F7",X"CF",X"3F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"3E",X"BE",X"BE",X"38",X"F8",X"24",X"60",X"30",X"18",X"0C",X"1C",X"18",X"38",X"F0",X"E0",X"90",
		X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"FC",X"FC",X"FC",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F9",X"C7",X"3F",X"FF",X"FF",X"FF",X"7F",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"7C",X"7F",X"77",X"77",X"77",X"37",X"37",X"17",X"0F",X"0F",X"02",X"03",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"1B",X"99",X"CF",X"E1",X"F3",X"FF",X"FF",X"F7",X"CF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"7F",X"BF",X"9F",X"7F",X"07",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",
		X"07",X"0F",X"FF",X"FE",X"FE",X"FC",X"F8",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"BF",X"9F",X"79",X"83",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"93",X"21",X"00",X"00",X"80",X"80",X"C0",X"E3",X"FF",X"FF",X"FF",
		X"38",X"3C",X"78",X"D9",X"8B",X"09",X"28",X"18",X"1C",X"4C",X"CC",X"8C",X"5C",X"F8",X"F0",X"00",
		X"0F",X"07",X"03",X"03",X"01",X"01",X"C2",X"23",X"03",X"87",X"C7",X"2E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"DC",X"FC",X"FC",X"FC",X"F8",X"F0",X"F3",X"E7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"E0",X"E0",
		X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"01",X"00",X"00",X"03",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"03",X"21",X"40",X"E4",X"F8",
		X"1C",X"3E",X"7C",X"D9",X"8B",X"09",X"28",X"18",X"9C",X"CC",X"8C",X"0C",X"5C",X"F8",X"F0",X"80",
		X"01",X"07",X"1F",X"7F",X"FF",X"FD",X"F9",X"71",X"31",X"E1",X"01",X"01",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"1E",X"1E",X"1F",X"1F",X"0F",X"37",X"3F",X"1E",X"1E",X"0F",X"0F",X"0F",X"07",X"07",
		X"03",X"33",X"4B",X"0F",X"17",X"25",X"0A",X"13",X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"D8",X"D8",X"DC",X"5C",X"7C",X"7C",X"78",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"F0",X"F9",X"FB",X"FB",X"FB",X"FF",X"FF",X"7F",X"7E",X"7E",X"7E",X"7C",X"3C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"F0",X"FC",X"FE",X"0E",X"FC",X"F0",X"FE",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"D0",X"F8",
		X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"04",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"0F",X"0F",X"0F",X"3F",X"3F",
		X"1F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"A0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"08",X"0C",X"5C",X"7F",X"3F",X"0F",X"03",X"03",X"01",X"01",X"18",X"18",X"10",X"88",
		X"3C",X"22",X"02",X"22",X"62",X"86",X"10",X"41",X"C0",X"E0",X"C0",X"E0",X"E0",X"10",X"00",X"00",
		X"E0",X"F0",X"30",X"30",X"F0",X"E0",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"8E",X"07",X"07",X"00",X"80",X"FE",X"FE",X"BE",X"BF",
		X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",X"F8",X"70",X"00",X"00",
		X"82",X"C0",X"60",X"60",X"20",X"10",X"80",X"80",X"22",X"23",X"47",X"0E",X"1E",X"FE",X"DE",X"8C",
		X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",X"03",X"1F",X"3F",X"3F",X"7F",X"FA",X"F8",X"70",X"20",
		X"00",X"00",X"00",X"20",X"30",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"20",X"30",X"10",X"18",X"18",
		X"00",X"00",X"00",X"10",X"18",X"0C",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",
		X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",
		X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"07",X"01",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"03",
		X"C7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",
		X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"E7",X"F7",X"7E",X"7E",X"3E",X"3C",X"1C",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",
		X"80",X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"CF",X"C3",X"41",X"40",X"40",X"40",X"40",X"C1",
		X"40",X"40",X"C0",X"F0",X"F0",X"C0",X"C0",X"E0",X"70",X"30",X"30",X"B0",X"B0",X"E0",X"C0",X"80",
		X"80",X"C0",X"E0",X"B0",X"B0",X"30",X"30",X"B0",X"B0",X"E0",X"C0",X"80",X"80",X"C0",X"E0",X"B0",
		X"00",X"00",X"01",X"03",X"07",X"07",X"8F",X"CF",X"DE",X"FE",X"FC",X"7F",X"7F",X"3C",X"30",X"00",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"B8",X"70",X"E0",
		X"FF",X"FF",X"FE",X"FC",X"FE",X"FC",X"FE",X"FF",X"FF",X"2E",X"63",X"30",X"84",X"86",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"70",X"38",X"F8",X"F0",X"C0",X"00",X"00",X"00",
		X"01",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"07",X"1F",X"1F",X"1F",X"0C",X"0C",X"02",X"00",
		X"31",X"70",X"F9",X"F9",X"9B",X"1B",X"1B",X"1B",X"1F",X"1F",X"1F",X"1F",X"0C",X"0C",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"70",X"38",X"F8",X"F0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"70",X"F9",X"F9",X"DB",X"DB",X"DB",X"DB",X"DF",X"DF",X"5F",X"1F",X"0C",X"0C",X"02",X"00",
		X"00",X"41",X"2B",X"13",X"43",X"41",X"81",X"50",X"21",X"83",X"C3",X"7F",X"3C",X"00",X"00",X"00",
		X"F8",X"1C",X"1D",X"0F",X"0F",X"87",X"03",X"0C",X"4D",X"1F",X"BF",X"3F",X"37",X"BD",X"1C",X"08",
		X"1C",X"0E",X"07",X"0F",X"07",X"07",X"0E",X"9E",X"FC",X"FE",X"FE",X"CC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"38",X"4C",X"76",X"B6",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B6",X"76",X"76",X"74",
		X"6C",X"68",X"58",X"50",X"A0",X"40",X"00",X"C0",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"03",X"47",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"00",X"80",X"C0",X"F0",X"E0",X"C0",X"84",X"10",X"10",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"03",X"07",X"0F",
		X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"EF",X"8F",X"07",X"07",
		X"03",X"03",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"0F",
		X"38",X"70",X"F0",X"E3",X"E7",X"C5",X"87",X"07",X"06",X"08",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"C0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"0E",X"0E",X"11",X"00",X"00",X"14",X"14",X"21",X"00",X"01",X"03",X"01",X"00",
		X"FE",X"A7",X"03",X"47",X"3F",X"3F",X"1F",X"19",X"83",X"06",X"2C",X"4C",X"8D",X"2F",X"07",X"02",
		X"00",X"00",X"18",X"BC",X"FC",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"00",
		X"E0",X"F0",X"F0",X"00",X"00",X"FC",X"FC",X"F8",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"C0",
		X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"F0",X"F0",X"F0",X"30",X"38",X"18",X"18",X"18",X"3C",X"33",X"07",X"1F",X"3F",X"7F",X"3F",
		X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",
		X"00",X"0D",X"9F",X"CF",X"84",X"A0",X"90",X"08",X"12",X"0B",X"07",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"06",X"06",X"09",X"00",X"0A",X"0A",X"08",X"11",X"00",X"07",X"0F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0B",X"09",X"06",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"83",X"CF",X"DF",X"9F",X"3F",
		X"7F",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"01",X"00",X"F0",X"7E",X"3F",X"F3",X"03",X"07",X"07",X"0E",X"1F",X"07",X"07",
		X"7F",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"07",X"07",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"10",X"70",X"7C",X"6F",X"76",X"31",X"3B",X"2A",X"00",
		X"22",X"21",X"65",X"26",X"24",X"14",X"04",X"0B",X"10",X"01",X"00",X"07",X"0F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"80",X"D0",X"F0",X"E0",X"E0",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"06",
		X"18",X"30",X"36",X"66",X"E9",X"C0",X"83",X"08",X"10",X"01",X"00",X"07",X"0F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"0E",X"07",X"0F",X"07",X"07",X"0E",X"9E",X"FC",X"FE",X"FE",X"CC",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",
		X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"F4",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",
		X"00",X"F0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"DC",X"C0",X"80",X"00",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"1C",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"FF",X"03",X"06",X"06",X"08",X"18",X"18",X"20",X"20",X"60",X"80",X"C0",X"E0",X"C0",X"80",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"F8",X"8C",X"06",X"02",X"02",X"06",X"8C",X"F8",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"8C",X"06",X"02",X"02",X"06",X"8C",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"80",X"84",X"8C",X"8C",X"C4",X"C0",X"E2",X"FE",X"FC",X"FC",X"FC",
		X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"1F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"C0",X"C0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",
		X"F8",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1E",X"BF",X"FF",X"DF",X"FE",X"FE",X"FC",X"F8",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"20",X"20",
		X"A8",X"70",X"00",X"00",X"00",X"00",X"00",X"50",X"28",X"28",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",X"0F",X"07",X"07",X"0F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"F0",X"F0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"9F",X"3F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"9F",X"9F",X"8F",X"87",X"C3",X"47",X"02",X"00",X"00",
		X"00",X"70",X"70",X"F8",X"FA",X"12",X"84",X"20",X"20",X"40",X"21",X"2B",X"1F",X"0F",X"0C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"70",X"38",X"38",X"1C",X"0E",X"0E",X"3E",X"FC",
		X"F0",X"60",X"40",X"00",X"02",X"01",X"83",X"87",X"87",X"83",X"C3",X"77",X"7E",X"FE",X"5C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"87",X"C7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"F0",X"1C",X"1E",X"0E",
		X"0E",X"07",X"07",X"C7",X"E3",X"E2",X"C0",X"18",X"3F",X"3E",X"7E",X"7F",X"3F",X"39",X"78",X"F0",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"06",X"02",X"06",X"0E",X"0E",X"0E",
		X"0E",X"7C",X"FC",X"FC",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"3C",X"79",X"79",X"F3",X"E7",X"CF",X"9F",X"9F",X"1F",
		X"3F",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"78",X"3C",X"0C",X"86",X"C3",X"71",X"0D",X"1E",X"3E",
		X"3E",X"3F",X"1E",X"1E",X"3F",X"FF",X"F1",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"82",X"D0",X"50",X"12",X"00",X"00",X"A0",X"26",X"7E",X"FF",X"FE",X"7C",
		X"00",X"00",X"80",X"80",X"A0",X"A0",X"C0",X"C0",X"02",X"02",X"0A",X"07",X"02",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"40",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"3F",X"3F",X"7F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"9F",X"8F",X"87",X"C3",X"CC",X"D0",X"F0",X"C1",X"0C",X"12",X"21",X"21",
		X"20",X"19",X"25",X"47",X"84",X"C2",X"80",X"01",X"01",X"23",X"27",X"7C",X"94",X"14",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"FE",X"FE",X"FC",X"F8",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"01",X"00",X"43",X"60",X"A3",X"00",X"02",X"00",X"00",X"C0",
		X"F3",X"DF",X"AF",X"EF",X"DF",X"9F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"05",X"02",X"0A",
		X"12",X"E4",X"48",X"A0",X"70",X"40",X"24",X"18",X"03",X"07",X"1B",X"03",X"03",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"F8",X"80",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"08",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"14",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"0E",X"15",X"84",
		X"84",X"84",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"C7",X"8F",X"9F",X"BF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"D8",X"08",X"08",X"18",X"19",X"1F",X"1F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"01",X"03",X"33",X"4E",X"04",X"87",X"80",X"9F",
		X"1C",X"1A",X"8A",X"1F",X"3F",X"7F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"82",X"0A",X"04",X"84",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"1F",X"3F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"0F",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",
		X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"03",X"00",X"01",X"01",X"01",X"08",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",X"A0",X"A0",X"A0",X"A0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"39",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"B8",X"00",X"00",X"03",X"01",X"09",X"0C",X"0C",X"1C",X"1C",X"1E",
		X"1E",X"3C",X"3C",X"3F",X"3F",X"BF",X"3F",X"3F",X"9F",X"0F",X"03",X"00",X"01",X"01",X"01",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"CE",X"1E",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",
		X"0F",X"0E",X"01",X"07",X"0F",X"03",X"03",X"37",X"67",X"53",X"13",X"0B",X"03",X"03",X"03",X"07",
		X"07",X"67",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"01",X"01",X"01",X"08",
		X"14",X"04",X"04",X"08",X"40",X"41",X"43",X"43",X"43",X"E3",X"E3",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"C0",X"C0",X"80",X"80",X"00",X"80",X"80",
		X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"08",X"10",X"08",X"0A",X"34",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"EE",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"7F",X"7F",X"39",X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"01",
		X"01",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"01",X"B9",
		X"3F",X"3F",X"3F",X"37",X"33",X"31",X"38",X"18",X"0C",X"02",X"00",X"00",X"00",X"01",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"1B",X"DE",X"F6",X"FC",X"FC",X"FC",
		X"7C",X"18",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"3C",X"FC",X"FC",X"FC",X"FE",X"BF",X"1F",X"1F",X"0F",X"0F",X"07",X"03",
		X"03",X"03",X"03",X"07",X"03",X"01",X"00",X"40",X"03",X"06",X"05",X"08",X"1C",X"1E",X"3F",X"FF",
		X"7F",X"7F",X"7F",X"7F",X"77",X"73",X"31",X"38",X"18",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"D0",X"B0",X"E0",X"E0",X"E0",X"80",X"C0",X"80",X"C0",
		X"C0",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"10",X"10",
		X"10",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"EF",X"8F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",
		X"03",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"BF",
		X"FF",X"FF",X"FF",X"F7",X"F3",X"31",X"38",X"18",X"0C",X"02",X"00",X"00",X"00",X"01",X"03",X"03",
		X"02",X"3C",X"44",X"89",X"81",X"81",X"80",X"80",X"80",X"C0",X"C1",X"00",X"18",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"14",X"34",X"3C",X"A8",X"F8",X"F8",X"F0",X"F0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"60",X"20",X"10",X"10",X"00",X"00",
		X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"7F",X"7F",X"6F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"FC",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",
		X"07",X"03",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"3F",X"BF",
		X"7F",X"7F",X"7F",X"7F",X"77",X"73",X"31",X"38",X"18",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"0F",X"07",X"06",X"06",X"0E",X"0E",X"1F",X"1F",X"1F",X"1F",X"3F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",
		X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3E",X"FE",X"FF",X"EF",X"FF",
		X"DF",X"0F",X"03",X"03",X"07",X"03",X"02",X"02",X"06",X"06",X"0F",X"0F",X"0F",X"1F",X"1F",X"7F",
		X"7F",X"3F",X"7F",X"7F",X"7F",X"77",X"73",X"31",X"38",X"18",X"0C",X"02",X"00",X"00",X"00",X"00",
		X"41",X"02",X"3C",X"44",X"89",X"80",X"81",X"80",X"80",X"80",X"C0",X"C1",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
