library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_graphx_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_graphx_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"68",X"78",X"5A",X"87",X"0D",X"A2",X"2A",X"22",X"66",X"66",X"EE",X"EE",X"66",X"66",X"66",
		X"F0",X"E0",X"3C",X"28",X"0F",X"69",X"E1",X"F0",X"C3",X"87",X"00",X"FF",X"FF",X"00",X"96",X"00",
		X"C1",X"2D",X"C3",X"0B",X"1E",X"D2",X"A1",X"2D",X"69",X"0F",X"00",X"FF",X"FF",X"00",X"78",X"00",
		X"F0",X"F0",X"C1",X"B0",X"2D",X"0B",X"45",X"45",X"44",X"66",X"66",X"77",X"77",X"66",X"66",X"66",
		X"F0",X"F0",X"34",X"F0",X"F0",X"E0",X"F0",X"34",X"F0",X"78",X"B0",X"F0",X"92",X"34",X"F0",X"F0",
		X"F0",X"F0",X"16",X"F0",X"F0",X"D0",X"F0",X"92",X"F0",X"E0",X"F0",X"92",X"F0",X"F0",X"34",X"F0",
		X"78",X"F0",X"78",X"F0",X"92",X"34",X"D0",X"F0",X"F0",X"F0",X"92",X"C1",X"F0",X"F0",X"F0",X"F0",
		X"D0",X"F0",X"E0",X"34",X"92",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"92",X"F0",X"E0",X"F0",X"F0",
		X"03",X"90",X"08",X"87",X"41",X"0F",X"0B",X"2D",X"07",X"02",X"08",X"41",X"09",X"0D",X"0F",X"0A",
		X"0E",X"0A",X"01",X"00",X"0C",X"0C",X"0F",X"43",X"94",X"0B",X"03",X"A1",X"07",X"03",X"28",X"05",
		X"07",X"0F",X"C2",X"07",X"03",X"04",X"02",X"41",X"02",X"01",X"09",X"08",X"0E",X"43",X"0E",X"09",
		X"0B",X"03",X"00",X"10",X"08",X"48",X"02",X"0F",X"09",X"03",X"25",X"4B",X"09",X"09",X"08",X"0E",
		X"83",X"07",X"0F",X"07",X"83",X"0F",X"0F",X"2C",X"41",X"41",X"29",X"29",X"0F",X"07",X"03",X"01",
		X"07",X"70",X"0F",X"1C",X"49",X"83",X"41",X"20",X"0F",X"07",X"0D",X"07",X"02",X"03",X"02",X"00",
		X"1C",X"0F",X"83",X"0F",X"0B",X"0A",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"02",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"EF",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"BF",X"FF",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"CF",X"FF",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"3F",X"FF",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0F",X"8F",X"AD",X"AD",X"0F",X"5E",X"2D",X"8F",X"4F",X"DE",X"9E",X"AF",X"8F",X"5E",X"8F",X"4B",
		X"3F",X"6F",X"5F",X"2F",X"BF",X"2F",X"BF",X"1F",X"2F",X"5F",X"AF",X"6F",X"BF",X"5F",X"AF",X"1F",
		X"0F",X"2F",X"2F",X"0F",X"0F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",X"4F",X"0F",X"0F",
		X"0F",X"1F",X"2F",X"1F",X"0F",X"0F",X"0F",X"1F",X"1F",X"4F",X"0F",X"0F",X"2F",X"0F",X"0F",X"2F",
		X"1E",X"3C",X"96",X"5A",X"38",X"34",X"1E",X"3C",X"34",X"1E",X"50",X"F0",X"3C",X"D2",X"34",X"F0",
		X"DF",X"AF",X"4F",X"CF",X"8F",X"8F",X"5E",X"8E",X"0F",X"0D",X"4B",X"2D",X"50",X"F0",X"F0",X"D0",
		X"8F",X"1F",X"2F",X"2F",X"0F",X"4F",X"0F",X"AF",X"BF",X"EF",X"1E",X"0F",X"D2",X"A0",X"F0",X"F0",
		X"0F",X"4F",X"8F",X"9F",X"4F",X"CF",X"2F",X"CF",X"EF",X"3F",X"4F",X"CF",X"0F",X"0F",X"58",X"F0",
		X"0F",X"4A",X"0C",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A5",X"4B",X"0D",X"87",X"07",X"0B",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"5A",X"4B",X"0F",X"09",X"86",X"0F",X"0B",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1C",X"29",X"1C",X"4B",X"A5",X"1A",X"06",X"04",X"0F",X"0F",X"07",X"0E",X"0C",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"EF",X"DF",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"BF",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"FF",X"CF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"3F",
		X"4F",X"2F",X"0F",X"0F",X"2F",X"2F",X"9F",X"1F",X"2F",X"0F",X"0F",X"0F",X"4F",X"2F",X"0F",X"8F",
		X"0F",X"1F",X"8F",X"0F",X"9F",X"0F",X"0F",X"8F",X"0F",X"AF",X"0F",X"1F",X"8F",X"4F",X"0F",X"1F",
		X"0F",X"9F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"0F",X"0F",X"0F",X"4F",X"8F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"87",X"97",X"0F",X"4B",X"A7",X"87",X"0F",X"0F",X"A7",X"0F",
		X"4F",X"8F",X"0F",X"2F",X"8F",X"5F",X"1F",X"8F",X"4F",X"2F",X"1F",X"0F",X"0F",X"1F",X"0F",X"C1",
		X"0F",X"CF",X"1F",X"2F",X"CF",X"0F",X"BF",X"1F",X"1F",X"2F",X"0F",X"0F",X"0F",X"60",X"06",X"F0",
		X"0F",X"0F",X"1F",X"0F",X"4F",X"1F",X"0F",X"3F",X"2F",X"0B",X"07",X"07",X"0B",X"C1",X"F0",X"F0",
		X"87",X"85",X"87",X"B7",X"07",X"D3",X"43",X"C3",X"A1",X"C2",X"C1",X"F0",X"E0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"1F",X"8F",X"0F",X"0F",X"0F",X"4F",X"4F",X"1F",X"AF",X"6F",X"FF",X"1F",X"2D",X"B0",
		X"CF",X"0F",X"8F",X"0F",X"0F",X"0F",X"8F",X"8F",X"2F",X"4F",X"FF",X"4F",X"87",X"0A",X"61",X"F0",
		X"0F",X"0F",X"4F",X"8F",X"0F",X"4F",X"0F",X"4F",X"8F",X"3F",X"5F",X"BF",X"9F",X"1C",X"0D",X"E0",
		X"0F",X"0F",X"4F",X"0F",X"0F",X"2F",X"1F",X"8F",X"0F",X"2F",X"1F",X"6F",X"BF",X"4F",X"8F",X"94",
		X"0F",X"0F",X"0F",X"2F",X"0F",X"8F",X"0F",X"0F",X"1F",X"0F",X"4F",X"8F",X"1F",X"4F",X"4F",X"0F",
		X"2F",X"8F",X"1F",X"2F",X"0F",X"0F",X"0F",X"1F",X"4F",X"AF",X"2F",X"8F",X"4F",X"2F",X"4F",X"1F",
		X"0F",X"4F",X"4F",X"0F",X"1F",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"8F",X"1F",X"0F",
		X"0F",X"2F",X"4F",X"2F",X"0F",X"1F",X"0F",X"2F",X"2F",X"8F",X"0F",X"0F",X"4F",X"0F",X"0F",X"4F",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0C",X"08",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0D",X"0F",X"0F",X"0D",X"05",X"03",X"0E",X"0E",X"09",X"0B",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"07",X"0F",X"0F",X"0E",X"0D",X"09",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"01",X"07",X"02",X"03",X"07",X"03",X"01",X"00",X"00",X"00",
		X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"EE",X"EE",X"66",X"66",X"22",X"2A",X"A2",X"0D",X"87",X"5A",X"78",X"68",X"F0",
		X"00",X"96",X"00",X"FF",X"FF",X"00",X"87",X"C3",X"F0",X"E1",X"69",X"0F",X"28",X"3C",X"E0",X"F0",
		X"00",X"78",X"00",X"FF",X"FF",X"00",X"0F",X"69",X"2D",X"A1",X"D2",X"1E",X"0B",X"C3",X"2D",X"C1",
		X"66",X"66",X"66",X"77",X"77",X"66",X"66",X"44",X"45",X"45",X"0B",X"2D",X"B0",X"C1",X"F0",X"F0",
		X"F0",X"F0",X"34",X"92",X"F0",X"B0",X"78",X"F0",X"34",X"F0",X"E0",X"F0",X"F0",X"34",X"F0",X"F0",
		X"F0",X"34",X"F0",X"F0",X"92",X"F0",X"E0",X"F0",X"92",X"F0",X"D0",X"F0",X"F0",X"16",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"C1",X"92",X"F0",X"F0",X"F0",X"D0",X"34",X"92",X"F0",X"78",X"F0",X"78",
		X"F0",X"F0",X"E0",X"F0",X"92",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"92",X"34",X"E0",X"F0",X"D0",
		X"0A",X"0F",X"0D",X"09",X"41",X"08",X"02",X"07",X"2D",X"0B",X"0F",X"41",X"87",X"08",X"90",X"03",
		X"05",X"28",X"03",X"07",X"A1",X"03",X"0B",X"94",X"43",X"0F",X"0C",X"0C",X"00",X"01",X"0A",X"0E",
		X"09",X"0E",X"43",X"0E",X"08",X"09",X"01",X"02",X"41",X"02",X"04",X"03",X"07",X"C2",X"0F",X"07",
		X"0E",X"08",X"09",X"09",X"4B",X"25",X"03",X"09",X"0F",X"02",X"48",X"08",X"10",X"00",X"03",X"0B",
		X"01",X"03",X"07",X"0F",X"29",X"29",X"41",X"41",X"2C",X"0F",X"0F",X"83",X"07",X"0F",X"07",X"83",
		X"00",X"02",X"03",X"02",X"07",X"0D",X"07",X"0F",X"20",X"41",X"83",X"49",X"1C",X"0F",X"70",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"0A",X"0B",X"0F",X"83",X"0F",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"02",X"07",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"EF",X"DF",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"BF",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"FF",X"CF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"3F",
		X"4B",X"8F",X"5E",X"8F",X"AF",X"9E",X"DE",X"4F",X"8F",X"2D",X"5E",X"0F",X"AD",X"AD",X"8F",X"0F",
		X"1F",X"AF",X"5F",X"BF",X"6F",X"AF",X"5F",X"2F",X"1F",X"BF",X"2F",X"BF",X"2F",X"5F",X"6F",X"3F",
		X"0F",X"0F",X"4F",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"0F",X"0F",X"2F",X"2F",X"0F",
		X"2F",X"0F",X"0F",X"2F",X"0F",X"0F",X"4F",X"1F",X"1F",X"0F",X"0F",X"0F",X"1F",X"2F",X"1F",X"0F",
		X"F0",X"34",X"D2",X"3C",X"F0",X"50",X"1E",X"34",X"3C",X"1E",X"34",X"38",X"5A",X"96",X"3C",X"1E",
		X"D0",X"F0",X"F0",X"50",X"2D",X"4B",X"0D",X"0F",X"8E",X"5E",X"8F",X"8F",X"CF",X"4F",X"AF",X"DF",
		X"F0",X"F0",X"A0",X"D2",X"0F",X"1E",X"EF",X"BF",X"AF",X"0F",X"4F",X"0F",X"2F",X"2F",X"1F",X"8F",
		X"F0",X"58",X"0F",X"0F",X"CF",X"4F",X"3F",X"EF",X"CF",X"2F",X"CF",X"4F",X"9F",X"8F",X"4F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"0C",X"4A",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0B",X"07",X"87",X"0D",X"4B",X"A5",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"0B",X"0F",X"86",X"09",X"0F",X"4B",X"5A",X"0F",
		X"00",X"00",X"0C",X"0E",X"07",X"0F",X"0F",X"04",X"06",X"1A",X"A5",X"4B",X"1C",X"29",X"1C",X"0F",
		X"DF",X"EF",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"BF",X"FF",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"CF",X"FF",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"3F",X"FF",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"8F",X"0F",X"2F",X"4F",X"0F",X"0F",X"0F",X"2F",X"1F",X"9F",X"2F",X"2F",X"0F",X"0F",X"2F",X"4F",
		X"1F",X"0F",X"4F",X"8F",X"1F",X"0F",X"AF",X"0F",X"8F",X"0F",X"0F",X"9F",X"0F",X"8F",X"1F",X"0F",
		X"0F",X"8F",X"4F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",X"9F",X"0F",
		X"0F",X"A7",X"0F",X"0F",X"87",X"A7",X"4B",X"0F",X"97",X"87",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"C1",X"0F",X"1F",X"0F",X"0F",X"1F",X"2F",X"4F",X"8F",X"1F",X"5F",X"8F",X"2F",X"0F",X"8F",X"4F",
		X"F0",X"06",X"60",X"0F",X"0F",X"0F",X"2F",X"1F",X"1F",X"BF",X"0F",X"CF",X"2F",X"1F",X"CF",X"0F",
		X"F0",X"F0",X"C1",X"0B",X"07",X"07",X"0B",X"2F",X"3F",X"0F",X"1F",X"4F",X"0F",X"1F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"E0",X"F0",X"C1",X"C2",X"A1",X"C3",X"43",X"D3",X"07",X"B7",X"87",X"85",X"87",
		X"B0",X"2D",X"1F",X"FF",X"6F",X"AF",X"1F",X"4F",X"4F",X"0F",X"0F",X"0F",X"8F",X"1F",X"0F",X"0F",
		X"F0",X"61",X"0A",X"87",X"4F",X"FF",X"4F",X"2F",X"8F",X"8F",X"0F",X"0F",X"0F",X"8F",X"0F",X"CF",
		X"E0",X"0D",X"1C",X"9F",X"BF",X"5F",X"3F",X"8F",X"4F",X"0F",X"4F",X"0F",X"8F",X"4F",X"0F",X"0F",
		X"94",X"8F",X"4F",X"BF",X"6F",X"1F",X"2F",X"0F",X"8F",X"1F",X"2F",X"0F",X"0F",X"4F",X"0F",X"0F",
		X"0F",X"4F",X"4F",X"1F",X"8F",X"4F",X"0F",X"1F",X"0F",X"0F",X"8F",X"0F",X"2F",X"0F",X"0F",X"0F",
		X"1F",X"4F",X"2F",X"4F",X"8F",X"2F",X"AF",X"4F",X"1F",X"0F",X"0F",X"0F",X"2F",X"1F",X"8F",X"2F",
		X"0F",X"1F",X"8F",X"0F",X"4F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",X"1F",X"0F",X"4F",X"4F",X"0F",
		X"4F",X"0F",X"0F",X"4F",X"0F",X"0F",X"8F",X"2F",X"2F",X"0F",X"1F",X"0F",X"2F",X"4F",X"2F",X"0F",
		X"00",X"00",X"00",X"00",X"0C",X"08",X"00",X"08",X"0C",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0B",X"09",X"0E",X"0E",X"03",X"05",X"0D",X"0F",X"0F",X"0D",X"04",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"09",X"0D",X"0E",X"0F",X"0F",X"07",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"03",X"02",X"07",X"01",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
