library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_spr_bit3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_spr_bit3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"C0",X"D0",X"CC",X"C1",X"47",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"07",X"47",X"C1",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"3E",X"3E",X"3F",X"3F",X"1F",X"1F",X"1E",X"08",X"01",X"00",X"E0",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"30",X"00",X"7C",X"FC",X"F8",X"00",X"03",X"07",X"07",X"00",
		X"00",X"E0",X"E0",X"E0",X"00",X"01",X"08",X"1E",X"1F",X"1F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3E",
		X"00",X"07",X"07",X"03",X"00",X"F8",X"FC",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"38",X"08",X"00",X"E0",X"C0",X"01",X"01",X"C0",X"E0",X"E0",X"00",
		X"40",X"40",X"40",X"40",X"40",X"C0",X"40",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"7D",X"73",X"63",X"3C",X"00",X"00",X"00",
		X"07",X"07",X"07",X"01",X"60",X"C4",X"1C",X"1C",X"78",X"DA",X"5C",X"8F",X"07",X"01",X"01",X"00",
		X"C0",X"C1",X"C3",X"C7",X"07",X"07",X"62",X"10",X"00",X"C0",X"C0",X"E0",X"E7",X"FF",X"9F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"02",X"C2",X"F8",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"7D",X"73",X"63",X"3C",X"00",X"00",X"00",
		X"07",X"07",X"07",X"01",X"60",X"C4",X"1C",X"1C",X"78",X"DA",X"5C",X"8F",X"07",X"01",X"01",X"00",
		X"C2",X"83",X"87",X"8F",X"07",X"0F",X"46",X"24",X"00",X"C0",X"C0",X"E0",X"E7",X"FF",X"9F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"02",X"C2",X"F8",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"02",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"38",X"7C",X"F9",X"E3",X"C7",X"78",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"3C",X"C6",X"00",X"09",X"3F",X"74",X"D0",X"AA",X"6E",X"7C",X"7F",X"3F",X"1F",X"1C",X"07",
		X"00",X"10",X"00",X"C0",X"E0",X"80",X"00",X"00",X"02",X"03",X"41",X"31",X"D9",X"F8",X"3C",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"40",X"78",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"38",X"7C",X"F9",X"E3",X"C7",X"78",X"00",X"00",X"00",X"00",X"00",
		X"78",X"38",X"C4",X"00",X"09",X"3F",X"74",X"D0",X"AA",X"6E",X"7C",X"7F",X"3F",X"1D",X"1D",X"07",
		X"20",X"30",X"10",X"80",X"C0",X"80",X"00",X"00",X"02",X"03",X"41",X"31",X"D9",X"F8",X"3C",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"40",X"78",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",
		X"80",X"A4",X"FE",X"0E",X"1C",X"3C",X"7C",X"F8",X"F8",X"F8",X"F8",X"D0",X"90",X"50",X"C0",X"C0",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",
		X"30",X"A4",X"EE",X"0E",X"1C",X"3C",X"7C",X"F8",X"F8",X"F8",X"F8",X"D0",X"90",X"50",X"C0",X"C0",
		X"00",X"E0",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"7C",X"7C",X"3E",X"0E",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"5F",X"7E",X"29",X"07",X"E6",X"FE",X"E6",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"E6",X"FE",X"E6",X"07",X"29",X"7E",X"5F",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"FE",X"FF",
		X"5F",X"5F",X"7E",X"29",X"07",X"E6",X"FE",X"E6",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"E6",X"FE",X"E6",X"07",X"29",X"7E",X"5F",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"FC",X"FE",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"1F",X"1E",X"3C",X"3A",X"3F",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"1C",X"1C",X"0C",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"0F",X"07",X"0F",
		X"8B",X"0B",X"0F",X"07",X"05",X"00",X"82",X"E7",X"FB",X"FD",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"D8",X"E0",X"F0",X"F8",X"7C",X"3E",X"9E",X"8F",X"25",X"17",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"3E",X"DE",X"FD",X"FB",X"FB",X"F7",X"C7",X"83",X"80",X"03",X"05",X"85",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"8B",X"0B",X"0F",X"07",X"05",X"00",X"82",X"E7",X"FB",X"FD",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"D8",X"E0",X"F0",X"F8",X"7C",X"3C",X"9E",X"8E",X"2E",X"1C",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"07",X"07",X"03",X"01",X"00",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"C3",X"CF",X"FE",X"9C",X"3F",X"27",X"27",X"27",X"27",X"3F",X"9C",X"FE",X"CF",X"C3",X"01",
		X"00",X"20",X"70",X"70",X"20",X"F0",X"FE",X"FF",X"FF",X"FE",X"F0",X"20",X"70",X"70",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"06",X"0F",X"0E",X"1D",X"1D",X"1D",X"1D",X"0E",X"0F",X"06",X"40",X"40",X"00",
		X"00",X"00",X"20",X"78",X"D8",X"80",X"F8",X"7F",X"7F",X"F8",X"80",X"D8",X"78",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"33",X"33",X"13",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"A8",X"C8",X"B0",X"5F",X"5F",X"B0",X"C8",X"A8",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"62",X"F8",X"EF",X"F8",X"62",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"2F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"00",X"00",X"00",X"30",X"70",X"70",X"70",X"70",X"30",X"00",X"00",X"00",X"04",X"04",
		X"00",X"10",X"33",X"7F",X"77",X"EE",X"E8",X"E8",X"E9",X"EF",X"F7",X"7F",X"73",X"30",X"00",X"00",
		X"40",X"C0",X"D8",X"98",X"00",X"D0",X"FE",X"FE",X"FE",X"F0",X"00",X"98",X"D8",X"60",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"7F",X"7F",X"3F",X"00",X"00",
		X"1F",X"1F",X"0F",X"1B",X"10",X"10",X"90",X"B0",X"31",X"16",X"30",X"F8",X"D8",X"9C",X"1C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"C3",X"C3",X"C3",X"83",X"03",X"23",X"23",X"67",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6C",X"58",X"F0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",X"38",X"38",X"38",X"38",X"0C",X"86",X"C6",X"C3",
		X"00",X"00",X"00",X"00",X"30",X"58",X"E8",X"7C",X"5C",X"1E",X"5F",X"43",X"93",X"3B",X"32",X"36",
		X"3C",X"1E",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"30",X"30",X"A0",X"E0",X"40",X"40",X"40",X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"70",X"70",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"47",X"4F",
		X"F3",X"F3",X"F1",X"F1",X"61",X"01",X"01",X"03",X"0F",X"1F",X"3E",X"FC",X"FF",X"7F",X"39",X"00",
		X"C0",X"80",X"00",X"00",X"06",X"0C",X"0D",X"07",X"27",X"4F",X"07",X"73",X"FB",X"33",X"86",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"E1",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",
		X"60",X"E0",X"E4",X"64",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"78",X"78",X"78",X"70",X"70",X"70",X"70",X"70",X"33",X"30",X"00",X"07",X"1E",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"06",X"8C",X"F8",X"F0",X"C0",X"E6",X"F0",X"DC",X"4F",X"65",X"31",X"1F",X"0F",X"07",
		X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"D0",X"D0",X"F8",X"F0",X"E0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"30",X"F8",X"38",X"00",X"38",X"7C",X"7C",X"7C",X"7C",X"7C",X"39",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"F8",X"F8",
		X"F0",X"F0",X"70",X"38",X"7C",X"EF",X"E0",X"B0",X"B4",X"A2",X"A0",X"89",X"DD",X"FF",X"7E",X"3F",
		X"70",X"00",X"00",X"00",X"76",X"FE",X"3E",X"1C",X"18",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"01",X"01",X"18",X"3F",X"39",X"00",X"00",X"02",X"02",X"04",X"00",X"40",X"40",X"C0",X"E0",X"E0",
		X"C0",X"00",X"30",X"00",X"C0",X"E0",X"30",X"1C",X"1E",X"0E",X"70",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"3E",X"7E",X"70",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"32",X"7B",X"7B",X"7B",X"7F",X"7F",X"7E",X"3C",X"00",X"00",
		X"00",X"00",X"40",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"39",X"07",X"01",
		X"64",X"46",X"C2",X"82",X"02",X"02",X"02",X"02",X"02",X"46",X"4C",X"7C",X"F8",X"E0",X"80",X"E0",
		X"00",X"00",X"00",X"00",X"01",X"1C",X"38",X"38",X"18",X"08",X"0C",X"05",X"07",X"03",X"02",X"02",
		X"20",X"60",X"40",X"C0",X"C0",X"68",X"28",X"78",X"78",X"7D",X"BF",X"9F",X"1F",X"3E",X"3C",X"64",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"41",X"E2",X"E6",X"F6",X"7C",X"00",
		X"02",X"07",X"07",X"0E",X"6E",X"5C",X"DC",X"B8",X"BA",X"76",X"74",X"2C",X"08",X"18",X"10",X"30",
		X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"FB",X"DC",X"CC",X"EC",X"EC",X"EC",X"CC",X"D8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"87",X"C7",X"E7",X"E7",X"E7",X"E7",X"37",X"1F",X"08",X"03",X"07",X"07",
		X"40",X"13",X"FF",X"FF",X"FF",X"7F",X"3F",X"17",X"1F",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",
		X"78",X"F0",X"E0",X"C0",X"00",X"E0",X"FE",X"FE",X"FE",X"7C",X"F8",X"F0",X"60",X"00",X"00",X"00",
		X"00",X"C3",X"E7",X"FF",X"FF",X"7E",X"8D",X"DF",X"DF",X"F3",X"D0",X"D0",X"D8",X"4F",X"C7",X"C3",
		X"00",X"00",X"00",X"F8",X"0C",X"C6",X"E6",X"E6",X"C6",X"8E",X"1C",X"3C",X"F8",X"F0",X"EC",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1C",X"3C",X"3C",X"3C",X"38",X"38",X"38",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"15",X"37",X"3B",X"C3",X"E3",X"E3",X"C1",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"E3",X"F1",X"F8",X"FC",X"3E",X"9E",X"CF",X"E7",X"F7",X"F3",X"EB",X"63",X"33",X"1E",X"00",
		X"18",X"18",X"38",X"38",X"3C",X"7C",X"7C",X"7C",X"7E",X"3E",X"3E",X"1E",X"1F",X"1F",X"3F",X"3F",
		X"67",X"77",X"53",X"0B",X"23",X"33",X"1E",X"18",X"18",X"18",X"18",X"1C",X"3E",X"FF",X"FF",X"F7",
		X"03",X"07",X"0E",X"1E",X"1E",X"1E",X"1F",X"1E",X"1F",X"1F",X"6F",X"07",X"07",X"07",X"03",X"09",
		X"00",X"00",X"00",X"00",X"00",X"18",X"98",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"3E",X"9E",X"CF",
		X"38",X"38",X"38",X"38",X"38",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1E",X"1E",X"1F",X"0F",X"03",X"07",X"0F",X"0E",X"0D",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"38",
		X"00",X"00",X"00",X"01",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",
		X"67",X"4F",X"4F",X"7F",X"FF",X"07",X"00",X"99",X"FB",X"FF",X"FF",X"C7",X"03",X"02",X"00",X"00",
		X"20",X"80",X"C0",X"F0",X"FC",X"FE",X"7F",X"1F",X"86",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"C0",X"C3",X"BF",X"6F",X"F7",X"D7",X"E0",X"F0",X"E0",X"E0",X"84",X"18",X"3C",X"24",
		X"00",X"00",X"00",X"FC",X"FE",X"FE",X"CE",X"3C",X"70",X"00",X"00",X"00",X"00",X"20",X"70",X"70",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"C0",X"D0",X"CC",X"C1",X"43",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"03",X"43",X"C1",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"3E",X"3E",X"3F",X"3F",X"1F",X"1F",X"1E",X"08",X"01",X"00",X"E0",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"30",X"00",X"7C",X"FC",X"F8",X"00",X"03",X"03",X"03",X"00",
		X"00",X"F0",X"F0",X"E0",X"00",X"01",X"08",X"1E",X"1F",X"1F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3E",
		X"00",X"03",X"03",X"03",X"00",X"F8",X"FC",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"38",X"08",X"00",X"E0",X"C0",X"01",X"01",X"C0",X"F0",X"F0",X"00",
		X"40",X"40",X"40",X"40",X"40",X"C0",X"40",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"02",X"02",X"07",X"07",X"06",X"06",X"06",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0C",X"1C",X"1C",X"20",X"20",X"20",X"60",X"40",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"30",X"3C",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"60",X"F8",X"3C",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"E2",X"08",X"1E",X"3F",X"07",X"01",X"00",X"00",X"01",X"01",
		X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"38",X"00",X"00",X"00",X"08",X"1D",X"3C",X"3E",X"7E",X"7E",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",
		X"03",X"03",X"07",X"07",X"07",X"03",X"83",X"99",X"3C",X"00",X"00",X"C0",X"F0",X"78",X"18",X"00",
		X"E2",X"E2",X"E2",X"C6",X"C4",X"C4",X"84",X"0C",X"18",X"08",X"18",X"10",X"30",X"60",X"00",X"00",
		X"03",X"03",X"C1",X"F0",X"F8",X"38",X"09",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"00",X"C0",X"F0",X"70",X"00",X"00",X"82",X"C3",X"41",X"01",X"01",X"F1",X"F1",X"F3",X"F1",X"F3",
		X"0E",X"0E",X"0E",X"0E",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"09",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"90",X"FF",X"FF",X"00",
		X"0E",X"0C",X"0D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"0C",X"0C",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"38",X"7F",X"7F",X"FF",X"FF",X"7F",X"1F",
		X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0E",X"0E",X"0E",
		X"00",X"00",X"7F",X"FF",X"D0",X"00",X"00",X"0F",X"3F",X"1F",X"1F",X"5F",X"CF",X"C0",X"C0",X"00",
		X"07",X"07",X"07",X"03",X"00",X"06",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"20",X"00",X"C0",X"E5",X"0F",X"0E",X"04",X"00",X"03",X"3F",X"00",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",
		X"04",X"0E",X"0F",X"05",X"00",X"00",X"00",X"20",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"01",X"01",X"00",X"00",X"0E",X"1F",X"1F",X"1F",X"9F",X"0E",X"00",X"00",X"01",X"9F",X"BF",X"00",
		X"FE",X"FE",X"EE",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"1C",X"38",X"78",X"F8",X"F8",X"F0",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"0E",X"1F",X"9F",X"1F",X"1F",X"0E",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",
		X"38",X"1C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"EE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"31",X"38",X"1E",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"01",X"03",X"03",X"F3",X"E1",X"C0",X"30",X"F7",
		X"FF",X"FE",X"FE",X"FE",X"FE",X"7E",X"7E",X"36",X"86",X"C6",X"C6",X"CE",X"8C",X"18",X"78",X"F0",
		X"03",X"01",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"C6",X"86",X"36",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"E3",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"8C",X"CE",X"C6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"20",X"81",X"C5",X"18",X"18",X"00",X"3D",X"00",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"3E",X"1E",X"86",X"C6",X"C6",X"86",X"0C",X"18",X"F8",X"00",
		X"00",X"00",X"00",X"18",X"18",X"05",X"01",X"20",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"18",X"0C",X"86",X"C6",X"C6",X"86",X"1E",X"3E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"06",X"02",X"18",X"0E",X"00",X"00",X"03",X"00",
		X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",X"0E",X"02",X"32",X"32",X"02",X"06",X"0C",X"BC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"32",X"32",X"02",X"0E",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"02",X"0D",X"0D",X"C1",X"C3",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C3",X"C1",X"0D",X"0D",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"05",X"25",X"63",X"67",X"67",X"67",X"67",X"63",X"25",X"05",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"09",X"0B",X"0B",X"0B",X"0B",X"09",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",
		X"FF",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FD",X"FF",X"FF",X"FF",X"FF",X"03",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"FE",X"FC",X"00",X"00",
		X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FD",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"F8",
		X"00",X"00",X"FC",X"FE",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"70",X"3E",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1E",X"3E",X"70",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"40",X"00",X"00",X"00",X"80",X"20",X"84",X"10",X"42",X"90",X"05",X"20",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"12",X"40",X"08",X"21",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"20",X"05",X"90",X"42",X"10",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"21",X"08",X"40",X"12",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",
		X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"3F",X"7F",X"7F",X"3F",X"7F",X"FF",X"FF",X"7F",X"30",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"F8",X"78",X"30",
		X"06",X"8E",X"CE",X"CE",X"EE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"7C",X"18",
		X"0E",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"F6",X"F8",X"F8",X"78",X"30",
		X"38",X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"3C",X"3C",X"3C",X"3C",X"3C",X"78",X"70",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0C",X"0E",X"1E",X"3D",X"3F",X"17",X"0F",X"2F",X"3F",X"19",X"03",X"03",X"03",X"01",
		X"00",X"00",X"60",X"F0",X"70",X"F0",X"E0",X"E6",X"C7",X"B3",X"F0",X"F0",X"F8",X"F8",X"F0",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"E0",X"FF",X"FF",X"FF",X"E0",X"40",X"03",X"0F",X"1F",X"7F",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"3F",X"FE",X"F8",X"F0",X"C0",X"02",X"07",X"FF",X"FF",
		X"40",X"E0",X"F8",X"FC",X"FE",X"FF",X"EF",X"47",X"03",X"47",X"EF",X"FF",X"FE",X"FC",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"02",X"87",X"FF",X"FF",X"FF",X"87",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"70",X"E0",X"E0",X"70",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"30",X"60",X"21",X"61",X"61",X"21",X"60",X"30",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"70",X"E0",X"E0",X"70",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"30",X"60",X"21",X"61",X"61",X"21",X"60",X"30",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"84",X"C3",X"F1",X"F9",X"81",X"81",X"F9",X"F1",X"C3",X"84",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"87",X"8D",X"8D",X"87",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"E0",X"F0",X"CC",X"60",X"30",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"60",X"61",X"21",X"61",X"40",X"60",X"A0",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"70",X"88",X"80",X"F1",X"F9",X"F1",X"E3",X"03",X"87",X"0E",X"3C",X"C0",X"F0",X"70",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"80",X"80",X"86",X"0D",X"0D",X"07",X"03",X"FF",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"04",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C8",X"8C",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"38",X"34",X"1A",X"13",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"18",X"18",X"30",X"20",X"E0",X"A0",X"00",
		X"01",X"03",X"07",X"1F",X"7E",X"F8",X"E0",X"7F",X"7F",X"3E",X"73",X"61",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"00",X"06",X"0C",X"0D",X"07",X"E7",X"FF",X"FE",X"36",X"CC",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"C0",X"F8",X"FC",X"F8",X"71",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"38",X"34",X"12",X"13",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"18",X"18",X"30",X"20",X"E0",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"70",X"E0",X"E0",X"70",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"11",X"31",X"63",X"27",X"66",X"66",X"27",X"63",X"31",X"11",X"10",X"00",X"00",
		X"00",X"00",X"10",X"8C",X"87",X"C3",X"E3",X"03",X"03",X"E3",X"C3",X"87",X"8C",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"87",X"8D",X"8D",X"87",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"70",X"E0",X"E0",X"70",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"11",X"31",X"63",X"27",X"66",X"66",X"27",X"63",X"31",X"11",X"10",X"00",X"00",
		X"00",X"00",X"10",X"8C",X"83",X"C1",X"E1",X"01",X"01",X"E1",X"C1",X"83",X"8C",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"87",X"8D",X"8D",X"87",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"FF",X"C7",X"6C",X"3F",
		X"00",X"00",X"01",X"12",X"36",X"27",X"27",X"67",X"63",X"20",X"60",X"E0",X"B0",X"D1",X"C0",X"80",
		X"00",X"00",X"C0",X"20",X"00",X"C1",X"E1",X"C1",X"81",X"03",X"07",X"0F",X"8F",X"1E",X"30",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"86",X"8D",X"8D",X"87",X"07",X"0F",X"FF",X"FF",
		X"38",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"DF",X"DE",X"66",X"3B",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"98",X"CF",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"12",X"37",X"67",X"67",X"23",X"20",X"70",X"D0",X"80",
		X"0F",X"3F",X"FE",X"F8",X"C1",X"FF",X"7B",X"39",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"07",X"0F",X"7F",X"FF",X"FF",X"7B",X"9B",X"EE",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"00",X"C0",X"E1",X"C1",X"81",X"03",X"03",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"86",X"8C",X"8D",
		X"E7",X"FF",X"DE",X"67",X"39",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"98",X"CF",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"16",X"37",X"67",X"67",X"23",X"20",X"70",X"D0",X"80",
		X"0F",X"3F",X"FE",X"F8",X"C1",X"FF",X"7B",X"39",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"07",X"0F",X"7F",X"FF",X"FF",X"7B",X"9B",X"EE",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"00",X"C0",X"E0",X"C0",X"80",X"01",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"86",X"8C",X"8D",
		X"00",X"00",X"00",X"07",X"38",X"70",X"70",X"38",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"30",X"7C",X"3E",X"60",X"60",X"3E",X"7C",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"20",X"38",X"1E",X"0F",X"07",X"07",X"07",X"07",X"0F",X"1E",X"38",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0D",X"0D",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"70",X"E0",X"E0",X"70",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"30",X"7C",X"3E",X"60",X"60",X"3E",X"7C",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"60",X"78",X"3E",X"1F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3E",X"78",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0D",X"0D",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"FF",X"C7",X"6C",X"3F",X"00",X"00",X"00",
		X"1C",X"22",X"20",X"3C",X"7E",X"7C",X"38",X"60",X"F0",X"90",X"90",X"C0",X"80",X"00",X"00",X"00",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"1E",X"3C",X"78",X"30",X"3F",X"1C",X"38",X"30",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0D",X"0D",X"07",X"07",X"0F",X"7F",X"FF",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"7F",X"71",X"67",X"6F",X"66",X"30",X"1F",X"00",X"00",
		X"60",X"7C",X"3E",X"3C",X"78",X"50",X"C0",X"80",X"90",X"4C",X"6F",X"6F",X"C3",X"83",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",X"1E",X"3E",X"3C",X"7B",X"E3",X"FF",X"FF",X"FD",X"38",X"30",
		X"00",X"00",X"06",X"0C",X"0D",X"07",X"07",X"3F",X"FF",X"FF",X"FF",X"FB",X"33",X"86",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"71",X"FF",X"E3",X"CE",X"DE",X"CC",X"61",X"3F",X"00",
		X"60",X"7C",X"3E",X"3C",X"78",X"50",X"C0",X"80",X"10",X"0C",X"8F",X"CF",X"C7",X"83",X"00",X"00",
		X"07",X"07",X"07",X"07",X"0F",X"0F",X"1E",X"1E",X"1C",X"7B",X"E3",X"FF",X"FD",X"FC",X"38",X"30",
		X"00",X"00",X"06",X"0D",X"0D",X"07",X"07",X"3F",X"C7",X"7F",X"FF",X"F3",X"86",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"70",X"E0",X"E0",X"70",X"3E",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"11",X"30",X"20",X"61",X"61",X"01",X"41",X"E1",X"21",X"20",X"00",X"00",X"00",
		X"00",X"00",X"8C",X"C7",X"C3",X"F1",X"F9",X"81",X"81",X"F9",X"F1",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"86",X"8D",X"8D",X"87",X"83",X"FF",X"FC",X"00",X"00",X"00",X"00",
		X"08",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"D0",X"88",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"78",X"26",X"20",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"18",X"18",X"30",X"20",X"30",X"10",X"00",
		X"01",X"03",X"07",X"0F",X"3E",X"F8",X"E0",X"5F",X"7F",X"3B",X"71",X"60",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"06",X"0C",X"0D",X"07",X"E7",X"FF",X"3E",X"CC",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"C0",X"F8",X"FC",X"F8",X"71",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F8",X"3C",X"1F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"07",X"07",X"03",X"03",X"03",
		X"00",X"00",X"10",X"10",X"02",X"12",X"10",X"10",X"18",X"0C",X"07",X"0F",X"07",X"07",X"03",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"1C",X"0F",X"07",X"03",X"01",X"11",X"08",X"00",X"00",X"00",X"1C",X"1F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"00",X"18",X"1C",X"07",X"03",X"02",X"02",X"12",X"12",X"02",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"05",X"01",X"10",X"10",X"10",X"10",X"02",X"02",X"00",X"00",X"18",X"0C",X"06",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"0F",X"0F",X"0F",X"07",X"01",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"08",
		X"70",X"10",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E7",X"67",X"61",X"60",X"60",X"60",X"70",X"50",X"00",X"00",X"00",X"80",X"80",X"C0",X"F0",X"F0",
		X"80",X"F8",X"FC",X"FC",X"3C",X"1C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"20",X"00",X"00",X"04",X"86",X"C7",X"E7",X"E1",X"60",X"60",X"00",X"00",X"00",X"C4",X"E6",
		X"18",X"18",X"18",X"18",X"08",X"00",X"80",X"C0",X"F0",X"F8",X"3E",X"1F",X"07",X"03",X"00",X"00",
		X"80",X"E4",X"E6",X"67",X"67",X"23",X"03",X"43",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"61",
		X"03",X"01",X"00",X"00",X"00",X"30",X"38",X"3E",X"1F",X"07",X"03",X"00",X"00",X"00",X"18",X"18",
		X"60",X"70",X"F3",X"F3",X"33",X"23",X"20",X"60",X"60",X"60",X"60",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"FF",X"FF",X"7F",X"07",X"00",X"00",X"00",X"E0",X"20",X"03",X"03",X"03",
		X"00",X"00",X"00",X"80",X"A0",X"B0",X"B0",X"B0",X"30",X"30",X"70",X"70",X"70",X"70",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"20",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"70",X"70",X"60",X"20",X"00",X"00",X"40",X"E0",X"E0",X"E0",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"70",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"01",X"00",X"00",X"0C",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"04",X"04",
		X"04",X"80",X"80",X"30",X"38",X"0E",X"07",X"01",X"80",X"C0",X"C0",X"E0",X"F1",X"70",X"38",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"30",X"38",X"0C",X"04",X"00",X"00",X"30",X"38",X"0E",X"07",X"01",X"00",X"30",X"38",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"1E",X"0E",X"07",X"07",X"23",X"11",X"00",X"00",X"00",X"30",X"3C",X"3E",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E1",X"E1",X"E0",X"E0",X"E0",X"E0",X"60",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"F1",X"F9",X"39",X"19",X"09",X"01",X"C1",X"C1",X"41",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C1",X"C1",X"C1",X"C1",X"C1",X"F1",X"F9",X"39",X"19",X"09",X"01",X"C1",X"C1",X"C1",X"C1",X"C1",
		X"80",X"A0",X"B0",X"3C",X"3C",X"0E",X"07",X"01",X"00",X"00",X"10",X"18",X"18",X"18",X"08",X"00",
		X"00",X"00",X"00",X"01",X"81",X"C1",X"E1",X"F1",X"79",X"39",X"18",X"09",X"07",X"83",X"C3",X"C1",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FF",X"3F",X"1F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"83",X"83",X"13",X"13",X"83",X"82",X"C0",X"C0",X"FF",X"9F",X"03",X"03",X"03",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"63",X"73",X"63",X"63",X"61",X"61",X"23",X"13",X"03",X"03",X"00",X"C0",X"E3",X"3B",X"1F",X"07",
		X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",
		X"40",X"60",X"78",X"7C",X"7D",X"3D",X"0D",X"05",X"11",X"11",X"13",X"13",X"03",X"03",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
