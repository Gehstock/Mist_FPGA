library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity berzerk_program2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of berzerk_program2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"07",X"01",X"0B",X"3C",X"7E",X"C7",X"D7",X"C7",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",
		X"3C",X"7E",X"E3",X"EB",X"E3",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F1",
		X"F5",X"F1",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F8",X"FA",X"F8",X"7E",
		X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"FC",X"FD",X"FC",X"7E",X"3C",X"DB",X"7E",
		X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",
		X"0B",X"3C",X"7E",X"3F",X"BF",X"3F",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",
		X"1F",X"5F",X"1F",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"8F",X"AF",X"8F",
		X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F1",X"F5",X"F1",X"7E",X"3C",X"DB",
		X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F1",X"F5",X"F1",X"7E",X"3C",X"6D",X"FF",X"FE",X"36",
		X"01",X"0B",X"3C",X"7E",X"F1",X"F5",X"F1",X"7E",X"3C",X"B6",X"FF",X"7F",X"6C",X"01",X"0B",X"3C",
		X"7E",X"8F",X"AF",X"8F",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"8F",X"AF",
		X"8F",X"7E",X"3C",X"B6",X"FF",X"7F",X"6C",X"01",X"0B",X"3C",X"7E",X"8F",X"AF",X"8F",X"7E",X"3C",
		X"6D",X"FF",X"FE",X"36",X"01",X"0B",X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"FF",X"1F",X"F8",
		X"E7",X"01",X"0B",X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"1F",X"F8",X"FF",X"07",X"01",X"0B",
		X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"F8",X"FF",X"1F",X"E0",X"01",X"0B",X"3C",X"7E",X"FF",
		X"C7",X"D7",X"46",X"3C",X"FF",X"1F",X"F8",X"E7",X"01",X"0B",X"3C",X"7E",X"FF",X"C7",X"D7",X"46",
		X"3C",X"F8",X"FF",X"1F",X"E0",X"01",X"0B",X"3C",X"7E",X"FF",X"C7",X"D7",X"46",X"3C",X"1F",X"F8",
		X"FF",X"07",X"02",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"07",X"E0",X"0F",X"78",X"13",X"C8",X"0A",X"D0",X"03",X"40",X"33",X"CC",X"09",X"F0",
		X"02",X"48",X"1E",X"78",X"06",X"60",X"02",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"06",X"60",X"12",X"48",X"08",X"90",X"10",X"08",X"22",X"44",X"24",X"48",X"0A",X"90",
		X"13",X"60",X"08",X"18",X"14",X"20",X"02",X"40",X"06",X"60",X"02",X"13",X"00",X"00",X"02",X"00",
		X"00",X"20",X"01",X"08",X"10",X"00",X"02",X"40",X"20",X"12",X"08",X"01",X"80",X"20",X"08",X"82",
		X"40",X"02",X"04",X"10",X"21",X"00",X"08",X"04",X"20",X"02",X"04",X"08",X"20",X"20",X"10",X"08",
		X"18",X"0C",X"01",X"01",X"00",X"00",X"82",X"01",X"02",X"18",X"18",X"00",X"82",X"01",X"03",X"10",
		X"38",X"10",X"00",X"82",X"01",X"04",X"10",X"38",X"38",X"10",X"00",X"82",X"01",X"05",X"18",X"3C",
		X"3C",X"3C",X"18",X"00",X"82",X"01",X"06",X"38",X"7C",X"7C",X"7C",X"7C",X"38",X"00",X"82",X"01",
		X"07",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"1C",X"00",X"82",X"01",X"08",X"18",X"7E",X"5A",X"FF",
		X"FF",X"7E",X"7E",X"18",X"00",X"81",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",
		X"7E",X"18",X"80",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",X"7E",X"18",
		X"40",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",X"7E",X"18",X"01",X"0A",
		X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",X"7E",X"18",X"00",X"82",X"01",X"09",X"00",X"00",
		X"00",X"3C",X"5A",X"FF",X"FF",X"C3",X"7E",X"00",X"81",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",
		X"FF",X"C3",X"7E",X"7E",X"18",X"80",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"C3",
		X"7E",X"7E",X"18",X"40",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"C3",X"7E",X"7E",
		X"18",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"C3",X"7E",X"7E",X"18",X"00",X"81",X"01",
		X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"E7",X"5A",X"7E",X"18",X"80",X"80",X"01",X"0A",X"18",
		X"7E",X"7E",X"DB",X"FF",X"FF",X"E7",X"5A",X"7E",X"18",X"40",X"80",X"01",X"0A",X"18",X"7E",X"7E",
		X"DB",X"FF",X"FF",X"E7",X"5A",X"7E",X"18",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"E7",
		X"5A",X"7E",X"18",X"00",X"82",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"3C",X"5A",X"C3",X"FF",
		X"00",X"82",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"5A",X"FF",X"00",X"82",X"01",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"FF",X"00",X"82",X"01",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"10",X"18",X"18",X"00",X"3C",X"5A",X"5A",X"5A",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"18",X"01",X"10",X"18",X"18",X"00",X"3C",X"5A",
		X"9A",X"59",X"18",X"18",X"24",X"22",X"41",X"41",X"81",X"81",X"C0",X"01",X"10",X"00",X"18",X"18",
		X"00",X"3C",X"5C",X"5A",X"3A",X"18",X"18",X"14",X"12",X"F2",X"82",X"02",X"03",X"01",X"10",X"18",
		X"18",X"00",X"3C",X"3C",X"3C",X"1A",X"18",X"18",X"0C",X"0A",X"0F",X"78",X"48",X"08",X"0C",X"01",
		X"10",X"18",X"18",X"00",X"3C",X"5A",X"59",X"9A",X"18",X"18",X"24",X"44",X"82",X"82",X"81",X"81",
		X"03",X"01",X"10",X"00",X"18",X"18",X"00",X"3C",X"3A",X"3A",X"DC",X"18",X"18",X"28",X"48",X"4F",
		X"41",X"40",X"80",X"01",X"10",X"18",X"18",X"00",X"3C",X"3C",X"3C",X"58",X"18",X"18",X"30",X"50",
		X"F0",X"1E",X"12",X"10",X"30",X"01",X"10",X"00",X"18",X"18",X"00",X"3C",X"5A",X"5A",X"5A",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"3C",X"01",X"11",X"18",X"24",X"24",X"42",X"81",X"81",X"81",
		X"81",X"81",X"42",X"24",X"24",X"24",X"24",X"24",X"42",X"3C",X"01",X"11",X"18",X"24",X"24",X"7E",
		X"C3",X"A5",X"A5",X"A5",X"E7",X"66",X"24",X"24",X"24",X"24",X"66",X"42",X"3C",X"01",X"11",X"3C",
		X"3C",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"3C",X"3C",X"3C",X"7E",X"7E",X"7E",
		X"01",X"0F",X"18",X"19",X"02",X"1C",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"1C",X"01",X"0F",X"18",X"18",X"00",X"1F",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"18",X"18",X"1C",X"1A",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"3C",X"3C",X"3A",X"3A",X"3A",X"18",X"18",X"18",
		X"18",X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"3C",X"3C",X"5C",X"9C",X"1C",X"18",X"18",
		X"18",X"18",X"18",X"18",X"38",X"01",X"0F",X"18",X"18",X"00",X"F8",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"38",X"01",X"0F",X"98",X"58",X"20",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"38",X"01",X"0F",X"18",X"18",X"00",X"1D",X"1B",X"19",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"00",X"3E",X"41",X"5D",X"51",X"5D",X"41",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"00",X"10",X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"7F",
		X"14",X"7F",X"14",X"14",X"14",X"14",X"7F",X"54",X"54",X"7F",X"15",X"15",X"7F",X"14",X"20",X"51",
		X"22",X"04",X"08",X"10",X"22",X"45",X"02",X"00",X"18",X"24",X"28",X"10",X"29",X"46",X"46",X"39",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"10",X"10",X"10",X"10",X"10",
		X"08",X"04",X"10",X"08",X"04",X"04",X"04",X"04",X"04",X"08",X"10",X"00",X"00",X"08",X"2A",X"1C",
		X"1C",X"2A",X"08",X"00",X"00",X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",X"80",X"00",X"00",
		X"00",X"18",X"18",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"20",
		X"40",X"1C",X"22",X"41",X"41",X"41",X"41",X"41",X"22",X"1C",X"08",X"18",X"08",X"08",X"08",X"08",
		X"08",X"08",X"1C",X"3E",X"41",X"01",X"01",X"3E",X"40",X"40",X"40",X"7F",X"3E",X"41",X"01",X"01",
		X"1E",X"01",X"01",X"41",X"3E",X"02",X"06",X"0A",X"12",X"22",X"7F",X"02",X"02",X"02",X"7F",X"40",
		X"40",X"40",X"7E",X"01",X"01",X"41",X"3E",X"3E",X"41",X"40",X"40",X"7E",X"41",X"41",X"41",X"3E",
		X"7F",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"08",X"3E",X"41",X"41",X"41",X"3E",X"41",X"41",
		X"41",X"3E",X"3E",X"41",X"41",X"41",X"3F",X"01",X"01",X"41",X"3E",X"00",X"00",X"00",X"18",X"18",
		X"00",X"00",X"18",X"18",X"98",X"18",X"00",X"00",X"18",X"18",X"08",X"10",X"00",X"02",X"04",X"08",
		X"10",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"00",X"3E",X"00",X"3E",X"00",X"00",X"00",X"20",
		X"10",X"08",X"04",X"02",X"04",X"08",X"10",X"20",X"1C",X"22",X"02",X"02",X"04",X"08",X"08",X"00",
		X"08",X"3E",X"41",X"4F",X"49",X"49",X"4F",X"40",X"40",X"3F",X"3E",X"41",X"41",X"41",X"7F",X"41",
		X"41",X"41",X"41",X"7E",X"41",X"41",X"41",X"7E",X"41",X"41",X"41",X"7E",X"3E",X"41",X"40",X"40",
		X"40",X"40",X"40",X"41",X"3E",X"7E",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"7E",X"7F",X"40",
		X"40",X"40",X"7C",X"40",X"40",X"40",X"7F",X"7F",X"40",X"40",X"40",X"7C",X"40",X"40",X"40",X"40",
		X"3E",X"41",X"40",X"40",X"47",X"41",X"41",X"41",X"3F",X"41",X"41",X"41",X"41",X"7F",X"41",X"41",
		X"41",X"41",X"1C",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"1C",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"41",X"3E",X"41",X"42",X"44",X"48",X"50",X"68",X"44",X"42",X"41",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"7F",X"41",X"63",X"55",X"49",X"41",X"41",X"41",X"41",X"41",X"41",
		X"61",X"51",X"49",X"45",X"43",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"41",X"41",X"41",X"41",
		X"3E",X"7E",X"41",X"41",X"41",X"7E",X"40",X"40",X"40",X"40",X"3E",X"41",X"41",X"41",X"41",X"41",
		X"45",X"42",X"3D",X"7E",X"41",X"41",X"41",X"7E",X"48",X"44",X"42",X"41",X"3E",X"41",X"40",X"40",
		X"3E",X"01",X"01",X"41",X"3E",X"7F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"41",X"41",
		X"41",X"41",X"41",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"22",X"22",X"14",X"14",X"08",X"08",
		X"41",X"41",X"41",X"41",X"41",X"49",X"55",X"63",X"41",X"41",X"41",X"22",X"14",X"08",X"14",X"22",
		X"41",X"41",X"41",X"41",X"22",X"14",X"08",X"08",X"08",X"08",X"08",X"7F",X"01",X"02",X"04",X"08",
		X"10",X"20",X"40",X"7F",X"3C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"3C",X"00",X"00",X"40",
		X"20",X"10",X"08",X"04",X"02",X"01",X"3C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"3C",X"08",
		X"14",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"18",X"18",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"46",X"42",
		X"42",X"46",X"3A",X"40",X"40",X"40",X"5C",X"62",X"42",X"42",X"62",X"5C",X"00",X"00",X"00",X"3C",
		X"42",X"40",X"40",X"42",X"3C",X"02",X"02",X"02",X"3A",X"46",X"42",X"42",X"46",X"3A",X"00",X"00",
		X"00",X"3C",X"42",X"7E",X"40",X"40",X"3C",X"0C",X"12",X"10",X"10",X"38",X"10",X"10",X"10",X"10",
		X"BA",X"46",X"42",X"42",X"46",X"3A",X"02",X"42",X"3C",X"40",X"40",X"40",X"7C",X"42",X"42",X"42",
		X"42",X"42",X"00",X"08",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"84",X"04",X"04",X"04",X"04",
		X"04",X"04",X"44",X"38",X"40",X"40",X"40",X"44",X"48",X"50",X"70",X"48",X"44",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"76",X"49",X"49",X"49",X"49",X"49",X"00",
		X"00",X"00",X"7C",X"42",X"42",X"42",X"42",X"42",X"00",X"00",X"00",X"3C",X"42",X"42",X"42",X"42",
		X"3C",X"DC",X"62",X"42",X"42",X"62",X"5C",X"40",X"40",X"40",X"BA",X"46",X"42",X"42",X"46",X"3A",
		X"02",X"02",X"02",X"00",X"00",X"00",X"5C",X"62",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"3C",
		X"42",X"30",X"0C",X"42",X"3C",X"00",X"10",X"10",X"7C",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"42",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"28",X"10",
		X"00",X"00",X"00",X"41",X"41",X"41",X"49",X"49",X"36",X"00",X"00",X"00",X"42",X"24",X"18",X"18",
		X"24",X"42",X"C2",X"42",X"42",X"42",X"46",X"3A",X"02",X"42",X"3C",X"00",X"00",X"00",X"7E",X"04",
		X"08",X"10",X"20",X"7E",X"0C",X"10",X"10",X"10",X"20",X"10",X"10",X"10",X"0C",X"08",X"08",X"08",
		X"00",X"00",X"08",X"08",X"08",X"00",X"18",X"04",X"04",X"04",X"02",X"04",X"04",X"04",X"18",X"08",
		X"00",X"1C",X"2A",X"08",X"08",X"14",X"22",X"00",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",
		X"55",X"08",X"00",X"1C",X"2A",X"08",X"08",X"14",X"22",X"00",X"02",X"28",X"00",X"0F",X"00",X"3F",
		X"00",X"FF",X"01",X"FF",X"03",X"FF",X"07",X"FF",X"0F",X"FF",X"1F",X"FF",X"1F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"3F",X"FF",X"3F",X"FF",X"1F",X"FF",X"1F",X"FF",X"0F",X"FF",
		X"07",X"FF",X"03",X"FF",X"01",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"0F",X"02",X"28",X"F0",X"00",
		X"FC",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"C0",X"FF",X"E0",X"FF",X"F0",X"FF",X"F8",X"FF",X"F8",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FC",X"FF",X"FC",X"FF",X"F8",X"FF",X"F8",
		X"FF",X"F0",X"FF",X"E0",X"FF",X"C0",X"FF",X"80",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"01",X"0C",
		X"20",X"30",X"18",X"0C",X"06",X"03",X"70",X"F8",X"C8",X"C8",X"F8",X"70",X"01",X"0C",X"04",X"0C",
		X"18",X"30",X"60",X"C0",X"0E",X"1F",X"13",X"13",X"1F",X"0E",X"02",X"07",X"00",X"03",X"00",X"1F",
		X"00",X"3C",X"00",X"60",X"00",X"C0",X"01",X"80",X"01",X"00",X"02",X"07",X"C0",X"00",X"F8",X"00",
		X"3C",X"00",X"06",X"00",X"03",X"00",X"01",X"80",X"00",X"80",X"02",X"07",X"01",X"00",X"01",X"80",
		X"00",X"C0",X"00",X"60",X"00",X"3C",X"00",X"1F",X"00",X"03",X"02",X"07",X"00",X"80",X"01",X"80",
		X"03",X"00",X"06",X"00",X"3C",X"00",X"F8",X"00",X"C0",X"00",X"02",X"02",X"FF",X"FF",X"FF",X"FF",
		X"02",X"08",X"00",X"30",X"00",X"78",X"00",X"CC",X"01",X"86",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"F0",X"02",X"08",X"0C",X"00",X"1E",X"00",X"33",X"00",X"61",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"C0",X"01",X"0B",X"F8",X"F8",X"98",X"68",X"68",X"08",X"68",X"68",X"68",X"F8",
		X"F8",X"02",X"06",X"00",X"00",X"FF",X"00",X"02",X"80",X"07",X"80",X"02",X"80",X"FF",X"00",X"02",
		X"06",X"60",X"00",X"FF",X"00",X"05",X"80",X"02",X"80",X"05",X"80",X"FF",X"00",X"02",X"06",X"06",
		X"00",X"FF",X"00",X"02",X"80",X"07",X"80",X"02",X"80",X"FF",X"00",X"02",X"06",X"00",X"00",X"FF",
		X"60",X"05",X"B0",X"02",X"80",X"05",X"80",X"FF",X"00",X"02",X"06",X"00",X"00",X"FF",X"00",X"02",
		X"B0",X"07",X"98",X"02",X"80",X"FF",X"00",X"02",X"06",X"00",X"00",X"FF",X"00",X"05",X"80",X"02",
		X"80",X"05",X"98",X"FF",X"0C",X"02",X"08",X"00",X"00",X"FF",X"00",X"02",X"80",X"07",X"80",X"02",
		X"80",X"FF",X"00",X"00",X"0C",X"00",X"06",X"02",X"06",X"00",X"00",X"FF",X"00",X"05",X"80",X"02",
		X"80",X"05",X"80",X"FF",X"00",X"01",X"17",X"30",X"78",X"FC",X"FC",X"FC",X"8C",X"B4",X"B4",X"8C",
		X"B4",X"B4",X"8C",X"FC",X"FC",X"78",X"30",X"30",X"78",X"30",X"34",X"3F",X"1F",X"04",X"02",X"1D",
		X"3F",X"FC",X"1F",X"F8",X"0F",X"F0",X"07",X"E0",X"FF",X"FF",X"80",X"01",X"93",X"29",X"AA",X"B9",
		X"BB",X"39",X"AA",X"A9",X"AA",X"A9",X"80",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"09",X"00",X"00",X"00",X"00",
		X"C0",X"40",X"40",X"40",X"78",X"01",X"08",X"00",X"00",X"00",X"00",X"C0",X"40",X"40",X"78",X"01",
		X"05",X"00",X"00",X"00",X"00",X"F8",X"01",X"05",X"00",X"78",X"40",X"40",X"C0",X"01",X"05",X"78",
		X"40",X"40",X"40",X"C0",X"01",X"05",X"04",X"04",X"FC",X"04",X"04",X"01",X"05",X"02",X"0C",X"74",
		X"84",X"08",X"01",X"05",X"02",X"1A",X"24",X"C8",X"08",X"01",X"05",X"09",X"12",X"24",X"48",X"90",
		X"01",X"05",X"10",X"13",X"24",X"58",X"40",X"01",X"05",X"10",X"21",X"2E",X"30",X"40",X"01",X"05",
		X"20",X"20",X"3F",X"20",X"20",X"01",X"05",X"40",X"30",X"2E",X"21",X"10",X"01",X"05",X"40",X"58",
		X"24",X"13",X"10",X"01",X"05",X"90",X"48",X"24",X"12",X"09",X"01",X"05",X"08",X"C8",X"24",X"1A",
		X"02",X"01",X"05",X"08",X"84",X"74",X"0C",X"02",X"01",X"01",X"5A",X"01",X"02",X"FF",X"5A",X"01",
		X"03",X"7E",X"FF",X"5A",X"01",X"04",X"DB",X"7E",X"FF",X"5A",X"01",X"05",X"3C",X"DB",X"7E",X"FF",
		X"5A",X"01",X"06",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"07",X"FF",X"7E",X"3C",X"DB",X"7E",
		X"FF",X"5A",X"01",X"08",X"EF",X"FF",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"09",X"FF",X"EF",
		X"FF",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0A",X"7E",X"FF",X"EF",X"FF",X"7E",X"3C",X"DB",
		X"7E",X"FF",X"5A",X"01",X"10",X"38",X"54",X"7C",X"28",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",
		X"10",X"38",X"28",X"28",X"6C",X"01",X"10",X"38",X"54",X"7C",X"28",X"38",X"10",X"7C",X"92",X"BA",
		X"90",X"38",X"10",X"38",X"28",X"68",X"0C",X"01",X"10",X"38",X"54",X"7C",X"28",X"38",X"10",X"7C",
		X"92",X"BA",X"12",X"38",X"10",X"38",X"28",X"2C",X"60",X"01",X"10",X"38",X"7C",X"7C",X"38",X"38",
		X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"38",X"28",X"28",X"6C",X"01",X"10",X"38",X"7C",X"7C",
		X"38",X"38",X"10",X"7C",X"92",X"BA",X"12",X"38",X"10",X"38",X"28",X"2C",X"60",X"01",X"10",X"38",
		X"7C",X"7C",X"38",X"38",X"10",X"7C",X"92",X"BA",X"90",X"38",X"10",X"38",X"28",X"68",X"0C",X"01",
		X"10",X"38",X"74",X"7C",X"30",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"38",X"28",X"28",
		X"3C",X"01",X"10",X"38",X"74",X"7C",X"30",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"7C",
		X"44",X"44",X"66",X"01",X"10",X"38",X"74",X"7C",X"30",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",
		X"10",X"10",X"10",X"10",X"18",X"01",X"10",X"38",X"5C",X"7C",X"18",X"38",X"10",X"7C",X"92",X"BA",
		X"92",X"38",X"10",X"38",X"28",X"28",X"78",X"01",X"10",X"38",X"5C",X"7C",X"18",X"38",X"10",X"7C",
		X"92",X"BA",X"92",X"38",X"10",X"7C",X"44",X"44",X"CC",X"01",X"10",X"38",X"5C",X"7C",X"18",X"38",
		X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"10",X"10",X"10",X"30",X"02",X"1E",X"80",X"00",X"80",
		X"00",X"80",X"00",X"80",X"07",X"80",X"08",X"80",X"10",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"40",X"40",X"40",X"40",X"20",X"80",X"1F",X"00",X"02",X"1E",X"00",X"01",X"00",X"01",X"00",
		X"01",X"E0",X"01",X"10",X"01",X"08",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",
		X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",
		X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"02",
		X"02",X"02",X"02",X"01",X"04",X"00",X"F8",X"01",X"08",X"3C",X"00",X"FF",X"FF",X"FF",X"7E",X"7E",
		X"3C",X"02",X"04",X"0F",X"FF",X"08",X"01",X"08",X"01",X"0F",X"FF",X"02",X"04",X"0F",X"FF",X"08",
		X"01",X"09",X"F9",X"0F",X"FF",X"02",X"06",X"0F",X"FF",X"08",X"01",X"0B",X"FD",X"0F",X"FF",X"01",
		X"F8",X"00",X"F0",X"02",X"08",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"03",X"FC",X"03",
		X"FC",X"01",X"F8",X"00",X"F0",X"02",X"0A",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"07",
		X"BE",X"07",X"BE",X"03",X"FC",X"03",X"FC",X"01",X"F8",X"00",X"F0",X"02",X"0C",X"0F",X"FF",X"08",
		X"01",X"0F",X"BF",X"0F",X"BF",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"03",X"FC",X"03",
		X"FC",X"01",X"F8",X"00",X"F0",X"02",X"0E",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"07",
		X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"03",X"FC",X"03",X"FC",X"01",
		X"F8",X"00",X"F0",X"02",X"0F",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"07",X"BE",X"07",
		X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"03",X"FC",X"03",X"FC",X"01",
		X"F8",X"00",X"F0",X"02",X"0C",X"1E",X"00",X"33",X"00",X"73",X"80",X"73",X"80",X"F3",X"C0",X"FF",
		X"C0",X"FF",X"C0",X"F3",X"C0",X"73",X"80",X"73",X"80",X"33",X"00",X"1E",X"00",X"02",X"0C",X"1E",
		X"00",X"3F",X"00",X"4F",X"80",X"67",X"80",X"E7",X"C0",X"FF",X"C0",X"FF",X"C0",X"F9",X"C0",X"79",
		X"80",X"7C",X"80",X"3F",X"00",X"1E",X"00",X"02",X"0C",X"1E",X"00",X"3F",X"00",X"7F",X"80",X"7F",
		X"80",X"FF",X"C0",X"8C",X"40",X"8C",X"40",X"FF",X"C0",X"7F",X"80",X"7F",X"80",X"3F",X"00",X"1E",
		X"00",X"02",X"0C",X"1E",X"00",X"3F",X"00",X"7C",X"80",X"79",X"80",X"F9",X"C0",X"FF",X"C0",X"FF",
		X"C0",X"E7",X"C0",X"67",X"80",X"4F",X"80",X"3F",X"00",X"1E",X"00",X"02",X"08",X"FF",X"F0",X"CF",
		X"30",X"B6",X"D0",X"BE",X"D0",X"A6",X"D0",X"B6",X"D0",X"C7",X"30",X"FF",X"F0",X"02",X"08",X"FF",
		X"F0",X"CE",X"30",X"B7",X"70",X"BF",X"70",X"A7",X"70",X"B7",X"70",X"C6",X"30",X"FF",X"F0",X"02",
		X"08",X"FF",X"F0",X"BB",X"B0",X"D7",X"30",X"EF",X"B0",X"EF",X"B0",X"D7",X"B0",X"BB",X"10",X"FF",
		X"F0",X"02",X"08",X"FF",X"F0",X"BA",X"10",X"D6",X"F0",X"EE",X"30",X"EF",X"D0",X"EF",X"D0",X"EE",
		X"30",X"FF",X"F0",X"01",X"10",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"18",X"18",X"3C",
		X"18",X"18",X"3C",X"18",X"18",X"01",X"08",X"3C",X"18",X"18",X"3C",X"18",X"18",X"3C",X"18",X"02",
		X"08",X"0E",X"00",X"01",X"C0",X"00",X"30",X"00",X"20",X"00",X"40",X"00",X"30",X"00",X"0C",X"00",
		X"03",X"02",X"08",X"0E",X"00",X"01",X"C0",X"00",X"30",X"00",X"70",X"00",X"C0",X"00",X"30",X"00",
		X"0C",X"00",X"03",X"02",X"08",X"00",X"00",X"0F",X"80",X"00",X"60",X"00",X"80",X"01",X"80",X"00",
		X"60",X"00",X"18",X"00",X"07",X"02",X"08",X"00",X"00",X"00",X"00",X"0E",X"00",X"01",X"C0",X"00",
		X"60",X"00",X"E0",X"00",X"1C",X"00",X"07",X"02",X"08",X"00",X"00",X"0C",X"00",X"03",X"80",X"00",
		X"70",X"00",X"20",X"00",X"40",X"00",X"38",X"00",X"07",X"02",X"08",X"00",X"00",X"00",X"01",X"00",
		X"C6",X"00",X"A8",X"01",X"30",X"02",X"00",X"04",X"00",X"08",X"00",X"02",X"08",X"00",X"01",X"00",
		X"02",X"00",X"64",X"00",X"98",X"01",X"00",X"02",X"00",X"04",X"00",X"08",X"00",X"02",X"08",X"00",
		X"00",X"00",X"03",X"00",X"0C",X"00",X"10",X"00",X"E0",X"03",X"00",X"04",X"00",X"08",X"00",X"02",
		X"08",X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"80",X"00",X"30",X"01",X"C0",X"0E",X"00",X"00",
		X"00",X"02",X"08",X"00",X"03",X"00",X"0E",X"00",X"18",X"00",X"D0",X"01",X"B0",X"02",X"00",X"04",
		X"00",X"08",X"00",X"02",X"08",X"00",X"00",X"00",X"07",X"00",X"8C",X"00",X"C8",X"01",X"B0",X"02",
		X"10",X"04",X"00",X"08",X"00",X"02",X"02",X"FF",X"F8",X"FF",X"F8",X"02",X"02",X"FF",X"F0",X"FF",
		X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
