library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_8L is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_8L is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"BF",X"BB",X"FE",X"EF",X"FB",X"E9",X"FE",X"FF",X"ED",X"AA",X"FA",X"FA",X"EF",X"B3",X"FF",
		X"BF",X"F2",X"AF",X"EB",X"EE",X"FA",X"F9",X"00",X"BA",X"FE",X"AB",X"EF",X"BF",X"FE",X"FF",X"00",
		X"BB",X"FA",X"FE",X"AB",X"FF",X"EF",X"DA",X"EB",X"BC",X"EA",X"7F",X"BB",X"BF",X"BE",X"EF",X"EB",
		X"BD",X"3A",X"BE",X"EB",X"EE",X"FF",X"A0",X"00",X"BA",X"FF",X"EF",X"EE",X"BF",X"A3",X"01",X"00",
		X"C0",X"00",X"00",X"80",X"C0",X"80",X"80",X"80",X"00",X"01",X"00",X"01",X"06",X"05",X"00",X"00",
		X"80",X"00",X"00",X"80",X"80",X"80",X"C0",X"F4",X"01",X"01",X"07",X"00",X"00",X"06",X"07",X"0D",
		X"80",X"80",X"C0",X"00",X"80",X"80",X"C0",X"C0",X"0B",X"37",X"3A",X"CE",X"3F",X"05",X"03",X"BF",
		X"80",X"80",X"00",X"01",X"80",X"80",X"80",X"80",X"0A",X"7B",X"6F",X"4F",X"B6",X"FD",X"2B",X"01",
		X"38",X"68",X"5C",X"BC",X"EC",X"AE",X"4E",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F6",X"76",X"73",X"D3",X"D9",X"F9",X"B8",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"00",X"80",X"80",X"C0",X"80",X"80",X"01",X"01",X"0E",X"04",X"03",X"00",X"01",X"00",
		X"C0",X"C0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"03",X"07",X"02",X"05",X"01",X"00",X"03",
		X"FE",X"F8",X"7C",X"B8",X"90",X"80",X"C1",X"1A",X"7F",X"FF",X"7F",X"3F",X"1F",X"D9",X"E2",X"F1",
		X"37",X"5F",X"BD",X"FF",X"5F",X"13",X"F0",X"FE",X"F9",X"BE",X"FF",X"E4",X"D9",X"F3",X"E7",X"37",
		X"F4",X"F0",X"E5",X"EA",X"DF",X"FC",X"FE",X"BB",X"FB",X"F4",X"E3",X"F3",X"FB",X"1F",X"3F",X"9F",
		X"07",X"EF",X"CD",X"A3",X"F3",X"F8",X"FC",X"F4",X"EE",X"D8",X"B8",X"B1",X"6D",X"7A",X"FD",X"FF",
		X"FB",X"BF",X"BB",X"FE",X"EF",X"FB",X"E9",X"FE",X"FF",X"ED",X"AA",X"FA",X"FA",X"EF",X"B3",X"FF",
		X"BF",X"F2",X"AF",X"EB",X"EE",X"BA",X"B9",X"BF",X"BA",X"FE",X"AB",X"EF",X"BF",X"FE",X"FB",X"AA",
		X"BF",X"EE",X"AA",X"EF",X"3B",X"9F",X"FA",X"B9",X"FA",X"7F",X"FA",X"E8",X"FA",X"BF",X"FF",X"FB",
		X"EE",X"EE",X"F3",X"BF",X"CE",X"AB",X"EE",X"BE",X"EF",X"CA",X"EE",X"FF",X"BE",X"FB",X"BF",X"FB",
		X"77",X"8D",X"87",X"CD",X"C6",X"E4",X"AC",X"F8",X"FC",X"E8",X"61",X"01",X"00",X"01",X"00",X"01",
		X"F0",X"D0",X"E0",X"E0",X"C0",X"80",X"40",X"80",X"01",X"03",X"03",X"03",X"00",X"03",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"36",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"80",X"FF",X"FF",X"C0",X"40",X"80",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"C0",X"40",X"80",X"FF",X"FF",X"C0",X"40",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"80",X"FF",X"FF",X"C0",X"40",X"80",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FC",X"FE",X"FE",X"E0",X"C0",X"C0",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",
		X"F0",X"E0",X"00",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F8",X"F0",X"00",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"C0",X"C0",X"D8",X"FC",X"FE",X"FE",X"E0",X"C0",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"C0",X"C0",X"C0",X"D0",X"F0",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"3F",X"3F",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"FF",X"C0",X"40",X"80",X"FF",X"FF",X"C0",X"40",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"80",X"FF",X"FF",X"C0",X"40",X"80",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"C0",X"40",X"80",X"FF",X"FF",X"C0",X"40",X"80",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"C0",X"40",X"80",X"FF",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"80",X"FF",X"FF",X"FF",X"FF",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"80",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"37",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"80",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"BF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"7F",X"7F",X"3F",X"3B",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"27",X"37",X"17",X"17",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"05",X"06",X"02",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"80",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"3F",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"10",X"A5",X"01",X"00",X"11",X"00",X"08",X"BF",X"52",X"29",X"06",X"F0",X"36",X"5C",X"23",
		X"A0",X"82",X"10",X"09",X"80",X"00",X"22",X"04",X"55",X"02",X"58",X"82",X"40",X"21",X"0A",X"26",
		X"FF",X"91",X"00",X"4A",X"91",X"00",X"10",X"50",X"FF",X"C4",X"4D",X"84",X"02",X"00",X"AC",X"00",
		X"81",X"72",X"1C",X"27",X"54",X"11",X"00",X"28",X"8C",X"08",X"80",X"A2",X"C4",X"74",X"9F",X"83",
		X"FF",X"30",X"0A",X"31",X"00",X"B8",X"15",X"80",X"FF",X"94",X"20",X"52",X"22",X"10",X"14",X"40",
		X"54",X"11",X"49",X"10",X"00",X"14",X"30",X"30",X"B1",X"10",X"40",X"90",X"0A",X"15",X"20",X"30",
		X"FF",X"99",X"52",X"04",X"1C",X"30",X"10",X"2A",X"28",X"14",X"00",X"44",X"40",X"08",X"00",X"20",
		X"14",X"82",X"08",X"92",X"70",X"19",X"10",X"90",X"80",X"24",X"04",X"90",X"50",X"08",X"00",X"62",
		X"00",X"02",X"00",X"0A",X"24",X"80",X"00",X"80",X"20",X"12",X"4A",X"28",X"8C",X"12",X"9A",X"43",
		X"01",X"08",X"12",X"00",X"A0",X"00",X"00",X"01",X"00",X"3A",X"80",X"10",X"53",X"02",X"29",X"0B",
		X"88",X"41",X"28",X"10",X"48",X"4D",X"02",X"08",X"84",X"04",X"80",X"00",X"0C",X"84",X"80",X"05",
		X"85",X"08",X"50",X"00",X"48",X"40",X"09",X"50",X"80",X"C0",X"A4",X"00",X"0C",X"04",X"0A",X"14",
		X"D0",X"30",X"5E",X"43",X"00",X"00",X"10",X"18",X"42",X"04",X"40",X"41",X"A8",X"70",X"08",X"4F",
		X"40",X"8A",X"10",X"14",X"21",X"B1",X"04",X"30",X"03",X"D0",X"80",X"42",X"24",X"40",X"40",X"21",
		X"14",X"10",X"00",X"90",X"04",X"D0",X"09",X"30",X"20",X"02",X"80",X"50",X"02",X"00",X"42",X"10",
		X"F0",X"72",X"34",X"77",X"09",X"12",X"91",X"30",X"10",X"08",X"80",X"02",X"80",X"18",X"00",X"48",
		X"08",X"00",X"20",X"00",X"44",X"80",X"00",X"02",X"80",X"02",X"44",X"20",X"52",X"00",X"09",X"83",
		X"00",X"00",X"00",X"08",X"20",X"00",X"82",X"80",X"00",X"44",X"00",X"02",X"0A",X"10",X"81",X"06",
		X"64",X"88",X"04",X"40",X"08",X"48",X"04",X"02",X"09",X"86",X"01",X"54",X"80",X"04",X"44",X"82",
		X"48",X"88",X"01",X"00",X"4A",X"04",X"49",X"80",X"A4",X"10",X"0D",X"84",X"94",X"20",X"04",X"84",
		X"90",X"4C",X"20",X"30",X"18",X"04",X"93",X"10",X"28",X"30",X"40",X"61",X"02",X"60",X"20",X"14",
		X"00",X"30",X"04",X"38",X"14",X"00",X"80",X"58",X"C0",X"60",X"22",X"14",X"A0",X"26",X"42",X"23",
		X"80",X"18",X"10",X"24",X"28",X"81",X"09",X"42",X"80",X"05",X"0A",X"1B",X"99",X"1B",X"D9",X"FC",
		X"01",X"02",X"29",X"07",X"84",X"04",X"23",X"01",X"7E",X"73",X"68",X"BC",X"4E",X"39",X"B4",X"DE",
		X"21",X"10",X"00",X"00",X"84",X"00",X"40",X"08",X"25",X"00",X"12",X"44",X"10",X"21",X"04",X"00",
		X"00",X"00",X"02",X"00",X"24",X"01",X"00",X"40",X"89",X"08",X"02",X"20",X"05",X"01",X"04",X"50",
		X"20",X"80",X"40",X"00",X"23",X"08",X"84",X"18",X"A5",X"00",X"14",X"82",X"00",X"84",X"04",X"00",
		X"02",X"20",X"00",X"20",X"00",X"C2",X"08",X"02",X"88",X"40",X"0D",X"00",X"80",X"46",X"01",X"01",
		X"00",X"98",X"52",X"20",X"00",X"92",X"18",X"09",X"B0",X"00",X"40",X"64",X"02",X"20",X"D0",X"08",
		X"14",X"10",X"26",X"41",X"90",X"08",X"10",X"08",X"24",X"22",X"60",X"11",X"80",X"E1",X"4A",X"A1",
		X"A4",X"0A",X"04",X"83",X"03",X"44",X"0E",X"03",X"F0",X"EE",X"3C",X"B0",X"EC",X"58",X"F6",X"BD",
		X"81",X"8E",X"81",X"43",X"34",X"0D",X"87",X"03",X"C7",X"EE",X"38",X"E0",X"DE",X"FC",X"C8",X"B7",
		X"02",X"00",X"80",X"10",X"00",X"00",X"80",X"00",X"12",X"00",X"00",X"00",X"21",X"10",X"04",X"01",
		X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"44",X"10",X"00",X"08",X"02",X"00",X"41",X"04",X"00",
		X"04",X"A4",X"00",X"02",X"11",X"04",X"00",X"20",X"48",X"22",X"84",X"90",X"04",X"11",X"94",X"08",
		X"0A",X"02",X"80",X"24",X"00",X"20",X"40",X"09",X"00",X"34",X"46",X"00",X"8A",X"54",X"89",X"61",
		X"90",X"B2",X"00",X"14",X"88",X"01",X"10",X"12",X"20",X"10",X"2E",X"A8",X"44",X"46",X"22",X"21",
		X"00",X"A0",X"90",X"0C",X"14",X"13",X"04",X"30",X"10",X"21",X"B4",X"01",X"21",X"40",X"22",X"24",
		X"84",X"03",X"01",X"24",X"71",X"8F",X"0B",X"CA",X"3C",X"38",X"8B",X"D6",X"EC",X"7D",X"AB",X"EE",
		X"07",X"43",X"31",X"0C",X"87",X"03",X"23",X"86",X"F0",X"D8",X"B7",X"F8",X"EC",X"D6",X"90",X"78",
		X"00",X"80",X"00",X"00",X"00",X"80",X"08",X"00",X"01",X"12",X"80",X"01",X"24",X"82",X"08",X"01",
		X"80",X"00",X"00",X"08",X"42",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"01",X"00",X"00",X"08",
		X"02",X"08",X"51",X"00",X"2A",X"02",X"00",X"90",X"64",X"02",X"14",X"20",X"86",X"08",X"81",X"14",
		X"00",X"02",X"40",X"0C",X"80",X"01",X"04",X"19",X"62",X"01",X"82",X"0A",X"84",X"10",X"05",X"92",
		X"15",X"A2",X"10",X"01",X"70",X"10",X"A0",X"01",X"A0",X"00",X"46",X"60",X"A0",X"08",X"31",X"20",
		X"14",X"40",X"10",X"00",X"00",X"11",X"72",X"08",X"28",X"12",X"24",X"80",X"2A",X"21",X"51",X"29",
		X"50",X"A1",X"00",X"50",X"89",X"21",X"02",X"50",X"F5",X"78",X"B8",X"74",X"8E",X"30",X"F3",X"EE",
		X"80",X"18",X"21",X"80",X"51",X"21",X"12",X"62",X"14",X"30",X"F0",X"E4",X"CA",X"BD",X"FA",X"A0",
		X"00",X"80",X"00",X"80",X"00",X"02",X"80",X"00",X"24",X"00",X"00",X"02",X"00",X"08",X"00",X"41",
		X"04",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"10",X"08",X"01",X"01",X"04",
		X"04",X"40",X"08",X"20",X"01",X"40",X"02",X"00",X"00",X"10",X"82",X"00",X"00",X"04",X"42",X"00",
		X"08",X"00",X"00",X"00",X"20",X"00",X"02",X"00",X"40",X"02",X"88",X"00",X"00",X"11",X"02",X"80",
		X"0A",X"90",X"01",X"80",X"50",X"00",X"00",X"22",X"23",X"10",X"22",X"04",X"48",X"A3",X"00",X"08",
		X"41",X"14",X"02",X"00",X"10",X"20",X"02",X"04",X"52",X"10",X"22",X"02",X"95",X"00",X"04",X"0A",
		X"86",X"A0",X"50",X"93",X"A7",X"01",X"00",X"56",X"FF",X"3E",X"FC",X"78",X"6B",X"B6",X"F8",X"7C",
		X"03",X"01",X"A0",X"40",X"10",X"04",X"11",X"A1",X"38",X"FB",X"D6",X"3C",X"78",X"FB",X"D7",X"7E",
		X"FB",X"FF",X"FB",X"FE",X"EF",X"FB",X"E9",X"FE",X"FF",X"ED",X"AA",X"FA",X"FE",X"EF",X"B7",X"FF",
		X"FF",X"F2",X"EF",X"EB",X"EE",X"FA",X"F9",X"FF",X"BA",X"FE",X"AF",X"EF",X"BB",X"FE",X"FB",X"AA",
		X"FF",X"EE",X"EA",X"EF",X"FB",X"FF",X"FA",X"F9",X"FA",X"7F",X"FA",X"EB",X"FA",X"BF",X"FF",X"FB",
		X"EE",X"EE",X"F3",X"FF",X"CE",X"EB",X"EE",X"FE",X"EF",X"CA",X"EE",X"FF",X"BE",X"FB",X"BF",X"FB",
		X"BB",X"FA",X"FE",X"EB",X"FF",X"FF",X"FA",X"EB",X"BC",X"EA",X"7F",X"BB",X"BF",X"BE",X"EF",X"EB",
		X"BD",X"FE",X"BE",X"EB",X"EE",X"FF",X"BA",X"EE",X"BA",X"FF",X"EF",X"EE",X"BB",X"AF",X"EA",X"FA",
		X"FB",X"BF",X"FB",X"FE",X"EF",X"FB",X"E9",X"FE",X"FF",X"ED",X"AA",X"FA",X"FA",X"EF",X"B3",X"FF",
		X"BF",X"F2",X"EF",X"EB",X"EE",X"FA",X"FB",X"E0",X"BA",X"FE",X"AB",X"EF",X"BF",X"FE",X"FB",X"00",
		X"AF",X"4C",X"6B",X"B6",X"9D",X"C7",X"CB",X"3C",X"2D",X"16",X"AC",X"1F",X"8E",X"E8",X"5E",X"2D",
		X"56",X"B8",X"1F",X"74",X"38",X"8E",X"37",X"09",X"98",X"3E",X"6B",X"9E",X"26",X"74",X"DB",X"1E",
		X"03",X"07",X"08",X"10",X"0F",X"47",X"0A",X"3C",X"FC",X"68",X"BE",X"9D",X"C2",X"26",X"7B",X"8E",
		X"5F",X"0E",X"11",X"BB",X"7E",X"2C",X"55",X"BF",X"04",X"EF",X"DA",X"2D",X"0E",X"F4",X"86",X"67",
		X"AF",X"76",X"B8",X"1D",X"47",X"61",X"0C",X"15",X"BE",X"C4",X"62",X"F9",X"62",X"86",X"FB",X"B6",
		X"88",X"6E",X"11",X"BB",X"7E",X"25",X"07",X"3B",X"45",X"E8",X"B2",X"3C",X"DA",X"F4",X"86",X"77",
		X"33",X"C4",X"6B",X"B6",X"9D",X"47",X"CB",X"3C",X"2D",X"16",X"AD",X"1F",X"8E",X"E8",X"5E",X"2D",
		X"56",X"B8",X"1F",X"74",X"38",X"8E",X"37",X"09",X"98",X"3E",X"6B",X"9E",X"26",X"74",X"DB",X"1E",
		X"29",X"D4",X"6B",X"B7",X"1E",X"35",X"EB",X"3F",X"3D",X"96",X"E4",X"28",X"1C",X"C0",X"78",X"C8",
		X"58",X"B6",X"1E",X"70",X"6C",X"FF",X"74",X"09",X"F2",X"30",X"C0",X"B0",X"7C",X"70",X"DF",X"16",
		X"00",X"00",X"00",X"02",X"02",X"08",X"07",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"60",X"B0",
		X"00",X"07",X"08",X"02",X"04",X"01",X"02",X"00",X"A0",X"10",X"50",X"A0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"24",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"05",X"38",X"02",X"05",X"02",X"08",X"10",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"04",X"1C",X"1C",X"1C",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"04",X"1C",X"1C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"EF",X"AF",X"AF",X"AF",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"2F",X"2F",X"2F",X"AF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"05",X"05",X"01",X"08",X"08",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"08",X"08",X"09",X"09",X"09",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",
		X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"FF",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"FF",
		X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",
		X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"FF",X"FF",X"CC",X"CC",X"FF",X"CC",X"CC",X"FF",X"FF",
		X"FF",X"7F",X"33",X"19",X"0C",X"06",X"03",X"01",X"FF",X"FF",X"33",X"99",X"CC",X"66",X"33",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"66",X"33",X"19",X"0C",X"06",X"03",X"01",
		X"FF",X"FF",X"33",X"99",X"CC",X"66",X"33",X"99",X"FF",X"FF",X"33",X"99",X"CC",X"66",X"33",X"99",
		X"CC",X"66",X"33",X"99",X"CC",X"66",X"33",X"FF",X"CC",X"66",X"33",X"99",X"CC",X"66",X"33",X"FF",
		X"FF",X"FF",X"33",X"FF",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"33",X"FF",X"CC",X"CC",X"CC",X"FF",
		X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",
		X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",
		X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",X"CC",X"CC",X"CC",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"92",X"92",X"92",X"92",X"92",X"FF",X"FF",X"FF",X"49",X"49",X"49",X"49",X"49",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"49",X"49",X"49",X"49",X"49",X"49",X"49",X"49",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"1F",X"00",X"11",X"0A",X"04",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"1F",X"04",X"55",X"5F",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"5F",X"55",X"55",X"10",X"1F",X"10",X"10",X"00",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"49",X"49",X"49",X"49",X"49",X"49",X"49",X"49",
		X"92",X"92",X"92",X"92",X"92",X"FF",X"FF",X"FF",X"49",X"49",X"49",X"49",X"49",X"FF",X"FF",X"FF",
		X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"47",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C0",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"00",X"00",X"7E",X"7E",X"7E",X"7F",X"7E",X"7E",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"7F",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"00",X"C4",X"C4",X"C4",X"C4",X"C0",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"47",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"B3",X"F3",X"B3",X"FF",X"B3",X"F3",X"F3",X"33",X"33",X"33",X"33",X"FF",X"33",X"33",X"33",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"FF",X"33",X"33",X"33",X"38",X"38",X"38",X"3F",X"F8",X"38",X"38",X"38",
		X"FF",X"33",X"33",X"33",X"FF",X"33",X"33",X"33",X"F8",X"38",X"38",X"3F",X"F8",X"38",X"38",X"38",
		X"FF",X"33",X"33",X"33",X"FF",X"33",X"33",X"33",X"F8",X"38",X"38",X"3F",X"F8",X"38",X"38",X"38",
		X"FF",X"B3",X"F3",X"B3",X"FF",X"B3",X"F3",X"B3",X"FF",X"33",X"33",X"33",X"FF",X"33",X"33",X"33",
		X"FF",X"B3",X"F3",X"B3",X"FF",X"B3",X"F3",X"B3",X"FF",X"33",X"33",X"33",X"FF",X"33",X"33",X"33",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"EF",X"8F",X"1F",X"3F",X"3F",X"7F",X"FF",X"7F",
		X"80",X"82",X"C1",X"83",X"81",X"00",X"8B",X"19",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"7C",X"79",X"73",X"BF",X"7F",X"3F",X"3F",X"FF",X"DF",X"DF",X"9F",
		X"4F",X"7E",X"78",X"74",X"60",X"78",X"70",X"64",X"9F",X"0F",X"1F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"1C",X"3A",X"3C",X"3C",X"7C",X"3E",X"3C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"3C",X"3E",X"3C",X"3C",X"34",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"3E",X"9E",X"8E",X"1F",X"FE",X"AF",X"9F",X"BF",
		X"00",X"00",X"00",X"00",X"43",X"C7",X"C7",X"CF",X"00",X"00",X"00",X"0C",X"1E",X"7E",X"FE",X"BE",
		X"CF",X"DF",X"47",X"43",X"40",X"21",X"47",X"7F",X"BE",X"BE",X"CE",X"9F",X"BE",X"BE",X"9E",X"9E",
		X"76",X"66",X"EF",X"EF",X"FF",X"FF",X"FF",X"FC",X"37",X"73",X"79",X"7C",X"7E",X"FE",X"FE",X"FC",
		X"F0",X"FC",X"FE",X"FF",X"FE",X"FF",X"7F",X"7F",X"00",X"0E",X"3F",X"7F",X"3F",X"1F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"02",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"06",X"02",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"0F",X"03",X"01",X"00",X"01",X"00",X"01",
		X"3F",X"9F",X"8E",X"9F",X"BF",X"BF",X"9F",X"FF",X"8E",X"1E",X"9E",X"5E",X"3E",X"BE",X"FE",X"FE",
		X"D7",X"DB",X"DB",X"F3",X"DB",X"B3",X"CB",X"DB",X"FC",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7C",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"2F",X"37",X"1F",X"B7",X"B7",X"3F",X"9B",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"00",X"00",X"03",X"BF",X"1F",X"8E",X"80",X"00",X"2C",X"FE",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0B",X"0F",X"1F",X"3F",X"3F",X"03",X"FC",X"F0",
		X"01",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"0E",X"0E",X"04",X"00",X"00",X"00",X"00",X"01",
		X"FE",X"FF",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"02",X"EC",X"FE",X"3F",X"1F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"30",X"30",X"38",X"3C",X"38",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",
		X"30",X"30",X"38",X"38",X"BD",X"FD",X"FD",X"FD",X"78",X"78",X"78",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"3F",X"3F",X"5F",X"5F",X"FF",
		X"00",X"01",X"01",X"03",X"03",X"07",X"1F",X"7F",X"EF",X"EF",X"FF",X"FF",X"FF",X"EF",X"FF",X"E7",
		X"3F",X"7F",X"71",X"70",X"60",X"28",X"2E",X"7D",X"FE",X"FE",X"FF",X"0F",X"03",X"01",X"00",X"00",
		X"7D",X"6F",X"67",X"73",X"73",X"7D",X"7C",X"7E",X"C1",X"C1",X"E1",X"C1",X"E1",X"F9",X"F9",X"FC",
		X"38",X"30",X"30",X"30",X"20",X"20",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"0D",X"1D",X"0D",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"FB",X"FF",X"7F",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"20",X"10",X"08",
		X"F2",X"F1",X"F8",X"FE",X"FE",X"F7",X"F7",X"FF",X"07",X"07",X"0F",X"0E",X"2E",X"2E",X"7F",X"7E",
		X"FF",X"FB",X"FB",X"FD",X"FF",X"05",X"06",X"06",X"FF",X"FF",X"FF",X"FF",X"1F",X"4F",X"AB",X"FF",
		X"FD",X"FD",X"FE",X"FE",X"FE",X"FF",X"FF",X"7F",X"F8",X"F8",X"F8",X"F8",X"F0",X"70",X"70",X"60",
		X"7E",X"78",X"E0",X"80",X"C0",X"80",X"C0",X"80",X"18",X"70",X"80",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"07",X"3F",X"7F",X"3F",X"01",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"7F",X"FF",X"FF",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"77",X"13",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"E7",X"E7",X"E3",X"E1",X"E1",
		X"FF",X"3F",X"0D",X"81",X"41",X"47",X"CF",X"CF",X"E1",X"E0",X"F3",X"A7",X"33",X"3F",X"7F",X"FF",
		X"76",X"66",X"62",X"63",X"71",X"78",X"7F",X"7F",X"1C",X"1C",X"08",X"80",X"20",X"28",X"F8",X"F0",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"F8",X"F8",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"16",X"1E",X"0A",X"15",X"0B",X"1F",X"2B",X"1F",
		X"02",X"07",X"0F",X"0F",X"0F",X"3F",X"3F",X"3F",X"17",X"2F",X"1B",X"2F",X"3F",X"3F",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"03",X"C1",X"70",X"1C",X"07",X"01",X"00",X"61",X"01",X"F0",X"00",X"00",X"00",X"80",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"F0",X"1E",X"03",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"81",X"E1",X"1D",X"03",
		X"E9",X"FF",X"EF",X"CE",X"C8",X"C0",X"C0",X"C0",X"FF",X"F9",X"80",X"00",X"00",X"00",X"00",X"02",
		X"C0",X"C0",X"80",X"81",X"82",X"1D",X"52",X"6A",X"0F",X"04",X"6A",X"4A",X"15",X"5A",X"AD",X"DA",
		X"DF",X"EF",X"7F",X"1F",X"0F",X"07",X"03",X"01",X"FD",X"FB",X"FF",X"FD",X"FD",X"FB",X"FF",X"FD",
		X"C1",X"F8",X"5E",X"A7",X"2B",X"55",X"6D",X"92",X"FF",X"FF",X"FB",X"FE",X"FE",X"FC",X"FD",X"FF",
		X"FC",X"FE",X"FE",X"FF",X"F6",X"FD",X"F4",X"F4",X"DF",X"DF",X"DF",X"DF",X"BF",X"9F",X"BF",X"BF",
		X"F0",X"F2",X"F5",X"E8",X"E2",X"F3",X"7B",X"7B",X"BF",X"9F",X"9F",X"5F",X"EF",X"6E",X"6E",X"B6",
		X"9F",X"9F",X"8F",X"8F",X"BF",X"9F",X"BF",X"9F",X"F0",X"F0",X"F8",X"F4",X"F0",X"F8",X"FC",X"F8",
		X"9F",X"BF",X"BE",X"9E",X"82",X"FF",X"FE",X"FE",X"E8",X"F0",X"F0",X"73",X"E7",X"F7",X"F3",X"FB",
		X"37",X"6E",X"6E",X"7C",X"5C",X"FE",X"FE",X"FD",X"FF",X"7F",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",
		X"F9",X"F9",X"FB",X"F9",X"FB",X"F3",X"F7",X"EF",X"FD",X"FF",X"EF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"14",X"03",X"4A",
		X"00",X"01",X"01",X"03",X"09",X"00",X"05",X"50",X"22",X"28",X"22",X"64",X"20",X"89",X"A2",X"CA",
		X"85",X"10",X"44",X"A5",X"0C",X"44",X"91",X"00",X"3F",X"7F",X"1F",X"1F",X"4F",X"57",X"63",X"41",
		X"24",X"84",X"84",X"A9",X"04",X"A0",X"62",X"24",X"42",X"14",X"84",X"05",X"08",X"44",X"C4",X"69",
		X"7B",X"7B",X"79",X"BD",X"FD",X"DF",X"DF",X"C3",X"36",X"17",X"0E",X"9B",X"03",X"87",X"87",X"83",
		X"F7",X"73",X"BB",X"3B",X"BB",X"1D",X"4F",X"97",X"01",X"80",X"D0",X"F6",X"F7",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"FF",X"87",X"E7",X"E7",X"E7",X"F8",X"F8",X"F8",X"FC",X"FE",X"FC",X"F8",X"E1",
		X"F3",X"F9",X"68",X"84",X"C0",X"F0",X"E0",X"FF",X"E3",X"CF",X"87",X"C3",X"49",X"26",X"27",X"83",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"04",X"06",X"10",X"15",
		X"00",X"00",X"01",X"05",X"05",X"05",X"15",X"56",X"54",X"5E",X"14",X"44",X"54",X"72",X"55",X"55",
		X"52",X"85",X"52",X"22",X"4B",X"C4",X"40",X"54",X"50",X"12",X"15",X"80",X"15",X"98",X"25",X"92",
		X"24",X"41",X"44",X"82",X"54",X"44",X"44",X"8A",X"80",X"0C",X"45",X"94",X"90",X"91",X"44",X"81",
		X"91",X"07",X"63",X"07",X"13",X"A3",X"27",X"47",X"74",X"F4",X"F5",X"3B",X"9F",X"99",X"98",X"D8",
		X"47",X"93",X"23",X"8B",X"23",X"21",X"2D",X"43",X"DE",X"FE",X"DE",X"FC",X"FC",X"FC",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"F8",X"FE",X"FF",X"FF",X"FF",X"43",X"33",X"38",X"3F",X"3F",X"3F",X"07",X"0F",
		X"FC",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"9F",X"9F",X"87",X"9D",X"85",X"8D",X"BD",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"05",X"0D",X"15",
		X"00",X"00",X"00",X"05",X"0C",X"1E",X"3E",X"3F",X"11",X"4C",X"05",X"C7",X"61",X"11",X"54",X"D5",
		X"51",X"5D",X"55",X"75",X"75",X"56",X"55",X"91",X"55",X"35",X"55",X"55",X"57",X"55",X"54",X"5D",
		X"55",X"45",X"0D",X"15",X"55",X"51",X"56",X"75",X"15",X"50",X"B5",X"C5",X"47",X"55",X"55",X"5D",
		X"0D",X"51",X"01",X"09",X"83",X"21",X"29",X"20",X"FF",X"DF",X"DF",X"DF",X"FF",X"FF",X"EF",X"EE",
		X"42",X"92",X"06",X"24",X"00",X"88",X"20",X"A2",X"E4",X"69",X"6C",X"7E",X"76",X"B6",X"B7",X"17",
		X"F3",X"E3",X"C3",X"E3",X"E3",X"83",X"01",X"01",X"85",X"83",X"81",X"83",X"87",X"9F",X"C3",X"C1",
		X"00",X"90",X"C0",X"C0",X"F4",X"F0",X"F0",X"DC",X"E1",X"E1",X"FD",X"F9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"5F",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3B",X"7B",X"DB",X"D9",X"FC",X"3E",X"3E",X"5A",X"DA",X"DA",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"C6",X"D5",X"CD",X"C9",X"D4",X"C5",X"CA",X"CE",
		X"EF",X"DF",X"5F",X"7F",X"DF",X"DD",X"DD",X"DC",X"85",X"89",X"85",X"8E",X"8D",X"C5",X"E1",X"F1",
		X"0A",X"41",X"53",X"02",X"24",X"82",X"02",X"52",X"27",X"17",X"11",X"58",X"01",X"94",X"20",X"02",
		X"40",X"88",X"42",X"62",X"40",X"08",X"90",X"42",X"90",X"31",X"10",X"90",X"16",X"03",X"42",X"12",
		X"DF",X"5F",X"50",X"40",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"C3",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"05",X"0D",X"15",X"37",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"25",X"3D",X"1D",X"0D",X"07",X"03",X"01",
		X"FB",X"FB",X"7B",X"7D",X"5D",X"59",X"5B",X"DB",X"B7",X"BF",X"B7",X"B7",X"BD",X"BD",X"DF",X"DF",
		X"FB",X"DA",X"DE",X"FA",X"EB",X"BB",X"AF",X"AB",X"DE",X"DE",X"DD",X"FD",X"FD",X"7D",X"7F",X"7F",
		X"DD",X"ED",X"DD",X"D9",X"DB",X"53",X"57",X"5E",X"F5",X"F1",X"E1",X"FA",X"F5",X"F3",X"F0",X"F1",
		X"7E",X"5F",X"4F",X"5B",X"5D",X"DE",X"DD",X"FB",X"F9",X"78",X"5C",X"7D",X"F4",X"FD",X"F1",X"71",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EB",X"7F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"6F",X"6F",X"6B",X"6B",X"EE",X"FE",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"D7",X"D6",X"D6",X"DE",X"FF",X"F7",X"F7",X"D5",X"59",X"79",X"79",X"E1",X"C6",X"C5",X"C1",X"40",
		X"C4",X"C4",X"C1",X"C4",X"C1",X"C9",X"41",X"01",X"51",X"19",X"59",X"15",X"74",X"40",X"16",X"54",
		X"1C",X"0D",X"03",X"01",X"00",X"00",X"00",X"00",X"D5",X"54",X"13",X"7D",X"D5",X"45",X"34",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"51",X"1D",X"75",X"D5",X"56",X"57",X"55",X"55",X"65",X"53",X"17",X"13",X"5B",X"57",X"57",X"D7",
		X"65",X"11",X"15",X"55",X"15",X"14",X"0D",X"01",X"46",X"5D",X"54",X"55",X"B8",X"58",X"58",X"52",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B8",X"54",X"48",X"58",X"05",X"08",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"82",X"2A",X"02",X"49",X"9A",X"21",X"22",X"21",X"08",X"88",X"1B",X"48",X"4C",X"49",X"28",
		X"AA",X"02",X"22",X"08",X"02",X"04",X"01",X"00",X"40",X"08",X"B0",X"62",X"28",X"28",X"88",X"26",
		X"59",X"49",X"7B",X"68",X"C8",X"48",X"E0",X"C4",X"FE",X"FE",X"7E",X"FF",X"7E",X"7F",X"3E",X"0F",
		X"A5",X"C9",X"DD",X"DF",X"CF",X"87",X"8F",X"DF",X"06",X"3F",X"FF",X"FD",X"FC",X"FE",X"7E",X"FE",
		X"DD",X"D9",X"D9",X"D8",X"DC",X"DC",X"D8",X"CC",X"FF",X"FF",X"DF",X"FF",X"FE",X"FE",X"DE",X"EE",
		X"88",X"9C",X"C8",X"CC",X"E4",X"E4",X"E0",X"E8",X"E5",X"FC",X"4E",X"5C",X"EE",X"5E",X"CE",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"30",X"30",X"3B",X"1B",X"FD",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"28",X"FF",X"FF",X"FF",X"FF",X"00",X"40",X"30",X"3B",X"FD",X"FD",X"FD",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"E0",X"FC",X"E7",X"FF",X"E6",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",
		X"01",X"00",X"03",X"87",X"0F",X"3F",X"FF",X"FF",X"F0",X"FC",X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"04",X"03",X"3F",X"FF",X"FF",X"FF",X"7E",X"1C",X"80",X"FF",X"3F",X"FF",X"3F",X"F8",X"8C",X"8F",
		X"04",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"8F",X"FF",X"FF",X"8F",X"8F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"F8",X"F0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F0",X"F8",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F8",X"04",X"04",X"0F",
		X"FE",X"FF",X"FF",X"F7",X"FB",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"00",X"40",X"F0",X"FA",X"FE",X"00",X"3F",X"FF",X"00",X"0A",X"77",X"BF",X"FC",X"01",X"FF",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"FF",
		X"00",X"00",X"80",X"60",X"00",X"E0",X"98",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FB",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"D0",X"F4",X"FB",X"FF",X"FF",X"FF",
		X"20",X"FF",X"20",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",X"00",X"FD",X"FD",X"FC",X"FC",X"F8",X"F8",X"F0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"03",X"0F",X"0F",X"03",X"23",X"2F",X"FD",X"FD",X"FD",X"FC",X"FC",X"FC",X"F8",X"F0",
		X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"FF",X"E7",X"C0",X"40",X"40",X"40",X"40",X"C0",
		X"01",X"07",X"1F",X"3F",X"7F",X"FF",X"FF",X"FE",X"80",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0E",X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"03",X"0E",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F8",
		X"FF",X"FF",X"00",X"00",X"00",X"FC",X"04",X"04",X"FF",X"FF",X"8F",X"8F",X"FF",X"07",X"07",X"07",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"E0",X"E0",X"FF",X"7F",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",
		X"55",X"55",X"55",X"55",X"D5",X"D5",X"7F",X"7F",X"57",X"57",X"57",X"57",X"57",X"56",X"FE",X"FE",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FB",X"07",X"1F",X"1F",X"07",X"07",X"1F",X"DF",
		X"8F",X"8F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"FF",X"F8",X"C0",X"C6",X"C6",X"06",X"3E",X"3C",
		X"D0",X"10",X"50",X"10",X"50",X"10",X"50",X"10",X"01",X"03",X"02",X"03",X"00",X"03",X"02",X"03",
		X"50",X"1F",X"D0",X"50",X"D0",X"50",X"D0",X"41",X"00",X"FF",X"00",X"00",X"00",X"7C",X"7F",X"FF",
		X"00",X"F7",X"17",X"F7",X"07",X"F7",X"17",X"F7",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"FF",X"07",X"07",X"07",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F0",X"F8",X"FC",X"F8",X"F8",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FC",X"F8",X"FC",X"FC",X"FE",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0F",X"0F",X"1F",X"7F",X"3F",X"8F",X"E3",
		X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FE",X"FF",X"7F",X"1F",X"0F",X"03",X"00",
		X"FC",X"F8",X"F0",X"E0",X"C0",X"E0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"7E",X"3F",X"8F",X"E3",X"F9",X"FC",X"FE",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"78",
		X"3F",X"38",X"38",X"7F",X"70",X"70",X"7F",X"38",X"FC",X"7C",X"7C",X"FC",X"7C",X"7C",X"FC",X"7C",
		X"38",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"7C",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0F",X"0E",X"2E",X"6E",X"EE",X"EE",X"EE",X"EF",X"EF",
		X"1F",X"3F",X"7F",X"E1",X"E1",X"FF",X"E1",X"E1",X"EF",X"EE",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",
		X"00",X"01",X"11",X"01",X"0F",X"8F",X"0E",X"7C",X"38",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"0E",X"EF",X"6F",X"61",X"1D",X"0D",X"8C",X"8F",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"38",X"BC",
		X"FE",X"FF",X"00",X"01",X"00",X"01",X"00",X"01",X"07",X"8F",X"3F",X"BC",X"18",X"B8",X"38",X"98",
		X"00",X"01",X"00",X"01",X"00",X"01",X"FE",X"FF",X"38",X"B8",X"18",X"BC",X"3F",X"8F",X"07",X"FF",
		X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"FF",X"3F",X"07",X"00",X"02",X"02",X"3F",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"0E",X"00",X"00",X"03",X"FF",X"0F",X"03",X"00",
		X"FF",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"07",X"3F",X"FF",X"FF",X"FC",X"FC",X"38",X"1F",X"E0",X"F7",X"F7",X"F7",X"00",X"00",X"00",
		X"00",X"F3",X"E7",X"8F",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FC",X"F8",X"F1",X"07",X"3F",X"1F",
		X"00",X"FF",X"FE",X"F8",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"1F",X"01",X"3E",X"7E",X"FD",
		X"F1",X"03",X"F3",X"F7",X"F7",X"F7",X"F7",X"F3",X"FB",X"F7",X"EF",X"DF",X"DE",X"FC",X"F9",X"F3",
		X"00",X"00",X"00",X"3F",X"21",X"00",X"30",X"30",X"0F",X"00",X"00",X"7C",X"44",X"00",X"60",X"60",
		X"30",X"B0",X"B0",X"30",X"30",X"FF",X"FF",X"0E",X"60",X"60",X"60",X"60",X"60",X"FF",X"FF",X"1C",
		X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"BF",X"DF",X"BE",X"86",X"F6",X"F6",X"F0",X"FF",X"FF",X"FF",
		X"DF",X"CF",X"CF",X"CF",X"CF",X"F7",X"F7",X"37",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C4",X"84",
		X"50",X"D0",X"50",X"D0",X"50",X"DF",X"10",X"50",X"7F",X"7D",X"00",X"00",X"00",X"FF",X"00",X"03",
		X"10",X"50",X"10",X"50",X"10",X"50",X"00",X"7F",X"02",X"03",X"00",X"03",X"02",X"00",X"01",X"FF",
		X"FF",X"FF",X"07",X"07",X"07",X"FF",X"05",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"B5",X"20",X"00",
		X"14",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"F4",X"F8",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"81",X"80",X"80",X"80",X"00",X"00",X"00",X"E7",X"C6",X"C6",X"63",X"31",X"38",X"3C",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0C",X"0C",X"0E",X"0E",X"FF",X"7F",X"7F",X"1C",X"18",X"18",X"1C",X"1C",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"37",X"36",X"35",X"37",X"37",X"F7",X"F7",X"FF",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7B",X"3B",X"07",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"E5",X"E4",X"3F",X"36",X"F8",X"F0",X"C0",X"30",X"00",X"00",
		X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"1C",X"78",X"F4",X"F8",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
