library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity time_pilot_char_grphx is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of time_pilot_char_grphx is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",X"E1",X"F0",X"F0",X"E1",X"C3",X"87",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"78",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"F0",X"E1",X"C3",X"87",
		X"00",X"00",X"00",X"FF",X"FF",X"11",X"11",X"11",X"00",X"00",X"00",X"FF",X"FF",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"99",X"99",X"66",X"00",X"00",X"00",X"10",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"31",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"EE",X"77",X"99",X"99",X"66",X"00",X"00",
		X"00",X"00",X"66",X"F9",X"F9",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"CC",X"EE",X"77",X"F9",X"F9",X"66",X"00",X"00",
		X"11",X"32",X"74",X"74",X"75",X"32",X"01",X"00",X"CC",X"E2",X"E5",X"E9",X"E1",X"C2",X"0C",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"11",X"11",X"11",X"FF",X"FF",X"11",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"11",X"11",X"11",X"FF",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"88",X"88",X"88",X"FF",X"FF",X"88",X"88",X"88",
		X"00",X"00",X"00",X"FF",X"FF",X"11",X"11",X"11",X"00",X"00",X"00",X"FF",X"FF",X"88",X"88",X"88",
		X"11",X"11",X"11",X"FF",X"FF",X"11",X"11",X"11",X"88",X"88",X"88",X"FF",X"FF",X"88",X"88",X"88",
		X"00",X"00",X"00",X"FF",X"FF",X"11",X"11",X"11",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",
		X"11",X"11",X"11",X"FF",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"FF",X"FF",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"F0",X"D2",X"A0",X"E1",X"B0",X"E2",X"70",X"90",X"42",X"02",X"7F",X"B7",X"74",X"59",X"20",
		X"00",X"49",X"A4",X"CE",X"AA",X"0C",X"B4",X"50",X"A0",X"F0",X"70",X"B8",X"70",X"D0",X"F8",X"60",
		X"70",X"F0",X"D0",X"F2",X"A4",X"93",X"35",X"7B",X"E0",X"70",X"F0",X"B2",X"58",X"24",X"82",X"ED",
		X"37",X"73",X"39",X"46",X"90",X"F2",X"F0",X"70",X"CF",X"CE",X"89",X"A8",X"42",X"F8",X"F0",X"E0",
		X"00",X"01",X"03",X"F7",X"F7",X"01",X"03",X"00",X"08",X"0C",X"0E",X"FF",X"FF",X"0C",X"0E",X"00",
		X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"80",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"80",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"A4",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"A4",
		X"70",X"F0",X"F0",X"FF",X"F0",X"70",X"70",X"77",X"E0",X"F0",X"F0",X"FF",X"F0",X"E0",X"E0",X"EE",
		X"70",X"70",X"70",X"70",X"F0",X"0F",X"F0",X"70",X"E0",X"E0",X"E0",X"E0",X"F0",X"0F",X"F0",X"E0",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"1E",X"3C",X"78",X"F0",X"F0",X"78",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",
		X"1E",X"3C",X"78",X"F0",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",X"E1",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"03",X"07",X"3F",X"3F",X"07",X"03",X"00",X"00",X"10",X"38",X"FC",X"FC",X"38",X"10",
		X"70",X"F0",X"F7",X"FF",X"FF",X"FF",X"FF",X"F7",X"80",X"C0",X"E8",X"FC",X"FC",X"FC",X"FC",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"3F",X"3F",X"37",X"33",X"70",X"F0",X"00",X"08",X"0C",X"0C",X"08",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"30",X"10",X"00",X"00",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"70",X"E8",X"FC",X"FC",X"FC",X"FC",X"EC",X"C8",X"80",
		X"33",X"33",X"33",X"37",X"3F",X"3F",X"07",X"03",X"00",X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",
		X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F0",X"C3",X"E1",X"87",X"F0",X"87",X"A5",X"A5",
		X"F0",X"3C",X"F0",X"F0",X"F0",X"B4",X"B4",X"3C",X"F7",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"FC",X"FC",X"FC",X"F8",X"F0",X"F0",X"F0",X"88",X"F0",X"F0",X"F0",X"96",X"A5",X"B4",X"F0",X"00",
		X"F0",X"B4",X"F0",X"F0",X"3C",X"F0",X"F0",X"00",X"F3",X"F3",X"F3",X"F1",X"F0",X"F0",X"F0",X"11",
		X"07",X"03",X"01",X"30",X"71",X"71",X"30",X"10",X"0F",X"0F",X"0F",X"0F",X"CF",X"CB",X"C1",X"80",
		X"00",X"30",X"70",X"F3",X"E3",X"43",X"07",X"07",X"00",X"00",X"80",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"0C",X"00",X"08",X"0C",X"2C",X"7C",X"FC",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"EE",X"CC",X"88",X"B8",X"F8",X"F0",X"F0",X"F0",
		X"77",X"33",X"11",X"D1",X"F1",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",
		X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"0C",X"0C",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"30",X"43",X"87",X"87",X"87",X"87",X"43",X"30",X"C0",X"2C",X"1E",X"1E",X"1E",X"1E",X"2C",X"C0",
		X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"78",X"78",X"78",X"78",X"78",X"78",X"0F",X"0F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"0F",
		X"0F",X"08",X"08",X"78",X"78",X"78",X"78",X"0F",X"0F",X"01",X"01",X"E1",X"E1",X"E1",X"E1",X"0F",
		X"0F",X"08",X"08",X"08",X"78",X"78",X"78",X"0F",X"0F",X"01",X"01",X"01",X"E1",X"E1",X"E1",X"0F",
		X"0F",X"08",X"08",X"08",X"08",X"08",X"78",X"0F",X"0F",X"01",X"01",X"01",X"01",X"01",X"E1",X"0F",
		X"00",X"10",X"54",X"12",X"F1",X"12",X"54",X"10",X"00",X"00",X"44",X"08",X"E0",X"08",X"44",X"00",
		X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"12",X"34",X"79",X"79",X"34",X"12",X"01",X"08",X"84",X"C2",X"E9",X"E9",X"C2",X"84",X"08",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0E",X"0E",X"E0",X"0E",X"0E",X"0F",X"0F",X"0F",X"44",X"66",X"77",X"66",X"44",X"0F",
		X"0F",X"0F",X"66",X"66",X"66",X"66",X"66",X"0F",X"0F",X"0F",X"07",X"07",X"70",X"07",X"07",X"0F",
		X"0C",X"3F",X"3F",X"0C",X"0C",X"0F",X"0F",X"0F",X"01",X"EF",X"EF",X"01",X"01",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0C",X"0C",X"3F",X"1D",X"0C",X"87",X"87",X"87",X"01",X"01",X"EF",X"CD",X"89",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"87",X"87",X"87",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"99",X"99",X"66",X"00",X"00",X"00",X"10",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"31",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"EE",X"77",X"99",X"99",X"66",X"00",X"00",
		X"00",X"00",X"66",X"F9",X"F9",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"CC",X"EE",X"77",X"F9",X"F9",X"66",X"00",X"00",
		X"11",X"32",X"74",X"74",X"75",X"32",X"01",X"00",X"CC",X"E2",X"E5",X"E9",X"E1",X"C2",X"0C",X"00",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"F0",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"F0",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"87",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"87",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"87",X"87",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0E",X"E0",X"0E",X"0F",X"0F",X"0F",X"2F",X"03",X"41",X"B4",X"12",X"A3",X"0F",
		X"0F",X"0F",X"4C",X"04",X"A0",X"0A",X"4C",X"0F",X"0F",X"0F",X"0F",X"07",X"70",X"07",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"1C",X"0F",X"1D",X"87",X"87",X"87",X"03",X"41",X"05",X"83",X"C3",
		X"0E",X"1D",X"0F",X"1C",X"0E",X"0F",X"0F",X"0F",X"C3",X"85",X"C3",X"41",X"03",X"87",X"87",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0E",X"E0",X"0E",X"0F",X"0F",X"0F",X"0F",X"45",X"44",X"44",X"44",X"45",X"0F",
		X"0F",X"0F",X"0C",X"88",X"88",X"88",X"0C",X"0F",X"0F",X"0F",X"0F",X"07",X"70",X"07",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"3F",X"0C",X"0E",X"87",X"87",X"87",X"03",X"01",X"EF",X"01",X"03",
		X"1F",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",X"0F",X"CF",X"03",X"01",X"01",X"03",X"87",X"87",X"87",
		X"0F",X"0F",X"0E",X"0E",X"E0",X"0E",X"0E",X"0F",X"0F",X"0F",X"66",X"66",X"66",X"66",X"66",X"0F",
		X"0F",X"0F",X"22",X"66",X"EE",X"66",X"22",X"0F",X"0F",X"0F",X"07",X"07",X"70",X"07",X"07",X"0F",
		X"0F",X"0F",X"0F",X"0C",X"0C",X"3F",X"3F",X"0C",X"87",X"87",X"87",X"01",X"01",X"EF",X"EF",X"01",
		X"0C",X"1D",X"3F",X"0C",X"0C",X"0F",X"0F",X"0F",X"89",X"CD",X"EF",X"01",X"01",X"87",X"87",X"87",
		X"00",X"00",X"03",X"07",X"3F",X"3F",X"07",X"03",X"00",X"00",X"10",X"38",X"FC",X"FC",X"38",X"10",
		X"0F",X"3C",X"0F",X"2D",X"E1",X"2D",X"0F",X"3C",X"0F",X"C3",X"4B",X"4B",X"78",X"4B",X"4B",X"C3",
		X"0F",X"0F",X"0F",X"0F",X"2D",X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",X"A5",X"B4",X"A5",X"2D",X"0F",
		X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"3F",X"3F",X"37",X"33",X"70",X"F0",X"00",X"08",X"0C",X"0C",X"08",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"30",X"10",X"00",X"00",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"70",X"E8",X"FC",X"FC",X"FC",X"FC",X"EC",X"C8",X"80",
		X"33",X"33",X"33",X"37",X"3F",X"3F",X"07",X"03",X"00",X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",
		X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F0",X"C3",X"E1",X"87",X"F0",X"87",X"A5",X"A5",
		X"F0",X"3C",X"F0",X"F0",X"F0",X"B4",X"B4",X"3C",X"F7",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"FC",X"FC",X"FC",X"F8",X"F0",X"F0",X"F0",X"88",X"F0",X"F0",X"F0",X"96",X"A5",X"B4",X"F0",X"00",
		X"F0",X"B4",X"F0",X"F0",X"3C",X"F0",X"F0",X"00",X"F3",X"F3",X"F3",X"F1",X"F0",X"F0",X"F0",X"11",
		X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"25",X"21",X"01",X"08",X"48",X"86",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"2D",X"2D",X"2D",
		X"0F",X"0F",X"0F",X"F0",X"07",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"EE",X"CC",X"88",X"B8",X"F8",X"F0",X"F0",X"F0",
		X"77",X"33",X"11",X"D1",X"F1",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",
		X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CE",X"9C",X"99",X"98",X"99",X"99",X"C9",X"FF",X"37",X"93",X"19",X"11",X"F9",X"F9",X"19",X"FF",
		X"8C",X"99",X"99",X"89",X"99",X"99",X"8C",X"FF",X"33",X"99",X"9F",X"3F",X"9F",X"99",X"33",X"FF",
		X"88",X"99",X"99",X"98",X"99",X"99",X"88",X"FF",X"71",X"3F",X"9F",X"97",X"9F",X"3F",X"71",X"FF",
		X"8C",X"99",X"99",X"89",X"99",X"99",X"9C",X"FF",X"13",X"F9",X"FF",X"71",X"F9",X"F9",X"F3",X"FF",
		X"9C",X"9E",X"9E",X"8E",X"9E",X"9E",X"9C",X"FF",X"93",X"97",X"97",X"17",X"97",X"97",X"93",X"FF",
		X"E9",X"F9",X"F8",X"F8",X"F8",X"99",X"C9",X"FF",X"19",X"33",X"37",X"3F",X"37",X"33",X"79",X"FF",
		X"99",X"98",X"98",X"99",X"99",X"99",X"89",X"FF",X"FC",X"F8",X"F0",X"F4",X"FC",X"FC",X"1C",X"FF",
		X"9C",X"89",X"89",X"89",X"99",X"99",X"9C",X"FF",X"93",X"99",X"19",X"19",X"19",X"99",X"93",X"FF",
		X"8C",X"99",X"99",X"89",X"99",X"9C",X"9F",X"FF",X"33",X"99",X"99",X"39",X"F9",X"F3",X"F1",X"FF",
		X"8C",X"99",X"99",X"8C",X"8F",X"99",X"9C",X"FF",X"33",X"99",X"9F",X"33",X"79",X"39",X"93",X"FF",
		X"89",X"E9",X"E9",X"E9",X"E9",X"E9",X"EC",X"FF",X"19",X"79",X"79",X"79",X"79",X"79",X"73",X"FF",
		X"99",X"99",X"99",X"99",X"98",X"C8",X"E9",X"FF",X"9C",X"9C",X"9C",X"94",X"90",X"38",X"7C",X"FF",
		X"99",X"99",X"C9",X"EC",X"CE",X"9E",X"9E",X"FF",X"99",X"99",X"39",X"73",X"37",X"97",X"97",X"FF",
		X"8C",X"FC",X"FC",X"EC",X"CC",X"9C",X"8C",X"FF",X"13",X"9F",X"3F",X"7F",X"FF",X"FF",X"13",X"FF",
		X"FC",X"EF",X"CF",X"0F",X"CF",X"9F",X"0C",X"FF",X"13",X"F3",X"F3",X"13",X"F3",X"F3",X"03",X"FF",
		X"FF",X"EE",X"CC",X"88",X"E8",X"EC",X"EE",X"EF",X"FF",X"7F",X"3F",X"10",X"70",X"7F",X"7F",X"7F",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FF",X"F7",X"F7",X"F7",X"F7",X"FF",X"FF",X"F7",X"FF",
		X"99",X"99",X"90",X"F9",X"F0",X"F9",X"F9",X"FF",X"99",X"99",X"90",X"F9",X"F0",X"F9",X"F9",X"FF",
		X"E9",X"C9",X"9F",X"CE",X"FC",X"89",X"EB",X"FF",X"7D",X"19",X"F3",X"37",X"9F",X"39",X"79",X"FF",
		X"CF",X"9F",X"CE",X"CF",X"9F",X"9F",X"CF",X"FF",X"39",X"93",X"37",X"7F",X"8F",X"9F",X"0F",X"FF",
		X"FC",X"EE",X"CF",X"CF",X"CF",X"EE",X"FC",X"FF",X"3F",X"77",X"F3",X"F3",X"F3",X"77",X"3F",X"FF",
		X"FF",X"9E",X"CE",X"08",X"CE",X"9E",X"FF",X"FF",X"FF",X"97",X"37",X"01",X"37",X"97",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F8",X"FF",X"EF",X"EF",X"CF",X"FF",X"FF",X"FF",X"F1",X"FF",X"7F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"EC",X"E9",X"FF",X"FF",X"FC",X"F9",X"F3",X"F7",X"7F",X"7F",X"FF",
		X"CE",X"9E",X"9C",X"8E",X"9E",X"9E",X"C8",X"FF",X"37",X"97",X"17",X"97",X"97",X"97",X"31",X"FF",
		X"CC",X"99",X"FF",X"FE",X"CF",X"99",X"8C",X"FF",X"33",X"99",X"99",X"33",X"F9",X"F9",X"13",X"FF",
		X"F8",X"F9",X"E8",X"9F",X"8F",X"F9",X"FC",X"FF",X"91",X"1F",X"13",X"99",X"09",X"99",X"93",X"FF",
		X"C8",X"99",X"9F",X"8E",X"9E",X"9E",X"CE",X"FF",X"31",X"99",X"F3",X"37",X"97",X"97",X"37",X"FF",
		X"CC",X"99",X"99",X"CC",X"9F",X"99",X"CC",X"FF",X"33",X"99",X"99",X"31",X"99",X"99",X"33",X"FF",
		X"FF",X"FF",X"EE",X"FF",X"FF",X"EE",X"FE",X"FC",X"FF",X"FF",X"77",X"FF",X"FF",X"77",X"F7",X"FF",
		X"FF",X"EF",X"C8",X"9F",X"C8",X"EF",X"FF",X"FF",X"1F",X"7F",X"F1",X"FF",X"F1",X"7F",X"1F",X"FF",
		X"8C",X"E9",X"FF",X"FF",X"FE",X"EF",X"8E",X"FF",X"F3",X"79",X"39",X"93",X"37",X"7F",X"F7",X"FF",
		X"FF",X"FE",X"FC",X"08",X"08",X"FE",X"FC",X"FF",X"F7",X"F3",X"F1",X"00",X"00",X"F3",X"F1",X"FF",
		X"EF",X"EF",X"EF",X"E0",X"E0",X"EF",X"EF",X"EF",X"7F",X"7F",X"7F",X"70",X"70",X"7F",X"7F",X"7F",
		X"FF",X"F0",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"FC",X"0C",X"0C",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F1",X"F0",X"FC",X"FE",X"FE",X"3F",X"3F",X"3F",X"3F",X"3F",X"37",X"37",X"37",
		X"EE",X"EE",X"EC",X"F0",X"F1",X"FF",X"FF",X"FF",X"77",X"77",X"37",X"0F",X"8F",X"FF",X"FF",X"FF",
		X"33",X"31",X"38",X"3C",X"3E",X"3F",X"0F",X"0F",X"FF",X"FF",X"FF",X"F7",X"F3",X"F1",X"08",X"0C",
		X"F0",X"F0",X"F3",X"E3",X"C3",X"83",X"13",X"33",X"C0",X"80",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"0F",X"0C",X"F8",X"F8",X"F8",X"F8",X"FC",X"FF",X"0F",X"03",X"C1",X"C1",X"C1",X"C1",X"C3",X"CF",
		X"FC",X"F8",X"F8",X"F8",X"FC",X"0E",X"0F",X"FF",X"F9",X"F0",X"F0",X"F0",X"F1",X"03",X"07",X"FF",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9E",X"9E",X"9E",X"FF",X"FF",X"FF",X"F8",X"F0",X"F3",X"F7",X"F7",
		X"3F",X"1C",X"88",X"C9",X"C9",X"88",X"1C",X"3F",X"CF",X"83",X"11",X"39",X"39",X"11",X"83",X"CF",
		X"EF",X"EF",X"9F",X"9F",X"EF",X"EF",X"CF",X"FF",X"79",X"79",X"99",X"99",X"79",X"79",X"39",X"F9",
		X"FE",X"EE",X"CE",X"80",X"C0",X"EE",X"FE",X"FE",X"77",X"37",X"17",X"00",X"10",X"37",X"77",X"F7",
		X"3E",X"3E",X"CE",X"CE",X"3E",X"3E",X"CE",X"CE",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"F0",X"F8",X"FC",X"CE",X"8F",X"CF",X"CF",X"FF",X"F0",X"F0",X"C0",X"10",X"90",X"98",X"9C",X"FE",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",
		X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",
		X"3F",X"3F",X"CF",X"CF",X"3F",X"3F",X"CF",X"CF",X"3C",X"3C",X"CC",X"CC",X"3C",X"3C",X"CC",X"CC",
		X"F0",X"F0",X"F0",X"F0",X"30",X"31",X"C3",X"C7",X"F0",X"F1",X"F3",X"F7",X"3F",X"3F",X"CF",X"CF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"C7",X"C7",X"C7",X"C0",X"C0",X"C7",X"C7",X"C7",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F0",X"00",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"EF",X"E0",X"E0",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"70",X"70",
		X"FE",X"FE",X"FE",X"E0",X"E0",X"EF",X"EF",X"EF",X"F7",X"F7",X"F7",X"00",X"00",X"7F",X"7F",X"7F",
		X"FE",X"FE",X"FE",X"00",X"00",X"EE",X"EE",X"EE",X"F7",X"F7",X"F7",X"07",X"07",X"77",X"77",X"77",
		X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"77",X"0F",X"0B",X"78",X"7F",X"67",X"30",X"00",X"C2",X"62",X"62",X"62",X"6E",X"6C",X"C0",
		X"00",X"33",X"77",X"DD",X"DD",X"77",X"33",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"66",X"FF",X"99",X"99",X"FF",X"FF",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"44",X"CC",X"88",X"88",X"FF",X"77",X"00",X"00",X"44",X"66",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"33",X"77",X"CC",X"88",X"FF",X"FF",X"00",X"00",X"88",X"CC",X"66",X"22",X"EE",X"EE",X"00",
		X"00",X"88",X"88",X"99",X"99",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"88",X"88",X"99",X"99",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"55",X"DD",X"99",X"88",X"FF",X"77",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"FF",X"FF",X"11",X"11",X"FF",X"FF",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"88",X"FF",X"FF",X"88",X"00",X"00",X"00",X"00",X"22",X"EE",X"EE",X"22",X"00",X"00",
		X"00",X"88",X"FF",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"22",X"66",X"44",X"00",
		X"00",X"88",X"CC",X"66",X"33",X"FF",X"FF",X"00",X"00",X"22",X"66",X"CC",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"FF",X"FF",X"66",X"33",X"66",X"FF",X"FF",X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"FF",X"FF",X"33",X"77",X"FF",X"FF",X"00",X"00",X"EE",X"EE",X"88",X"00",X"EE",X"EE",X"00",
		X"00",X"77",X"FF",X"88",X"88",X"FF",X"77",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"66",X"FF",X"99",X"99",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"77",X"FF",X"88",X"88",X"FF",X"77",X"00",X"00",X"AA",X"EE",X"66",X"44",X"CC",X"88",X"00",
		X"00",X"66",X"FF",X"99",X"99",X"FF",X"FF",X"00",X"00",X"22",X"66",X"CC",X"88",X"EE",X"EE",X"00",
		X"00",X"44",X"DD",X"99",X"99",X"FF",X"66",X"00",X"00",X"CC",X"EE",X"22",X"22",X"66",X"44",X"00",
		X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"88",X"CC",X"66",X"66",X"CC",X"88",X"00",
		X"FF",X"FF",X"00",X"11",X"00",X"FF",X"FF",X"00",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",
		X"00",X"CC",X"EE",X"33",X"33",X"EE",X"CC",X"00",X"00",X"66",X"EE",X"88",X"88",X"EE",X"66",X"00",
		X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",
		X"00",X"CC",X"EE",X"BB",X"99",X"88",X"88",X"00",X"00",X"22",X"22",X"22",X"AA",X"EE",X"66",X"00",
		X"00",X"00",X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",X"00",X"22",X"22",X"EE",X"EE",X"00",X"00",
		X"00",X"99",X"99",X"99",X"77",X"33",X"11",X"11",X"22",X"22",X"22",X"22",X"AA",X"EE",X"66",X"22",
		X"00",X"00",X"FF",X"FF",X"88",X"88",X"00",X"00",X"00",X"00",X"EE",X"EE",X"22",X"22",X"00",X"00",
		X"00",X"11",X"33",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"77",X"33",X"11",X"00",X"88",X"88",X"88",X"88",X"EE",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"FF",X"FF",X"22",X"22",X"FF",X"FF",X"22",X"88",X"EE",X"EE",X"88",X"88",X"EE",X"EE",X"88",
		X"00",X"44",X"55",X"DD",X"DD",X"77",X"22",X"00",X"00",X"88",X"CC",X"66",X"66",X"44",X"44",X"00",
		X"00",X"CC",X"66",X"33",X"11",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"88",X"CC",X"66",X"00",
		X"00",X"44",X"EE",X"BB",X"BB",X"FF",X"44",X"00",X"AA",X"EE",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"88",X"CC",X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CC",X"77",X"33",X"00",X"00",X"00",X"00",X"22",X"66",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"33",X"77",X"CC",X"88",X"00",X"00",X"00",X"00",X"88",X"CC",X"66",X"22",X"00",X"00",
		X"11",X"55",X"77",X"33",X"33",X"77",X"55",X"11",X"00",X"44",X"CC",X"88",X"88",X"CC",X"44",X"00",
		X"00",X"11",X"11",X"77",X"77",X"11",X"11",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",X"11",X"00",X"00",
		X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"44",X"66",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"66",X"22",X"00",
		X"00",X"77",X"FF",X"AA",X"99",X"FF",X"77",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"22",X"00",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",
		X"00",X"66",X"FF",X"99",X"88",X"CC",X"44",X"00",X"00",X"22",X"22",X"22",X"AA",X"EE",X"66",X"00",
		X"00",X"66",X"FF",X"99",X"99",X"CC",X"44",X"00",X"00",X"CC",X"EE",X"22",X"22",X"66",X"44",X"00",
		X"00",X"FF",X"FF",X"66",X"22",X"11",X"11",X"00",X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",
		X"00",X"99",X"BB",X"AA",X"AA",X"EE",X"EE",X"00",X"00",X"CC",X"EE",X"22",X"22",X"66",X"44",X"00",
		X"00",X"44",X"DD",X"99",X"99",X"FF",X"77",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"CC",X"EE",X"BB",X"99",X"CC",X"CC",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",
		X"00",X"66",X"FF",X"99",X"99",X"FF",X"66",X"00",X"00",X"CC",X"EE",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"77",X"FF",X"99",X"99",X"FF",X"66",X"00",X"00",X"CC",X"EE",X"22",X"22",X"66",X"44",X"00",
		X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",X"11",X"00",X"00",
		X"00",X"88",X"88",X"CC",X"66",X"33",X"11",X"00",X"00",X"22",X"22",X"66",X"CC",X"88",X"00",X"00",
		X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",
		X"00",X"11",X"33",X"66",X"CC",X"88",X"88",X"00",X"00",X"00",X"88",X"CC",X"66",X"22",X"22",X"00",
		X"00",X"66",X"FF",X"99",X"88",X"CC",X"44",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"70",X"D0",X"80",X"D0",X"F0",X"00",X"00",X"00",X"00",X"80",X"80",X"F0",X"F0",X"00",
		X"00",X"00",X"60",X"C0",X"C0",X"F0",X"70",X"00",X"00",X"00",X"60",X"30",X"30",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"70",X"90",X"F0",X"F0",X"00",X"00",X"00",X"E0",X"B0",X"10",X"B0",X"F0",X"00",
		X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"90",X"90",X"90",X"F0",X"00",
		X"00",X"00",X"00",X"70",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"F0",X"90",X"90",X"10",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"70",X"00",X"00",X"00",X"00",X"80",X"E0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"40",X"40",X"40",X"70",X"00",X"00",X"00",X"00",X"F0",X"90",X"90",X"90",X"00",
		X"00",X"00",X"00",X"40",X"40",X"40",X"70",X"00",X"00",X"00",X"00",X"F0",X"90",X"90",X"F0",X"00",
		X"00",X"00",X"00",X"70",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"00",X"00",
		X"00",X"00",X"00",X"70",X"40",X"40",X"70",X"00",X"00",X"00",X"00",X"F0",X"90",X"90",X"F0",X"00",
		X"00",X"00",X"00",X"70",X"40",X"40",X"70",X"00",X"00",X"00",X"00",X"F0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"40",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"10",X"00",
		X"00",X"00",X"F0",X"90",X"90",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"F0",X"90",X"90",X"F0",X"10",X"00",X"F0",X"F0",X"10",X"10",X"10",X"10",X"F0",X"00",
		X"33",X"44",X"88",X"8A",X"8A",X"89",X"44",X"33",X"CC",X"22",X"11",X"15",X"15",X"19",X"22",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
