library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity time_pilot_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of time_pilot_prog is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"B1",X"07",X"FF",X"FF",X"FF",X"33",X"4B",X"85",X"6F",X"30",X"01",X"24",X"7E",X"C9",X"4F",
		X"87",X"DF",X"5E",X"23",X"56",X"23",X"C9",X"4E",X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"41",
		X"7B",X"D6",X"20",X"5F",X"D0",X"15",X"C9",X"4D",X"7B",X"C6",X"20",X"5F",X"D0",X"14",X"C9",X"49",
		X"E1",X"D7",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"E5",X"26",X"AC",X"3A",X"B2",X"A9",X"6F",X"CB",
		X"7E",X"28",X"0A",X"72",X"2C",X"73",X"2C",X"7D",X"E6",X"3F",X"32",X"B2",X"A9",X"E1",X"C9",X"0F",
		X"A7",X"11",X"ED",X"77",X"68",X"D7",X"34",X"F1",X"D7",X"A5",X"3B",X"7C",X"FD",X"3B",X"7D",X"F1",
		X"DC",X"A5",X"8C",X"57",X"34",X"B9",X"C3",X"D8",X"00",X"32",X"00",X"C2",X"21",X"11",X"B4",X"06",
		X"30",X"36",X"00",X"23",X"10",X"FB",X"32",X"00",X"C2",X"21",X"10",X"B4",X"06",X"30",X"36",X"00",
		X"23",X"10",X"FB",X"32",X"00",X"C2",X"21",X"00",X"A8",X"11",X"01",X"A8",X"01",X"FF",X"07",X"36",
		X"00",X"ED",X"B0",X"32",X"00",X"C2",X"06",X"00",X"21",X"D8",X"00",X"AF",X"86",X"23",X"10",X"FC",
		X"D6",X"87",X"C4",X"D8",X"00",X"C3",X"66",X"58",X"32",X"00",X"C3",X"32",X"00",X"C2",X"C3",X"93",
		X"0B",X"21",X"20",X"A4",X"0E",X"0E",X"11",X"20",X"00",X"19",X"06",X"10",X"CD",X"C7",X"00",X"23",
		X"23",X"10",X"F9",X"0D",X"20",X"F0",X"C9",X"E5",X"36",X"56",X"23",X"36",X"83",X"11",X"1F",X"00",
		X"19",X"36",X"C7",X"23",X"36",X"EF",X"E1",X"C9",X"F5",X"C5",X"D5",X"E5",X"08",X"D9",X"F5",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"65",X"03",X"CD",X"86",X"52",X"AF",X"32",X"00",X"C3",
		X"32",X"00",X"C2",X"3C",X"32",X"87",X"A9",X"3A",X"32",X"AD",X"A7",X"28",X"09",X"3A",X"C2",X"A9",
		X"A7",X"20",X"03",X"32",X"87",X"A9",X"3A",X"87",X"A9",X"32",X"02",X"C3",X"3A",X"00",X"C2",X"2F",
		X"32",X"AD",X"A9",X"3A",X"00",X"C3",X"2F",X"32",X"AE",X"A9",X"3A",X"20",X"C3",X"2F",X"32",X"AF",
		X"A9",X"3A",X"40",X"C3",X"2F",X"32",X"B0",X"A9",X"3A",X"60",X"C3",X"2F",X"32",X"B1",X"A9",X"21",
		X"80",X"A9",X"34",X"21",X"CE",X"A9",X"7E",X"3C",X"27",X"77",X"21",X"17",X"A8",X"7E",X"A7",X"28",
		X"01",X"35",X"21",X"12",X"A8",X"7E",X"A7",X"28",X"01",X"35",X"21",X"F4",X"A8",X"7E",X"A7",X"28",
		X"01",X"35",X"CD",X"BE",X"48",X"21",X"74",X"01",X"E5",X"3A",X"AB",X"A9",X"E6",X"03",X"F7",X"C2",
		X"15",X"51",X"16",X"FE",X"17",X"1F",X"0F",X"6F",X"A6",X"14",X"88",X"57",X"A5",X"BF",X"34",X"D7",
		X"F1",X"96",X"F1",X"B9",X"CD",X"D4",X"55",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"D9",
		X"08",X"E1",X"D1",X"C1",X"3A",X"00",X"16",X"32",X"00",X"C3",X"F1",X"C9",X"87",X"30",X"01",X"24",
		X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"23",X"C9",X"21",X"00",X"A4",X"22",X"89",X"A9",
		X"3E",X"20",X"32",X"88",X"A9",X"06",X"F0",X"21",X"A5",X"4B",X"AF",X"86",X"23",X"10",X"FC",X"D6",
		X"11",X"C4",X"67",X"01",X"C9",X"21",X"04",X"A4",X"22",X"89",X"A9",X"3A",X"CD",X"0C",X"32",X"88",
		X"A9",X"C9",X"2A",X"89",X"A9",X"06",X"20",X"11",X"20",X"00",X"36",X"F1",X"CB",X"94",X"36",X"10",
		X"CB",X"D4",X"19",X"10",X"F5",X"2A",X"89",X"A9",X"23",X"22",X"89",X"A9",X"21",X"88",X"A9",X"35",
		X"C9",X"AF",X"32",X"E2",X"A9",X"2A",X"45",X"0D",X"22",X"E3",X"A9",X"2A",X"0C",X"28",X"22",X"E5",
		X"A9",X"06",X"00",X"21",X"33",X"0E",X"AF",X"86",X"23",X"10",X"FC",X"D6",X"FD",X"C4",X"69",X"00",
		X"C9",X"CD",X"6F",X"02",X"2A",X"F5",X"32",X"ED",X"4B",X"E3",X"A9",X"A7",X"ED",X"42",X"29",X"29",
		X"29",X"29",X"3E",X"00",X"DE",X"00",X"6C",X"67",X"22",X"E7",X"A9",X"2A",X"45",X"0B",X"ED",X"4B",
		X"E5",X"A9",X"A7",X"ED",X"42",X"29",X"29",X"29",X"29",X"3E",X"00",X"DE",X"00",X"6C",X"67",X"22",
		X"E9",X"A9",X"2A",X"E3",X"A9",X"ED",X"4B",X"E7",X"A9",X"09",X"22",X"E3",X"A9",X"2A",X"E5",X"A9",
		X"ED",X"4B",X"E9",X"A9",X"09",X"22",X"E5",X"A9",X"CD",X"6F",X"02",X"ED",X"5B",X"B2",X"14",X"A7",
		X"ED",X"52",X"C2",X"32",X"02",X"21",X"E2",X"A9",X"34",X"7E",X"21",X"90",X"02",X"D7",X"21",X"E3",
		X"A9",X"36",X"00",X"23",X"73",X"21",X"E5",X"A9",X"36",X"00",X"23",X"72",X"7B",X"A7",X"C9",X"3A",
		X"E4",X"A9",X"87",X"87",X"87",X"6F",X"26",X"00",X"29",X"29",X"3A",X"E6",X"A9",X"85",X"6F",X"3E",
		X"A4",X"84",X"67",X"3A",X"0B",X"AD",X"77",X"CB",X"94",X"3A",X"0C",X"AD",X"77",X"CB",X"D4",X"C9",
		X"10",X"04",X"11",X"04",X"12",X"04",X"13",X"04",X"14",X"04",X"15",X"04",X"16",X"04",X"17",X"04",
		X"18",X"04",X"19",X"04",X"1A",X"04",X"1B",X"04",X"1C",X"04",X"1D",X"04",X"1D",X"05",X"1D",X"06",
		X"1D",X"07",X"1D",X"08",X"1D",X"09",X"1D",X"0A",X"1D",X"0B",X"1D",X"0C",X"1D",X"0D",X"1D",X"0E",
		X"1D",X"0F",X"1D",X"10",X"1D",X"11",X"1D",X"12",X"1D",X"13",X"1D",X"14",X"1D",X"15",X"1D",X"16",
		X"1D",X"17",X"1D",X"18",X"1D",X"19",X"1D",X"1A",X"1D",X"1B",X"1D",X"1C",X"1D",X"1D",X"1D",X"1E",
		X"1C",X"1E",X"1B",X"1E",X"1A",X"1E",X"19",X"1E",X"18",X"1E",X"17",X"1E",X"16",X"1E",X"15",X"1E",
		X"14",X"1E",X"13",X"1E",X"12",X"1E",X"11",X"1E",X"10",X"1E",X"0F",X"1E",X"0E",X"1E",X"0D",X"1E",
		X"0C",X"1E",X"0B",X"1E",X"0A",X"1E",X"09",X"1E",X"08",X"1E",X"07",X"1E",X"06",X"1E",X"05",X"1E",
		X"04",X"1E",X"03",X"1E",X"02",X"1E",X"02",X"1D",X"02",X"1C",X"02",X"1B",X"02",X"1A",X"02",X"19",
		X"02",X"18",X"02",X"17",X"02",X"16",X"02",X"15",X"02",X"14",X"02",X"13",X"02",X"12",X"02",X"11",
		X"02",X"10",X"02",X"0F",X"02",X"0E",X"02",X"0D",X"02",X"0C",X"02",X"0B",X"02",X"0A",X"02",X"09",
		X"02",X"08",X"02",X"07",X"02",X"06",X"02",X"05",X"02",X"04",X"03",X"04",X"04",X"04",X"05",X"04",
		X"06",X"04",X"07",X"04",X"08",X"04",X"09",X"04",X"0A",X"04",X"0B",X"04",X"0C",X"04",X"0D",X"04",
		X"0E",X"04",X"0F",X"04",X"00",X"21",X"30",X"AA",X"11",X"10",X"B0",X"3A",X"87",X"A9",X"A7",X"CA",
		X"56",X"05",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"21",X"10",
		X"AA",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",
		X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",
		X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",
		X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",
		X"A0",X"21",X"36",X"AA",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",
		X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"21",X"60",X"AA",X"11",X"10",X"B4",X"ED",X"A0",
		X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",
		X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"21",X"40",X"AA",X"ED",X"A0",X"7E",X"C6",
		X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",
		X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",
		X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",
		X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",
		X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",
		X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",
		X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",
		X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",
		X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"21",X"66",X"AA",X"ED",
		X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",
		X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",
		X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0E",X"2F",X"12",X"2C",X"1C",X"3A",X"AB",X"A9",X"FE",
		X"03",X"C0",X"3A",X"AC",X"A9",X"21",X"32",X"08",X"BE",X"D8",X"FE",X"08",X"D0",X"3A",X"11",X"B4",
		X"C6",X"80",X"38",X"0A",X"32",X"11",X"B4",X"21",X"10",X"B0",X"7E",X"C6",X"80",X"77",X"3A",X"13",
		X"B4",X"C6",X"80",X"38",X"0A",X"32",X"13",X"B4",X"21",X"12",X"B0",X"7E",X"C6",X"80",X"77",X"3A",
		X"15",X"B4",X"C6",X"80",X"38",X"0A",X"32",X"15",X"B4",X"21",X"14",X"B0",X"7E",X"C6",X"80",X"77",
		X"3A",X"37",X"B4",X"C6",X"80",X"38",X"0A",X"32",X"37",X"B4",X"21",X"36",X"B0",X"7E",X"C6",X"80",
		X"77",X"3A",X"39",X"B4",X"C6",X"80",X"38",X"0A",X"32",X"39",X"B4",X"21",X"38",X"B0",X"7E",X"C6",
		X"80",X"77",X"3A",X"3B",X"B4",X"C6",X"80",X"38",X"0A",X"32",X"3B",X"B4",X"21",X"3A",X"B0",X"7E",
		X"C6",X"80",X"77",X"3A",X"3D",X"B4",X"C6",X"80",X"38",X"0A",X"32",X"3D",X"B4",X"21",X"3C",X"B0",
		X"7E",X"C6",X"80",X"77",X"3A",X"3F",X"B4",X"C6",X"80",X"38",X"0A",X"32",X"3F",X"B4",X"21",X"3E",
		X"B0",X"7E",X"C6",X"80",X"77",X"C9",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",
		X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",
		X"A0",X"21",X"10",X"AA",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",
		X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",
		X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",
		X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",
		X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",
		X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",
		X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",
		X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",
		X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",
		X"2C",X"1C",X"ED",X"A0",X"21",X"36",X"AA",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",
		X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",
		X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",X"2C",X"1C",X"ED",X"A0",X"7E",X"C6",X"0F",X"2F",X"12",
		X"2C",X"1C",X"ED",X"A0",X"21",X"60",X"AA",X"11",X"10",X"B4",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",
		X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",
		X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"21",X"40",X"AA",X"7E",X"EE",
		X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",
		X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",
		X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",
		X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",
		X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",
		X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",
		X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",
		X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",
		X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",
		X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",
		X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"21",X"66",
		X"AA",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",
		X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",
		X"2C",X"1C",X"7E",X"EE",X"C0",X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"7E",X"EE",X"C0",
		X"12",X"2C",X"1C",X"7E",X"3C",X"12",X"2C",X"1C",X"C3",X"BC",X"04",X"06",X"00",X"21",X"A0",X"4A",
		X"AF",X"86",X"23",X"10",X"FC",X"D6",X"B8",X"C2",X"FA",X"08",X"3A",X"0C",X"AD",X"FE",X"05",X"F5",
		X"3E",X"05",X"32",X"0C",X"AD",X"3E",X"F1",X"32",X"0B",X"AD",X"CD",X"E1",X"01",X"F1",X"CC",X"1A",
		X"0F",X"C3",X"1A",X"0F",X"06",X"00",X"21",X"99",X"4C",X"97",X"AE",X"23",X"10",X"FC",X"C6",X"95",
		X"C4",X"11",X"0F",X"3A",X"30",X"AD",X"A7",X"28",X"17",X"ED",X"5B",X"5B",X"12",X"3A",X"32",X"AD",
		X"A7",X"28",X"01",X"1C",X"FF",X"3A",X"0E",X"AD",X"A7",X"28",X"05",X"16",X"07",X"FF",X"18",X"04",
		X"11",X"02",X"02",X"FF",X"CD",X"09",X"08",X"CD",X"F0",X"19",X"C3",X"1A",X"0F",X"47",X"C3",X"03",
		X"53",X"3A",X"00",X"60",X"FE",X"55",X"CA",X"00",X"60",X"31",X"00",X"B0",X"32",X"00",X"C2",X"21",
		X"00",X"C3",X"06",X"08",X"36",X"00",X"23",X"10",X"FB",X"3A",X"4B",X"2D",X"32",X"08",X"C3",X"C3",
		X"69",X"00",X"21",X"9F",X"A7",X"11",X"E0",X"FF",X"06",X"0E",X"36",X"F1",X"CB",X"94",X"36",X"16",
		X"CB",X"D4",X"19",X"10",X"F5",X"C9",X"CD",X"06",X"0B",X"CD",X"39",X"0B",X"21",X"1C",X"A6",X"11",
		X"FE",X"AB",X"CD",X"FC",X"1A",X"3A",X"AE",X"A9",X"CB",X"5F",X"C2",X"15",X"32",X"3A",X"86",X"A9",
		X"3D",X"C8",X"11",X"19",X"01",X"FF",X"C3",X"1A",X"0F",X"3A",X"04",X"AD",X"87",X"47",X"87",X"87",
		X"80",X"21",X"7C",X"08",X"DF",X"46",X"23",X"4E",X"23",X"3A",X"02",X"AD",X"5F",X"E6",X"07",X"CF",
		X"08",X"7B",X"21",X"9F",X"A7",X"11",X"E0",X"FF",X"0F",X"0F",X"E6",X"1F",X"28",X"0A",X"70",X"19",
		X"3D",X"28",X"05",X"71",X"19",X"3D",X"20",X"F6",X"08",X"77",X"19",X"36",X"F1",X"C9",X"CD",X"39",
		X"0B",X"CD",X"06",X"0B",X"11",X"00",X"01",X"06",X"02",X"FF",X"1C",X"10",X"FC",X"1C",X"06",X"05",
		X"FF",X"1C",X"10",X"FC",X"1E",X"14",X"FF",X"1C",X"FF",X"21",X"6A",X"17",X"06",X"18",X"AF",X"AE",
		X"2C",X"10",X"FC",X"D6",X"C9",X"C2",X"FA",X"08",X"C3",X"1A",X"0F",X"BC",X"A6",X"10",X"30",X"F1",
		X"7C",X"68",X"3B",X"A5",X"38",X"FD",X"F1",X"96",X"5D",X"17",X"9B",X"B9",X"4C",X"4F",X"F1",X"41",
		X"72",X"A6",X"F1",X"8D",X"E2",X"FB",X"37",X"A7",X"F1",X"AB",X"31",X"07",X"F1",X"5A",X"75",X"85",
		X"D9",X"1B",X"F1",X"C1",X"E1",X"FA",X"F1",X"B3",X"A0",X"47",X"7B",X"78",X"F1",X"04",X"05",X"C2",
		X"F1",X"DE",X"F9",X"BB",X"93",X"AC",X"F1",X"36",X"06",X"4B",X"F1",X"EE",X"D3",X"D4",X"21",X"5E",
		X"33",X"06",X"1E",X"C9",X"CD",X"01",X"02",X"C0",X"06",X"00",X"21",X"80",X"48",X"97",X"AE",X"23",
		X"10",X"FC",X"C6",X"D0",X"C2",X"D9",X"00",X"11",X"13",X"01",X"FF",X"1E",X"00",X"FF",X"1E",X"14",
		X"FF",X"1C",X"FF",X"1E",X"0C",X"FF",X"CD",X"DC",X"4B",X"21",X"95",X"A9",X"AF",X"06",X"05",X"77",
		X"23",X"10",X"FC",X"36",X"03",X"ED",X"5B",X"93",X"A9",X"3A",X"99",X"A9",X"21",X"C7",X"12",X"CF",
		X"12",X"CB",X"92",X"1A",X"32",X"90",X"A9",X"C3",X"1A",X"0F",X"4B",X"01",X"4A",X"01",X"49",X"01",
		X"48",X"01",X"47",X"01",X"46",X"01",X"45",X"01",X"40",X"01",X"3E",X"01",X"3C",X"01",X"3A",X"01",
		X"38",X"01",X"32",X"01",X"2F",X"01",X"2D",X"01",X"27",X"01",X"24",X"01",X"21",X"01",X"1E",X"01",
		X"18",X"01",X"15",X"01",X"12",X"01",X"0C",X"01",X"09",X"01",X"06",X"01",X"00",X"01",X"FD",X"00",
		X"FA",X"00",X"F7",X"00",X"F1",X"00",X"EE",X"00",X"EB",X"00",X"E5",X"00",X"E2",X"00",X"DE",X"00",
		X"D8",X"00",X"D5",X"00",X"D1",X"00",X"CA",X"00",X"C6",X"00",X"C3",X"00",X"BC",X"00",X"B6",X"00",
		X"AE",X"00",X"A9",X"00",X"9F",X"00",X"9C",X"00",X"93",X"00",X"8A",X"00",X"84",X"00",X"7B",X"00",
		X"71",X"00",X"6B",X"00",X"61",X"00",X"57",X"00",X"50",X"00",X"45",X"00",X"3B",X"00",X"34",X"00",
		X"29",X"00",X"1E",X"00",X"13",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"F8",X"FF",X"ED",X"FF",
		X"00",X"00",X"D7",X"FF",X"CC",X"FF",X"C5",X"FF",X"BB",X"FF",X"B0",X"FF",X"A9",X"FF",X"9F",X"FF",
		X"95",X"FF",X"8F",X"FF",X"85",X"FF",X"7C",X"FF",X"76",X"FF",X"6D",X"FF",X"64",X"FF",X"61",X"FF",
		X"64",X"FF",X"52",X"FF",X"4A",X"FF",X"44",X"FF",X"3D",X"FF",X"3A",X"FF",X"36",X"FF",X"2F",X"FF",
		X"2B",X"FF",X"28",X"FF",X"22",X"FF",X"1E",X"FF",X"1B",X"FF",X"15",X"FF",X"12",X"FF",X"0F",X"FF",
		X"0F",X"FF",X"06",X"FF",X"03",X"FF",X"00",X"FF",X"FA",X"FE",X"F7",X"FE",X"F4",X"FE",X"EE",X"FE",
		X"EB",X"FE",X"E8",X"FE",X"E2",X"FE",X"DF",X"FE",X"DC",X"FE",X"D9",X"FE",X"D3",X"FE",X"D1",X"FE",
		X"CE",X"FE",X"C8",X"FE",X"C6",X"FE",X"C4",X"FE",X"C2",X"FE",X"C0",X"FE",X"BB",X"FE",X"BA",X"FE",
		X"B9",X"FE",X"B8",X"FE",X"B7",X"FE",X"B6",X"FE",X"B5",X"FE",X"B5",X"FE",X"B6",X"FE",X"B7",X"FE",
		X"B8",X"FE",X"B9",X"FE",X"BA",X"FE",X"BB",X"FE",X"C0",X"FE",X"C2",X"FE",X"C4",X"FE",X"C6",X"FE",
		X"C8",X"FE",X"CE",X"FE",X"D1",X"FE",X"D3",X"FE",X"D9",X"FE",X"DC",X"FE",X"DF",X"FE",X"E2",X"FE",
		X"E8",X"FE",X"EB",X"FE",X"EE",X"FE",X"F4",X"FE",X"F7",X"FE",X"FA",X"FE",X"00",X"FF",X"03",X"FF",
		X"06",X"FF",X"09",X"FF",X"0F",X"FF",X"12",X"FF",X"15",X"FF",X"1B",X"FF",X"1E",X"FF",X"22",X"FF",
		X"28",X"FF",X"2B",X"FF",X"2F",X"FF",X"36",X"FF",X"3A",X"FF",X"3D",X"FF",X"44",X"FF",X"4A",X"FF",
		X"52",X"FF",X"57",X"FF",X"61",X"FF",X"64",X"FF",X"6D",X"FF",X"76",X"FF",X"7C",X"FF",X"85",X"FF",
		X"8F",X"FF",X"95",X"FF",X"9F",X"FF",X"A9",X"FF",X"B0",X"FF",X"BB",X"FF",X"C5",X"FF",X"CC",X"FF",
		X"D7",X"FF",X"E2",X"FF",X"ED",X"FF",X"F8",X"FF",X"00",X"00",X"00",X"00",X"08",X"00",X"13",X"00",
		X"1E",X"00",X"29",X"00",X"34",X"00",X"3B",X"00",X"45",X"00",X"50",X"00",X"57",X"00",X"61",X"00",
		X"6B",X"00",X"71",X"00",X"7B",X"00",X"84",X"00",X"8A",X"00",X"93",X"00",X"9C",X"00",X"9F",X"00",
		X"9F",X"00",X"AE",X"00",X"B6",X"00",X"BC",X"00",X"C3",X"00",X"C6",X"00",X"CA",X"00",X"D1",X"00",
		X"D5",X"00",X"D8",X"00",X"DE",X"00",X"E2",X"00",X"E5",X"00",X"EB",X"00",X"EE",X"00",X"F1",X"00",
		X"EE",X"00",X"FA",X"00",X"FD",X"00",X"00",X"01",X"06",X"01",X"09",X"01",X"0C",X"01",X"12",X"01",
		X"15",X"01",X"18",X"01",X"1E",X"01",X"21",X"01",X"24",X"01",X"27",X"01",X"2D",X"01",X"2F",X"01",
		X"27",X"01",X"38",X"01",X"3A",X"01",X"3C",X"01",X"3E",X"01",X"40",X"01",X"45",X"01",X"46",X"01",
		X"47",X"01",X"48",X"01",X"49",X"01",X"4A",X"01",X"4B",X"01",X"77",X"A6",X"13",X"ED",X"DC",X"A5",
		X"7D",X"34",X"F1",X"F1",X"F1",X"B9",X"FD",X"21",X"10",X"AA",X"06",X"04",X"0E",X"04",X"16",X"A0",
		X"1E",X"D8",X"FD",X"72",X"31",X"FD",X"73",X"00",X"FD",X"71",X"01",X"FD",X"36",X"30",X"6C",X"FD",
		X"23",X"FD",X"23",X"0C",X"7A",X"D6",X"10",X"57",X"10",X"E8",X"C9",X"21",X"41",X"AA",X"11",X"02",
		X"00",X"06",X"04",X"AF",X"77",X"19",X"10",X"FC",X"C9",X"3A",X"80",X"A9",X"CB",X"47",X"28",X"06",
		X"11",X"00",X"01",X"C3",X"38",X"00",X"11",X"1F",X"01",X"C3",X"38",X"00",X"AF",X"86",X"23",X"10",
		X"FC",X"B9",X"C8",X"C9",X"AF",X"AE",X"23",X"10",X"FC",X"B9",X"C8",X"C3",X"00",X"00",X"AF",X"86",
		X"23",X"0D",X"28",X"02",X"18",X"F9",X"CB",X"47",X"C8",X"C3",X"00",X"00",X"21",X"06",X"0B",X"06",
		X"24",X"0E",X"00",X"7E",X"91",X"23",X"10",X"FB",X"EB",X"BE",X"C9",X"0F",X"A7",X"13",X"88",X"0D",
		X"ED",X"C4",X"F1",X"ED",X"DC",X"A5",X"D7",X"DC",X"F1",X"8C",X"0D",X"DC",X"DC",X"68",X"3B",X"B9",
		X"C3",X"93",X"0B",X"26",X"AC",X"3A",X"B3",X"A9",X"6F",X"7E",X"07",X"DA",X"90",X"0B",X"4E",X"36",
		X"FF",X"23",X"46",X"36",X"FF",X"23",X"7D",X"E6",X"3F",X"32",X"B3",X"A9",X"79",X"E6",X"0F",X"21",
		X"BC",X"0B",X"CD",X"8C",X"01",X"78",X"21",X"90",X"0B",X"E5",X"EB",X"E9",X"DD",X"0B",X"F2",X"0B",
		X"0F",X"0C",X"39",X"0C",X"90",X"0C",X"72",X"4D",X"D7",X"0D",X"AC",X"0E",X"DC",X"0B",X"DC",X"0B",
		X"21",X"34",X"23",X"0C",X"DC",X"0B",X"DC",X"0B",X"DC",X"0B",X"DC",X"0B",X"C9",X"21",X"50",X"0C",
		X"CD",X"8C",X"01",X"EB",X"5E",X"23",X"56",X"23",X"23",X"7E",X"FE",X"B9",X"C8",X"12",X"23",X"E7",
		X"18",X"F7",X"21",X"50",X"0C",X"CD",X"8C",X"01",X"EB",X"5E",X"23",X"56",X"23",X"4E",X"23",X"7E",
		X"FE",X"B9",X"C8",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"23",X"E7",X"C3",X"FF",X"0B",X"21",
		X"50",X"0C",X"CD",X"8C",X"01",X"EB",X"5E",X"23",X"56",X"23",X"23",X"3A",X"0C",X"AD",X"E6",X"0F",
		X"4F",X"18",X"DC",X"21",X"50",X"0C",X"CD",X"8C",X"01",X"EB",X"5E",X"23",X"56",X"23",X"23",X"3A",
		X"0C",X"AD",X"C6",X"0A",X"E6",X"0F",X"4F",X"18",X"C6",X"21",X"50",X"0C",X"CD",X"8C",X"01",X"EB",
		X"5E",X"23",X"56",X"23",X"23",X"7E",X"FE",X"B9",X"C8",X"3E",X"F1",X"12",X"23",X"E7",X"18",X"F5",
		X"6B",X"08",X"73",X"16",X"7F",X"30",X"1D",X"58",X"FA",X"49",X"D6",X"15",X"4C",X"58",X"09",X"25",
		X"CA",X"15",X"67",X"01",X"42",X"4E",X"10",X"18",X"CE",X"48",X"A4",X"1B",X"FA",X"0A",X"31",X"24",
		X"3B",X"12",X"9B",X"45",X"A4",X"2C",X"4F",X"00",X"9E",X"31",X"6E",X"29",X"7B",X"0B",X"5C",X"34",
		X"D2",X"3E",X"48",X"33",X"49",X"0F",X"14",X"4C",X"54",X"59",X"ED",X"55",X"D8",X"23",X"00",X"49",
		X"4F",X"06",X"00",X"3A",X"30",X"AD",X"A7",X"CA",X"E8",X"0C",X"79",X"A7",X"CA",X"E9",X"0C",X"21",
		X"27",X"0D",X"09",X"09",X"09",X"11",X"33",X"AD",X"3A",X"32",X"AD",X"A7",X"28",X"03",X"11",X"36",
		X"AD",X"1A",X"86",X"27",X"12",X"13",X"23",X"1A",X"8E",X"27",X"12",X"13",X"23",X"1A",X"8E",X"27",
		X"12",X"21",X"8D",X"A9",X"01",X"03",X"00",X"1A",X"BE",X"38",X"0F",X"20",X"07",X"1B",X"2B",X"0D",
		X"20",X"F5",X"18",X"06",X"EB",X"ED",X"B8",X"CD",X"6B",X"0D",X"3A",X"32",X"AD",X"A7",X"20",X"05",
		X"CD",X"57",X"0D",X"18",X"03",X"CD",X"61",X"0D",X"C9",X"3A",X"31",X"AD",X"A7",X"20",X"1B",X"3A",
		X"31",X"0B",X"CD",X"F2",X"0B",X"CD",X"57",X"0D",X"3A",X"C6",X"15",X"CD",X"39",X"0C",X"11",X"01",
		X"A5",X"06",X"06",X"3E",X"F1",X"12",X"E7",X"10",X"FA",X"C9",X"3E",X"06",X"CD",X"F2",X"0B",X"CD",
		X"57",X"0D",X"3E",X"07",X"CD",X"F2",X"0B",X"CD",X"61",X"0D",X"C9",X"3C",X"A2",X"C7",X"AC",X"7C",
		X"A2",X"43",X"AB",X"FC",X"A1",X"BE",X"AC",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",
		X"00",X"03",X"00",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"06",X"00",X"00",X"07",X"00",X"00",
		X"08",X"00",X"00",X"09",X"00",X"00",X"10",X"00",X"00",X"15",X"00",X"00",X"20",X"00",X"00",X"30",
		X"00",X"00",X"40",X"00",X"00",X"50",X"00",X"11",X"81",X"A7",X"21",X"35",X"AD",X"0E",X"10",X"18",
		X"12",X"11",X"01",X"A5",X"21",X"38",X"AD",X"0E",X"10",X"18",X"08",X"11",X"41",X"A6",X"21",X"8D",
		X"A9",X"0E",X"10",X"06",X"00",X"CD",X"A0",X"0D",X"2B",X"CD",X"A0",X"0D",X"2B",X"CD",X"81",X"0D",
		X"C9",X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"90",X"0D",X"E7",X"7E",X"CD",X"90",X"0D",X"E7",X"C9",
		X"E6",X"0F",X"E5",X"21",X"CC",X"0D",X"CF",X"E1",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"C9",
		X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"AF",X"0D",X"E7",X"7E",X"CD",X"AF",X"0D",X"E7",X"C9",X"E6",
		X"0F",X"28",X"03",X"04",X"18",X"08",X"3A",X"46",X"32",X"04",X"05",X"28",X"01",X"AF",X"E5",X"21",
		X"CC",X"0D",X"CF",X"E1",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"C9",X"13",X"96",X"9B",X"CD",
		X"F3",X"7F",X"65",X"02",X"17",X"5D",X"F1",X"11",X"63",X"A4",X"FE",X"64",X"38",X"02",X"3E",X"63",
		X"D9",X"06",X"00",X"D6",X"1E",X"38",X"03",X"04",X"18",X"F9",X"C6",X"1E",X"0E",X"00",X"D6",X"0A",
		X"38",X"03",X"0C",X"18",X"F9",X"C6",X"0A",X"16",X"00",X"D6",X"05",X"38",X"03",X"14",X"18",X"F9",
		X"C6",X"05",X"5F",X"D9",X"D9",X"7B",X"D9",X"A7",X"28",X"0C",X"06",X"01",X"0E",X"13",X"08",X"CD",
		X"8D",X"0E",X"08",X"3D",X"20",X"F8",X"D9",X"7A",X"D9",X"A7",X"28",X"0C",X"06",X"32",X"0E",X"11",
		X"08",X"CD",X"9C",X"0E",X"08",X"3D",X"20",X"F8",X"D9",X"79",X"D9",X"A7",X"28",X"0C",X"06",X"CE",
		X"0E",X"16",X"08",X"CD",X"70",X"0E",X"08",X"3D",X"20",X"F8",X"D9",X"78",X"D9",X"A7",X"28",X"0C",
		X"06",X"23",X"0E",X"11",X"08",X"CD",X"70",X"0E",X"08",X"3D",X"20",X"F8",X"01",X"10",X"F1",X"21",
		X"DD",X"59",X"19",X"38",X"05",X"CD",X"8D",X"0E",X"18",X"F5",X"AF",X"2A",X"A0",X"00",X"ED",X"5B",
		X"A3",X"00",X"ED",X"4B",X"9D",X"00",X"19",X"09",X"85",X"84",X"D6",X"69",X"C2",X"00",X"00",X"C9",
		X"78",X"3C",X"12",X"3D",X"1B",X"12",X"EF",X"78",X"C6",X"02",X"12",X"3C",X"13",X"12",X"21",X"00",
		X"FC",X"19",X"EF",X"71",X"2B",X"71",X"EB",X"E7",X"EB",X"71",X"23",X"71",X"C9",X"EB",X"70",X"2B",
		X"36",X"F1",X"CB",X"94",X"71",X"23",X"71",X"CB",X"D4",X"EB",X"EF",X"C9",X"EB",X"04",X"70",X"05",
		X"2B",X"70",X"CB",X"94",X"71",X"23",X"71",X"CB",X"D4",X"EB",X"EF",X"C9",X"3A",X"01",X"AD",X"FE",
		X"64",X"D0",X"3E",X"0E",X"CD",X"0F",X"0C",X"EF",X"EF",X"21",X"01",X"AD",X"06",X"01",X"3A",X"0C",
		X"AD",X"4F",X"C5",X"0E",X"00",X"7E",X"D6",X"0A",X"38",X"03",X"0C",X"18",X"F9",X"C6",X"0A",X"08",
		X"79",X"C1",X"CD",X"EB",X"0E",X"E7",X"08",X"CD",X"EB",X"0E",X"E7",X"11",X"48",X"17",X"01",X"8C",
		X"10",X"1A",X"81",X"4F",X"13",X"10",X"FA",X"C2",X"09",X"25",X"C9",X"E6",X"0F",X"28",X"10",X"06",
		X"00",X"E5",X"21",X"06",X"0F",X"CF",X"E1",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"C9",X"78",
		X"A7",X"28",X"EE",X"05",X"EF",X"C9",X"E3",X"49",X"A8",X"64",X"27",X"AE",X"42",X"B0",X"D5",X"86",
		X"F1",X"21",X"AB",X"A9",X"34",X"AF",X"32",X"AC",X"A9",X"C9",X"21",X"AC",X"A9",X"34",X"C9",X"21",
		X"54",X"0F",X"E5",X"3A",X"AC",X"A9",X"E6",X"0F",X"F7",X"B1",X"27",X"5E",X"33",X"D7",X"5B",X"75",
		X"4C",X"74",X"07",X"AF",X"16",X"94",X"56",X"99",X"11",X"0B",X"33",X"B4",X"08",X"C3",X"18",X"E2",
		X"12",X"FB",X"12",X"0F",X"4A",X"23",X"13",X"B5",X"15",X"73",X"A6",X"14",X"7E",X"29",X"F8",X"96",
		X"5D",X"96",X"13",X"B9",X"3A",X"30",X"AD",X"A7",X"C0",X"3A",X"86",X"A9",X"A7",X"20",X"11",X"3A",
		X"C0",X"A9",X"A7",X"C8",X"3A",X"AE",X"A9",X"E6",X"18",X"C8",X"CD",X"B6",X"15",X"C3",X"90",X"16",
		X"AF",X"32",X"AC",X"A9",X"3A",X"36",X"17",X"32",X"AB",X"A9",X"C9",X"87",X"87",X"21",X"6A",X"18",
		X"11",X"D3",X"A9",X"DF",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"C9",X"F1",X"01",X"F1",
		X"02",X"F1",X"03",X"F1",X"04",X"F1",X"05",X"3A",X"11",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"11",X"B4",X"3A",
		X"10",X"B0",X"C6",X"80",X"32",X"10",X"B0",X"3A",X"13",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"13",X"B4",X"3A",
		X"12",X"B0",X"C6",X"80",X"32",X"12",X"B0",X"3A",X"15",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"15",X"B4",X"3A",
		X"14",X"B0",X"C6",X"80",X"32",X"14",X"B0",X"3A",X"37",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"37",X"B4",X"3A",
		X"36",X"B0",X"C6",X"80",X"32",X"36",X"B0",X"3A",X"39",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"39",X"B4",X"3A",
		X"38",X"B0",X"C6",X"80",X"32",X"38",X"B0",X"3A",X"3B",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"3B",X"B4",X"3A",
		X"3A",X"B0",X"C6",X"80",X"32",X"3A",X"B0",X"3A",X"3D",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"3D",X"B4",X"3A",
		X"3C",X"B0",X"C6",X"80",X"32",X"3C",X"B0",X"3A",X"3F",X"B4",X"CB",X"7F",X"28",X"19",X"4F",X"3A",
		X"00",X"C0",X"81",X"30",X"12",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"3F",X"B4",X"3A",
		X"3E",X"B0",X"C6",X"80",X"32",X"3E",X"B0",X"C9",X"3A",X"11",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"11",X"B4",
		X"3A",X"10",X"B0",X"C6",X"80",X"32",X"10",X"B0",X"3A",X"13",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"13",X"B4",
		X"3A",X"12",X"B0",X"C6",X"80",X"32",X"12",X"B0",X"3A",X"15",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"15",X"B4",
		X"3A",X"14",X"B0",X"C6",X"80",X"32",X"14",X"B0",X"3A",X"37",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"37",X"B4",
		X"3A",X"36",X"B0",X"C6",X"80",X"32",X"36",X"B0",X"3A",X"39",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"39",X"B4",
		X"3A",X"38",X"B0",X"C6",X"80",X"32",X"38",X"B0",X"3A",X"3B",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"3B",X"B4",
		X"3A",X"3A",X"B0",X"C6",X"80",X"32",X"3A",X"B0",X"3A",X"3D",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"3D",X"B4",
		X"3A",X"3C",X"B0",X"C6",X"80",X"32",X"3C",X"B0",X"3A",X"3F",X"B4",X"CB",X"7F",X"28",X"19",X"4F",
		X"3A",X"00",X"C0",X"81",X"30",X"F2",X"23",X"23",X"2B",X"2B",X"79",X"E6",X"7F",X"32",X"3F",X"B4",
		X"3A",X"3E",X"B0",X"C6",X"80",X"32",X"3E",X"B0",X"C9",X"CD",X"B4",X"31",X"CD",X"DF",X"1E",X"CD",
		X"E3",X"23",X"CD",X"AF",X"36",X"CD",X"97",X"0F",X"CD",X"B3",X"47",X"CD",X"B7",X"43",X"CD",X"A1",
		X"28",X"CD",X"97",X"0F",X"CD",X"BC",X"2C",X"CD",X"D6",X"40",X"CD",X"97",X"0F",X"CD",X"5F",X"3B",
		X"CD",X"DA",X"3D",X"CD",X"36",X"3E",X"CD",X"97",X"0F",X"CD",X"EA",X"3F",X"CD",X"4F",X"4E",X"CD",
		X"B8",X"40",X"CD",X"97",X"0F",X"CD",X"DE",X"4D",X"CD",X"05",X"52",X"CD",X"3A",X"4D",X"CD",X"09",
		X"08",X"CD",X"98",X"10",X"3A",X"00",X"A8",X"3C",X"CA",X"71",X"12",X"3D",X"C0",X"CD",X"B6",X"15",
		X"3A",X"C6",X"AC",X"A7",X"C4",X"B8",X"2D",X"CD",X"34",X"56",X"21",X"00",X"AD",X"35",X"F5",X"3A",
		X"32",X"AD",X"A7",X"11",X"10",X"AD",X"28",X"03",X"11",X"20",X"AD",X"21",X"00",X"AD",X"01",X"10",
		X"00",X"ED",X"B0",X"F1",X"28",X"3D",X"3A",X"32",X"AD",X"A7",X"21",X"20",X"AD",X"28",X"03",X"21",
		X"10",X"AD",X"7E",X"A7",X"28",X"09",X"3A",X"32",X"AD",X"3C",X"E6",X"01",X"32",X"32",X"AD",X"3E",
		X"5A",X"32",X"EB",X"A9",X"3A",X"52",X"4B",X"32",X"AC",X"A9",X"C9",X"18",X"A7",X"13",X"A5",X"3B",
		X"87",X"F1",X"34",X"0E",X"34",X"D7",X"BF",X"F1",X"7F",X"13",X"13",X"13",X"13",X"F1",X"88",X"DC",
		X"ED",X"11",X"B9",X"3A",X"30",X"AD",X"A7",X"CA",X"FB",X"12",X"11",X"09",X"02",X"3A",X"32",X"AD",
		X"A7",X"28",X"01",X"1C",X"FF",X"11",X"0B",X"0A",X"FF",X"3E",X"B4",X"32",X"EB",X"A9",X"C3",X"1A",
		X"0F",X"3A",X"02",X"AD",X"A7",X"C0",X"3A",X"C6",X"AC",X"A7",X"C8",X"21",X"10",X"A8",X"11",X"10",
		X"00",X"06",X"0F",X"7E",X"A7",X"C0",X"19",X"10",X"FA",X"CD",X"34",X"56",X"3A",X"30",X"AD",X"A7",
		X"28",X"29",X"21",X"43",X"AA",X"06",X"17",X"AF",X"77",X"2C",X"2C",X"10",X"FB",X"CD",X"B8",X"2D",
		X"3A",X"32",X"AD",X"A7",X"11",X"10",X"AD",X"28",X"03",X"11",X"20",X"AD",X"21",X"00",X"AD",X"01",
		X"10",X"00",X"ED",X"B0",X"3A",X"35",X"4A",X"32",X"AC",X"A9",X"C9",X"3A",X"D1",X"07",X"32",X"C6",
		X"AC",X"CD",X"B6",X"15",X"C3",X"FB",X"12",X"74",X"B1",X"CC",X"EC",X"5C",X"16",X"39",X"50",X"67",
		X"21",X"7A",X"C5",X"F7",X"BE",X"54",X"80",X"2F",X"5F",X"9F",X"6D",X"44",X"B8",X"E7",X"BD",X"89",
		X"59",X"1A",X"21",X"EB",X"A9",X"35",X"C0",X"3A",X"32",X"AD",X"A7",X"21",X"20",X"AD",X"28",X"03",
		X"21",X"10",X"AD",X"7E",X"A7",X"C2",X"26",X"12",X"C3",X"1A",X"0F",X"AF",X"32",X"30",X"AD",X"32",
		X"AC",X"A9",X"32",X"32",X"AD",X"3A",X"D3",X"16",X"32",X"AB",X"A9",X"3A",X"01",X"49",X"2A",X"02",
		X"49",X"DF",X"AC",X"D6",X"9B",X"32",X"AC",X"A9",X"C9",X"11",X"E0",X"FF",X"06",X"0D",X"77",X"19",
		X"10",X"FC",X"C9",X"3A",X"80",X"A9",X"E6",X"02",X"C0",X"3A",X"F0",X"A9",X"A7",X"20",X"04",X"CD",
		X"67",X"13",X"C9",X"3D",X"20",X"07",X"CD",X"67",X"13",X"CD",X"2A",X"14",X"C9",X"3D",X"20",X"07",
		X"CD",X"93",X"13",X"CD",X"C5",X"14",X"C9",X"3D",X"20",X"04",X"CD",X"C5",X"14",X"C9",X"3D",X"20",
		X"04",X"CD",X"CC",X"13",X"C9",X"3E",X"5A",X"32",X"EB",X"A9",X"CD",X"B6",X"15",X"CD",X"75",X"4C",
		X"3A",X"50",X"27",X"32",X"AC",X"A9",X"C9",X"3A",X"F1",X"A9",X"FE",X"08",X"20",X"08",X"3E",X"01",
		X"32",X"F0",X"A9",X"CD",X"11",X"58",X"3A",X"F1",X"A9",X"E6",X"01",X"3E",X"3E",X"28",X"02",X"3E",
		X"00",X"47",X"3A",X"40",X"AA",X"E6",X"C0",X"80",X"32",X"40",X"AA",X"3A",X"F1",X"A9",X"3C",X"32",
		X"F1",X"A9",X"C9",X"3A",X"F3",X"A9",X"A7",X"20",X"09",X"3E",X"03",X"32",X"F0",X"A9",X"3E",X"3F",
		X"18",X"18",X"E6",X"04",X"20",X"04",X"3E",X"3F",X"18",X"10",X"3D",X"20",X"04",X"3E",X"36",X"18",
		X"09",X"3D",X"20",X"04",X"3E",X"3E",X"18",X"02",X"3E",X"37",X"47",X"3A",X"40",X"AA",X"E6",X"C0",
		X"80",X"32",X"40",X"AA",X"3A",X"F3",X"A9",X"3D",X"32",X"F3",X"A9",X"C9",X"3E",X"05",X"32",X"F0",
		X"A9",X"3A",X"32",X"AD",X"A7",X"3A",X"1C",X"AD",X"47",X"28",X"04",X"3A",X"2C",X"AD",X"47",X"3A",
		X"87",X"A9",X"A7",X"78",X"28",X"22",X"21",X"44",X"A0",X"11",X"45",X"A0",X"D9",X"06",X"1C",X"D9",
		X"01",X"1A",X"00",X"77",X"ED",X"B0",X"11",X"06",X"00",X"19",X"54",X"5D",X"13",X"D9",X"10",X"EF",
		X"3A",X"F6",X"A9",X"3D",X"32",X"F6",X"A9",X"C9",X"21",X"BE",X"A3",X"11",X"BD",X"A3",X"D9",X"06",
		X"1C",X"D9",X"01",X"1A",X"00",X"77",X"ED",X"B8",X"11",X"FA",X"FF",X"19",X"54",X"5D",X"1B",X"D9",
		X"10",X"EF",X"3A",X"F6",X"A9",X"3D",X"32",X"F6",X"A9",X"C9",X"3A",X"F2",X"A9",X"CB",X"47",X"28",
		X"6C",X"2A",X"F7",X"A9",X"7E",X"FE",X"FF",X"20",X"12",X"3E",X"00",X"32",X"F2",X"A9",X"3E",X"02",
		X"32",X"F0",X"A9",X"2A",X"F7",X"A9",X"2B",X"22",X"F7",X"A9",X"C9",X"CD",X"63",X"15",X"2A",X"F7",
		X"A9",X"7E",X"E6",X"01",X"23",X"22",X"F7",X"A9",X"28",X"0F",X"11",X"20",X"00",X"21",X"F0",X"A5",
		X"34",X"19",X"34",X"21",X"F2",X"A5",X"34",X"19",X"34",X"2A",X"F7",X"A9",X"7E",X"E6",X"01",X"23",
		X"22",X"F7",X"A9",X"28",X"09",X"11",X"20",X"00",X"21",X"F1",X"A5",X"34",X"19",X"34",X"0E",X"02",
		X"11",X"D1",X"A5",X"CD",X"9D",X"4A",X"2A",X"F7",X"A9",X"11",X"F3",X"FF",X"19",X"22",X"F7",X"A9",
		X"0E",X"00",X"11",X"31",X"A6",X"CD",X"9D",X"4A",X"CD",X"8C",X"15",X"18",X"20",X"3E",X"F1",X"21",
		X"B1",X"A7",X"CD",X"19",X"13",X"21",X"D1",X"A5",X"CD",X"19",X"13",X"21",X"10",X"A6",X"77",X"19",
		X"77",X"21",X"11",X"A6",X"77",X"19",X"77",X"21",X"12",X"A6",X"77",X"19",X"77",X"3A",X"F2",X"A9",
		X"3D",X"32",X"F2",X"A9",X"C9",X"3A",X"F4",X"A9",X"CB",X"47",X"28",X"6F",X"2A",X"F7",X"A9",X"7E",
		X"E6",X"FE",X"28",X"15",X"3E",X"00",X"32",X"F4",X"A9",X"3E",X"04",X"32",X"F0",X"A9",X"CD",X"E4",
		X"56",X"2A",X"F7",X"A9",X"23",X"22",X"F7",X"A9",X"C9",X"CD",X"63",X"15",X"0E",X"01",X"11",X"51",
		X"A4",X"CD",X"9D",X"4A",X"2A",X"F7",X"A9",X"11",X"0D",X"00",X"19",X"22",X"F7",X"A9",X"0E",X"03",
		X"11",X"B1",X"A7",X"CD",X"9D",X"4A",X"2A",X"F7",X"A9",X"7E",X"E6",X"01",X"2B",X"22",X"F7",X"A9",
		X"28",X"09",X"11",X"20",X"00",X"21",X"F1",X"A5",X"35",X"19",X"35",X"2A",X"F7",X"A9",X"7E",X"E6",
		X"01",X"2B",X"22",X"F7",X"A9",X"28",X"0F",X"11",X"20",X"00",X"21",X"F0",X"A5",X"35",X"19",X"35",
		X"21",X"F2",X"A5",X"35",X"19",X"35",X"CD",X"8C",X"15",X"18",X"20",X"3E",X"F1",X"21",X"B1",X"A7",
		X"CD",X"19",X"13",X"21",X"D1",X"A5",X"CD",X"19",X"13",X"21",X"10",X"A6",X"77",X"19",X"77",X"21",
		X"11",X"A6",X"77",X"19",X"77",X"21",X"12",X"A6",X"77",X"19",X"77",X"3A",X"F4",X"A9",X"3D",X"32",
		X"F4",X"A9",X"C9",X"11",X"00",X"A4",X"21",X"51",X"A4",X"01",X"20",X"00",X"D9",X"06",X"1C",X"D9",
		X"1A",X"77",X"13",X"09",X"D9",X"10",X"F8",X"D9",X"21",X"F0",X"A5",X"1A",X"77",X"09",X"13",X"1A",
		X"77",X"13",X"21",X"F2",X"A5",X"1A",X"77",X"09",X"13",X"1A",X"77",X"C9",X"11",X"00",X"A4",X"21",
		X"51",X"A4",X"01",X"20",X"00",X"D9",X"06",X"1C",X"D9",X"7E",X"12",X"13",X"09",X"D9",X"10",X"F8",
		X"D9",X"21",X"F0",X"A5",X"7E",X"12",X"09",X"13",X"7E",X"12",X"13",X"21",X"F2",X"A5",X"7E",X"12",
		X"09",X"13",X"7E",X"12",X"C9",X"C9",X"21",X"41",X"AA",X"06",X"18",X"AF",X"77",X"2C",X"2C",X"10",
		X"FB",X"C9",X"3A",X"AC",X"A9",X"E6",X"07",X"F7",X"E2",X"15",X"5F",X"A5",X"13",X"77",X"D7",X"34",
		X"87",X"FD",X"DC",X"B9",X"FE",X"15",X"60",X"A6",X"14",X"C4",X"FD",X"10",X"ED",X"77",X"68",X"D7",
		X"34",X"B9",X"CD",X"9A",X"01",X"3A",X"49",X"17",X"32",X"AC",X"A9",X"0E",X"00",X"21",X"48",X"56",
		X"3A",X"AB",X"A9",X"96",X"23",X"0D",X"20",X"FB",X"EE",X"4E",X"32",X"AB",X"A9",X"C9",X"CD",X"C2",
		X"01",X"C0",X"11",X"05",X"01",X"FF",X"1C",X"FF",X"1C",X"FF",X"11",X"01",X"06",X"FF",X"3E",X"13",
		X"32",X"01",X"A7",X"32",X"E1",X"A6",X"21",X"3F",X"16",X"06",X"06",X"5E",X"23",X"56",X"23",X"7E",
		X"12",X"13",X"EB",X"36",X"05",X"EB",X"23",X"10",X"F2",X"CD",X"6B",X"0D",X"3E",X"01",X"32",X"AB",
		X"A9",X"3C",X"32",X"AC",X"A9",X"3A",X"C0",X"A9",X"A7",X"C8",X"11",X"0D",X"01",X"FF",X"C9",X"FB",
		X"AD",X"FD",X"39",X"AD",X"68",X"43",X"AB",X"7C",X"FE",X"AB",X"A5",X"BE",X"AC",X"38",X"C7",X"AC",
		X"3B",X"21",X"7B",X"16",X"E5",X"3A",X"AC",X"A9",X"F7",X"4B",X"07",X"34",X"17",X"3F",X"2D",X"3E",
		X"08",X"48",X"17",X"6A",X"17",X"8C",X"17",X"B9",X"17",X"52",X"32",X"E2",X"17",X"19",X"4B",X"FB",
		X"17",X"30",X"27",X"26",X"A6",X"13",X"88",X"57",X"A5",X"BF",X"B9",X"3A",X"86",X"A9",X"A7",X"C2",
		X"11",X"0F",X"3A",X"C0",X"A9",X"A7",X"C8",X"3A",X"AE",X"A9",X"E6",X"18",X"C8",X"CD",X"B6",X"15",
		X"3A",X"AE",X"A9",X"CB",X"67",X"20",X"05",X"CB",X"5F",X"20",X"7E",X"C9",X"3E",X"FF",X"32",X"30",
		X"AD",X"32",X"31",X"AD",X"3A",X"C1",X"A9",X"32",X"10",X"AD",X"32",X"20",X"AD",X"18",X"7B",X"06",
		X"00",X"21",X"9F",X"4D",X"3A",X"AB",X"A9",X"96",X"23",X"10",X"FC",X"EE",X"A2",X"32",X"AB",X"A9",
		X"CD",X"97",X"0F",X"CD",X"DF",X"1E",X"CD",X"97",X"0F",X"CD",X"BC",X"2C",X"CD",X"98",X"10",X"3A",
		X"80",X"A9",X"E6",X"01",X"28",X"1C",X"21",X"EB",X"A9",X"35",X"20",X"16",X"11",X"09",X"03",X"FF",
		X"1E",X"0E",X"FF",X"1E",X"1A",X"FF",X"AF",X"32",X"0E",X"AD",X"3E",X"2A",X"32",X"EB",X"A9",X"C3",
		X"1A",X"0F",X"3A",X"0E",X"AD",X"A7",X"C8",X"3A",X"80",X"A9",X"E6",X"0F",X"28",X"09",X"FE",X"05",
		X"28",X"09",X"FE",X"0A",X"28",X"09",X"C9",X"16",X"02",X"18",X"06",X"16",X"0A",X"18",X"02",X"16",
		X"0B",X"3A",X"04",X"AD",X"C6",X"1A",X"5F",X"FF",X"C9",X"AF",X"32",X"31",X"AD",X"32",X"20",X"AD",
		X"3D",X"32",X"30",X"AD",X"3A",X"C1",X"A9",X"32",X"10",X"AD",X"3E",X"03",X"32",X"AB",X"A9",X"AF",
		X"32",X"AC",X"A9",X"C9",X"CD",X"01",X"02",X"C0",X"21",X"48",X"17",X"06",X"22",X"AF",X"96",X"23",
		X"10",X"FC",X"32",X"17",X"A8",X"C3",X"1A",X"0F",X"CD",X"06",X"0B",X"CD",X"39",X"0B",X"21",X"EB",
		X"A9",X"35",X"C0",X"21",X"3C",X"A6",X"11",X"C7",X"AC",X"7E",X"12",X"13",X"CB",X"94",X"7E",X"12",
		X"11",X"03",X"03",X"FF",X"1C",X"FF",X"C3",X"1A",X"0F",X"31",X"CD",X"DA",X"19",X"3A",X"7C",X"A6",
		X"FE",X"7C",X"C2",X"9B",X"45",X"11",X"13",X"01",X"FF",X"CD",X"DC",X"4B",X"21",X"DC",X"A5",X"11",
		X"FB",X"AD",X"7E",X"12",X"13",X"CB",X"94",X"7E",X"12",X"C3",X"1A",X"0F",X"CD",X"06",X"0B",X"CD",
		X"39",X"0B",X"21",X"EB",X"A9",X"35",X"C0",X"CD",X"DA",X"19",X"3A",X"B3",X"47",X"C6",X"02",X"6F",
		X"C6",X"6A",X"67",X"7E",X"FE",X"3B",X"C2",X"CA",X"15",X"21",X"7C",X"A6",X"11",X"43",X"AB",X"7E",
		X"12",X"13",X"CB",X"94",X"7E",X"12",X"C3",X"1A",X"0F",X"3A",X"0D",X"59",X"4F",X"3A",X"40",X"4A",
		X"21",X"06",X"0B",X"06",X"33",X"86",X"23",X"10",X"FC",X"FE",X"EF",X"CA",X"1A",X"0F",X"3A",X"89",
		X"4C",X"32",X"08",X"C3",X"21",X"5C",X"A6",X"11",X"39",X"AD",X"7E",X"12",X"13",X"CB",X"94",X"7E",
		X"12",X"C9",X"3E",X"FF",X"32",X"3F",X"AA",X"11",X"B9",X"17",X"0E",X"08",X"CD",X"D9",X"4B",X"3A",
		X"C0",X"27",X"CD",X"1E",X"29",X"32",X"6F",X"AA",X"C3",X"1A",X"0F",X"C3",X"1A",X"0F",X"21",X"1D",
		X"18",X"E5",X"3A",X"AC",X"A9",X"F7",X"1E",X"18",X"DB",X"2C",X"30",X"18",X"E6",X"07",X"8A",X"18",
		X"72",X"A6",X"14",X"7D",X"A5",X"38",X"34",X"F1",X"68",X"0E",X"34",X"D7",X"B9",X"C9",X"CD",X"B6",
		X"15",X"21",X"FC",X"A5",X"11",X"BE",X"AC",X"CD",X"FC",X"1A",X"CD",X"B5",X"01",X"C3",X"1A",X"0F",
		X"CD",X"06",X"0B",X"CD",X"39",X"0B",X"11",X"01",X"01",X"FF",X"1E",X"14",X"FF",X"1C",X"FF",X"1E",
		X"0F",X"3A",X"C3",X"A9",X"A7",X"28",X"02",X"1C",X"1C",X"FF",X"1C",X"FF",X"1E",X"16",X"FF",X"1E",
		X"00",X"FF",X"3A",X"86",X"A9",X"FE",X"02",X"30",X"07",X"11",X"17",X"01",X"FF",X"C3",X"1A",X"0F",
		X"11",X"19",X"01",X"FF",X"CD",X"1A",X"0F",X"C3",X"1A",X"0F",X"00",X"02",X"06",X"0D",X"00",X"03",
		X"07",X"0C",X"00",X"04",X"08",X"0B",X"02",X"06",X"0A",X"0A",X"04",X"08",X"0C",X"09",X"07",X"0A",
		X"0D",X"07",X"0B",X"0D",X"0E",X"05",X"0F",X"0F",X"0F",X"05",X"CD",X"06",X"0B",X"CD",X"39",X"0B",
		X"3A",X"AE",X"A9",X"CB",X"67",X"C2",X"9E",X"18",X"CB",X"5F",X"C2",X"15",X"32",X"C9",X"CD",X"2B",
		X"0B",X"3E",X"FF",X"32",X"30",X"AD",X"32",X"31",X"AD",X"3A",X"C1",X"A9",X"32",X"10",X"AD",X"32",
		X"20",X"AD",X"CD",X"0E",X"46",X"21",X"86",X"A9",X"7E",X"D6",X"02",X"27",X"77",X"CD",X"FB",X"4A",
		X"C3",X"2A",X"17",X"3A",X"80",X"A9",X"E6",X"01",X"C2",X"84",X"19",X"CD",X"D1",X"1E",X"21",X"95",
		X"A9",X"0F",X"CB",X"16",X"23",X"0F",X"CB",X"16",X"23",X"0F",X"0F",X"0F",X"CB",X"16",X"23",X"0F",
		X"CB",X"16",X"7E",X"E6",X"07",X"3D",X"28",X"3B",X"2B",X"7E",X"E6",X"07",X"3D",X"28",X"34",X"2B",
		X"7E",X"FE",X"FF",X"CC",X"80",X"19",X"E6",X"07",X"3D",X"28",X"1B",X"2B",X"7E",X"FE",X"7F",X"CC",
		X"80",X"19",X"E6",X"07",X"3D",X"28",X"02",X"18",X"5A",X"21",X"99",X"A9",X"35",X"7E",X"FE",X"80",
		X"38",X"3C",X"36",X"1A",X"18",X"38",X"21",X"99",X"A9",X"34",X"7E",X"FE",X"1B",X"38",X"2F",X"36",
		X"00",X"18",X"2B",X"3A",X"99",X"A9",X"21",X"C7",X"12",X"CF",X"2A",X"91",X"A9",X"ED",X"5B",X"93",
		X"A9",X"12",X"77",X"3A",X"90",X"A9",X"CB",X"92",X"12",X"CB",X"D2",X"E7",X"23",X"22",X"91",X"A9",
		X"ED",X"53",X"93",X"A9",X"21",X"9A",X"A9",X"35",X"28",X"2B",X"AF",X"32",X"99",X"A9",X"ED",X"5B",
		X"93",X"A9",X"3A",X"99",X"A9",X"21",X"C7",X"12",X"CF",X"12",X"CB",X"92",X"3E",X"10",X"12",X"AF",
		X"32",X"9C",X"A9",X"3A",X"80",X"A9",X"E6",X"07",X"20",X"30",X"21",X"EB",X"A9",X"35",X"20",X"2A",
		X"2A",X"93",X"A9",X"36",X"F1",X"3E",X"3C",X"32",X"EB",X"A9",X"CD",X"34",X"56",X"C3",X"1A",X"0F",
		X"36",X"00",X"AF",X"C9",X"21",X"9C",X"A9",X"34",X"2A",X"93",X"A9",X"CB",X"94",X"3A",X"9C",X"A9",
		X"CB",X"67",X"28",X"04",X"36",X"14",X"18",X"02",X"36",X"10",X"21",X"20",X"AD",X"3A",X"10",X"AD",
		X"B6",X"C0",X"3A",X"C0",X"A9",X"A7",X"20",X"26",X"3A",X"86",X"A9",X"FE",X"01",X"D8",X"28",X"10",
		X"3A",X"AE",X"A9",X"E6",X"18",X"C8",X"FE",X"08",X"28",X"0E",X"CD",X"B6",X"15",X"C3",X"9E",X"18",
		X"3A",X"AE",X"A9",X"E6",X"18",X"FE",X"08",X"C0",X"CD",X"B6",X"15",X"C3",X"15",X"32",X"3A",X"AE",
		X"A9",X"E6",X"18",X"C8",X"CD",X"B6",X"15",X"C3",X"90",X"16",X"21",X"BC",X"A2",X"06",X"0D",X"7E",
		X"FE",X"10",X"28",X"05",X"FE",X"05",X"C2",X"FA",X"49",X"11",X"E0",X"FF",X"19",X"10",X"F0",X"C9",
		X"21",X"00",X"00",X"22",X"08",X"A8",X"22",X"0A",X"A8",X"22",X"06",X"AD",X"AF",X"32",X"0D",X"AD",
		X"32",X"F7",X"A8",X"32",X"05",X"AD",X"3A",X"D6",X"A9",X"32",X"D7",X"A9",X"3A",X"0A",X"AD",X"32",
		X"C0",X"AC",X"AF",X"32",X"81",X"AA",X"32",X"C6",X"AC",X"3E",X"80",X"32",X"02",X"A8",X"AF",X"32",
		X"01",X"A8",X"3E",X"FF",X"32",X"00",X"A8",X"3E",X"78",X"32",X"41",X"AA",X"3E",X"84",X"32",X"10",
		X"AA",X"CD",X"AF",X"20",X"CD",X"55",X"27",X"DD",X"21",X"C0",X"A8",X"FD",X"21",X"28",X"AA",X"CD",
		X"0D",X"3C",X"06",X"07",X"DD",X"21",X"50",X"A8",X"FD",X"21",X"1A",X"AA",X"DD",X"21",X"E0",X"A8",
		X"FD",X"21",X"2C",X"AA",X"CD",X"FB",X"3D",X"DD",X"21",X"F0",X"A8",X"FD",X"21",X"2E",X"AA",X"CD",
		X"AD",X"48",X"CD",X"DE",X"2B",X"11",X"10",X"00",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"10",X"F2",
		X"CD",X"E4",X"1A",X"FD",X"21",X"28",X"AA",X"FD",X"36",X"00",X"00",X"FD",X"36",X"02",X"00",X"FD",
		X"36",X"04",X"00",X"FD",X"36",X"06",X"00",X"FD",X"36",X"31",X"00",X"FD",X"36",X"33",X"00",X"FD",
		X"36",X"35",X"00",X"FD",X"36",X"37",X"00",X"CD",X"A5",X"30",X"3A",X"04",X"AD",X"07",X"07",X"07",
		X"07",X"E6",X"F0",X"47",X"3A",X"C0",X"AC",X"80",X"21",X"04",X"1B",X"D7",X"1A",X"32",X"44",X"A8",
		X"13",X"1A",X"32",X"37",X"A8",X"13",X"1A",X"32",X"27",X"A8",X"13",X"1A",X"32",X"17",X"A8",X"32",
		X"14",X"A8",X"13",X"1A",X"32",X"C1",X"AC",X"13",X"1A",X"32",X"C4",X"AC",X"13",X"1A",X"32",X"C6",
		X"A8",X"13",X"1A",X"32",X"D6",X"A8",X"13",X"1A",X"32",X"E6",X"A8",X"13",X"1A",X"32",X"F4",X"A8",
		X"32",X"F6",X"A8",X"C9",X"DD",X"21",X"10",X"A8",X"3E",X"01",X"06",X"17",X"11",X"10",X"00",X"DD",
		X"36",X"00",X"00",X"DD",X"77",X"0F",X"3C",X"DD",X"19",X"10",X"F4",X"C9",X"7E",X"12",X"13",X"CB",
		X"94",X"7E",X"12",X"C9",X"B1",X"1B",X"BB",X"1B",X"C5",X"1B",X"CF",X"1B",X"D9",X"1B",X"E3",X"1B",
		X"ED",X"1B",X"F7",X"1B",X"01",X"1C",X"0B",X"1C",X"15",X"1C",X"1F",X"1C",X"29",X"1C",X"33",X"1C",
		X"3D",X"1C",X"47",X"1C",X"51",X"1C",X"5B",X"1C",X"65",X"1C",X"6F",X"1C",X"79",X"1C",X"83",X"1C",
		X"8D",X"1C",X"97",X"1C",X"A1",X"1C",X"AB",X"1C",X"B5",X"1C",X"BF",X"1C",X"C9",X"1C",X"D3",X"1C",
		X"DD",X"1C",X"E7",X"1C",X"F1",X"1C",X"FB",X"1C",X"05",X"1D",X"0F",X"1D",X"19",X"1D",X"23",X"1D",
		X"2D",X"1D",X"37",X"1D",X"41",X"1D",X"4B",X"1D",X"55",X"1D",X"5F",X"1D",X"69",X"1D",X"73",X"1D",
		X"7D",X"1D",X"87",X"1D",X"91",X"1D",X"9B",X"1D",X"A5",X"1D",X"AF",X"1D",X"B9",X"1D",X"C3",X"1D",
		X"CD",X"1D",X"D7",X"1D",X"E1",X"1D",X"EB",X"1D",X"F5",X"1D",X"FF",X"1D",X"09",X"1E",X"13",X"1E",
		X"1D",X"1E",X"27",X"1E",X"31",X"1E",X"3B",X"1E",X"45",X"1E",X"4F",X"1E",X"59",X"1E",X"63",X"1E",
		X"6D",X"1E",X"77",X"1E",X"81",X"1E",X"8B",X"1E",X"95",X"1E",X"9F",X"1E",X"A9",X"1E",X"B3",X"1E",
		X"BD",X"1E",X"C7",X"1E",X"5F",X"A5",X"13",X"00",X"D7",X"34",X"34",X"F1",X"88",X"57",X"A5",X"BF",
		X"B9",X"00",X"20",X"50",X"3C",X"04",X"50",X"00",X"50",X"18",X"5A",X"01",X"20",X"4E",X"3C",X"04",
		X"50",X"00",X"4E",X"18",X"54",X"01",X"28",X"4C",X"32",X"05",X"60",X"01",X"4C",X"1C",X"4E",X"02",
		X"28",X"48",X"28",X"05",X"60",X"01",X"48",X"1C",X"48",X"02",X"30",X"46",X"1E",X"06",X"70",X"01",
		X"46",X"1C",X"42",X"03",X"30",X"44",X"1E",X"06",X"70",X"02",X"44",X"20",X"3C",X"03",X"38",X"42",
		X"1E",X"06",X"80",X"02",X"42",X"20",X"36",X"03",X"38",X"40",X"1E",X"06",X"80",X"02",X"40",X"20",
		X"30",X"04",X"40",X"3F",X"1E",X"07",X"90",X"03",X"3F",X"24",X"2A",X"04",X"40",X"3E",X"1E",X"07",
		X"90",X"03",X"3E",X"24",X"24",X"04",X"40",X"3D",X"1E",X"07",X"A0",X"03",X"3D",X"24",X"1E",X"04",
		X"40",X"3C",X"1E",X"07",X"B0",X"03",X"3C",X"28",X"1E",X"04",X"48",X"3B",X"1E",X"07",X"C0",X"03",
		X"3B",X"28",X"1E",X"04",X"48",X"3A",X"1E",X"07",X"D0",X"03",X"3A",X"2C",X"1E",X"04",X"48",X"39",
		X"1E",X"07",X"E0",X"03",X"39",X"30",X"1E",X"04",X"48",X"38",X"19",X"07",X"F0",X"03",X"38",X"30",
		X"19",X"01",X"28",X"48",X"32",X"05",X"50",X"01",X"5C",X"00",X"1E",X"01",X"28",X"48",X"28",X"05",
		X"50",X"01",X"5A",X"00",X"1E",X"02",X"30",X"48",X"1E",X"05",X"60",X"01",X"58",X"00",X"1E",X"02",
		X"30",X"48",X"1E",X"06",X"60",X"01",X"56",X"00",X"1E",X"02",X"30",X"48",X"1E",X"06",X"70",X"02",
		X"54",X"00",X"1E",X"03",X"38",X"40",X"1E",X"06",X"70",X"02",X"52",X"00",X"1E",X"03",X"38",X"40",
		X"1E",X"06",X"80",X"02",X"50",X"00",X"1E",X"03",X"38",X"40",X"1E",X"06",X"80",X"02",X"4C",X"00",
		X"1E",X"04",X"40",X"40",X"1E",X"07",X"90",X"02",X"4C",X"00",X"1E",X"04",X"40",X"40",X"1E",X"07",
		X"90",X"02",X"48",X"00",X"1E",X"04",X"48",X"38",X"1E",X"07",X"A0",X"02",X"48",X"00",X"1E",X"04",
		X"48",X"38",X"1E",X"07",X"B0",X"02",X"48",X"00",X"1E",X"04",X"48",X"38",X"1E",X"07",X"C0",X"02",
		X"48",X"00",X"1E",X"04",X"48",X"38",X"1E",X"07",X"D0",X"02",X"48",X"00",X"1E",X"04",X"50",X"38",
		X"1E",X"07",X"E0",X"02",X"48",X"00",X"1E",X"04",X"58",X"30",X"19",X"07",X"F0",X"02",X"48",X"00",
		X"19",X"01",X"20",X"50",X"32",X"03",X"50",X"01",X"50",X"08",X"1E",X"01",X"20",X"50",X"28",X"04",
		X"50",X"01",X"50",X"08",X"1E",X"01",X"20",X"50",X"1E",X"04",X"60",X"01",X"50",X"0C",X"1E",X"01",
		X"28",X"50",X"1E",X"04",X"60",X"02",X"50",X"0C",X"1E",X"01",X"28",X"48",X"1E",X"05",X"70",X"02",
		X"48",X"10",X"1E",X"01",X"28",X"48",X"1E",X"05",X"80",X"02",X"48",X"10",X"1E",X"01",X"30",X"48",
		X"1E",X"05",X"90",X"03",X"48",X"14",X"1E",X"01",X"30",X"48",X"1E",X"06",X"A0",X"03",X"48",X"14",
		X"1E",X"02",X"30",X"40",X"1E",X"06",X"B0",X"03",X"40",X"18",X"1E",X"02",X"38",X"40",X"1E",X"06",
		X"C0",X"03",X"40",X"18",X"1E",X"02",X"38",X"40",X"1E",X"06",X"D0",X"03",X"40",X"18",X"1E",X"02",
		X"38",X"40",X"1E",X"06",X"D0",X"03",X"40",X"18",X"1E",X"02",X"40",X"38",X"1E",X"06",X"E0",X"03",
		X"38",X"18",X"1E",X"02",X"48",X"38",X"1E",X"06",X"E0",X"03",X"38",X"18",X"1E",X"02",X"50",X"38",
		X"1E",X"06",X"F0",X"03",X"38",X"18",X"1E",X"03",X"58",X"30",X"19",X"07",X"F0",X"03",X"30",X"18",
		X"19",X"01",X"20",X"50",X"1E",X"04",X"60",X"01",X"50",X"00",X"1E",X"01",X"20",X"50",X"1E",X"04",
		X"70",X"01",X"50",X"00",X"1E",X"01",X"28",X"50",X"1E",X"04",X"80",X"01",X"50",X"00",X"1E",X"01",
		X"28",X"50",X"1E",X"05",X"90",X"02",X"50",X"00",X"1E",X"01",X"30",X"48",X"1E",X"05",X"A0",X"02",
		X"48",X"00",X"1E",X"01",X"30",X"48",X"1E",X"05",X"B0",X"02",X"48",X"00",X"1E",X"01",X"38",X"48",
		X"1E",X"05",X"C0",X"03",X"48",X"00",X"1E",X"01",X"38",X"48",X"1E",X"06",X"D0",X"03",X"48",X"00",
		X"1E",X"01",X"40",X"40",X"1E",X"06",X"E0",X"03",X"40",X"00",X"1E",X"01",X"40",X"40",X"1E",X"06",
		X"F0",X"03",X"40",X"00",X"1E",X"01",X"48",X"40",X"1E",X"06",X"F0",X"03",X"40",X"00",X"1E",X"01",
		X"48",X"40",X"1E",X"06",X"F0",X"03",X"40",X"00",X"1E",X"01",X"50",X"38",X"1E",X"06",X"F0",X"03",
		X"38",X"00",X"1E",X"01",X"50",X"38",X"1E",X"06",X"F0",X"03",X"38",X"00",X"1E",X"01",X"58",X"38",
		X"1E",X"06",X"F0",X"03",X"38",X"00",X"1E",X"01",X"58",X"30",X"19",X"06",X"F0",X"03",X"30",X"00",
		X"19",X"01",X"20",X"50",X"5A",X"03",X"00",X"01",X"58",X"3C",X"64",X"01",X"20",X"50",X"5A",X"03",
		X"10",X"01",X"54",X"46",X"5A",X"01",X"28",X"50",X"50",X"04",X"20",X"01",X"52",X"50",X"50",X"01",
		X"28",X"50",X"46",X"04",X"30",X"02",X"50",X"5A",X"46",X"01",X"30",X"48",X"46",X"04",X"40",X"02",
		X"4E",X"64",X"46",X"01",X"30",X"48",X"3C",X"05",X"50",X"02",X"4B",X"6E",X"3C",X"01",X"38",X"48",
		X"3C",X"05",X"60",X"03",X"48",X"78",X"3C",X"01",X"38",X"40",X"32",X"05",X"70",X"03",X"46",X"82",
		X"3C",X"01",X"40",X"40",X"32",X"05",X"80",X"03",X"44",X"8C",X"32",X"01",X"40",X"40",X"28",X"05",
		X"90",X"03",X"44",X"96",X"32",X"01",X"48",X"40",X"28",X"05",X"A0",X"03",X"42",X"A0",X"32",X"01",
		X"48",X"3C",X"1E",X"05",X"B0",X"03",X"42",X"AA",X"28",X"01",X"50",X"3C",X"1E",X"05",X"C0",X"03",
		X"40",X"B4",X"28",X"01",X"50",X"3C",X"1E",X"05",X"D0",X"03",X"3C",X"BE",X"28",X"01",X"58",X"38",
		X"1E",X"05",X"E0",X"03",X"38",X"C8",X"1E",X"01",X"58",X"30",X"19",X"05",X"F0",X"03",X"34",X"D2",
		X"19",X"3A",X"87",X"A9",X"A7",X"21",X"AF",X"A9",X"20",X"03",X"21",X"B0",X"A9",X"7E",X"C9",X"DD",
		X"21",X"00",X"A8",X"FD",X"21",X"10",X"AA",X"3A",X"00",X"A8",X"A7",X"C8",X"3C",X"C2",X"10",X"20",
		X"3A",X"30",X"AD",X"A7",X"CA",X"4B",X"21",X"CD",X"D1",X"1E",X"E6",X"0F",X"20",X"03",X"C3",X"42",
		X"1F",X"21",X"2E",X"1F",X"CF",X"47",X"3A",X"02",X"A8",X"90",X"CA",X"42",X"1F",X"4F",X"3A",X"04",
		X"AD",X"E6",X"0F",X"FE",X"03",X"30",X"04",X"16",X"03",X"18",X"02",X"16",X"04",X"79",X"C6",X"01",
		X"FE",X"03",X"DA",X"3E",X"1F",X"79",X"FE",X"80",X"D2",X"6F",X"1F",X"C3",X"68",X"1F",X"00",X"00",
		X"80",X"00",X"C0",X"E0",X"A0",X"00",X"40",X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"78",X"32",
		X"02",X"A8",X"21",X"55",X"1F",X"E5",X"3A",X"04",X"AD",X"A7",X"CA",X"4E",X"59",X"FE",X"03",X"DA",
		X"65",X"59",X"C3",X"6B",X"59",X"AF",X"67",X"6F",X"ED",X"52",X"22",X"08",X"A8",X"AF",X"67",X"6F",
		X"ED",X"42",X"22",X"0A",X"A8",X"C3",X"AF",X"20",X"92",X"80",X"32",X"02",X"A8",X"18",X"D3",X"82",
		X"80",X"32",X"02",X"A8",X"18",X"CC",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"DD",X"F1",X"F1",
		X"F1",X"F1",X"F0",X"F1",X"F1",X"F1",X"F1",X"C3",X"F1",X"F1",X"F1",X"F1",X"EA",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"B7",X"F1",X"F1",X"F1",X"F1",X"4D",X"F1",X"F1",X"F1",X"E5",
		X"2D",X"6E",X"F1",X"F1",X"5E",X"61",X"E6",X"F1",X"F1",X"F1",X"B2",X"F1",X"F1",X"F1",X"F1",X"53",
		X"F1",X"F1",X"F1",X"F1",X"95",X"F1",X"F1",X"F1",X"45",X"CA",X"F1",X"F1",X"F1",X"C6",X"2C",X"97",
		X"F1",X"F1",X"81",X"69",X"1E",X"F1",X"F1",X"BC",X"A1",X"60",X"F1",X"F1",X"F4",X"EB",X"F1",X"F1",
		X"F1",X"F1",X"48",X"F1",X"F1",X"F1",X"E0",X"63",X"35",X"F1",X"F1",X"AA",X"B4",X"8A",X"F1",X"F1",
		X"51",X"E9",X"F6",X"F1",X"F1",X"82",X"92",X"98",X"F1",X"F1",X"F1",X"46",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"19",X"DF",X"78",X"C9",
		X"DD",X"7E",X"00",X"FE",X"B4",X"38",X"29",X"DD",X"36",X"00",X"B4",X"FD",X"36",X"01",X"FF",X"3A",
		X"04",X"AD",X"FE",X"02",X"D4",X"79",X"56",X"CD",X"D2",X"56",X"3A",X"FE",X"AB",X"FE",X"A5",X"C2",
		X"63",X"20",X"11",X"FF",X"AB",X"1A",X"FE",X"05",X"CA",X"40",X"20",X"FE",X"10",X"C2",X"63",X"20",
		X"DD",X"35",X"00",X"DD",X"7E",X"00",X"FE",X"B3",X"28",X"1C",X"FE",X"AB",X"28",X"1D",X"FE",X"A3",
		X"28",X"1E",X"FE",X"9B",X"28",X"1F",X"FE",X"93",X"28",X"20",X"FE",X"8B",X"28",X"21",X"FE",X"83",
		X"28",X"22",X"C9",X"C3",X"2E",X"1F",X"11",X"76",X"1F",X"18",X"1E",X"11",X"94",X"1F",X"18",X"19",
		X"11",X"B2",X"1F",X"18",X"14",X"11",X"D0",X"1F",X"18",X"0F",X"11",X"D0",X"1F",X"18",X"0A",X"11",
		X"B2",X"1F",X"18",X"05",X"11",X"EE",X"1F",X"18",X"00",X"21",X"AF",X"A5",X"06",X"C1",X"3A",X"04",
		X"AD",X"80",X"4F",X"D9",X"3A",X"7A",X"33",X"47",X"D9",X"3A",X"02",X"49",X"47",X"1A",X"77",X"CB",
		X"94",X"71",X"CB",X"D4",X"23",X"13",X"10",X"F5",X"3E",X"1B",X"DF",X"D9",X"10",X"EA",X"C9",X"DD",
		X"21",X"00",X"A8",X"11",X"20",X"00",X"3A",X"02",X"A8",X"C6",X"04",X"0F",X"0F",X"0F",X"E6",X"1F",
		X"21",X"CE",X"20",X"DF",X"7E",X"32",X"11",X"AA",X"19",X"7E",X"32",X"40",X"AA",X"C9",X"F0",X"F1",
		X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"E8",X"F7",X"F6",X"F5",X"F4",X"F3",X"F2",X"F1",X"F0",X"EF",
		X"EE",X"ED",X"EC",X"EB",X"EA",X"E9",X"E8",X"E9",X"EA",X"EB",X"EC",X"ED",X"EE",X"EF",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"21",X"F3",
		X"AD",X"EB",X"3A",X"14",X"AD",X"A7",X"28",X"28",X"FE",X"03",X"28",X"24",X"FE",X"01",X"28",X"25",
		X"21",X"FA",X"22",X"7E",X"3C",X"32",X"F2",X"AD",X"EB",X"73",X"2C",X"72",X"21",X"FB",X"AD",X"7E",
		X"FE",X"FD",X"C2",X"3D",X"21",X"23",X"7E",X"FE",X"10",X"C8",X"FE",X"05",X"C8",X"C3",X"51",X"22",
		X"21",X"8C",X"21",X"18",X"DE",X"21",X"51",X"22",X"18",X"D9",X"C9",X"21",X"F2",X"AD",X"7E",X"47",
		X"E6",X"3F",X"28",X"07",X"3D",X"28",X"04",X"05",X"70",X"18",X"0F",X"23",X"5E",X"23",X"56",X"13",
		X"72",X"2B",X"73",X"EB",X"7E",X"1B",X"3C",X"12",X"18",X"E1",X"78",X"D9",X"07",X"07",X"E6",X"03",
		X"CA",X"42",X"1F",X"3D",X"28",X"0B",X"3A",X"02",X"A8",X"C6",X"03",X"32",X"02",X"A8",X"C3",X"42",
		X"1F",X"3A",X"02",X"A8",X"D6",X"03",X"32",X"02",X"A8",X"C3",X"42",X"1F",X"3C",X"3C",X"3C",X"3C",
		X"0B",X"95",X"03",X"66",X"95",X"7C",X"59",X"8D",X"4B",X"8E",X"4A",X"02",X"8B",X"1A",X"55",X"0E",
		X"8A",X"7C",X"4E",X"05",X"8A",X"0B",X"86",X"46",X"03",X"4A",X"0D",X"7C",X"5A",X"36",X"AB",X"08",
		X"55",X"08",X"56",X"01",X"4A",X"05",X"56",X"03",X"7C",X"4D",X"BC",X"83",X"0A",X"4B",X"07",X"BC",
		X"81",X"72",X"02",X"56",X"02",X"6A",X"01",X"95",X"3B",X"88",X"53",X"03",X"BC",X"95",X"46",X"0B",
		X"95",X"04",X"A0",X"0C",X"4A",X"02",X"56",X"03",X"55",X"01",X"95",X"03",X"4A",X"04",X"8A",X"02",
		X"4A",X"02",X"8A",X"29",X"8B",X"06",X"4B",X"16",X"4A",X"01",X"95",X"0D",X"88",X"53",X"01",X"6A",
		X"0F",X"8A",X"08",X"8B",X"0D",X"4B",X"08",X"8B",X"07",X"55",X"02",X"69",X"89",X"03",X"4B",X"01",
		X"7C",X"6F",X"05",X"8B",X"4B",X"0D",X"8B",X"01",X"4E",X"83",X"01",X"8B",X"0F",X"55",X"05",X"A2",
		X"42",X"10",X"60",X"26",X"4B",X"02",X"8B",X"08",X"4B",X"05",X"8F",X"4F",X"01",X"95",X"17",X"4A",
		X"0E",X"8A",X"04",X"A0",X"1B",X"8B",X"11",X"4B",X"0A",X"52",X"97",X"4D",X"8F",X"47",X"06",X"8B",
		X"02",X"55",X"03",X"9D",X"67",X"8A",X"0A",X"56",X"05",X"8B",X"02",X"48",X"88",X"03",X"55",X"09",
		X"60",X"03",X"76",X"13",X"8B",X"24",X"4B",X"2F",X"8B",X"05",X"8B",X"08",X"8A",X"15",X"96",X"3C",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"0A",X"95",X"60",X"04",X"9E",X"53",X"0D",X"8B",X"02",X"4B",X"0F",
		X"93",X"53",X"07",X"A9",X"54",X"0A",X"96",X"03",X"60",X"0F",X"8A",X"23",X"48",X"B9",X"02",X"82",
		X"59",X"9F",X"59",X"01",X"8B",X"22",X"AB",X"02",X"4B",X"02",X"8B",X"07",X"55",X"AC",X"42",X"01",
		X"50",X"90",X"02",X"55",X"35",X"90",X"50",X"04",X"92",X"5B",X"89",X"1F",X"48",X"88",X"05",X"8C",
		X"42",X"05",X"4A",X"3C",X"0C",X"46",X"86",X"3C",X"04",X"93",X"5E",X"06",X"4B",X"09",X"4A",X"0A",
		X"7C",X"7C",X"6F",X"BC",X"01",X"8B",X"07",X"92",X"48",X"07",X"88",X"7C",X"7C",X"45",X"11",X"90",
		X"50",X"01",X"8B",X"07",X"4B",X"0C",X"8B",X"0A",X"76",X"AB",X"12",X"87",X"47",X"18",X"8B",X"03",
		X"8A",X"02",X"96",X"08",X"4B",X"02",X"8B",X"07",X"95",X"3C",X"3C",X"17",X"55",X"3C",X"05",X"56",
		X"20",X"7C",X"44",X"06",X"67",X"BC",X"4D",X"8E",X"0C",X"56",X"02",X"4A",X"1A",X"4B",X"39",X"55",
		X"25",X"56",X"20",X"55",X"0B",X"4B",X"03",X"60",X"06",X"4A",X"03",X"41",X"01",X"BC",X"9F",X"50",
		X"04",X"96",X"0F",X"4B",X"07",X"8B",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"02",X"90",
		X"45",X"02",X"4B",X"02",X"48",X"88",X"07",X"8A",X"55",X"01",X"4A",X"01",X"58",X"82",X"03",X"8A",
		X"5F",X"01",X"60",X"07",X"B2",X"52",X"03",X"46",X"86",X"1E",X"49",X"89",X"08",X"4B",X"01",X"94",
		X"49",X"05",X"8A",X"4A",X"3C",X"3C",X"0A",X"BC",X"84",X"11",X"53",X"88",X"01",X"4A",X"0B",X"6B",
		X"06",X"4B",X"24",X"4A",X"11",X"56",X"08",X"4A",X"0E",X"4B",X"07",X"55",X"07",X"4B",X"07",X"7C",
		X"72",X"8E",X"01",X"AF",X"44",X"02",X"56",X"8B",X"04",X"5A",X"85",X"02",X"8A",X"02",X"90",X"45",
		X"09",X"8B",X"01",X"48",X"89",X"41",X"02",X"4B",X"05",X"B5",X"10",X"4D",X"83",X"03",X"B5",X"4B",
		X"03",X"A0",X"07",X"72",X"88",X"08",X"4B",X"01",X"50",X"85",X"03",X"8B",X"02",X"55",X"05",X"95",
		X"06",X"60",X"06",X"55",X"01",X"4B",X"09",X"48",X"8F",X"47",X"03",X"4B",X"01",X"96",X"07",X"8A",
		X"05",X"6A",X"18",X"4B",X"0A",X"8B",X"06",X"8A",X"02",X"44",X"84",X"06",X"8B",X"08",X"8B",X"14",
		X"BC",X"84",X"03",X"59",X"83",X"02",X"8B",X"03",X"60",X"08",X"8B",X"05",X"7C",X"5A",X"01",X"B6",
		X"0A",X"48",X"95",X"4D",X"01",X"8A",X"09",X"51",X"BC",X"85",X"65",X"2D",X"6B",X"01",X"95",X"4D",
		X"83",X"02",X"8A",X"4A",X"01",X"8B",X"02",X"72",X"85",X"53",X"01",X"95",X"02",X"8B",X"06",X"95",
		X"03",X"8B",X"01",X"8A",X"01",X"4A",X"07",X"95",X"01",X"6B",X"03",X"97",X"41",X"05",X"4B",X"0B",
		X"48",X"88",X"05",X"60",X"3C",X"3C",X"3C",X"3C",X"73",X"A6",X"14",X"7E",X"29",X"F8",X"9B",X"13",
		X"13",X"96",X"B9",X"3A",X"00",X"A8",X"3C",X"C2",X"96",X"24",X"3A",X"C6",X"AC",X"A7",X"C2",X"96",
		X"24",X"CD",X"D1",X"1E",X"07",X"07",X"07",X"07",X"21",X"8E",X"A9",X"CB",X"16",X"7E",X"E6",X"03",
		X"FE",X"01",X"21",X"81",X"AA",X"20",X"02",X"36",X"03",X"3A",X"30",X"AD",X"A7",X"28",X"05",X"7E",
		X"A7",X"CA",X"96",X"24",X"23",X"7E",X"A7",X"C2",X"96",X"24",X"DD",X"21",X"80",X"AA",X"06",X"06",
		X"DD",X"7E",X"00",X"A7",X"28",X"23",X"ED",X"5B",X"46",X"0D",X"DD",X"19",X"10",X"F2",X"C3",X"96",
		X"24",X"16",X"A7",X"13",X"96",X"ED",X"DC",X"F1",X"8C",X"68",X"3B",X"0D",X"ED",X"F1",X"96",X"13",
		X"13",X"13",X"13",X"F1",X"88",X"DC",X"ED",X"11",X"B9",X"CD",X"7E",X"56",X"AF",X"67",X"6F",X"ED",
		X"4B",X"08",X"A8",X"ED",X"42",X"29",X"29",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"AF",X"67",X"6F",
		X"ED",X"4B",X"0A",X"A8",X"ED",X"42",X"29",X"29",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"3A",X"02",
		X"A8",X"C6",X"04",X"0F",X"0F",X"0F",X"E6",X"1F",X"21",X"71",X"27",X"CD",X"8C",X"01",X"DD",X"35",
		X"00",X"DD",X"36",X"03",X"00",X"DD",X"73",X"04",X"DD",X"36",X"05",X"00",X"DD",X"72",X"06",X"21",
		X"81",X"AA",X"35",X"23",X"36",X"06",X"3A",X"82",X"AA",X"A7",X"28",X"04",X"3D",X"32",X"82",X"AA",
		X"DD",X"21",X"80",X"AA",X"06",X"06",X"D9",X"DD",X"7E",X"00",X"A7",X"28",X"46",X"3C",X"20",X"4C",
		X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"ED",X"5B",X"08",X"A8",X"19",X"DD",X"56",X"04",X"DD",X"5E",
		X"03",X"19",X"7C",X"C6",X"10",X"FE",X"10",X"DA",X"FC",X"24",X"DD",X"74",X"04",X"DD",X"75",X"03",
		X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"ED",X"5B",X"0A",X"A8",X"19",X"DD",X"56",X"06",X"DD",X"5E",
		X"05",X"19",X"7C",X"C6",X"08",X"FE",X"18",X"DA",X"FC",X"24",X"DD",X"74",X"06",X"DD",X"75",X"05",
		X"CD",X"37",X"53",X"11",X"10",X"00",X"DD",X"19",X"D9",X"10",X"AB",X"C9",X"AF",X"DD",X"77",X"00",
		X"DD",X"77",X"04",X"DD",X"77",X"06",X"C3",X"F3",X"24",X"E0",X"A4",X"14",X"9B",X"10",X"0D",X"88",
		X"B9",X"21",X"00",X"AC",X"06",X"40",X"36",X"FF",X"23",X"10",X"FB",X"CD",X"67",X"4B",X"32",X"00",
		X"C2",X"CD",X"A5",X"4B",X"32",X"00",X"C2",X"CD",X"6A",X"52",X"32",X"00",X"C2",X"C3",X"AA",X"52",
		X"19",X"01",X"18",X"01",X"17",X"01",X"16",X"01",X"15",X"01",X"14",X"01",X"13",X"01",X"10",X"01",
		X"0E",X"01",X"0C",X"01",X"0A",X"01",X"08",X"01",X"04",X"01",X"01",X"01",X"FF",X"00",X"FB",X"00",
		X"F8",X"00",X"F5",X"00",X"F2",X"00",X"EE",X"00",X"EB",X"00",X"E8",X"00",X"E4",X"00",X"E1",X"00",
		X"DE",X"00",X"DA",X"00",X"D7",X"00",X"D4",X"00",X"D1",X"00",X"CD",X"00",X"CA",X"00",X"C7",X"00",
		X"C3",X"00",X"C0",X"00",X"BC",X"00",X"B8",X"00",X"B5",X"00",X"B1",X"00",X"AC",X"00",X"A8",X"00",
		X"A5",X"00",X"A0",X"00",X"9A",X"00",X"94",X"00",X"8F",X"00",X"87",X"00",X"84",X"00",X"7D",X"00",
		X"76",X"00",X"70",X"00",X"69",X"00",X"61",X"00",X"5B",X"00",X"53",X"00",X"4B",X"00",X"44",X"00",
		X"3B",X"00",X"33",X"00",X"2C",X"00",X"23",X"00",X"1A",X"00",X"11",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"FF",X"EF",X"FF",X"00",X"00",X"DD",X"FF",X"D4",X"FF",X"CD",X"FF",X"C5",X"FF",
		X"BC",X"FF",X"B5",X"FF",X"AD",X"FF",X"A5",X"FF",X"9F",X"FF",X"97",X"FF",X"90",X"FF",X"8A",X"FF",
		X"83",X"FF",X"7C",X"FF",X"79",X"FF",X"7C",X"FF",X"6C",X"FF",X"66",X"FF",X"60",X"FF",X"5B",X"FF",
		X"58",X"FF",X"54",X"FF",X"4F",X"FF",X"4B",X"FF",X"48",X"FF",X"44",X"FF",X"40",X"FF",X"3D",X"FF",
		X"39",X"FF",X"36",X"FF",X"33",X"FF",X"33",X"FF",X"2C",X"FF",X"29",X"FF",X"26",X"FF",X"22",X"FF",
		X"1F",X"FF",X"1C",X"FF",X"18",X"FF",X"15",X"FF",X"12",X"FF",X"0E",X"FF",X"0B",X"FF",X"08",X"FF",
		X"05",X"FF",X"01",X"FF",X"FF",X"FE",X"FC",X"FE",X"F8",X"FE",X"F6",X"FE",X"F4",X"FE",X"F2",X"FE",
		X"F0",X"FE",X"ED",X"FE",X"EC",X"FE",X"EB",X"FE",X"EA",X"FE",X"E9",X"FE",X"E8",X"FE",X"E7",X"FE",
		X"E7",X"FE",X"E8",X"FE",X"E9",X"FE",X"EA",X"FE",X"EB",X"FE",X"EC",X"FE",X"ED",X"FE",X"F0",X"FE",
		X"F2",X"FE",X"F4",X"FE",X"F6",X"FE",X"F8",X"FE",X"FC",X"FE",X"FF",X"FE",X"01",X"FF",X"05",X"FF",
		X"08",X"FF",X"0B",X"FF",X"0E",X"FF",X"12",X"FF",X"15",X"FF",X"18",X"FF",X"1C",X"FF",X"1F",X"FF",
		X"22",X"FF",X"26",X"FF",X"29",X"FF",X"2C",X"FF",X"2F",X"FF",X"33",X"FF",X"36",X"FF",X"39",X"FF",
		X"3D",X"FF",X"40",X"FF",X"44",X"FF",X"48",X"FF",X"4B",X"FF",X"4F",X"FF",X"54",X"FF",X"58",X"FF",
		X"5B",X"FF",X"60",X"FF",X"66",X"FF",X"6C",X"FF",X"71",X"FF",X"79",X"FF",X"7C",X"FF",X"83",X"FF",
		X"8A",X"FF",X"90",X"FF",X"97",X"FF",X"9F",X"FF",X"A5",X"FF",X"AD",X"FF",X"B5",X"FF",X"BC",X"FF",
		X"C5",X"FF",X"CD",X"FF",X"D4",X"FF",X"DD",X"FF",X"E6",X"FF",X"EF",X"FF",X"F8",X"FF",X"00",X"00",
		X"00",X"00",X"08",X"00",X"11",X"00",X"1A",X"00",X"23",X"00",X"2C",X"00",X"33",X"00",X"3B",X"00",
		X"44",X"00",X"4B",X"00",X"53",X"00",X"5B",X"00",X"61",X"00",X"69",X"00",X"70",X"00",X"76",X"00",
		X"7D",X"00",X"84",X"00",X"87",X"00",X"87",X"00",X"94",X"00",X"9A",X"00",X"A0",X"00",X"A5",X"00",
		X"A8",X"00",X"AC",X"00",X"B1",X"00",X"B5",X"00",X"B8",X"00",X"BC",X"00",X"C0",X"00",X"C3",X"00",
		X"C7",X"00",X"CA",X"00",X"CD",X"00",X"CA",X"00",X"D4",X"00",X"D7",X"00",X"DA",X"00",X"DE",X"00",
		X"E1",X"00",X"E4",X"00",X"E8",X"00",X"EB",X"00",X"EE",X"00",X"F2",X"00",X"F5",X"00",X"F8",X"00",
		X"FB",X"00",X"FF",X"00",X"01",X"01",X"FB",X"00",X"08",X"01",X"0A",X"01",X"0C",X"01",X"0E",X"01",
		X"10",X"01",X"13",X"01",X"14",X"01",X"15",X"01",X"16",X"01",X"17",X"01",X"18",X"01",X"19",X"01",
		X"3A",X"6F",X"AA",X"FE",X"76",X"C2",X"30",X"25",X"CD",X"2B",X"0B",X"CD",X"0E",X"21",X"AF",X"32",
		X"31",X"AD",X"32",X"20",X"AD",X"32",X"30",X"AD",X"32",X"AC",X"A9",X"3C",X"32",X"10",X"AD",X"3E",
		X"03",X"32",X"AB",X"A9",X"C9",X"DD",X"21",X"80",X"AA",X"21",X"6E",X"27",X"3A",X"61",X"08",X"5F",
		X"3A",X"01",X"5C",X"57",X"06",X"06",X"DD",X"77",X"00",X"DD",X"77",X"04",X"DD",X"19",X"10",X"F6",
		X"C9",X"7E",X"84",X"7E",X"85",X"7E",X"86",X"7D",X"87",X"7C",X"88",X"7B",X"89",X"7A",X"8A",X"79",
		X"8A",X"78",X"8A",X"77",X"8A",X"76",X"8A",X"75",X"89",X"74",X"88",X"73",X"87",X"72",X"86",X"72",
		X"85",X"72",X"84",X"72",X"83",X"72",X"82",X"73",X"81",X"74",X"80",X"75",X"7F",X"76",X"7E",X"77",
		X"7E",X"78",X"7E",X"79",X"7E",X"7A",X"7E",X"7B",X"7F",X"7C",X"80",X"7D",X"81",X"7E",X"82",X"7E",
		X"83",X"CD",X"34",X"58",X"3E",X"78",X"32",X"64",X"AC",X"3E",X"84",X"32",X"65",X"AC",X"21",X"00",
		X"00",X"22",X"16",X"AD",X"22",X"26",X"AD",X"3A",X"CD",X"A9",X"32",X"12",X"AD",X"32",X"22",X"AD",
		X"AF",X"32",X"14",X"AD",X"32",X"24",X"AD",X"32",X"32",X"AD",X"32",X"13",X"AD",X"32",X"23",X"AD",
		X"32",X"1D",X"AD",X"32",X"2D",X"AD",X"32",X"0C",X"AD",X"3C",X"32",X"11",X"AD",X"32",X"21",X"AD",
		X"32",X"1E",X"AD",X"32",X"2E",X"AD",X"3A",X"30",X"AD",X"A7",X"28",X"39",X"AF",X"67",X"6F",X"32",
		X"33",X"AD",X"22",X"34",X"AD",X"32",X"36",X"AD",X"22",X"37",X"AD",X"11",X"00",X"04",X"FF",X"3A",
		X"C4",X"A9",X"CD",X"7B",X"0F",X"06",X"00",X"21",X"50",X"15",X"97",X"AE",X"23",X"10",X"FC",X"C6",
		X"01",X"32",X"08",X"C3",X"3A",X"D3",X"A9",X"32",X"1A",X"AD",X"32",X"2A",X"AD",X"3E",X"96",X"32",
		X"EB",X"A9",X"C3",X"1A",X"0F",X"21",X"D0",X"A9",X"7E",X"3C",X"FE",X"04",X"38",X"02",X"3E",X"01",
		X"77",X"32",X"14",X"AD",X"3C",X"32",X"11",X"AD",X"AF",X"32",X"80",X"A9",X"32",X"CE",X"A9",X"32",
		X"CF",X"A9",X"CD",X"67",X"4B",X"21",X"80",X"AA",X"11",X"81",X"AA",X"36",X"00",X"01",X"5F",X"00",
		X"ED",X"B0",X"21",X"00",X"A8",X"11",X"01",X"A8",X"36",X"00",X"01",X"7F",X"01",X"ED",X"B0",X"3E",
		X"02",X"CD",X"7B",X"0F",X"3A",X"D3",X"A9",X"32",X"1A",X"AD",X"32",X"2A",X"AD",X"0E",X"00",X"21",
		X"10",X"33",X"3A",X"AB",X"A9",X"96",X"23",X"0D",X"20",X"FB",X"EE",X"90",X"32",X"AB",X"A9",X"21",
		X"74",X"AC",X"06",X"10",X"36",X"80",X"23",X"10",X"FB",X"3E",X"5A",X"32",X"EB",X"A9",X"C3",X"1A",
		X"0F",X"CD",X"B7",X"28",X"CD",X"C2",X"28",X"CD",X"CD",X"28",X"CD",X"D8",X"28",X"CD",X"E3",X"28",
		X"CD",X"EE",X"28",X"CD",X"FE",X"28",X"C9",X"DD",X"21",X"50",X"A8",X"FD",X"21",X"1A",X"AA",X"C3",
		X"0E",X"29",X"DD",X"21",X"60",X"A8",X"FD",X"21",X"1C",X"AA",X"C3",X"0E",X"29",X"DD",X"21",X"70",
		X"A8",X"FD",X"21",X"1E",X"AA",X"C3",X"0E",X"29",X"DD",X"21",X"80",X"A8",X"FD",X"21",X"20",X"AA",
		X"C3",X"0E",X"29",X"DD",X"21",X"90",X"A8",X"FD",X"21",X"22",X"AA",X"C3",X"0E",X"29",X"3A",X"0D",
		X"AD",X"A7",X"C0",X"DD",X"21",X"A0",X"A8",X"FD",X"21",X"24",X"AA",X"C3",X"0E",X"29",X"3A",X"0D",
		X"AD",X"A7",X"C0",X"DD",X"21",X"B0",X"A8",X"FD",X"21",X"26",X"AA",X"C3",X"0E",X"29",X"3A",X"04",
		X"AD",X"E6",X"07",X"F7",X"27",X"29",X"4C",X"29",X"84",X"29",X"B0",X"29",X"D5",X"29",X"86",X"EB",
		X"4E",X"EB",X"23",X"13",X"10",X"F8",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"3C",X"28",X"07",X"3C",
		X"CA",X"52",X"2B",X"C3",X"93",X"2B",X"CD",X"EF",X"2B",X"CD",X"40",X"58",X"CD",X"83",X"2B",X"DA",
		X"DE",X"2B",X"CD",X"D6",X"3E",X"CD",X"3C",X"2A",X"CD",X"43",X"42",X"C9",X"DD",X"7E",X"00",X"A7",
		X"C8",X"3C",X"28",X"07",X"3C",X"CA",X"52",X"2B",X"C3",X"93",X"2B",X"CD",X"EF",X"2B",X"CD",X"54",
		X"58",X"CD",X"83",X"2B",X"DA",X"DE",X"2B",X"CD",X"D6",X"3E",X"CD",X"47",X"2A",X"C9",X"09",X"A7",
		X"32",X"82",X"6E",X"58",X"B5",X"77",X"E4",X"E8",X"EC",X"9D",X"CB",X"4F",X"55",X"FE",X"A3",X"31",
		X"81",X"5B",X"9A",X"B9",X"DD",X"7E",X"00",X"A7",X"C8",X"3C",X"28",X"07",X"3C",X"CA",X"52",X"2B",
		X"C3",X"93",X"2B",X"3A",X"80",X"A9",X"E6",X"03",X"FE",X"03",X"DC",X"EF",X"2B",X"CD",X"40",X"58",
		X"CD",X"83",X"2B",X"DA",X"DE",X"2B",X"CD",X"D6",X"3E",X"CD",X"97",X"2A",X"CD",X"43",X"42",X"C9",
		X"DD",X"7E",X"00",X"A7",X"C8",X"3C",X"28",X"07",X"3C",X"CA",X"52",X"2B",X"C3",X"93",X"2B",X"CD",
		X"EF",X"2B",X"CD",X"A4",X"58",X"CD",X"83",X"2B",X"DA",X"DE",X"2B",X"CD",X"D6",X"3E",X"CD",X"FC",
		X"2A",X"CD",X"43",X"42",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"3C",X"28",X"07",X"3C",X"CA",X"52",
		X"2B",X"C3",X"93",X"2B",X"CD",X"F7",X"29",X"CD",X"83",X"2B",X"DA",X"DE",X"2B",X"CD",X"38",X"2B",
		X"CD",X"D6",X"3E",X"CD",X"43",X"42",X"C9",X"3E",X"78",X"FD",X"96",X"31",X"C6",X"48",X"FE",X"90",
		X"38",X"1A",X"3E",X"84",X"FD",X"96",X"31",X"C6",X"48",X"FE",X"90",X"38",X"0F",X"CD",X"EF",X"2B",
		X"3A",X"80",X"A9",X"0F",X"E6",X"01",X"CA",X"AA",X"58",X"C3",X"60",X"58",X"AF",X"32",X"04",X"AD",
		X"CD",X"EF",X"2B",X"3E",X"04",X"32",X"04",X"AD",X"18",X"E6",X"DD",X"7E",X"04",X"3D",X"CA",X"93",
		X"2B",X"DD",X"77",X"04",X"DD",X"36",X"00",X"FF",X"CD",X"BA",X"2B",X"C9",X"CD",X"57",X"2A",X"FD",
		X"71",X"30",X"78",X"FD",X"77",X"01",X"C9",X"CD",X"57",X"2A",X"79",X"C6",X"35",X"FD",X"77",X"30",
		X"78",X"C6",X"10",X"FD",X"77",X"01",X"C9",X"11",X"10",X"00",X"DD",X"7E",X"02",X"C6",X"08",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"21",X"77",X"2A",X"DF",X"46",X"19",X"4E",X"3A",X"80",X"A9",X"CB",
		X"4F",X"C8",X"78",X"C6",X"08",X"47",X"C9",X"0C",X"0D",X"0E",X"0F",X"08",X"0F",X"0E",X"0D",X"0C",
		X"0B",X"0A",X"09",X"08",X"09",X"0A",X"0B",X"41",X"41",X"41",X"41",X"81",X"C1",X"C1",X"C1",X"C1",
		X"C1",X"C1",X"C1",X"41",X"41",X"41",X"41",X"DD",X"7E",X"02",X"C6",X"04",X"E6",X"F8",X"0F",X"0F",
		X"E6",X"3F",X"21",X"BC",X"2A",X"DF",X"46",X"3A",X"80",X"A9",X"E6",X"02",X"20",X"0A",X"80",X"FD",
		X"77",X"01",X"23",X"7E",X"FD",X"77",X"30",X"C9",X"3E",X"08",X"18",X"F2",X"80",X"DC",X"80",X"DC",
		X"80",X"DC",X"80",X"DC",X"81",X"DC",X"81",X"DC",X"82",X"DC",X"83",X"DC",X"84",X"5C",X"84",X"5C",
		X"83",X"5C",X"82",X"5C",X"81",X"5C",X"81",X"5C",X"80",X"5C",X"80",X"5C",X"80",X"5C",X"80",X"5C",
		X"80",X"5C",X"80",X"5C",X"81",X"5C",X"81",X"5C",X"82",X"5C",X"83",X"5C",X"84",X"DC",X"84",X"DC",
		X"83",X"DC",X"82",X"DC",X"81",X"DC",X"81",X"DC",X"80",X"DC",X"80",X"DC",X"11",X"10",X"00",X"DD",
		X"7E",X"02",X"C6",X"08",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"21",X"18",X"2B",X"DF",X"7E",X"FD",
		X"77",X"01",X"19",X"7E",X"FD",X"77",X"30",X"C9",X"2C",X"2D",X"2E",X"2F",X"28",X"2F",X"2E",X"2D",
		X"2C",X"2B",X"2A",X"29",X"28",X"29",X"2A",X"2B",X"5B",X"5B",X"5B",X"5B",X"9B",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"5B",X"5B",X"5B",X"5B",X"3A",X"80",X"A9",X"0F",X"0F",X"E6",X"03",X"C6",
		X"D8",X"47",X"DD",X"7E",X"04",X"D6",X"01",X"87",X"87",X"80",X"FD",X"77",X"01",X"FD",X"36",X"30",
		X"61",X"C9",X"DD",X"35",X"0E",X"28",X"01",X"C9",X"DD",X"34",X"00",X"DD",X"36",X"0E",X"80",X"C9",
		X"FD",X"66",X"31",X"DD",X"6E",X"03",X"ED",X"5B",X"08",X"A8",X"19",X"FD",X"74",X"31",X"DD",X"75",
		X"03",X"FD",X"66",X"00",X"DD",X"6E",X"05",X"ED",X"5B",X"0A",X"A8",X"19",X"FD",X"74",X"00",X"DD",
		X"75",X"05",X"C9",X"FD",X"7E",X"31",X"C6",X"09",X"FE",X"03",X"D8",X"FD",X"7E",X"00",X"D6",X"03",
		X"FE",X"03",X"C9",X"DD",X"7E",X"00",X"FE",X"F0",X"CA",X"AC",X"2B",X"FE",X"3C",X"CC",X"BA",X"2B",
		X"D2",X"B4",X"2B",X"DD",X"35",X"00",X"28",X"36",X"CD",X"22",X"2C",X"C9",X"DD",X"36",X"00",X"3B",
		X"CD",X"BA",X"2B",X"C9",X"DD",X"35",X"00",X"C3",X"40",X"58",X"CD",X"83",X"56",X"21",X"02",X"AD",
		X"7E",X"A7",X"28",X"01",X"35",X"DD",X"7E",X"0E",X"CB",X"7F",X"C8",X"3A",X"12",X"A8",X"A7",X"C8",
		X"21",X"11",X"A8",X"35",X"C0",X"DD",X"7E",X"0F",X"C6",X"80",X"32",X"21",X"A8",X"C9",X"AF",X"DD",
		X"77",X"00",X"DD",X"77",X"03",X"DD",X"77",X"05",X"FD",X"77",X"00",X"FD",X"77",X"31",X"C9",X"DD",
		X"7E",X"01",X"DD",X"96",X"02",X"4F",X"C6",X"02",X"FE",X"04",X"D8",X"DD",X"46",X"02",X"79",X"FE",
		X"80",X"30",X"0C",X"21",X"1D",X"2C",X"3A",X"04",X"AD",X"CF",X"80",X"DD",X"77",X"02",X"C9",X"21",
		X"1D",X"2C",X"3A",X"04",X"AD",X"CF",X"90",X"ED",X"44",X"DD",X"77",X"02",X"C9",X"01",X"01",X"02",
		X"02",X"05",X"21",X"31",X"2C",X"E5",X"DD",X"7E",X"00",X"FE",X"20",X"D2",X"B4",X"2B",X"C3",X"60",
		X"2B",X"DD",X"7E",X"00",X"FE",X"2A",X"D2",X"71",X"2C",X"FE",X"0A",X"30",X"45",X"3A",X"21",X"A8",
		X"CB",X"7F",X"CA",X"DE",X"2B",X"3A",X"21",X"A8",X"CB",X"BF",X"DD",X"BE",X"0F",X"C2",X"DE",X"2B",
		X"3A",X"80",X"A9",X"E6",X"07",X"28",X"03",X"DD",X"34",X"00",X"FD",X"36",X"01",X"FC",X"FD",X"36",
		X"30",X"6C",X"DD",X"7E",X"00",X"FE",X"01",X"C0",X"11",X"0C",X"04",X"FF",X"AF",X"32",X"21",X"A8",
		X"C9",X"FD",X"7E",X"30",X"4F",X"E6",X"C0",X"47",X"3A",X"80",X"A9",X"E6",X"0F",X"80",X"FD",X"77",
		X"30",X"C9",X"D6",X"0A",X"0F",X"E6",X"0F",X"47",X"21",X"94",X"2C",X"CF",X"FD",X"77",X"01",X"FD",
		X"36",X"30",X"3C",X"C9",X"FF",X"FF",X"7D",X"7D",X"7E",X"7E",X"7D",X"7D",X"5B",X"5B",X"5A",X"5A",
		X"59",X"59",X"58",X"58",X"18",X"A7",X"13",X"A5",X"3B",X"87",X"F1",X"34",X"0E",X"34",X"D7",X"BF",
		X"F1",X"65",X"13",X"13",X"13",X"13",X"F1",X"88",X"DC",X"ED",X"11",X"B9",X"DD",X"21",X"00",X"A9",
		X"FD",X"21",X"30",X"AA",X"3A",X"04",X"AD",X"A7",X"28",X"2B",X"FE",X"04",X"28",X"34",X"CD",X"21",
		X"2D",X"CD",X"36",X"2D",X"CD",X"36",X"2D",X"CD",X"68",X"2D",X"C9",X"CD",X"C2",X"01",X"C0",X"01",
		X"04",X"00",X"21",X"80",X"49",X"97",X"AE",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C6",X"BD",X"C2",
		X"11",X"0F",X"C3",X"1A",X"0F",X"CD",X"15",X"2D",X"CD",X"36",X"2D",X"CD",X"36",X"2D",X"CD",X"68",
		X"2D",X"C9",X"CD",X"2D",X"2D",X"CD",X"2D",X"2D",X"CD",X"62",X"2D",X"CD",X"62",X"2D",X"CD",X"68",
		X"2D",X"CD",X"68",X"2D",X"C9",X"CD",X"6E",X"2D",X"CD",X"58",X"30",X"CD",X"58",X"30",X"C3",X"9B",
		X"30",X"CD",X"6E",X"2D",X"CD",X"58",X"30",X"CD",X"8A",X"30",X"C3",X"9B",X"30",X"CD",X"6E",X"2D",
		X"CD",X"58",X"30",X"C3",X"9B",X"30",X"CD",X"93",X"2D",X"CD",X"58",X"30",X"C3",X"9B",X"30",X"3A",
		X"C0",X"A9",X"A7",X"C2",X"1A",X"0F",X"CD",X"FB",X"4A",X"11",X"08",X"01",X"FF",X"3A",X"17",X"A8",
		X"A7",X"C2",X"3E",X"2E",X"CD",X"06",X"0B",X"CD",X"39",X"0B",X"21",X"6B",X"08",X"06",X"14",X"C3",
		X"E8",X"43",X"CD",X"93",X"2D",X"C3",X"9B",X"30",X"CD",X"F4",X"2D",X"C3",X"9B",X"30",X"FD",X"56",
		X"31",X"DD",X"5E",X"03",X"2A",X"08",X"A8",X"CD",X"31",X"2E",X"FD",X"74",X"31",X"DD",X"75",X"03",
		X"FD",X"56",X"00",X"DD",X"5E",X"05",X"2A",X"0A",X"A8",X"CD",X"31",X"2E",X"FD",X"74",X"00",X"DD",
		X"75",X"05",X"C9",X"FD",X"56",X"31",X"DD",X"5E",X"03",X"2A",X"08",X"A8",X"CD",X"3E",X"30",X"FD",
		X"74",X"31",X"DD",X"75",X"03",X"FD",X"56",X"00",X"DD",X"5E",X"05",X"2A",X"0A",X"A8",X"CD",X"3E",
		X"30",X"FD",X"74",X"00",X"DD",X"75",X"05",X"C9",X"21",X"01",X"AD",X"34",X"21",X"04",X"AD",X"7E",
		X"3C",X"FE",X"05",X"38",X"01",X"AF",X"77",X"3A",X"01",X"AD",X"FE",X"06",X"38",X"09",X"FE",X"0B",
		X"38",X"0A",X"3A",X"D5",X"A9",X"18",X"08",X"3A",X"D3",X"A9",X"18",X"03",X"3A",X"D4",X"A9",X"32",
		X"0A",X"AD",X"3A",X"CD",X"A9",X"32",X"02",X"AD",X"AF",X"32",X"0D",X"AD",X"32",X"C6",X"AC",X"3D",
		X"32",X"0E",X"AD",X"C9",X"FD",X"56",X"31",X"DD",X"5E",X"03",X"2A",X"08",X"A8",X"CD",X"4D",X"30",
		X"FD",X"74",X"31",X"DD",X"75",X"03",X"FD",X"56",X"00",X"DD",X"5E",X"05",X"2A",X"0A",X"A8",X"CD",
		X"4D",X"30",X"FD",X"74",X"00",X"DD",X"75",X"05",X"C9",X"32",X"C1",X"A9",X"79",X"0F",X"0F",X"4F",
		X"E6",X"01",X"32",X"C2",X"A9",X"79",X"0F",X"4F",X"E6",X"01",X"32",X"C3",X"A9",X"79",X"C3",X"A8",
		X"49",X"44",X"4D",X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"09",X"19",X"C9",X"32",X"01",
		X"31",X"01",X"30",X"01",X"2F",X"01",X"2E",X"01",X"2D",X"01",X"2C",X"01",X"28",X"01",X"26",X"01",
		X"24",X"01",X"22",X"01",X"20",X"01",X"1B",X"01",X"18",X"01",X"16",X"01",X"11",X"01",X"0E",X"01",
		X"0B",X"01",X"08",X"01",X"03",X"01",X"00",X"01",X"FD",X"00",X"F8",X"00",X"F5",X"00",X"F2",X"00",
		X"ED",X"00",X"EA",X"00",X"E7",X"00",X"E4",X"00",X"DF",X"00",X"DC",X"00",X"D9",X"00",X"D4",X"00",
		X"D1",X"00",X"CD",X"00",X"C8",X"00",X"C5",X"00",X"C1",X"00",X"BB",X"00",X"B7",X"00",X"B4",X"00",
		X"AE",X"00",X"A8",X"00",X"A1",X"00",X"9C",X"00",X"93",X"00",X"90",X"00",X"88",X"00",X"80",X"00",
		X"7A",X"00",X"72",X"00",X"69",X"00",X"63",X"00",X"5A",X"00",X"51",X"00",X"4A",X"00",X"40",X"00",
		X"37",X"00",X"30",X"00",X"26",X"00",X"1C",X"00",X"12",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FF",X"EE",X"FF",X"00",X"00",X"DA",X"FF",X"D0",X"FF",X"C9",X"FF",X"C0",X"FF",X"B6",X"FF",
		X"AF",X"FF",X"A6",X"FF",X"9D",X"FF",X"97",X"FF",X"8E",X"FF",X"86",X"FF",X"80",X"FF",X"78",X"FF",
		X"70",X"FF",X"6D",X"FF",X"70",X"FF",X"5F",X"FF",X"58",X"FF",X"52",X"FF",X"4C",X"FF",X"49",X"FF",
		X"45",X"FF",X"3F",X"FF",X"3B",X"FF",X"38",X"FF",X"33",X"FF",X"2F",X"FF",X"2C",X"FF",X"27",X"FF",
		X"24",X"FF",X"21",X"FF",X"21",X"FF",X"19",X"FF",X"16",X"FF",X"13",X"FF",X"0E",X"FF",X"0B",X"FF",
		X"08",X"FF",X"03",X"FF",X"00",X"FF",X"FD",X"FE",X"F8",X"FE",X"F5",X"FE",X"F2",X"FE",X"EF",X"FE",
		X"EA",X"FE",X"E8",X"FE",X"E5",X"FE",X"E0",X"FE",X"DE",X"FE",X"DC",X"FE",X"DA",X"FE",X"D8",X"FE",
		X"D4",X"FE",X"D3",X"FE",X"D2",X"FE",X"D1",X"FE",X"D0",X"FE",X"CF",X"FE",X"CE",X"FE",X"CE",X"FE",
		X"CF",X"FE",X"D0",X"FE",X"D1",X"FE",X"D2",X"FE",X"D3",X"FE",X"D4",X"FE",X"D8",X"FE",X"DA",X"FE",
		X"DC",X"FE",X"DE",X"FE",X"E0",X"FE",X"E5",X"FE",X"E8",X"FE",X"EA",X"FE",X"EF",X"FE",X"F2",X"FE",
		X"F5",X"FE",X"F8",X"FE",X"FD",X"FE",X"00",X"FF",X"03",X"FF",X"08",X"FF",X"0B",X"FF",X"0E",X"FF",
		X"13",X"FF",X"16",X"FF",X"19",X"FF",X"1C",X"FF",X"21",X"FF",X"24",X"FF",X"27",X"FF",X"2C",X"FF",
		X"2F",X"FF",X"33",X"FF",X"38",X"FF",X"3B",X"FF",X"3F",X"FF",X"45",X"FF",X"49",X"FF",X"4C",X"FF",
		X"52",X"FF",X"58",X"FF",X"5F",X"FF",X"64",X"FF",X"6D",X"FF",X"70",X"FF",X"78",X"FF",X"80",X"FF",
		X"86",X"FF",X"8E",X"FF",X"97",X"FF",X"9D",X"FF",X"A6",X"FF",X"AF",X"FF",X"B6",X"FF",X"C0",X"FF",
		X"C9",X"FF",X"D0",X"FF",X"DA",X"FF",X"E4",X"FF",X"EE",X"FF",X"F8",X"FF",X"00",X"00",X"00",X"00",
		X"08",X"00",X"12",X"00",X"1C",X"00",X"26",X"00",X"30",X"00",X"37",X"00",X"40",X"00",X"4A",X"00",
		X"51",X"00",X"5A",X"00",X"63",X"00",X"69",X"00",X"72",X"00",X"7A",X"00",X"80",X"00",X"88",X"00",
		X"90",X"00",X"93",X"00",X"93",X"00",X"A1",X"00",X"A8",X"00",X"AE",X"00",X"B4",X"00",X"B7",X"00",
		X"BB",X"00",X"C1",X"00",X"C5",X"00",X"C8",X"00",X"CD",X"00",X"D1",X"00",X"D4",X"00",X"D9",X"00",
		X"DC",X"00",X"DF",X"00",X"DC",X"00",X"E7",X"00",X"EA",X"00",X"ED",X"00",X"F2",X"00",X"F5",X"00",
		X"F8",X"00",X"FD",X"00",X"00",X"01",X"03",X"01",X"08",X"01",X"0B",X"01",X"0E",X"01",X"11",X"01",
		X"16",X"01",X"18",X"01",X"11",X"01",X"20",X"01",X"22",X"01",X"24",X"01",X"26",X"01",X"28",X"01",
		X"2C",X"01",X"2D",X"01",X"2E",X"01",X"2F",X"01",X"30",X"01",X"31",X"01",X"32",X"01",X"44",X"4D",
		X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"A7",X"ED",X"42",X"19",X"C9",X"44",X"4D",X"CB",
		X"28",X"CB",X"19",X"A7",X"ED",X"42",X"19",X"C9",X"FD",X"46",X"31",X"FD",X"4E",X"00",X"3E",X"10",
		X"80",X"FD",X"77",X"33",X"FD",X"71",X"02",X"C3",X"9B",X"30",X"FD",X"46",X"31",X"FD",X"4E",X"00",
		X"26",X"08",X"2E",X"6E",X"7E",X"81",X"FD",X"70",X"33",X"FD",X"77",X"02",X"C3",X"9B",X"30",X"73",
		X"A6",X"10",X"F1",X"D7",X"34",X"A5",X"87",X"BF",X"F1",X"B9",X"FD",X"46",X"31",X"FD",X"4E",X"00",
		X"26",X"F0",X"2E",X"10",X"09",X"FD",X"74",X"33",X"FD",X"75",X"02",X"11",X"10",X"00",X"DD",X"19",
		X"FD",X"23",X"FD",X"23",X"C9",X"21",X"6B",X"08",X"0E",X"22",X"06",X"10",X"CD",X"4C",X"0B",X"3A",
		X"04",X"AD",X"87",X"87",X"87",X"4F",X"21",X"76",X"31",X"DF",X"11",X"31",X"AA",X"06",X"08",X"7E",
		X"12",X"23",X"13",X"13",X"10",X"F9",X"3A",X"04",X"AD",X"FE",X"04",X"4F",X"CA",X"56",X"31",X"3E",
		X"CC",X"21",X"60",X"AA",X"11",X"02",X"00",X"06",X"08",X"77",X"19",X"10",X"FC",X"79",X"FE",X"04",
		X"DA",X"17",X"31",X"21",X"C7",X"AC",X"7E",X"FE",X"3B",X"C2",X"5B",X"31",X"23",X"7E",X"FE",X"05",
		X"CA",X"F8",X"30",X"FE",X"10",X"C2",X"5B",X"31",X"06",X"08",X"FD",X"21",X"30",X"AA",X"21",X"5E",
		X"31",X"7E",X"FD",X"77",X"31",X"23",X"7E",X"FD",X"77",X"00",X"23",X"FD",X"23",X"FD",X"23",X"10",
		X"F0",X"C3",X"BC",X"2C",X"C3",X"7F",X"30",X"21",X"39",X"AD",X"7E",X"FE",X"68",X"C2",X"14",X"31",
		X"23",X"7E",X"FE",X"10",X"CA",X"2C",X"31",X"FE",X"05",X"C2",X"14",X"31",X"21",X"6E",X"31",X"06",
		X"04",X"FD",X"21",X"30",X"AA",X"7E",X"FD",X"77",X"31",X"C6",X"10",X"FD",X"77",X"33",X"23",X"7E",
		X"FD",X"77",X"00",X"FD",X"77",X"02",X"23",X"11",X"10",X"00",X"DD",X"19",X"11",X"04",X"00",X"FD",
		X"19",X"10",X"E2",X"C3",X"BC",X"2C",X"3E",X"28",X"C3",X"D1",X"30",X"C3",X"76",X"31",X"40",X"68",
		X"38",X"62",X"60",X"70",X"68",X"D8",X"88",X"58",X"99",X"B0",X"37",X"43",X"CF",X"78",X"20",X"D0",
		X"50",X"60",X"A0",X"A0",X"D0",X"60",X"60",X"68",X"61",X"60",X"61",X"62",X"63",X"5C",X"74",X"75",
		X"76",X"60",X"61",X"64",X"65",X"5D",X"77",X"78",X"79",X"66",X"67",X"64",X"65",X"5E",X"7A",X"7B",
		X"7C",X"60",X"61",X"62",X"63",X"5F",X"31",X"30",X"33",X"32",X"85",X"86",X"87",X"85",X"08",X"A7",
		X"32",X"CA",X"7E",X"C8",X"FF",X"5F",X"93",X"FB",X"C4",X"AF",X"D8",X"2A",X"6C",X"E1",X"7A",X"42",
		X"BD",X"B0",X"5A",X"B9",X"3A",X"05",X"AD",X"4F",X"E6",X"F0",X"28",X"0D",X"FE",X"30",X"C2",X"6C",
		X"32",X"3A",X"03",X"49",X"FE",X"30",X"C2",X"C9",X"31",X"79",X"E6",X"0F",X"FE",X"07",X"D0",X"DD",
		X"21",X"50",X"A8",X"FD",X"21",X"1A",X"AA",X"87",X"4F",X"06",X"00",X"FD",X"09",X"87",X"87",X"87",
		X"4F",X"DD",X"09",X"DD",X"7E",X"00",X"3C",X"C0",X"CD",X"3A",X"32",X"DD",X"7E",X"08",X"FE",X"10",
		X"C8",X"FE",X"11",X"28",X"0C",X"87",X"21",X"65",X"AC",X"DF",X"CD",X"B8",X"33",X"DD",X"77",X"01",
		X"C9",X"21",X"65",X"AC",X"CD",X"B8",X"33",X"C6",X"80",X"DD",X"77",X"01",X"DD",X"36",X"08",X"10",
		X"DD",X"36",X"09",X"00",X"C9",X"CD",X"2B",X"0B",X"AF",X"32",X"31",X"AD",X"32",X"20",X"AD",X"3D",
		X"32",X"30",X"AD",X"3A",X"C1",X"A9",X"32",X"10",X"AD",X"21",X"86",X"A9",X"7E",X"D6",X"01",X"27",
		X"77",X"CD",X"FB",X"4A",X"CD",X"30",X"4B",X"C3",X"2A",X"17",X"DD",X"7E",X"09",X"A7",X"C8",X"3D",
		X"DD",X"77",X"09",X"4F",X"DD",X"7E",X"0A",X"21",X"38",X"34",X"D7",X"EB",X"79",X"CF",X"DD",X"77",
		X"08",X"C9",X"01",X"00",X"03",X"21",X"08",X"00",X"1E",X"00",X"7B",X"AE",X"23",X"0B",X"5F",X"79",
		X"B0",X"20",X"F7",X"3E",X"52",X"83",X"C2",X"11",X"0F",X"C3",X"1A",X"0F",X"79",X"E6",X"0F",X"FE",
		X"07",X"C0",X"DD",X"21",X"64",X"AC",X"3A",X"02",X"A8",X"C6",X"40",X"CD",X"D1",X"59",X"EB",X"29",
		X"29",X"29",X"7C",X"C6",X"78",X"DD",X"77",X"10",X"7C",X"ED",X"44",X"C6",X"78",X"DD",X"77",X"14",
		X"29",X"7C",X"C6",X"78",X"DD",X"77",X"12",X"7C",X"ED",X"44",X"C6",X"78",X"DD",X"77",X"16",X"60",
		X"69",X"29",X"29",X"29",X"7C",X"C6",X"84",X"DD",X"77",X"11",X"7C",X"ED",X"44",X"C6",X"84",X"DD",
		X"77",X"15",X"29",X"7C",X"C6",X"84",X"DD",X"77",X"13",X"7C",X"ED",X"44",X"C6",X"84",X"DD",X"77",
		X"17",X"3A",X"02",X"A8",X"CD",X"D1",X"59",X"EB",X"29",X"29",X"29",X"7C",X"C6",X"78",X"DD",X"77",
		X"18",X"29",X"7C",X"C6",X"78",X"DD",X"77",X"1A",X"60",X"69",X"29",X"29",X"29",X"7C",X"C6",X"84",
		X"DD",X"77",X"19",X"29",X"7C",X"C6",X"84",X"DD",X"77",X"1B",X"C9",X"32",X"00",X"C2",X"21",X"EB",
		X"A9",X"36",X"0C",X"01",X"00",X"00",X"10",X"FE",X"32",X"00",X"C2",X"0D",X"20",X"F8",X"35",X"20",
		X"F2",X"AF",X"CD",X"F8",X"55",X"3A",X"87",X"4C",X"C3",X"A8",X"00",X"21",X"EB",X"A9",X"35",X"C0",
		X"CD",X"C3",X"4C",X"D2",X"26",X"33",X"11",X"09",X"03",X"FF",X"1E",X"0B",X"FF",X"3A",X"43",X"08",
		X"32",X"AC",X"A9",X"C3",X"E7",X"12",X"CD",X"3A",X"58",X"3E",X"00",X"32",X"0C",X"AD",X"3E",X"F1",
		X"32",X"0B",X"AD",X"CD",X"E1",X"01",X"06",X"00",X"21",X"F1",X"01",X"AF",X"86",X"23",X"10",X"FC",
		X"D6",X"19",X"C4",X"11",X"0F",X"C3",X"1A",X"0F",X"11",X"A7",X"13",X"68",X"3B",X"34",X"F1",X"68",
		X"D7",X"F1",X"DC",X"0F",X"68",X"F1",X"88",X"57",X"A5",X"BF",X"34",X"D7",X"ED",X"B9",X"3A",X"AB",
		X"A9",X"21",X"8C",X"17",X"06",X"1E",X"86",X"23",X"10",X"FC",X"C6",X"2C",X"32",X"AB",X"A9",X"3A",
		X"32",X"AD",X"A7",X"11",X"1B",X"AD",X"3A",X"14",X"AD",X"28",X"06",X"11",X"2B",X"AD",X"3A",X"24",
		X"AD",X"87",X"21",X"8D",X"0F",X"CF",X"12",X"32",X"0B",X"AD",X"23",X"13",X"7E",X"12",X"21",X"0C",
		X"AD",X"BE",X"77",X"CC",X"1A",X"0F",X"CD",X"E1",X"01",X"C3",X"1A",X"0F",X"3A",X"32",X"AD",X"A7",
		X"11",X"1B",X"AD",X"3A",X"14",X"AD",X"28",X"06",X"11",X"2B",X"AD",X"3A",X"24",X"AD",X"87",X"21",
		X"8D",X"0F",X"DF",X"ED",X"A0",X"ED",X"A0",X"C9",X"0E",X"00",X"FD",X"46",X"31",X"5E",X"2D",X"7E",
		X"90",X"30",X"04",X"ED",X"44",X"CB",X"C1",X"57",X"FD",X"46",X"00",X"7B",X"90",X"30",X"04",X"ED",
		X"44",X"CB",X"C9",X"5F",X"08",X"7B",X"08",X"92",X"28",X"35",X"30",X"02",X"CB",X"D1",X"2E",X"00",
		X"CB",X"51",X"20",X"03",X"62",X"18",X"02",X"63",X"5A",X"06",X"08",X"AF",X"ED",X"6A",X"7C",X"38",
		X"03",X"BB",X"38",X"03",X"93",X"67",X"AF",X"3F",X"10",X"F2",X"45",X"79",X"21",X"15",X"34",X"DF",
		X"78",X"0F",X"0F",X"E6",X"1F",X"CB",X"6E",X"28",X"04",X"47",X"3E",X"1F",X"90",X"86",X"C9",X"21",
		X"1D",X"34",X"79",X"CF",X"C9",X"20",X"40",X"C0",X"A0",X"00",X"60",X"E0",X"80",X"20",X"60",X"E0",
		X"A0",X"21",X"50",X"0C",X"CD",X"8C",X"01",X"EB",X"5E",X"23",X"56",X"23",X"23",X"3A",X"0C",X"AD",
		X"C6",X"05",X"E6",X"0F",X"4F",X"C3",X"FF",X"0B",X"6F",X"34",X"8F",X"34",X"AF",X"34",X"CF",X"34",
		X"EF",X"34",X"0F",X"35",X"2F",X"35",X"4F",X"35",X"6F",X"35",X"8F",X"35",X"AF",X"35",X"CF",X"35",
		X"EF",X"35",X"0F",X"36",X"2F",X"36",X"4F",X"36",X"6F",X"36",X"8F",X"36",X"11",X"A7",X"13",X"68",
		X"3B",X"34",X"F1",X"88",X"57",X"A5",X"BF",X"34",X"D7",X"F1",X"68",X"3B",X"57",X"BF",X"B9",X"11",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"11",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0D",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0C",X"0D",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0C",X"0D",X"0D",X"11",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"10",X"10",X"10",X"11",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"10",X"10",X"10",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"11",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"10",X"10",X"10",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"10",X"10",X"10",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0D",X"10",X"10",X"10",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0D",X"10",X"10",X"10",X"3A",
		X"C6",X"AC",X"A7",X"C0",X"3A",X"04",X"AD",X"FE",X"04",X"CA",X"6E",X"38",X"21",X"05",X"AD",X"3A",
		X"06",X"AD",X"E6",X"0F",X"FE",X"07",X"CA",X"55",X"38",X"DA",X"BD",X"37",X"FE",X"09",X"DA",X"9F",
		X"37",X"7E",X"A7",X"C0",X"CD",X"4B",X"4B",X"0F",X"3A",X"04",X"AD",X"8F",X"21",X"C2",X"AC",X"36",
		X"FF",X"23",X"77",X"3A",X"02",X"A8",X"C6",X"08",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"21",X"D9",
		X"38",X"DF",X"4E",X"3A",X"C3",X"AC",X"87",X"87",X"87",X"87",X"21",X"7B",X"39",X"DF",X"EB",X"3A",
		X"C1",X"AC",X"47",X"3A",X"02",X"AD",X"A7",X"20",X"02",X"06",X"05",X"AF",X"32",X"11",X"A8",X"DD",
		X"21",X"50",X"A8",X"FD",X"21",X"1A",X"AA",X"DD",X"7E",X"00",X"A7",X"C2",X"68",X"37",X"1A",X"81",
		X"87",X"21",X"E9",X"38",X"CF",X"FD",X"77",X"31",X"23",X"7E",X"FD",X"77",X"00",X"3A",X"02",X"A8",
		X"C6",X"80",X"DD",X"77",X"01",X"DD",X"77",X"02",X"CD",X"2D",X"38",X"C6",X"09",X"DD",X"77",X"0A",
		X"13",X"1A",X"DD",X"77",X"0E",X"13",X"DD",X"36",X"03",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",
		X"09",X"20",X"D9",X"CD",X"3A",X"32",X"D9",X"DD",X"36",X"00",X"FE",X"DD",X"7E",X"0E",X"A7",X"20",
		X"03",X"DD",X"34",X"00",X"21",X"11",X"A8",X"34",X"EB",X"11",X"10",X"00",X"DD",X"19",X"FD",X"23",
		X"FD",X"23",X"EB",X"10",X"A2",X"AF",X"32",X"C2",X"AC",X"3E",X"E4",X"32",X"12",X"A8",X"21",X"11",
		X"A8",X"7E",X"FE",X"05",X"D2",X"17",X"58",X"21",X"C1",X"AC",X"BE",X"7E",X"32",X"11",X"A8",X"D2",
		X"17",X"58",X"C9",X"06",X"05",X"DD",X"21",X"90",X"A8",X"FD",X"21",X"22",X"AA",X"18",X"37",X"7E",
		X"A7",X"28",X"03",X"FE",X"30",X"C0",X"21",X"50",X"A8",X"11",X"10",X"00",X"01",X"00",X"07",X"7E",
		X"A7",X"28",X"01",X"0C",X"19",X"10",X"F8",X"79",X"FE",X"02",X"D0",X"18",X"07",X"7E",X"A7",X"28",
		X"03",X"FE",X"30",X"C0",X"3A",X"02",X"AD",X"A7",X"28",X"C9",X"3A",X"C1",X"AC",X"47",X"DD",X"21",
		X"B0",X"A8",X"FD",X"21",X"26",X"AA",X"DD",X"7E",X"00",X"A7",X"C2",X"47",X"38",X"DD",X"35",X"00",
		X"3A",X"02",X"A8",X"0F",X"0F",X"E6",X"3F",X"4F",X"CD",X"4B",X"4B",X"E6",X"0F",X"D6",X"08",X"81",
		X"E6",X"3F",X"21",X"FB",X"39",X"CF",X"87",X"87",X"21",X"3B",X"3A",X"CF",X"FD",X"77",X"31",X"23",
		X"7E",X"FD",X"77",X"00",X"3A",X"02",X"A8",X"C6",X"80",X"DD",X"77",X"01",X"DD",X"77",X"02",X"CD",
		X"2D",X"38",X"DD",X"77",X"0A",X"AF",X"32",X"C5",X"AC",X"DD",X"36",X"03",X"00",X"DD",X"36",X"05",
		X"00",X"DD",X"36",X"09",X"20",X"CD",X"3A",X"32",X"DD",X"36",X"0E",X"00",X"C9",X"CD",X"4B",X"4B",
		X"21",X"C4",X"AC",X"BE",X"30",X"0C",X"21",X"CF",X"A9",X"7E",X"3C",X"FE",X"05",X"38",X"01",X"AF",
		X"77",X"C9",X"E6",X"03",X"C6",X"05",X"C9",X"11",X"F0",X"FF",X"DD",X"19",X"FD",X"2B",X"FD",X"2B",
		X"05",X"C2",X"D6",X"37",X"C9",X"7E",X"A7",X"C0",X"DD",X"21",X"50",X"A8",X"11",X"10",X"00",X"06",
		X"05",X"DD",X"36",X"08",X"11",X"DD",X"36",X"09",X"00",X"DD",X"19",X"10",X"F4",X"C9",X"DD",X"21",
		X"50",X"A8",X"FD",X"21",X"1A",X"AA",X"3A",X"C1",X"AC",X"47",X"3A",X"0D",X"AD",X"A7",X"28",X"02",
		X"06",X"05",X"C5",X"DD",X"7E",X"00",X"A7",X"C2",X"C0",X"38",X"CD",X"4B",X"4B",X"E6",X"FC",X"21",
		X"3B",X"3A",X"CF",X"FD",X"77",X"31",X"23",X"7E",X"FD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",
		X"DD",X"77",X"02",X"3A",X"C1",X"AC",X"90",X"21",X"D2",X"38",X"CF",X"DD",X"77",X"0A",X"DD",X"36",
		X"09",X"20",X"CD",X"3A",X"32",X"DD",X"36",X"04",X"01",X"DD",X"36",X"0E",X"00",X"DD",X"35",X"00",
		X"11",X"10",X"00",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"C1",X"10",X"B6",X"3E",X"E4",X"32",X"12",
		X"A8",X"C9",X"0A",X"0B",X"0D",X"0E",X"0F",X"09",X"0C",X"08",X"0C",X"0F",X"13",X"16",X"1A",X"1D",
		X"21",X"24",X"28",X"2B",X"2F",X"33",X"37",X"3A",X"3D",X"F0",X"10",X"F0",X"20",X"F0",X"30",X"F0",
		X"40",X"F0",X"50",X"F0",X"60",X"F0",X"70",X"F0",X"80",X"F0",X"90",X"F0",X"A0",X"F0",X"B0",X"F0",
		X"C0",X"F0",X"D0",X"F0",X"E0",X"F0",X"F0",X"E0",X"F8",X"D0",X"F8",X"C0",X"F8",X"B0",X"F8",X"A0",
		X"F8",X"90",X"F8",X"80",X"F8",X"70",X"F8",X"60",X"F8",X"50",X"F8",X"40",X"F8",X"30",X"F8",X"20",
		X"F8",X"10",X"F8",X"00",X"F0",X"00",X"E0",X"00",X"D0",X"00",X"C0",X"00",X"B0",X"00",X"A0",X"00",
		X"90",X"00",X"80",X"00",X"70",X"00",X"60",X"00",X"50",X"00",X"40",X"00",X"30",X"00",X"20",X"00",
		X"10",X"10",X"10",X"20",X"10",X"30",X"10",X"40",X"10",X"50",X"10",X"60",X"10",X"70",X"10",X"80",
		X"10",X"90",X"10",X"A0",X"10",X"B0",X"10",X"C0",X"10",X"D0",X"10",X"E0",X"10",X"F0",X"10",X"F0",
		X"20",X"F0",X"30",X"F0",X"40",X"F0",X"50",X"F0",X"60",X"F0",X"70",X"F0",X"80",X"F0",X"90",X"F0",
		X"A0",X"F0",X"B0",X"F0",X"C0",X"F0",X"D0",X"F0",X"E0",X"F0",X"F0",X"00",X"01",X"01",X"11",X"FF",
		X"11",X"02",X"21",X"FE",X"21",X"03",X"31",X"FD",X"31",X"00",X"00",X"00",X"11",X"01",X"01",X"FF",
		X"01",X"02",X"11",X"FE",X"11",X"03",X"21",X"FD",X"21",X"00",X"00",X"00",X"01",X"02",X"11",X"FE",
		X"11",X"03",X"21",X"FD",X"21",X"04",X"31",X"FC",X"31",X"00",X"00",X"00",X"31",X"03",X"01",X"FD",
		X"01",X"04",X"11",X"FC",X"11",X"03",X"11",X"FD",X"11",X"00",X"00",X"00",X"01",X"03",X"01",X"FD",
		X"01",X"04",X"11",X"FC",X"11",X"05",X"21",X"FB",X"21",X"00",X"00",X"00",X"01",X"03",X"11",X"FD",
		X"11",X"00",X"21",X"03",X"21",X"FD",X"21",X"00",X"31",X"00",X"00",X"03",X"01",X"FD",X"01",X"03",
		X"11",X"FD",X"11",X"05",X"11",X"FB",X"11",X"00",X"29",X"00",X"00",X"00",X"01",X"03",X"11",X"FD",
		X"11",X"05",X"21",X"FB",X"21",X"03",X"31",X"FD",X"31",X"00",X"00",X"08",X"09",X"0A",X"0B",X"0C",
		X"0D",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",
		X"1B",X"1B",X"1C",X"1D",X"1E",X"1F",X"20",X"21",X"22",X"22",X"23",X"24",X"25",X"26",X"27",X"28",
		X"29",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",
		X"38",X"38",X"39",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"F0",X"10",X"60",X"00",X"F0",
		X"20",X"80",X"00",X"F0",X"30",X"80",X"00",X"F0",X"40",X"80",X"00",X"F0",X"50",X"80",X"00",X"F0",
		X"60",X"80",X"00",X"F0",X"70",X"80",X"00",X"F0",X"80",X"80",X"00",X"F0",X"90",X"80",X"00",X"F0",
		X"A0",X"80",X"00",X"F0",X"B0",X"80",X"00",X"F0",X"C0",X"80",X"00",X"F0",X"D0",X"80",X"00",X"F0",
		X"E0",X"80",X"00",X"F0",X"F0",X"A0",X"00",X"E0",X"F8",X"C0",X"00",X"D0",X"F8",X"C0",X"00",X"C0",
		X"F8",X"C0",X"00",X"B0",X"F8",X"C0",X"00",X"A0",X"F8",X"C0",X"00",X"90",X"F8",X"C0",X"00",X"80",
		X"F8",X"C0",X"00",X"70",X"F8",X"C0",X"00",X"60",X"F8",X"C0",X"00",X"50",X"F8",X"C0",X"00",X"40",
		X"F8",X"C0",X"00",X"30",X"F8",X"C0",X"00",X"20",X"F8",X"C0",X"00",X"10",X"F8",X"C0",X"00",X"00",
		X"F0",X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"10",X"20",X"00",X"10",X"10",X"40",X"00",X"20",
		X"10",X"40",X"00",X"30",X"10",X"40",X"00",X"40",X"10",X"40",X"00",X"50",X"10",X"40",X"00",X"60",
		X"10",X"40",X"00",X"70",X"10",X"40",X"00",X"80",X"10",X"40",X"00",X"90",X"10",X"40",X"00",X"A0",
		X"10",X"40",X"00",X"B0",X"10",X"40",X"00",X"C0",X"10",X"40",X"00",X"D0",X"10",X"40",X"00",X"E0",
		X"10",X"40",X"00",X"F0",X"10",X"60",X"00",X"F0",X"20",X"80",X"00",X"F0",X"30",X"80",X"00",X"F0",
		X"40",X"80",X"00",X"F0",X"50",X"80",X"00",X"F0",X"60",X"80",X"00",X"F0",X"70",X"80",X"00",X"F0",
		X"80",X"80",X"00",X"F0",X"90",X"80",X"00",X"F0",X"A0",X"80",X"00",X"F0",X"B0",X"80",X"00",X"F0",
		X"C0",X"80",X"00",X"F0",X"D0",X"80",X"00",X"F0",X"E0",X"80",X"00",X"F0",X"F0",X"A0",X"00",X"3A",
		X"04",X"AD",X"3D",X"C0",X"DD",X"21",X"C0",X"A8",X"FD",X"21",X"28",X"AA",X"DD",X"7E",X"00",X"A7",
		X"CA",X"25",X"3C",X"3C",X"C2",X"94",X"3B",X"CD",X"05",X"3E",X"FD",X"7E",X"31",X"C6",X"10",X"FD",
		X"77",X"33",X"FD",X"7E",X"00",X"FD",X"77",X"02",X"CD",X"C4",X"3C",X"DA",X"0D",X"3C",X"CD",X"E9",
		X"3C",X"C3",X"25",X"3D",X"3D",X"4F",X"21",X"DC",X"A8",X"7E",X"A7",X"CA",X"A9",X"3B",X"35",X"DD",
		X"36",X"00",X"FF",X"CD",X"83",X"56",X"C3",X"77",X"3B",X"79",X"FE",X"61",X"38",X"0F",X"DD",X"36",
		X"00",X"61",X"CD",X"83",X"56",X"FD",X"36",X"30",X"3D",X"FD",X"36",X"32",X"3D",X"DD",X"35",X"00",
		X"28",X"4B",X"CD",X"60",X"2B",X"FD",X"7E",X"31",X"C6",X"10",X"FD",X"77",X"33",X"FD",X"7E",X"00",
		X"FD",X"77",X"02",X"DD",X"7E",X"00",X"D6",X"40",X"CA",X"F1",X"3B",X"D8",X"4F",X"E6",X"07",X"C0",
		X"79",X"0F",X"0F",X"0F",X"3D",X"21",X"09",X"3C",X"CF",X"FD",X"77",X"03",X"3C",X"FD",X"77",X"01",
		X"C9",X"11",X"0B",X"04",X"FF",X"FD",X"36",X"03",X"FA",X"FD",X"36",X"01",X"FB",X"FD",X"36",X"30",
		X"6C",X"FD",X"36",X"32",X"6C",X"DD",X"35",X"00",X"C9",X"96",X"94",X"92",X"90",X"AF",X"DD",X"77",
		X"00",X"DD",X"77",X"10",X"FD",X"77",X"00",X"FD",X"77",X"31",X"32",X"5B",X"AA",X"32",X"2A",X"AA",
		X"DD",X"36",X"0E",X"80",X"C9",X"3A",X"80",X"A9",X"E6",X"01",X"C0",X"DD",X"35",X"0E",X"CA",X"32",
		X"3C",X"C9",X"3A",X"0D",X"AD",X"A7",X"C0",X"3A",X"02",X"A8",X"47",X"C6",X"08",X"E6",X"7F",X"FE",
		X"10",X"38",X"32",X"78",X"0F",X"0F",X"E6",X"3E",X"21",X"84",X"3C",X"CF",X"FD",X"77",X"31",X"23",
		X"7E",X"FD",X"77",X"00",X"78",X"C6",X"C0",X"E6",X"80",X"DD",X"77",X"02",X"CD",X"42",X"59",X"DD",
		X"73",X"0A",X"DD",X"72",X"0B",X"DD",X"71",X"0C",X"DD",X"70",X"0D",X"3E",X"03",X"32",X"DC",X"A8",
		X"DD",X"36",X"00",X"FF",X"C9",X"3A",X"80",X"A9",X"4F",X"3E",X"10",X"CB",X"59",X"20",X"02",X"ED",
		X"44",X"80",X"18",X"C0",X"EC",X"80",X"EC",X"88",X"EC",X"90",X"EC",X"A0",X"EC",X"B0",X"EC",X"C0",
		X"EC",X"D0",X"EC",X"E0",X"F0",X"EC",X"F0",X"EC",X"F0",X"E0",X"F0",X"D0",X"F0",X"C0",X"F0",X"B0",
		X"F0",X"A0",X"F0",X"90",X"F0",X"80",X"F0",X"78",X"F0",X"70",X"F0",X"60",X"F0",X"50",X"F0",X"40",
		X"F0",X"30",X"F0",X"28",X"F0",X"20",X"EC",X"20",X"EC",X"30",X"EC",X"40",X"EC",X"50",X"EC",X"60",
		X"EC",X"70",X"EC",X"78",X"DD",X"7E",X"02",X"C6",X"40",X"CB",X"7F",X"C2",X"D9",X"3C",X"FD",X"7E",
		X"31",X"C6",X"13",X"FE",X"03",X"D8",X"C3",X"E1",X"3C",X"FD",X"7E",X"31",X"C6",X"10",X"FE",X"03",
		X"D8",X"FD",X"7E",X"00",X"C6",X"02",X"FE",X"04",X"C9",X"3A",X"80",X"A9",X"E6",X"02",X"47",X"3A",
		X"DC",X"A8",X"4F",X"3E",X"03",X"91",X"87",X"87",X"C6",X"A0",X"80",X"4F",X"DD",X"7E",X"02",X"C6",
		X"40",X"FE",X"80",X"38",X"10",X"FD",X"71",X"01",X"0C",X"FD",X"71",X"03",X"FD",X"36",X"30",X"ED",
		X"FD",X"36",X"32",X"ED",X"C9",X"FD",X"71",X"03",X"0C",X"FD",X"71",X"01",X"FD",X"36",X"30",X"6D",
		X"FD",X"36",X"32",X"6D",X"C9",X"DD",X"7E",X"00",X"3C",X"C0",X"3A",X"F4",X"A8",X"A7",X"C0",X"3A",
		X"C6",X"A8",X"A7",X"C8",X"FE",X"01",X"CA",X"40",X"3D",X"3A",X"E0",X"A8",X"A7",X"CA",X"45",X"3D",
		X"3A",X"40",X"A8",X"A7",X"C0",X"06",X"02",X"3A",X"D6",X"A8",X"57",X"87",X"5F",X"3E",X"84",X"FD",
		X"96",X"00",X"82",X"BB",X"D2",X"6F",X"3D",X"3E",X"78",X"FD",X"96",X"31",X"82",X"BB",X"D2",X"6F",
		X"3D",X"D9",X"11",X"10",X"00",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"D9",X"10",X"DF",X"C9",X"CD",
		X"5F",X"56",X"21",X"7F",X"AC",X"CD",X"B8",X"33",X"67",X"3E",X"18",X"EB",X"21",X"D4",X"A8",X"34",
		X"46",X"CB",X"40",X"20",X"02",X"ED",X"44",X"EB",X"84",X"08",X"FD",X"46",X"31",X"FD",X"4E",X"00",
		X"3A",X"C6",X"A8",X"FE",X"01",X"CA",X"9F",X"3D",X"3A",X"E0",X"A8",X"A7",X"CA",X"CF",X"3D",X"DD",
		X"21",X"40",X"A8",X"FD",X"21",X"18",X"AA",X"FD",X"70",X"31",X"FD",X"71",X"00",X"08",X"CD",X"C5",
		X"59",X"DD",X"73",X"0A",X"DD",X"72",X"0B",X"DD",X"71",X"0C",X"DD",X"70",X"0D",X"FD",X"36",X"01",
		X"4D",X"FD",X"36",X"30",X"62",X"DD",X"35",X"00",X"3A",X"F6",X"A8",X"32",X"F4",X"A8",X"C9",X"DD",
		X"21",X"E0",X"A8",X"FD",X"21",X"2C",X"AA",X"C3",X"A7",X"3D",X"3A",X"04",X"AD",X"3D",X"C0",X"DD",
		X"21",X"E0",X"A8",X"FD",X"21",X"2C",X"AA",X"CD",X"EB",X"3D",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",
		X"3C",X"C2",X"FB",X"3D",X"CD",X"05",X"3E",X"CD",X"83",X"2B",X"D0",X"CD",X"AB",X"40",X"3A",X"F6",
		X"A8",X"DD",X"77",X"0E",X"C9",X"DD",X"66",X"0B",X"DD",X"6E",X"0A",X"ED",X"5B",X"08",X"A8",X"19",
		X"FD",X"56",X"31",X"DD",X"5E",X"03",X"19",X"FD",X"74",X"31",X"DD",X"75",X"03",X"DD",X"66",X"0D",
		X"DD",X"6E",X"0C",X"ED",X"5B",X"0A",X"A8",X"19",X"FD",X"56",X"00",X"DD",X"5E",X"05",X"19",X"FD",
		X"74",X"00",X"DD",X"75",X"05",X"C9",X"DD",X"21",X"10",X"A8",X"FD",X"21",X"12",X"AA",X"CD",X"63",
		X"3E",X"DD",X"21",X"20",X"A8",X"FD",X"21",X"14",X"AA",X"CD",X"63",X"3E",X"DD",X"21",X"30",X"A8",
		X"FD",X"21",X"16",X"AA",X"CD",X"63",X"3E",X"DD",X"21",X"40",X"A8",X"FD",X"21",X"18",X"AA",X"CD",
		X"63",X"3E",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"3C",X"C2",X"8E",X"3E",X"3A",X"04",X"AD",X"FE",
		X"04",X"CC",X"7E",X"3E",X"CD",X"05",X"3E",X"CD",X"83",X"2B",X"D0",X"C3",X"AB",X"40",X"3A",X"80",
		X"A9",X"0F",X"E6",X"07",X"C6",X"40",X"FD",X"77",X"01",X"FD",X"36",X"30",X"44",X"C9",X"3A",X"04",
		X"AD",X"FE",X"04",X"28",X"03",X"C3",X"AB",X"40",X"DD",X"7E",X"00",X"FE",X"01",X"CA",X"AB",X"40",
		X"DD",X"35",X"00",X"FE",X"3C",X"D4",X"CB",X"3E",X"CD",X"60",X"2B",X"DD",X"7E",X"00",X"FE",X"1C",
		X"D8",X"D6",X"1C",X"0F",X"0F",X"E6",X"07",X"21",X"C3",X"3E",X"CF",X"FD",X"77",X"01",X"FD",X"36",
		X"30",X"03",X"C9",X"FF",X"E6",X"E7",X"E7",X"E6",X"E6",X"E5",X"E4",X"DD",X"36",X"00",X"3B",X"C3",
		X"83",X"56",X"92",X"A6",X"14",X"B9",X"3A",X"80",X"A9",X"E6",X"07",X"C6",X"05",X"DD",X"BE",X"0F",
		X"C0",X"3A",X"17",X"A8",X"A7",X"C0",X"21",X"10",X"A8",X"11",X"12",X"AA",X"3A",X"44",X"A8",X"A7",
		X"C8",X"47",X"7E",X"A7",X"28",X"09",X"7D",X"C6",X"10",X"6F",X"1C",X"1C",X"10",X"F4",X"C9",X"22",
		X"91",X"A9",X"ED",X"53",X"93",X"A9",X"3A",X"27",X"A8",X"47",X"87",X"4F",X"3E",X"78",X"FD",X"96",
		X"31",X"80",X"B9",X"30",X"08",X"3E",X"84",X"FD",X"96",X"00",X"80",X"B9",X"D8",X"3A",X"37",X"A8",
		X"47",X"87",X"4F",X"3A",X"02",X"A8",X"DD",X"96",X"02",X"80",X"B9",X"D0",X"7A",X"FE",X"02",X"CA",
		X"9E",X"3F",X"21",X"7F",X"AC",X"CD",X"B8",X"33",X"4F",X"DD",X"96",X"02",X"C6",X"10",X"FE",X"20",
		X"D0",X"CD",X"93",X"3F",X"DD",X"E5",X"FD",X"E5",X"FD",X"56",X"31",X"FD",X"5E",X"00",X"DD",X"2A",
		X"91",X"A9",X"FD",X"2A",X"93",X"A9",X"FD",X"72",X"31",X"FD",X"73",X"00",X"3A",X"04",X"AD",X"A7",
		X"79",X"20",X"05",X"CD",X"CB",X"59",X"18",X"03",X"CD",X"D1",X"59",X"DD",X"73",X"0A",X"DD",X"72",
		X"0B",X"DD",X"71",X"0C",X"DD",X"70",X"0D",X"FD",X"7E",X"31",X"FD",X"7E",X"00",X"FD",X"36",X"01",
		X"4D",X"FD",X"36",X"30",X"62",X"3A",X"14",X"A8",X"32",X"17",X"A8",X"DD",X"35",X"00",X"FD",X"E1",
		X"DD",X"E1",X"C9",X"3A",X"04",X"AD",X"FE",X"03",X"DA",X"5F",X"56",X"C3",X"69",X"56",X"3A",X"E6",
		X"A8",X"47",X"87",X"4F",X"3E",X"84",X"FD",X"96",X"00",X"80",X"B9",X"D0",X"C3",X"32",X"3F",X"DD",
		X"7E",X"02",X"C6",X"08",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"21",X"CA",X"3F",X"CF",X"FD",X"77",
		X"01",X"11",X"10",X"00",X"19",X"7E",X"FD",X"77",X"30",X"C9",X"48",X"49",X"4A",X"4B",X"4C",X"4B",
		X"4A",X"49",X"48",X"49",X"4A",X"4B",X"4C",X"4B",X"4A",X"49",X"F4",X"B4",X"B4",X"B4",X"B4",X"34",
		X"34",X"34",X"34",X"74",X"74",X"74",X"74",X"F4",X"F4",X"F4",X"3A",X"04",X"AD",X"A7",X"C0",X"DD",
		X"21",X"C0",X"A8",X"FD",X"21",X"28",X"AA",X"06",X"03",X"DD",X"7E",X"00",X"A7",X"CA",X"0B",X"40",
		X"3C",X"20",X"05",X"CD",X"17",X"40",X"18",X"03",X"CD",X"6C",X"40",X"11",X"10",X"00",X"DD",X"19",
		X"FD",X"23",X"FD",X"23",X"10",X"E3",X"C9",X"FD",X"56",X"31",X"DD",X"5E",X"03",X"DD",X"7E",X"01",
		X"A7",X"28",X"05",X"21",X"80",X"FE",X"18",X"03",X"21",X"80",X"01",X"19",X"ED",X"5B",X"08",X"A8",
		X"19",X"FD",X"74",X"31",X"DD",X"75",X"03",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"11",X"09",X"00",
		X"19",X"DD",X"75",X"07",X"DD",X"74",X"08",X"FD",X"56",X"00",X"DD",X"5E",X"05",X"19",X"ED",X"5B",
		X"0A",X"A8",X"19",X"FD",X"74",X"00",X"DD",X"75",X"05",X"FD",X"7E",X"31",X"C6",X"10",X"FE",X"20",
		X"DA",X"AB",X"40",X"FD",X"7E",X"00",X"FE",X"F8",X"D2",X"AB",X"40",X"C9",X"DD",X"7E",X"00",X"FE",
		X"3C",X"D4",X"9D",X"40",X"DD",X"35",X"00",X"28",X"32",X"CD",X"60",X"2B",X"DD",X"7E",X"00",X"FE",
		X"1C",X"D8",X"D6",X"1C",X"0F",X"0F",X"E6",X"0F",X"21",X"94",X"40",X"CF",X"FD",X"77",X"01",X"FD",
		X"36",X"30",X"0E",X"C9",X"FF",X"9A",X"99",X"98",X"98",X"99",X"99",X"9A",X"9B",X"DD",X"36",X"00",
		X"3B",X"3A",X"04",X"AD",X"A7",X"CA",X"8E",X"56",X"C3",X"8E",X"56",X"DD",X"36",X"00",X"00",X"FD",
		X"36",X"00",X"00",X"FD",X"36",X"31",X"00",X"C9",X"3A",X"04",X"AD",X"FE",X"02",X"D8",X"3A",X"80",
		X"A9",X"E6",X"1F",X"C0",X"3A",X"C0",X"A8",X"3C",X"C8",X"3A",X"D0",X"A8",X"3C",X"C8",X"3A",X"E0",
		X"A8",X"3C",X"C8",X"C3",X"79",X"56",X"3A",X"04",X"AD",X"FE",X"02",X"D8",X"DD",X"21",X"C0",X"A8",
		X"FD",X"21",X"28",X"AA",X"3A",X"C6",X"A8",X"A7",X"C8",X"47",X"DD",X"7E",X"00",X"A7",X"CA",X"0B",
		X"41",X"3C",X"20",X"14",X"3A",X"04",X"AD",X"FE",X"04",X"CA",X"94",X"41",X"DD",X"7E",X"0E",X"A7",
		X"C2",X"8B",X"41",X"CD",X"17",X"41",X"18",X"03",X"CD",X"3C",X"41",X"11",X"10",X"00",X"DD",X"19",
		X"FD",X"23",X"FD",X"23",X"10",X"D4",X"C9",X"C5",X"3A",X"80",X"A9",X"E6",X"0F",X"DD",X"BE",X"0F",
		X"20",X"09",X"21",X"7F",X"AC",X"CD",X"B8",X"33",X"DD",X"77",X"01",X"CD",X"01",X"42",X"CD",X"AA",
		X"58",X"CD",X"AF",X"3F",X"C1",X"CD",X"83",X"2B",X"D0",X"C3",X"AB",X"40",X"DD",X"7E",X"00",X"FE",
		X"3C",X"D4",X"9D",X"40",X"CD",X"60",X"2B",X"DD",X"35",X"00",X"CA",X"AB",X"40",X"DD",X"7E",X"00",
		X"FE",X"1C",X"D8",X"D6",X"1C",X"0F",X"0F",X"E6",X"07",X"57",X"3A",X"04",X"AD",X"FE",X"04",X"30",
		X"15",X"21",X"6E",X"41",X"7A",X"CF",X"FD",X"77",X"01",X"FD",X"36",X"30",X"0D",X"C9",X"FF",X"9E",
		X"9F",X"9F",X"9E",X"9E",X"9D",X"9C",X"21",X"83",X"41",X"7A",X"CF",X"FD",X"77",X"01",X"FD",X"36",
		X"30",X"02",X"C9",X"FF",X"E2",X"E3",X"E3",X"E2",X"E2",X"E1",X"E0",X"CD",X"6C",X"3E",X"DD",X"35",
		X"0E",X"C3",X"0B",X"41",X"DD",X"7E",X"04",X"A7",X"CA",X"A4",X"41",X"DD",X"35",X"04",X"CD",X"B8",
		X"41",X"C3",X"0B",X"41",X"C5",X"CD",X"B6",X"58",X"CD",X"F1",X"41",X"CD",X"83",X"2B",X"C1",X"D2",
		X"0B",X"41",X"CD",X"AB",X"40",X"C3",X"0B",X"41",X"C5",X"3A",X"80",X"A9",X"E6",X"0F",X"20",X"1F",
		X"21",X"75",X"AC",X"DD",X"CB",X"0F",X"46",X"20",X"03",X"21",X"79",X"AC",X"CD",X"B8",X"33",X"47",
		X"7A",X"FE",X"10",X"30",X"07",X"08",X"FE",X"10",X"DC",X"EC",X"41",X"08",X"DD",X"70",X"01",X"CD",
		X"1F",X"42",X"CD",X"B6",X"58",X"CD",X"F1",X"41",X"C1",X"C3",X"83",X"2B",X"DD",X"36",X"04",X"00",
		X"C9",X"3A",X"80",X"A9",X"0F",X"E6",X"07",X"C6",X"50",X"FD",X"77",X"01",X"FD",X"36",X"30",X"0A",
		X"C9",X"DD",X"7E",X"01",X"DD",X"96",X"02",X"C6",X"01",X"FE",X"02",X"D8",X"FE",X"80",X"DD",X"7E",
		X"02",X"30",X"06",X"C6",X"01",X"DD",X"77",X"02",X"C9",X"D6",X"01",X"DD",X"77",X"02",X"C9",X"3A",
		X"80",X"A9",X"E6",X"03",X"C8",X"DD",X"7E",X"01",X"DD",X"96",X"02",X"C6",X"01",X"FE",X"02",X"D8",
		X"FE",X"80",X"DD",X"7E",X"02",X"30",X"06",X"C6",X"02",X"DD",X"77",X"02",X"C9",X"D6",X"02",X"DD",
		X"77",X"02",X"C9",X"3A",X"80",X"A9",X"E6",X"07",X"C6",X"05",X"DD",X"BE",X"0F",X"C0",X"21",X"F4",
		X"A8",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"21",X"C0",X"A8",X"11",X"28",X"AA",X"3A",X"C6",X"A8",
		X"A7",X"C8",X"47",X"7E",X"A7",X"CA",X"71",X"42",X"7D",X"C6",X"10",X"6F",X"13",X"13",X"10",X"F3",
		X"C9",X"22",X"91",X"A9",X"ED",X"53",X"93",X"A9",X"3A",X"D6",X"A8",X"57",X"87",X"4F",X"3E",X"78",
		X"FD",X"96",X"31",X"82",X"B9",X"30",X"08",X"3E",X"84",X"FD",X"96",X"00",X"82",X"B9",X"D8",X"DD",
		X"4E",X"02",X"3A",X"04",X"AD",X"A7",X"CA",X"9C",X"42",X"C3",X"B7",X"42",X"3A",X"E6",X"A8",X"57",
		X"87",X"4F",X"3E",X"84",X"FD",X"96",X"00",X"82",X"B9",X"D0",X"3E",X"78",X"FD",X"96",X"31",X"38",
		X"04",X"0E",X"00",X"18",X"02",X"0E",X"01",X"FD",X"56",X"31",X"DD",X"5E",X"03",X"FD",X"66",X"00",
		X"DD",X"6E",X"05",X"D9",X"DD",X"E5",X"FD",X"E5",X"DD",X"2A",X"91",X"A9",X"FD",X"2A",X"93",X"A9",
		X"D9",X"DD",X"73",X"03",X"FD",X"72",X"31",X"DD",X"75",X"05",X"FD",X"74",X"00",X"DD",X"71",X"01",
		X"3A",X"04",X"AD",X"FE",X"04",X"CA",X"AE",X"43",X"A7",X"C2",X"13",X"43",X"FD",X"36",X"01",X"4F",
		X"79",X"0F",X"CB",X"2F",X"E6",X"C0",X"C6",X"0B",X"FD",X"77",X"30",X"DD",X"36",X"07",X"00",X"DD",
		X"36",X"08",X"FF",X"DD",X"35",X"00",X"3A",X"F6",X"A8",X"32",X"F4",X"A8",X"FD",X"E1",X"DD",X"E1",
		X"C3",X"64",X"56",X"3A",X"04",X"AD",X"FE",X"03",X"CA",X"6F",X"43",X"D2",X"4C",X"43",X"21",X"7F",
		X"AC",X"CD",X"B8",X"33",X"DD",X"77",X"01",X"DD",X"7E",X"0F",X"0F",X"E6",X"80",X"C6",X"40",X"DD",
		X"86",X"01",X"DD",X"77",X"02",X"CD",X"AF",X"3F",X"DD",X"35",X"00",X"3A",X"F6",X"A8",X"32",X"F4",
		X"A8",X"DD",X"36",X"0E",X"00",X"FD",X"E1",X"DD",X"E1",X"C3",X"6E",X"56",X"21",X"7F",X"AC",X"CD",
		X"B8",X"33",X"DD",X"77",X"01",X"DD",X"77",X"02",X"CD",X"AF",X"3F",X"DD",X"35",X"00",X"3A",X"F6",
		X"A8",X"32",X"F4",X"A8",X"DD",X"36",X"0E",X"00",X"FD",X"E1",X"DD",X"E1",X"C3",X"74",X"56",X"C5",
		X"79",X"C6",X"40",X"E6",X"80",X"79",X"20",X"07",X"C6",X"1A",X"DD",X"77",X"02",X"18",X"05",X"D6",
		X"1A",X"DD",X"77",X"02",X"CD",X"8E",X"59",X"DD",X"73",X"0A",X"DD",X"72",X"0B",X"DD",X"71",X"0C",
		X"DD",X"70",X"0D",X"C1",X"DD",X"71",X"02",X"CD",X"AF",X"3F",X"DD",X"36",X"0E",X"20",X"DD",X"35",
		X"00",X"3A",X"F6",X"A8",X"32",X"F4",X"A8",X"FD",X"E1",X"DD",X"E1",X"C3",X"6E",X"56",X"3A",X"E6",
		X"A8",X"DD",X"77",X"04",X"C3",X"13",X"43",X"3A",X"C6",X"AC",X"3C",X"C8",X"3A",X"0D",X"AD",X"A7",
		X"20",X"2E",X"3A",X"80",X"A9",X"E6",X"07",X"FE",X"05",X"C0",X"DD",X"21",X"A0",X"A8",X"FD",X"21",
		X"24",X"AA",X"3A",X"02",X"AD",X"DD",X"B6",X"00",X"DD",X"B6",X"10",X"C0",X"3E",X"FF",X"32",X"0D",
		X"AD",X"DD",X"36",X"04",X"07",X"C3",X"DB",X"46",X"AF",X"86",X"23",X"10",X"FC",X"C3",X"AD",X"07",
		X"DD",X"21",X"A0",X"A8",X"FD",X"21",X"24",X"AA",X"DD",X"7E",X"00",X"A7",X"CA",X"35",X"45",X"3C",
		X"C2",X"40",X"45",X"DD",X"66",X"0C",X"DD",X"6E",X"0D",X"ED",X"5B",X"08",X"A8",X"19",X"FD",X"56",
		X"31",X"DD",X"5E",X"03",X"19",X"FD",X"74",X"31",X"DD",X"75",X"03",X"DD",X"66",X"1C",X"DD",X"6E",
		X"1D",X"ED",X"5B",X"0A",X"A8",X"19",X"FD",X"56",X"00",X"DD",X"5E",X"05",X"19",X"FD",X"74",X"00",
		X"DD",X"75",X"05",X"FD",X"7E",X"31",X"C6",X"10",X"FD",X"77",X"33",X"FD",X"7E",X"00",X"FD",X"77",
		X"02",X"CD",X"47",X"44",X"C3",X"F0",X"46",X"CD",X"C4",X"3C",X"DA",X"DB",X"46",X"3A",X"04",X"AD",
		X"57",X"FE",X"04",X"CA",X"A2",X"44",X"7A",X"87",X"87",X"87",X"87",X"47",X"3A",X"80",X"A9",X"E6",
		X"02",X"80",X"47",X"3E",X"07",X"DD",X"96",X"04",X"0F",X"E6",X"03",X"5F",X"87",X"87",X"80",X"21",
		X"F1",X"44",X"DF",X"46",X"23",X"4E",X"21",X"31",X"45",X"7A",X"DF",X"56",X"DD",X"7E",X"02",X"C6",
		X"40",X"FE",X"80",X"38",X"10",X"FD",X"70",X"01",X"FD",X"71",X"03",X"7A",X"C6",X"80",X"FD",X"77",
		X"30",X"FD",X"77",X"32",X"C9",X"FD",X"71",X"01",X"FD",X"70",X"03",X"FD",X"72",X"30",X"FD",X"72",
		X"32",X"C9",X"DD",X"7E",X"04",X"5F",X"FE",X"07",X"CA",X"BF",X"44",X"DD",X"34",X"06",X"DD",X"4E",
		X"06",X"CB",X"79",X"20",X"14",X"7B",X"C6",X"02",X"B9",X"30",X"04",X"DD",X"36",X"06",X"80",X"FD",
		X"36",X"30",X"70",X"FD",X"36",X"32",X"70",X"18",X"13",X"79",X"E6",X"7F",X"FE",X"03",X"38",X"04",
		X"DD",X"36",X"06",X"00",X"FD",X"36",X"30",X"51",X"FD",X"36",X"32",X"51",X"11",X"02",X"02",X"21",
		X"D5",X"D4",X"3A",X"80",X"A9",X"CB",X"57",X"20",X"01",X"19",X"FD",X"75",X"01",X"FD",X"74",X"03",
		X"C9",X"39",X"38",X"39",X"38",X"3B",X"3A",X"3D",X"3C",X"3B",X"3A",X"3D",X"3C",X"3D",X"3C",X"3F",
		X"3E",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",
		X"BF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C6",X"C7",X"C8",X"C9",X"C8",X"C9",X"CA",
		X"CB",X"CC",X"CD",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"CE",X"CF",X"D0",X"D1",X"D0",X"D1",X"D2",
		X"D3",X"E9",X"58",X"6F",X"6E",X"DD",X"7E",X"0E",X"A7",X"CA",X"63",X"46",X"DD",X"35",X"0E",X"C9",
		X"4F",X"DD",X"7E",X"04",X"A7",X"28",X"0D",X"DD",X"35",X"04",X"DD",X"36",X"00",X"FF",X"CD",X"83",
		X"56",X"C3",X"03",X"44",X"79",X"FE",X"F0",X"C2",X"B3",X"45",X"AF",X"32",X"DC",X"A8",X"CD",X"34",
		X"56",X"CD",X"D2",X"56",X"21",X"10",X"A8",X"11",X"10",X"00",X"06",X"0F",X"0E",X"14",X"7E",X"3C",
		X"20",X"22",X"71",X"D9",X"11",X"02",X"04",X"FF",X"D9",X"19",X"79",X"C6",X"0A",X"4F",X"10",X"EE",
		X"0E",X"3C",X"3E",X"FE",X"32",X"C6",X"AC",X"DD",X"36",X"00",X"E4",X"FD",X"36",X"30",X"3D",X"FD",
		X"36",X"32",X"3D",X"C9",X"3C",X"20",X"E2",X"36",X"00",X"18",X"DE",X"16",X"A7",X"13",X"96",X"ED",
		X"DC",X"F1",X"8C",X"68",X"3B",X"0D",X"ED",X"F1",X"9B",X"13",X"13",X"13",X"13",X"F1",X"88",X"DC",
		X"ED",X"11",X"B9",X"CD",X"60",X"2B",X"FD",X"7E",X"31",X"47",X"C6",X"13",X"FE",X"03",X"38",X"15",
		X"78",X"C6",X"10",X"FD",X"77",X"33",X"FD",X"7E",X"00",X"47",X"C6",X"08",X"FE",X"28",X"38",X"05",
		X"FD",X"70",X"02",X"18",X"08",X"FD",X"36",X"01",X"FF",X"FD",X"36",X"03",X"FF",X"DD",X"7E",X"00",
		X"FE",X"B4",X"28",X"3F",X"38",X"13",X"D6",X"B4",X"0F",X"0F",X"0F",X"3D",X"E6",X"07",X"21",X"1B",
		X"46",X"CF",X"FD",X"77",X"03",X"3C",X"FD",X"77",X"01",X"DD",X"35",X"00",X"CA",X"46",X"46",X"DD",
		X"7E",X"00",X"FE",X"5A",X"C0",X"FD",X"36",X"01",X"FF",X"FD",X"36",X"03",X"FF",X"C9",X"21",X"7C",
		X"A6",X"7E",X"4F",X"3A",X"43",X"AB",X"91",X"C2",X"43",X"46",X"C9",X"94",X"96",X"96",X"94",X"92",
		X"90",X"90",X"94",X"DD",X"35",X"00",X"FD",X"36",X"01",X"FE",X"FD",X"36",X"03",X"FD",X"FD",X"36",
		X"30",X"6C",X"FD",X"36",X"32",X"6C",X"3A",X"00",X"A8",X"3C",X"CC",X"0B",X"58",X"11",X"0D",X"04",
		X"C3",X"38",X"00",X"C3",X"1B",X"46",X"3E",X"FF",X"32",X"C6",X"AC",X"DD",X"36",X"00",X"00",X"21",
		X"43",X"AB",X"7E",X"FE",X"7C",X"C2",X"60",X"46",X"23",X"7E",X"FE",X"10",X"C8",X"FE",X"05",X"C8",
		X"C3",X"9B",X"45",X"3A",X"C6",X"AC",X"A7",X"C0",X"3A",X"02",X"A8",X"47",X"3A",X"80",X"A9",X"4F",
		X"3E",X"10",X"CB",X"59",X"20",X"02",X"ED",X"44",X"80",X"0F",X"0F",X"E6",X"3E",X"21",X"84",X"3C",
		X"CF",X"FD",X"77",X"31",X"23",X"7E",X"FD",X"77",X"00",X"78",X"C6",X"C0",X"E6",X"80",X"DD",X"77",
		X"02",X"CD",X"BA",X"46",X"DD",X"7E",X"04",X"FE",X"06",X"30",X"04",X"DD",X"36",X"04",X"05",X"DD",
		X"36",X"00",X"FF",X"C3",X"F7",X"57",X"3A",X"80",X"A9",X"4F",X"E6",X"1C",X"CB",X"41",X"20",X"02",
		X"ED",X"44",X"80",X"0F",X"0F",X"E6",X"3E",X"C3",X"7D",X"46",X"21",X"CE",X"46",X"E5",X"3A",X"04",
		X"AD",X"E6",X"07",X"F7",X"42",X"59",X"4E",X"59",X"4E",X"59",X"65",X"59",X"6B",X"59",X"DD",X"72",
		X"0C",X"DD",X"73",X"0D",X"DD",X"70",X"1C",X"DD",X"71",X"1D",X"C9",X"AF",X"DD",X"77",X"00",X"FD",
		X"77",X"00",X"FD",X"77",X"02",X"FD",X"77",X"31",X"FD",X"77",X"33",X"DD",X"36",X"0E",X"5F",X"C9",
		X"DD",X"7E",X"00",X"3C",X"C0",X"3A",X"17",X"A8",X"A7",X"C0",X"06",X"02",X"3A",X"27",X"A8",X"57",
		X"87",X"5F",X"FD",X"7E",X"00",X"C6",X"08",X"FE",X"28",X"38",X"1B",X"FD",X"7E",X"31",X"C6",X"10",
		X"FE",X"20",X"38",X"12",X"3E",X"84",X"FD",X"96",X"00",X"82",X"BB",X"30",X"17",X"3E",X"78",X"FD",
		X"96",X"31",X"82",X"BB",X"30",X"0E",X"D9",X"11",X"10",X"00",X"DD",X"19",X"FD",X"23",X"FD",X"23",
		X"D9",X"10",X"CF",X"C9",X"21",X"30",X"A8",X"D9",X"21",X"16",X"AA",X"06",X"02",X"D9",X"7E",X"A7",
		X"28",X"0A",X"11",X"10",X"00",X"19",X"D9",X"23",X"23",X"10",X"F2",X"C9",X"22",X"91",X"A9",X"D9",
		X"22",X"93",X"A9",X"CD",X"5F",X"56",X"21",X"7F",X"AC",X"CD",X"B8",X"33",X"67",X"EB",X"21",X"B4",
		X"A8",X"34",X"3E",X"18",X"CB",X"46",X"20",X"02",X"ED",X"44",X"EB",X"84",X"FD",X"46",X"31",X"FD",
		X"4E",X"00",X"DD",X"2A",X"91",X"A9",X"FD",X"2A",X"93",X"A9",X"DD",X"77",X"02",X"FD",X"70",X"31",
		X"FD",X"71",X"00",X"21",X"95",X"47",X"E5",X"3A",X"04",X"AD",X"F7",X"8E",X"59",X"8E",X"59",X"94",
		X"59",X"94",X"59",X"94",X"59",X"DD",X"73",X"0A",X"DD",X"72",X"0B",X"DD",X"71",X"0C",X"DD",X"70",
		X"0D",X"FD",X"36",X"01",X"4D",X"FD",X"36",X"30",X"62",X"DD",X"35",X"00",X"3A",X"14",X"A8",X"32",
		X"17",X"A8",X"C9",X"3A",X"04",X"AD",X"FE",X"04",X"C8",X"DD",X"21",X"F0",X"A8",X"FD",X"21",X"2E",
		X"AA",X"DD",X"7E",X"00",X"A7",X"CA",X"53",X"48",X"3C",X"C2",X"F2",X"47",X"CD",X"05",X"3E",X"CD",
		X"83",X"2B",X"DA",X"AD",X"48",X"3A",X"80",X"A9",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"21",X"EA",
		X"47",X"CF",X"FD",X"77",X"01",X"FD",X"36",X"30",X"75",X"C9",X"00",X"01",X"02",X"03",X"03",X"02",
		X"01",X"00",X"CD",X"60",X"2B",X"DD",X"7E",X"00",X"FE",X"10",X"CA",X"31",X"48",X"FE",X"3C",X"D2",
		X"09",X"48",X"DD",X"35",X"00",X"C0",X"C3",X"AD",X"48",X"DD",X"36",X"00",X"3B",X"CD",X"FF",X"57",
		X"DD",X"7E",X"07",X"FE",X"04",X"D2",X"24",X"48",X"21",X"2D",X"48",X"CF",X"FD",X"77",X"01",X"FD",
		X"36",X"30",X"6C",X"C9",X"FD",X"36",X"01",X"8F",X"FD",X"36",X"30",X"6C",X"C9",X"F9",X"FC",X"8D",
		X"8E",X"DD",X"35",X"00",X"DD",X"7E",X"07",X"DD",X"34",X"07",X"FE",X"04",X"D2",X"49",X"48",X"21",
		X"4F",X"48",X"DF",X"5E",X"16",X"04",X"C3",X"38",X"00",X"11",X"0F",X"04",X"C3",X"38",X"00",X"0A",
		X"0C",X"0D",X"0E",X"3A",X"0D",X"AD",X"A7",X"C0",X"3A",X"80",X"A9",X"E6",X"01",X"C8",X"DD",X"35",
		X"0E",X"C0",X"3A",X"02",X"A8",X"C6",X"08",X"0F",X"0F",X"0F",X"E6",X"1E",X"21",X"8D",X"48",X"CF",
		X"FD",X"77",X"31",X"23",X"7E",X"FD",X"77",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"00",
		X"DD",X"36",X"0C",X"40",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"00",X"FF",X"C9",X"F0",X"40",X"F0",
		X"80",X"F0",X"F8",X"60",X"F8",X"80",X"F8",X"A0",X"F8",X"10",X"F8",X"00",X"80",X"00",X"90",X"10",
		X"10",X"30",X"10",X"60",X"10",X"80",X"10",X"A0",X"10",X"C0",X"10",X"F0",X"28",X"DD",X"36",X"00",
		X"00",X"FD",X"36",X"00",X"00",X"FD",X"36",X"31",X"00",X"DD",X"36",X"0E",X"F0",X"C9",X"CD",X"E7",
		X"48",X"CD",X"41",X"49",X"CD",X"11",X"49",X"CD",X"84",X"49",X"CD",X"D6",X"49",X"C9",X"2C",X"A7",
		X"13",X"FD",X"3B",X"88",X"0D",X"DC",X"F1",X"BF",X"68",X"0D",X"D7",X"F1",X"FD",X"3B",X"FD",X"DC",
		X"FD",X"A5",X"57",X"ED",X"F1",X"52",X"B9",X"3A",X"AE",X"A9",X"0F",X"0F",X"0F",X"21",X"83",X"A9",
		X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"CD",X"F1",X"57",X"0E",X"01",X"C3",X"6E",X"49",
		X"BC",X"A6",X"05",X"30",X"F1",X"7C",X"68",X"3B",X"A5",X"38",X"FD",X"F1",X"96",X"5D",X"17",X"9B",
		X"B9",X"3A",X"AE",X"A9",X"21",X"CA",X"A9",X"0F",X"0F",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",
		X"C0",X"EB",X"CD",X"F1",X"57",X"21",X"82",X"A9",X"34",X"EB",X"23",X"7E",X"C6",X"10",X"77",X"47",
		X"23",X"7E",X"90",X"D0",X"7E",X"4F",X"E6",X"F0",X"C6",X"10",X"2B",X"ED",X"44",X"86",X"77",X"18",
		X"2D",X"3A",X"AE",X"A9",X"21",X"C7",X"A9",X"0F",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",
		X"EB",X"CD",X"F1",X"57",X"21",X"81",X"A9",X"34",X"EB",X"23",X"7E",X"C6",X"10",X"77",X"47",X"23",
		X"7E",X"90",X"D0",X"7E",X"4F",X"E6",X"F0",X"C6",X"10",X"2B",X"ED",X"44",X"86",X"77",X"3A",X"C0",
		X"A9",X"A7",X"20",X"10",X"79",X"E6",X"0F",X"21",X"86",X"A9",X"86",X"27",X"77",X"30",X"02",X"36",
		X"99",X"CD",X"FB",X"4A",X"3A",X"81",X"A9",X"A7",X"C8",X"21",X"84",X"A9",X"7E",X"A7",X"20",X"07",
		X"36",X"30",X"3C",X"32",X"0A",X"C3",X"C9",X"35",X"28",X"09",X"7E",X"FE",X"18",X"C0",X"AF",X"32",
		X"0A",X"C3",X"C9",X"21",X"81",X"A9",X"35",X"C9",X"0F",X"4F",X"E6",X"07",X"32",X"C4",X"A9",X"79",
		X"0F",X"0F",X"0F",X"E6",X"01",X"32",X"C6",X"A9",X"32",X"00",X"C2",X"3A",X"3E",X"0C",X"32",X"02",
		X"C3",X"CD",X"B1",X"00",X"06",X"00",X"21",X"DE",X"27",X"AF",X"86",X"23",X"10",X"FC",X"D6",X"C5",
		X"C4",X"D8",X"00",X"C3",X"EB",X"32",X"3A",X"82",X"A9",X"A7",X"C8",X"21",X"85",X"A9",X"7E",X"A7",
		X"20",X"07",X"36",X"30",X"3C",X"32",X"0C",X"C3",X"C9",X"35",X"28",X"09",X"7E",X"FE",X"18",X"C0",
		X"AF",X"32",X"0C",X"C3",X"C9",X"21",X"82",X"A9",X"35",X"C9",X"EE",X"A6",X"14",X"A5",X"3B",X"87",
		X"F1",X"DC",X"D7",X"BF",X"F1",X"DC",X"C4",X"FD",X"ED",X"F1",X"7D",X"A5",X"38",X"34",X"B9",X"3A",
		X"13",X"32",X"32",X"F0",X"A9",X"3E",X"00",X"32",X"F1",X"A9",X"3E",X"FF",X"32",X"F2",X"A9",X"3E",
		X"04",X"32",X"F3",X"A9",X"3E",X"FF",X"32",X"F4",X"A9",X"3E",X"08",X"32",X"F6",X"A9",X"21",X"F1",
		X"56",X"22",X"F7",X"A9",X"06",X"0D",X"21",X"00",X"A4",X"0E",X"14",X"71",X"23",X"10",X"FC",X"3E",
		X"00",X"77",X"23",X"77",X"23",X"06",X"0D",X"71",X"23",X"10",X"FC",X"3E",X"0E",X"06",X"04",X"77",
		X"23",X"10",X"FC",X"21",X"B1",X"A7",X"CB",X"94",X"3A",X"0C",X"AD",X"4F",X"3E",X"A0",X"81",X"CD",
		X"19",X"13",X"21",X"D1",X"A5",X"CB",X"94",X"3E",X"20",X"81",X"CD",X"19",X"13",X"21",X"10",X"A6",
		X"CB",X"94",X"3E",X"A0",X"81",X"77",X"19",X"3E",X"20",X"81",X"77",X"21",X"12",X"A6",X"CB",X"94",
		X"3E",X"E0",X"81",X"77",X"19",X"3E",X"60",X"81",X"77",X"21",X"11",X"A6",X"CB",X"94",X"3E",X"A0",
		X"81",X"77",X"19",X"3E",X"20",X"81",X"77",X"CD",X"9C",X"33",X"C3",X"1A",X"0F",X"06",X"0D",X"2A",
		X"F7",X"A9",X"7E",X"A7",X"EB",X"28",X"09",X"7E",X"3C",X"CB",X"41",X"28",X"02",X"3D",X"3D",X"77",
		X"CB",X"49",X"11",X"20",X"00",X"28",X"03",X"11",X"E0",X"FF",X"19",X"EB",X"2A",X"F7",X"A9",X"23",
		X"CB",X"41",X"28",X"02",X"2B",X"2B",X"22",X"F7",X"A9",X"10",X"D7",X"C9",X"3A",X"B1",X"A9",X"E6",
		X"0F",X"FE",X"0F",X"20",X"05",X"21",X"C0",X"A9",X"36",X"FF",X"21",X"95",X"4B",X"CF",X"32",X"C9",
		X"A9",X"3A",X"B1",X"A9",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"FE",X"0F",X"20",X"05",X"21",X"C0",
		X"A9",X"36",X"FF",X"21",X"95",X"4B",X"CF",X"32",X"CC",X"A9",X"C9",X"0E",X"10",X"11",X"7F",X"A4",
		X"21",X"86",X"A9",X"CD",X"81",X"0D",X"C9",X"2A",X"41",X"AB",X"7D",X"AC",X"2F",X"87",X"87",X"ED",
		X"6A",X"22",X"41",X"AB",X"ED",X"5F",X"85",X"AC",X"C9",X"11",X"CC",X"0B",X"01",X"89",X"00",X"3A",
		X"50",X"1A",X"67",X"1A",X"81",X"4F",X"13",X"10",X"FA",X"94",X"C4",X"11",X"0F",X"C3",X"1A",X"0F",
		X"21",X"1B",X"0D",X"06",X"03",X"5E",X"23",X"56",X"23",X"1A",X"08",X"3E",X"04",X"82",X"57",X"1A",
		X"5E",X"23",X"56",X"23",X"12",X"1C",X"08",X"12",X"10",X"EB",X"C9",X"D9",X"21",X"3F",X"AB",X"11",
		X"40",X"AB",X"01",X"10",X"00",X"ED",X"B8",X"21",X"40",X"AB",X"3A",X"37",X"AB",X"AE",X"32",X"30",
		X"AB",X"21",X"80",X"A9",X"86",X"D9",X"C9",X"21",X"84",X"4B",X"11",X"30",X"AB",X"01",X"11",X"00",
		X"ED",X"B0",X"DD",X"2A",X"6D",X"08",X"2A",X"70",X"08",X"DD",X"7D",X"DD",X"84",X"85",X"C6",X"44",
		X"C2",X"00",X"60",X"C9",X"FF",X"05",X"F6",X"80",X"32",X"17",X"9C",X"C9",X"DD",X"21",X"74",X"98",
		X"FD",X"BF",X"24",X"AE",X"46",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"11",X"13",X"15",X"21",
		X"22",X"24",X"31",X"33",X"01",X"21",X"B1",X"4B",X"11",X"08",X"AB",X"01",X"28",X"00",X"ED",X"B0",
		X"C9",X"00",X"00",X"00",X"01",X"7C",X"11",X"68",X"F1",X"01",X"00",X"88",X"00",X"3B",X"11",X"A5",
		X"F1",X"02",X"60",X"84",X"00",X"38",X"11",X"FD",X"F1",X"03",X"20",X"65",X"00",X"68",X"11",X"68",
		X"F1",X"04",X"00",X"43",X"00",X"BF",X"11",X"A5",X"F1",X"C3",X"AE",X"08",X"21",X"08",X"AB",X"11",
		X"11",X"A7",X"0E",X"14",X"CD",X"1F",X"4C",X"21",X"10",X"AB",X"11",X"13",X"A7",X"0E",X"16",X"CD",
		X"1F",X"4C",X"21",X"18",X"AB",X"11",X"15",X"A7",X"0E",X"12",X"CD",X"1F",X"4C",X"21",X"20",X"AB",
		X"11",X"17",X"A7",X"0E",X"15",X"CD",X"1F",X"4C",X"21",X"28",X"AB",X"11",X"19",X"A7",X"0E",X"13",
		X"CD",X"1F",X"4C",X"C9",X"73",X"A6",X"14",X"7E",X"29",X"F8",X"96",X"5D",X"F3",X"13",X"B9",X"E5",
		X"7E",X"87",X"86",X"21",X"B4",X"4C",X"CF",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"23",X"E7",
		X"7E",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"23",X"E7",X"7E",X"12",X"CB",X"92",X"79",X"12",
		X"CB",X"D2",X"21",X"80",X"FF",X"19",X"EB",X"E1",X"23",X"23",X"23",X"CD",X"73",X"0D",X"E5",X"21",
		X"A0",X"FF",X"19",X"EB",X"E1",X"23",X"23",X"23",X"7E",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",
		X"23",X"E7",X"7E",X"12",X"CB",X"92",X"79",X"12",X"CB",X"D2",X"23",X"E7",X"7E",X"12",X"CB",X"92",
		X"79",X"12",X"CB",X"D2",X"C9",X"CD",X"D2",X"07",X"3A",X"32",X"AD",X"A7",X"21",X"10",X"AD",X"28",
		X"03",X"21",X"20",X"AD",X"11",X"00",X"AD",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"30",X"AD",X"A7",
		X"CA",X"1A",X"0F",X"3A",X"01",X"AD",X"16",X"06",X"5F",X"FF",X"3A",X"00",X"AD",X"3D",X"16",X"05",
		X"5F",X"FF",X"06",X"00",X"21",X"50",X"5B",X"97",X"AE",X"23",X"10",X"FC",X"C6",X"FF",X"32",X"08",
		X"C3",X"C3",X"1A",X"0F",X"96",X"ED",X"DC",X"9B",X"3B",X"87",X"CD",X"D7",X"87",X"F3",X"DC",X"C4",
		X"7F",X"DC",X"C4",X"21",X"0B",X"AB",X"06",X"05",X"3A",X"32",X"AD",X"A7",X"11",X"35",X"AD",X"28",
		X"03",X"11",X"38",X"AD",X"E5",X"D5",X"CD",X"2B",X"4D",X"30",X"09",X"D1",X"E1",X"3E",X"08",X"CF",
		X"10",X"F2",X"37",X"C9",X"05",X"28",X"3F",X"21",X"27",X"AB",X"11",X"2F",X"AB",X"78",X"87",X"87",
		X"87",X"4F",X"06",X"00",X"ED",X"B8",X"EB",X"2B",X"36",X"F1",X"2B",X"36",X"F1",X"2B",X"36",X"F1",
		X"22",X"91",X"A9",X"2B",X"D1",X"01",X"03",X"00",X"EB",X"ED",X"B8",X"1A",X"E1",X"21",X"31",X"A5",
		X"87",X"CF",X"22",X"93",X"A9",X"21",X"08",X"AB",X"11",X"08",X"00",X"06",X"05",X"AF",X"77",X"19",
		X"3C",X"10",X"FB",X"37",X"3F",X"C9",X"21",X"2F",X"AB",X"18",X"CC",X"0E",X"03",X"1A",X"BE",X"D8",
		X"20",X"05",X"1B",X"2B",X"0D",X"20",X"F6",X"37",X"3F",X"C9",X"21",X"05",X"AD",X"CD",X"67",X"4D",
		X"D8",X"2C",X"CD",X"67",X"4D",X"38",X"04",X"2C",X"CD",X"67",X"4D",X"21",X"D7",X"A9",X"7E",X"A7",
		X"C8",X"35",X"C0",X"3A",X"D6",X"A9",X"77",X"3A",X"C0",X"AC",X"3C",X"FE",X"10",X"38",X"02",X"3E",
		X"0F",X"32",X"C0",X"AC",X"C3",X"9A",X"1A",X"7E",X"C6",X"01",X"27",X"77",X"FE",X"60",X"D8",X"36",
		X"00",X"C9",X"4F",X"3A",X"30",X"AD",X"A7",X"C8",X"11",X"83",X"A7",X"79",X"FE",X"07",X"38",X"02",
		X"3E",X"06",X"A7",X"28",X"0C",X"06",X"09",X"0E",X"18",X"08",X"CD",X"AF",X"4D",X"08",X"3D",X"20",
		X"F8",X"01",X"10",X"F1",X"21",X"DD",X"59",X"19",X"30",X"05",X"CD",X"CF",X"4D",X"18",X"F5",X"06",
		X"00",X"21",X"11",X"07",X"97",X"AE",X"23",X"10",X"FC",X"C6",X"19",X"C2",X"B1",X"4B",X"C9",X"78",
		X"C6",X"03",X"12",X"3D",X"1B",X"12",X"E7",X"78",X"12",X"3C",X"13",X"12",X"21",X"00",X"FC",X"19",
		X"E7",X"71",X"2B",X"71",X"7D",X"C6",X"20",X"6F",X"30",X"01",X"24",X"71",X"23",X"71",X"C9",X"EB",
		X"70",X"2B",X"36",X"F1",X"CB",X"94",X"71",X"23",X"71",X"CB",X"D4",X"EB",X"E7",X"C9",X"3A",X"30",
		X"AD",X"A7",X"C8",X"3A",X"C3",X"A9",X"E6",X"01",X"21",X"1B",X"4E",X"28",X"03",X"21",X"30",X"4E",
		X"4E",X"06",X"00",X"23",X"3A",X"32",X"AD",X"A7",X"3A",X"35",X"AD",X"28",X"03",X"3A",X"38",X"AD",
		X"ED",X"B1",X"21",X"03",X"AD",X"20",X"11",X"CB",X"46",X"C0",X"CB",X"C6",X"21",X"00",X"AD",X"7E",
		X"34",X"16",X"05",X"5F",X"FF",X"C3",X"05",X"58",X"CB",X"86",X"C9",X"14",X"01",X"06",X"11",X"16",
		X"21",X"26",X"31",X"36",X"41",X"46",X"51",X"56",X"61",X"66",X"71",X"76",X"81",X"86",X"91",X"96",
		X"11",X"02",X"08",X"14",X"20",X"26",X"32",X"38",X"44",X"50",X"56",X"62",X"68",X"74",X"80",X"86",
		X"92",X"98",X"6F",X"A6",X"14",X"88",X"57",X"A5",X"BF",X"34",X"D7",X"F1",X"9B",X"F1",X"B9",X"3A",
		X"04",X"AD",X"FE",X"04",X"CA",X"2A",X"4F",X"3D",X"CA",X"BC",X"4E",X"3A",X"80",X"A9",X"E6",X"01",
		X"C2",X"35",X"4F",X"CD",X"5D",X"4F",X"06",X"04",X"11",X"10",X"A8",X"FD",X"21",X"12",X"AA",X"2E",
		X"05",X"26",X"0B",X"CD",X"85",X"51",X"3A",X"0D",X"AD",X"A7",X"20",X"1B",X"06",X"07",X"2E",X"07",
		X"26",X"0F",X"CD",X"52",X"51",X"06",X"03",X"2E",X"06",X"26",X"0D",X"CD",X"21",X"51",X"06",X"01",
		X"2E",X"08",X"26",X"11",X"C3",X"B3",X"51",X"06",X"05",X"2E",X"07",X"26",X"0F",X"CD",X"52",X"51",
		X"CD",X"B1",X"50",X"06",X"03",X"11",X"C0",X"A8",X"FD",X"21",X"28",X"AA",X"2E",X"06",X"26",X"0D",
		X"CD",X"21",X"51",X"06",X"01",X"2E",X"08",X"26",X"11",X"C3",X"B3",X"51",X"3A",X"80",X"A9",X"E6",
		X"01",X"C2",X"35",X"4F",X"CD",X"7E",X"4F",X"06",X"04",X"11",X"10",X"A8",X"FD",X"21",X"12",X"AA",
		X"2E",X"05",X"26",X"0B",X"CD",X"85",X"51",X"3A",X"0D",X"AD",X"A7",X"20",X"25",X"06",X"07",X"2E",
		X"07",X"26",X"0F",X"CD",X"52",X"51",X"CD",X"7E",X"50",X"06",X"01",X"11",X"E0",X"A8",X"FD",X"21",
		X"2C",X"AA",X"2E",X"05",X"26",X"0B",X"CD",X"85",X"51",X"06",X"01",X"2E",X"08",X"26",X"11",X"C3",
		X"B3",X"51",X"06",X"05",X"2E",X"07",X"26",X"0F",X"CD",X"52",X"51",X"CD",X"B1",X"50",X"CD",X"7E",
		X"50",X"06",X"01",X"11",X"E0",X"A8",X"FD",X"21",X"2C",X"AA",X"2E",X"05",X"26",X"0B",X"CD",X"85",
		X"51",X"06",X"01",X"2E",X"08",X"26",X"11",X"C3",X"B3",X"51",X"3A",X"80",X"A9",X"E6",X"01",X"CA",
		X"63",X"4E",X"C3",X"32",X"50",X"3A",X"0D",X"AD",X"A7",X"C2",X"BF",X"4F",X"11",X"50",X"A8",X"FD",
		X"21",X"1A",X"AA",X"DD",X"21",X"80",X"AA",X"08",X"3E",X"07",X"47",X"08",X"0E",X"06",X"ED",X"53",
		X"93",X"A9",X"FD",X"22",X"91",X"A9",X"2E",X"07",X"26",X"0F",X"C3",X"11",X"52",X"11",X"C0",X"A8",
		X"FD",X"21",X"28",X"AA",X"DD",X"21",X"80",X"AA",X"08",X"3E",X"03",X"47",X"08",X"0E",X"06",X"ED",
		X"53",X"93",X"A9",X"FD",X"22",X"91",X"A9",X"2E",X"07",X"26",X"0F",X"C3",X"11",X"52",X"2E",X"06",
		X"26",X"0D",X"1E",X"17",X"16",X"1F",X"FD",X"21",X"80",X"AA",X"06",X"06",X"3A",X"C0",X"A8",X"3C",
		X"C0",X"FD",X"7E",X"00",X"3C",X"20",X"1F",X"3A",X"28",X"AA",X"FD",X"96",X"06",X"85",X"BC",X"30",
		X"15",X"3A",X"59",X"AA",X"FD",X"96",X"04",X"83",X"BA",X"30",X"0B",X"3E",X"F0",X"32",X"C0",X"A8",
		X"FD",X"77",X"00",X"CD",X"DE",X"51",X"FD",X"7D",X"C6",X"10",X"FD",X"6F",X"10",X"D3",X"C9",X"11",
		X"50",X"A8",X"FD",X"21",X"1A",X"AA",X"DD",X"21",X"80",X"AA",X"08",X"3E",X"05",X"47",X"08",X"0E",
		X"06",X"ED",X"53",X"93",X"A9",X"FD",X"22",X"91",X"A9",X"2E",X"07",X"26",X"0F",X"CD",X"11",X"52",
		X"3A",X"04",X"AD",X"A7",X"28",X"45",X"FE",X"04",X"28",X"41",X"2E",X"06",X"26",X"0D",X"1E",X"17",
		X"16",X"1F",X"FD",X"21",X"80",X"AA",X"06",X"06",X"3A",X"A0",X"A8",X"3C",X"C0",X"FD",X"7E",X"00",
		X"3C",X"20",X"1F",X"3A",X"24",X"AA",X"FD",X"96",X"06",X"85",X"BC",X"30",X"15",X"3A",X"55",X"AA",
		X"FD",X"96",X"04",X"83",X"BA",X"30",X"0B",X"3E",X"F0",X"32",X"A0",X"A8",X"FD",X"77",X"00",X"CD",
		X"DE",X"51",X"FD",X"7D",X"C6",X"10",X"FD",X"6F",X"10",X"D3",X"C9",X"2E",X"08",X"26",X"11",X"C3",
		X"EE",X"4F",X"3A",X"0D",X"AD",X"A7",X"C2",X"5A",X"50",X"11",X"10",X"A8",X"FD",X"21",X"12",X"AA",
		X"DD",X"21",X"80",X"AA",X"08",X"3E",X"0B",X"47",X"08",X"0E",X"06",X"ED",X"53",X"93",X"A9",X"FD",
		X"22",X"91",X"A9",X"2E",X"07",X"26",X"0F",X"C3",X"11",X"52",X"11",X"10",X"A8",X"FD",X"21",X"12",
		X"AA",X"DD",X"21",X"80",X"AA",X"08",X"3E",X"09",X"47",X"08",X"0E",X"06",X"ED",X"53",X"93",X"A9",
		X"FD",X"22",X"91",X"A9",X"2E",X"07",X"26",X"0F",X"CD",X"11",X"52",X"C3",X"E0",X"4F",X"DD",X"21",
		X"10",X"AA",X"3A",X"00",X"A8",X"3C",X"C0",X"3A",X"C0",X"A8",X"3C",X"C0",X"3A",X"28",X"AA",X"DD",
		X"96",X"00",X"C6",X"06",X"FE",X"0D",X"D0",X"3A",X"59",X"AA",X"DD",X"96",X"31",X"C6",X"18",X"FE",
		X"21",X"D0",X"3E",X"F0",X"32",X"00",X"A8",X"32",X"C0",X"A8",X"AF",X"32",X"DC",X"A8",X"C3",X"DE",
		X"51",X"3A",X"04",X"AD",X"A7",X"28",X"37",X"FE",X"04",X"28",X"33",X"DD",X"21",X"10",X"AA",X"3A",
		X"00",X"A8",X"3C",X"C0",X"3A",X"A0",X"A8",X"3C",X"C0",X"3A",X"24",X"AA",X"DD",X"96",X"00",X"C6",
		X"06",X"FE",X"0D",X"D0",X"3A",X"55",X"AA",X"DD",X"96",X"31",X"C6",X"19",X"FE",X"23",X"D0",X"3E",
		X"F0",X"32",X"00",X"A8",X"32",X"A0",X"A8",X"AF",X"32",X"A4",X"A8",X"C3",X"DE",X"51",X"DD",X"21",
		X"10",X"AA",X"3A",X"00",X"A8",X"3C",X"C0",X"3A",X"A0",X"A8",X"3C",X"C0",X"3A",X"24",X"AA",X"DD",
		X"96",X"00",X"C6",X"08",X"FE",X"11",X"D0",X"3A",X"55",X"AA",X"DD",X"96",X"31",X"C6",X"19",X"FE",
		X"23",X"D0",X"3E",X"F0",X"32",X"00",X"A8",X"32",X"A0",X"A8",X"AF",X"32",X"A4",X"A8",X"C3",X"DE",
		X"51",X"3A",X"00",X"A8",X"3C",X"C0",X"1A",X"3C",X"20",X"1D",X"3A",X"10",X"AA",X"FD",X"96",X"00",
		X"85",X"BC",X"30",X"13",X"3A",X"41",X"AA",X"FD",X"96",X"31",X"85",X"BC",X"30",X"09",X"3E",X"F0",
		X"32",X"00",X"A8",X"12",X"CD",X"DE",X"51",X"7B",X"C6",X"10",X"5F",X"FD",X"23",X"FD",X"23",X"10",
		X"D5",X"C9",X"3A",X"00",X"A8",X"3C",X"C0",X"1A",X"3C",X"20",X"1F",X"3A",X"10",X"AA",X"FD",X"96",
		X"00",X"85",X"BC",X"30",X"15",X"3A",X"41",X"AA",X"FD",X"96",X"31",X"C6",X"08",X"FE",X"11",X"30",
		X"09",X"3E",X"F0",X"32",X"00",X"A8",X"12",X"CD",X"DE",X"51",X"7B",X"C6",X"10",X"5F",X"FD",X"23",
		X"FD",X"23",X"10",X"D3",X"C9",X"3A",X"00",X"A8",X"3C",X"C0",X"1A",X"3C",X"20",X"1A",X"3A",X"10",
		X"AA",X"FD",X"96",X"00",X"85",X"BC",X"30",X"10",X"3A",X"41",X"AA",X"FD",X"96",X"31",X"85",X"BC",
		X"30",X"06",X"3E",X"F0",X"32",X"00",X"A8",X"12",X"7B",X"C6",X"10",X"5F",X"FD",X"23",X"FD",X"23",
		X"10",X"D8",X"C9",X"3A",X"00",X"A8",X"3C",X"C0",X"1A",X"3C",X"20",X"17",X"3A",X"10",X"AA",X"FD",
		X"96",X"00",X"85",X"BC",X"30",X"0D",X"3A",X"41",X"AA",X"FD",X"96",X"31",X"85",X"BC",X"30",X"03",
		X"3E",X"F0",X"12",X"7B",X"C6",X"10",X"5F",X"FD",X"23",X"FD",X"23",X"10",X"DB",X"C9",X"D5",X"3A",
		X"9D",X"A9",X"A7",X"28",X"15",X"3A",X"9E",X"A9",X"3C",X"32",X"9E",X"A9",X"E6",X"07",X"3C",X"5F",
		X"16",X"04",X"FF",X"D1",X"3E",X"1E",X"32",X"9D",X"A9",X"C9",X"11",X"01",X"04",X"FF",X"D1",X"3E",
		X"1E",X"32",X"9D",X"A9",X"C9",X"21",X"9D",X"A9",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"2C",X"77",
		X"C9",X"DD",X"7E",X"00",X"3C",X"20",X"3D",X"1A",X"3C",X"20",X"2F",X"FD",X"7E",X"00",X"C6",X"08",
		X"FE",X"19",X"38",X"26",X"FD",X"7E",X"31",X"C6",X"10",X"FE",X"11",X"38",X"1D",X"DD",X"7E",X"06",
		X"FD",X"96",X"00",X"85",X"BC",X"30",X"13",X"DD",X"7E",X"04",X"FD",X"96",X"31",X"85",X"BC",X"30",
		X"09",X"3E",X"F0",X"DD",X"77",X"00",X"12",X"CD",X"DE",X"51",X"7B",X"C6",X"10",X"5F",X"FD",X"23",
		X"FD",X"23",X"10",X"C3",X"FD",X"2A",X"91",X"A9",X"ED",X"5B",X"93",X"A9",X"08",X"47",X"08",X"DD",
		X"7D",X"C6",X"10",X"DD",X"6F",X"0D",X"C2",X"11",X"52",X"C9",X"21",X"84",X"AE",X"22",X"80",X"AE",
		X"21",X"04",X"AE",X"22",X"00",X"AE",X"C9",X"06",X"00",X"21",X"DE",X"27",X"AF",X"86",X"23",X"10",
		X"FC",X"D6",X"C5",X"C4",X"D4",X"53",X"CD",X"0E",X"53",X"CD",X"D2",X"52",X"3A",X"00",X"AE",X"FE",
		X"04",X"28",X"D7",X"4F",X"06",X"00",X"21",X"00",X"AE",X"11",X"80",X"AE",X"ED",X"B0",X"C6",X"80",
		X"32",X"80",X"AE",X"21",X"04",X"AE",X"22",X"00",X"AE",X"C9",X"3A",X"C9",X"08",X"32",X"8D",X"A9",
		X"3A",X"74",X"08",X"32",X"CD",X"A9",X"3A",X"60",X"C3",X"2F",X"32",X"B1",X"A9",X"CD",X"CC",X"4A",
		X"3A",X"00",X"C2",X"2F",X"4F",X"E6",X"03",X"C6",X"03",X"FE",X"06",X"20",X"02",X"3E",X"FF",X"C3",
		X"19",X"2E",X"3A",X"0C",X"AD",X"E6",X"0F",X"4F",X"2A",X"00",X"AE",X"7D",X"D6",X"04",X"C8",X"0F",
		X"0F",X"E6",X"1F",X"47",X"21",X"04",X"AE",X"5E",X"2C",X"56",X"2C",X"1A",X"E6",X"10",X"20",X"0E",
		X"7E",X"CB",X"D2",X"12",X"CB",X"92",X"2C",X"7E",X"2C",X"81",X"12",X"10",X"EA",X"C9",X"2C",X"2C",
		X"10",X"E5",X"C9",X"CD",X"0C",X"20",X"FE",X"67",X"C2",X"8D",X"0F",X"C3",X"1A",X"0F",X"2A",X"80",
		X"AE",X"7D",X"E6",X"7F",X"D6",X"04",X"C8",X"0F",X"0F",X"E6",X"1F",X"47",X"21",X"84",X"AE",X"5E",
		X"2C",X"56",X"2C",X"1A",X"E6",X"10",X"20",X"0A",X"2C",X"2C",X"CB",X"D2",X"3E",X"20",X"12",X"10",
		X"EE",X"C9",X"2C",X"2C",X"10",X"E9",X"C9",X"DD",X"7E",X"04",X"C6",X"07",X"47",X"16",X"28",X"07",
		X"CB",X"12",X"07",X"CB",X"12",X"E6",X"E0",X"5F",X"DD",X"7E",X"06",X"C6",X"07",X"4F",X"0F",X"0F",
		X"0F",X"E6",X"1F",X"83",X"5F",X"79",X"07",X"07",X"07",X"E6",X"38",X"4F",X"78",X"06",X"00",X"CB",
		X"57",X"28",X"01",X"04",X"0F",X"0F",X"E6",X"C0",X"81",X"4F",X"21",X"D4",X"53",X"09",X"7E",X"23",
		X"46",X"23",X"A7",X"28",X"10",X"E5",X"2A",X"00",X"AE",X"73",X"2C",X"72",X"2C",X"77",X"2C",X"70",
		X"2C",X"22",X"00",X"AE",X"E1",X"13",X"7E",X"23",X"46",X"23",X"A7",X"28",X"10",X"E5",X"2A",X"00",
		X"AE",X"73",X"2C",X"72",X"2C",X"77",X"2C",X"70",X"2C",X"22",X"00",X"AE",X"E1",X"7B",X"C6",X"1F",
		X"5F",X"30",X"01",X"14",X"7E",X"23",X"46",X"23",X"A7",X"28",X"10",X"E5",X"2A",X"00",X"AE",X"73",
		X"2C",X"72",X"2C",X"77",X"2C",X"70",X"2C",X"22",X"00",X"AE",X"E1",X"13",X"7E",X"23",X"46",X"23",
		X"A7",X"28",X"10",X"E5",X"2A",X"00",X"AE",X"73",X"2C",X"72",X"2C",X"77",X"2C",X"70",X"2C",X"22",
		X"00",X"AE",X"E1",X"C9",X"24",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"24",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"20",X"39",X"60",
		X"00",X"00",X"00",X"00",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B7",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B7",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"20",X"6D",X"60",
		X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2B",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"B1",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2B",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"20",X"8E",X"60",
		X"00",X"00",X"00",X"00",X"74",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4C",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"74",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"D5",X"20",X"D5",X"60",
		X"00",X"00",X"00",X"00",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2B",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"B1",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2B",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"A0",X"8E",X"E0",
		X"00",X"00",X"00",X"00",X"30",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B7",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B7",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"A0",X"6D",X"E0",
		X"00",X"00",X"00",X"00",X"24",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"24",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"A0",X"39",X"E0",
		X"00",X"00",X"00",X"00",X"3A",X"20",X"00",X"00",X"3A",X"A0",X"00",X"00",X"8F",X"20",X"00",X"00",
		X"8F",X"A0",X"00",X"00",X"70",X"20",X"00",X"00",X"70",X"A0",X"00",X"00",X"66",X"20",X"00",X"00",
		X"66",X"A0",X"00",X"00",X"70",X"60",X"00",X"00",X"70",X"E0",X"00",X"00",X"8F",X"60",X"00",X"00",
		X"8F",X"E0",X"00",X"00",X"3A",X"60",X"00",X"00",X"3A",X"E0",X"00",X"00",X"C7",X"20",X"C7",X"60",
		X"C7",X"A0",X"C7",X"E0",X"21",X"43",X"AC",X"7E",X"A7",X"C8",X"35",X"F5",X"23",X"7E",X"CD",X"F8",
		X"55",X"F1",X"C8",X"3D",X"06",X"00",X"4F",X"5D",X"54",X"23",X"ED",X"B0",X"C9",X"73",X"A6",X"14",
		X"7E",X"29",X"F8",X"96",X"5D",X"17",X"9B",X"B9",X"32",X"00",X"C0",X"3E",X"01",X"32",X"04",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"32",X"04",X"C3",X"C9",X"E5",X"F5",X"3A",X"30",
		X"AD",X"A7",X"20",X"16",X"F1",X"E1",X"C9",X"E5",X"F5",X"3A",X"30",X"AD",X"A7",X"20",X"0B",X"3A",
		X"C6",X"A9",X"A7",X"20",X"05",X"F1",X"E1",X"C9",X"E5",X"F5",X"21",X"43",X"AC",X"34",X"7E",X"CF",
		X"F1",X"77",X"E1",X"C9",X"3A",X"7C",X"16",X"CD",X"28",X"56",X"3A",X"9C",X"0A",X"CD",X"28",X"56",
		X"3A",X"84",X"14",X"CD",X"28",X"56",X"3A",X"78",X"0C",X"CD",X"28",X"56",X"3A",X"D3",X"07",X"CD",
		X"28",X"56",X"3A",X"B4",X"33",X"CD",X"28",X"56",X"3A",X"04",X"AD",X"C6",X"8C",X"18",X"C9",X"3A",
		X"A2",X"07",X"18",X"A8",X"3A",X"DE",X"16",X"18",X"A3",X"3A",X"9F",X"4C",X"18",X"9E",X"3A",X"D8",
		X"07",X"CD",X"0C",X"56",X"3A",X"6B",X"27",X"18",X"93",X"3A",X"FE",X"07",X"18",X"8E",X"3A",X"70",
		X"32",X"18",X"94",X"3A",X"A6",X"07",X"CD",X"17",X"56",X"3A",X"DA",X"4C",X"18",X"89",X"3A",X"87",
		X"2D",X"C3",X"0C",X"56",X"0E",X"00",X"21",X"31",X"08",X"3A",X"AB",X"A9",X"96",X"23",X"0D",X"20",
		X"FB",X"EE",X"C2",X"32",X"AB",X"A9",X"CD",X"97",X"0F",X"CD",X"DF",X"1E",X"CD",X"97",X"0F",X"CD",
		X"BC",X"2C",X"CD",X"E3",X"23",X"CD",X"98",X"10",X"21",X"EB",X"A9",X"35",X"C0",X"0E",X"00",X"21",
		X"A7",X"12",X"3A",X"AB",X"A9",X"96",X"23",X"0D",X"20",X"FB",X"EE",X"59",X"32",X"AB",X"A9",X"C3",
		X"1A",X"0F",X"3A",X"5B",X"0C",X"CD",X"0C",X"56",X"3A",X"55",X"08",X"CD",X"0C",X"56",X"3A",X"75",
		X"16",X"CD",X"0C",X"56",X"3A",X"CB",X"27",X"CD",X"17",X"56",X"3A",X"A0",X"33",X"C3",X"17",X"56",
		X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3A",X"2E",X"32",X"C3",X"28",X"56",X"3A",X"04",X"AD",X"C6",X"0C",X"C3",X"0C",X"56",X"3A",
		X"9B",X"07",X"C3",X"0C",X"56",X"3A",X"4E",X"2D",X"C3",X"0C",X"56",X"3A",X"EE",X"49",X"C3",X"0C",
		X"56",X"3A",X"A9",X"07",X"C3",X"0C",X"56",X"3A",X"3A",X"27",X"C3",X"0C",X"56",X"0C",X"A7",X"13",
		X"88",X"57",X"34",X"A5",X"ED",X"34",X"F1",X"87",X"34",X"88",X"68",X"ED",X"FD",X"DC",X"F1",X"77",
		X"68",X"FD",X"3B",X"B9",X"3A",X"67",X"17",X"C3",X"0C",X"56",X"3A",X"FA",X"18",X"C3",X"0C",X"56",
		X"21",X"D7",X"59",X"C3",X"BC",X"58",X"21",X"00",X"5C",X"C3",X"BC",X"58",X"60",X"A7",X"14",X"96",
		X"10",X"0D",X"88",X"B9",X"21",X"00",X"5E",X"C3",X"BC",X"58",X"21",X"30",X"25",X"C3",X"BC",X"58",
		X"21",X"3E",X"2E",X"C3",X"BC",X"58",X"2A",X"81",X"25",X"01",X"00",X"04",X"16",X"10",X"72",X"23",
		X"0B",X"79",X"B0",X"20",X"F9",X"32",X"00",X"C2",X"2A",X"37",X"4A",X"01",X"00",X"04",X"16",X"F1",
		X"72",X"23",X"0B",X"79",X"B0",X"20",X"F9",X"21",X"00",X"00",X"3A",X"00",X"00",X"86",X"23",X"08",
		X"7C",X"FE",X"60",X"30",X"06",X"08",X"32",X"00",X"C2",X"18",X"F2",X"08",X"D6",X"AF",X"C2",X"D7",
		X"59",X"C3",X"11",X"25",X"21",X"FA",X"08",X"C3",X"BC",X"58",X"21",X"D7",X"59",X"C3",X"FE",X"58",
		X"21",X"00",X"5C",X"C3",X"FE",X"58",X"21",X"00",X"5E",X"C3",X"FE",X"58",X"DD",X"7E",X"02",X"4F",
		X"87",X"30",X"01",X"24",X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"79",X"C6",X"C0",X"01",
		X"80",X"01",X"30",X"03",X"01",X"80",X"FF",X"09",X"46",X"2B",X"4E",X"2A",X"08",X"A8",X"19",X"DD",
		X"5E",X"03",X"FD",X"56",X"31",X"19",X"DD",X"75",X"03",X"FD",X"74",X"31",X"2A",X"0A",X"A8",X"09",
		X"DD",X"5E",X"05",X"FD",X"56",X"00",X"19",X"DD",X"75",X"05",X"FD",X"74",X"00",X"C9",X"DD",X"7E",
		X"02",X"4F",X"87",X"30",X"01",X"24",X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"79",X"C6",
		X"C0",X"01",X"80",X"01",X"30",X"03",X"01",X"80",X"FF",X"09",X"46",X"2B",X"4E",X"2A",X"08",X"A8",
		X"19",X"19",X"DD",X"5E",X"03",X"FD",X"56",X"31",X"19",X"DD",X"75",X"03",X"FD",X"74",X"31",X"2A",
		X"0A",X"A8",X"09",X"09",X"DD",X"5E",X"05",X"FD",X"56",X"00",X"19",X"DD",X"75",X"05",X"FD",X"74",
		X"00",X"C9",X"21",X"D7",X"59",X"C3",X"6E",X"59",X"21",X"00",X"5C",X"C3",X"6E",X"59",X"21",X"00",
		X"5E",X"C3",X"6E",X"59",X"73",X"A6",X"14",X"7E",X"29",X"F8",X"96",X"5D",X"02",X"13",X"B9",X"21",
		X"30",X"25",X"C3",X"6E",X"59",X"21",X"3E",X"2E",X"C3",X"6E",X"59",X"21",X"FA",X"08",X"DD",X"7E",
		X"02",X"4F",X"87",X"30",X"01",X"24",X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"79",X"C6",
		X"C0",X"01",X"80",X"01",X"30",X"03",X"01",X"80",X"FF",X"09",X"46",X"2B",X"4E",X"C9",X"21",X"D7",
		X"59",X"C3",X"9D",X"59",X"21",X"00",X"5C",X"C3",X"9D",X"59",X"21",X"00",X"5E",X"DD",X"7E",X"02",
		X"4F",X"87",X"30",X"01",X"24",X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"CB",X"23",X"CB",
		X"12",X"79",X"C6",X"C0",X"01",X"80",X"01",X"30",X"03",X"01",X"80",X"FF",X"09",X"46",X"2B",X"4E",
		X"CB",X"21",X"CB",X"10",X"C9",X"21",X"D7",X"59",X"C3",X"A0",X"59",X"21",X"00",X"5C",X"C3",X"A0",
		X"59",X"21",X"00",X"5E",X"C3",X"A0",X"59",X"CE",X"00",X"CD",X"00",X"CC",X"00",X"CB",X"00",X"CA",
		X"00",X"C9",X"00",X"C8",X"00",X"C8",X"00",X"C6",X"00",X"C4",X"00",X"C2",X"00",X"C0",X"00",X"BF",
		X"00",X"BC",X"00",X"BA",X"00",X"B9",X"00",X"B6",X"00",X"B3",X"00",X"B0",X"00",X"AF",X"00",X"AC",
		X"00",X"A9",X"00",X"A8",X"00",X"A5",X"00",X"A2",X"00",X"A1",X"00",X"9E",X"00",X"9B",X"00",X"98",
		X"00",X"97",X"00",X"94",X"00",X"91",X"00",X"90",X"00",X"8D",X"00",X"89",X"00",X"88",X"00",X"85",
		X"00",X"81",X"00",X"7F",X"00",X"7B",X"00",X"78",X"00",X"76",X"00",X"70",X"00",X"6D",X"00",X"68",
		X"00",X"63",X"00",X"60",X"00",X"5C",X"00",X"58",X"00",X"52",X"00",X"4E",X"00",X"49",X"00",X"43",
		X"00",X"3E",X"00",X"39",X"00",X"32",X"00",X"2C",X"00",X"27",X"00",X"20",X"00",X"1A",X"00",X"14",
		X"00",X"0E",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"F8",X"FF",X"F2",X"FF",X"00",X"00",X"E6",
		X"FF",X"E0",X"FF",X"D9",X"FF",X"D4",X"FF",X"CE",X"FF",X"C7",X"FF",X"C2",X"FF",X"BD",X"FF",X"B7",
		X"FF",X"B2",X"FF",X"AE",X"FF",X"A8",X"FF",X"A4",X"FF",X"A0",X"FF",X"9D",X"FF",X"A0",X"FF",X"93",
		X"FF",X"90",X"FF",X"8A",X"FF",X"88",X"FF",X"85",X"FF",X"81",X"FF",X"7F",X"FF",X"7B",X"FF",X"78",
		X"FF",X"77",X"FF",X"73",X"FF",X"70",X"FF",X"6F",X"FF",X"6C",X"FF",X"69",X"FF",X"69",X"FF",X"65",
		X"FF",X"62",X"FF",X"5F",X"FF",X"5E",X"FF",X"5B",X"FF",X"58",X"FF",X"57",X"FF",X"54",X"FF",X"51",
		X"FF",X"50",X"FF",X"4D",X"FF",X"4A",X"FF",X"47",X"FF",X"46",X"FF",X"44",X"FF",X"41",X"FF",X"40",
		X"FF",X"3E",X"FF",X"3C",X"FF",X"3A",X"FF",X"38",X"FF",X"38",X"FF",X"37",X"FF",X"36",X"FF",X"35",
		X"FF",X"34",X"FF",X"33",X"FF",X"32",X"FF",X"32",X"FF",X"33",X"FF",X"34",X"FF",X"35",X"FF",X"36",
		X"FF",X"37",X"FF",X"38",X"FF",X"38",X"FF",X"3A",X"FF",X"3C",X"FF",X"3E",X"FF",X"40",X"FF",X"41",
		X"FF",X"44",X"FF",X"46",X"FF",X"47",X"FF",X"4A",X"FF",X"4D",X"FF",X"50",X"FF",X"51",X"FF",X"54",
		X"FF",X"57",X"FF",X"58",X"FF",X"5B",X"FF",X"5E",X"FF",X"5F",X"FF",X"62",X"FF",X"65",X"FF",X"68",
		X"FF",X"69",X"FF",X"6C",X"FF",X"6F",X"FF",X"70",X"FF",X"73",X"FF",X"77",X"FF",X"78",X"FF",X"7B",
		X"FF",X"7F",X"FF",X"81",X"FF",X"85",X"FF",X"88",X"FF",X"8A",X"FF",X"90",X"FF",X"93",X"FF",X"98",
		X"FF",X"9D",X"FF",X"A0",X"FF",X"A4",X"FF",X"A8",X"FF",X"AE",X"FF",X"B2",X"FF",X"B7",X"FF",X"BD",
		X"FF",X"C2",X"FF",X"C7",X"FF",X"CE",X"FF",X"D4",X"FF",X"D9",X"FF",X"E0",X"FF",X"E6",X"FF",X"EC",
		X"FF",X"F2",X"FF",X"F8",X"FF",X"00",X"00",X"00",X"00",X"08",X"00",X"0E",X"00",X"14",X"00",X"1A",
		X"00",X"20",X"00",X"27",X"00",X"2C",X"00",X"32",X"00",X"39",X"00",X"3E",X"00",X"43",X"00",X"49",
		X"00",X"4E",X"00",X"52",X"00",X"58",X"00",X"5C",X"00",X"60",X"00",X"63",X"00",X"63",X"00",X"6D",
		X"00",X"70",X"00",X"76",X"00",X"78",X"00",X"7B",X"00",X"7F",X"00",X"81",X"00",X"85",X"00",X"88",
		X"00",X"89",X"00",X"8D",X"00",X"90",X"00",X"91",X"00",X"94",X"00",X"97",X"00",X"94",X"00",X"9B",
		X"00",X"9E",X"00",X"A1",X"00",X"A2",X"00",X"A5",X"00",X"A8",X"00",X"A9",X"00",X"AC",X"00",X"AF",
		X"00",X"B0",X"00",X"B3",X"00",X"B6",X"00",X"B9",X"00",X"BA",X"00",X"BC",X"00",X"B9",X"00",X"C0",
		X"00",X"C2",X"00",X"C4",X"00",X"C6",X"00",X"C8",X"00",X"C8",X"00",X"C9",X"00",X"CA",X"00",X"CB",
		X"00",X"CC",X"00",X"CD",X"00",X"CE",X"00",X"CD",X"D2",X"07",X"CD",X"01",X"02",X"C0",X"21",X"DD",
		X"0B",X"97",X"47",X"AE",X"23",X"10",X"FC",X"C6",X"E4",X"C4",X"11",X"0F",X"3A",X"AB",X"A9",X"21",
		X"34",X"17",X"06",X"14",X"86",X"23",X"10",X"FC",X"C6",X"77",X"32",X"AB",X"A9",X"C3",X"1A",X"0F",
		X"E7",X"00",X"E6",X"00",X"E5",X"00",X"E4",X"00",X"E3",X"00",X"E2",X"00",X"E1",X"00",X"E0",X"00",
		X"DE",X"00",X"DC",X"00",X"DA",X"00",X"D8",X"00",X"D6",X"00",X"D3",X"00",X"D1",X"00",X"CF",X"00",
		X"CC",X"00",X"C9",X"00",X"C6",X"00",X"C4",X"00",X"C1",X"00",X"BE",X"00",X"BC",X"00",X"B9",X"00",
		X"B6",X"00",X"B4",X"00",X"B1",X"00",X"AE",X"00",X"AB",X"00",X"A9",X"00",X"A6",X"00",X"A3",X"00",
		X"A1",X"00",X"9E",X"00",X"9A",X"00",X"98",X"00",X"95",X"00",X"91",X"00",X"8E",X"00",X"8A",X"00",
		X"87",X"00",X"84",X"00",X"7E",X"00",X"7A",X"00",X"75",X"00",X"6F",X"00",X"6C",X"00",X"67",X"00",
		X"62",X"00",X"5C",X"00",X"57",X"00",X"51",X"00",X"4B",X"00",X"45",X"00",X"3F",X"00",X"38",X"00",
		X"31",X"00",X"2B",X"00",X"24",X"00",X"1D",X"00",X"16",X"00",X"0F",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"FF",X"F1",X"FF",X"00",X"00",X"E3",X"FF",X"DC",X"FF",X"D5",X"FF",X"CF",X"FF",
		X"C8",X"FF",X"C1",X"FF",X"BB",X"FF",X"B5",X"FF",X"AF",X"FF",X"A9",X"FF",X"A4",X"FF",X"9E",X"FF",
		X"99",X"FF",X"94",X"FF",X"91",X"FF",X"94",X"FF",X"86",X"FF",X"82",X"FF",X"7C",X"FF",X"79",X"FF",
		X"76",X"FF",X"72",X"FF",X"6F",X"FF",X"6B",X"FF",X"68",X"FF",X"66",X"FF",X"62",X"FF",X"5F",X"FF",
		X"5D",X"FF",X"5A",X"FF",X"57",X"FF",X"57",X"FF",X"52",X"FF",X"4F",X"FF",X"4C",X"FF",X"4A",X"FF",
		X"47",X"FF",X"44",X"FF",X"42",X"FF",X"3F",X"FF",X"3C",X"FF",X"3A",X"FF",X"37",X"FF",X"34",X"FF",
		X"31",X"FF",X"2F",X"FF",X"2D",X"FF",X"2A",X"FF",X"28",X"FF",X"26",X"FF",X"24",X"FF",X"22",X"FF",
		X"20",X"FF",X"1F",X"FF",X"1E",X"FF",X"1D",X"FF",X"1C",X"FF",X"1B",X"FF",X"1A",X"FF",X"19",X"FF",
		X"19",X"FF",X"1A",X"FF",X"1B",X"FF",X"1C",X"FF",X"1D",X"FF",X"1E",X"FF",X"1F",X"FF",X"20",X"FF",
		X"22",X"FF",X"24",X"FF",X"26",X"FF",X"28",X"FF",X"2A",X"FF",X"2D",X"FF",X"2F",X"FF",X"31",X"FF",
		X"34",X"FF",X"37",X"FF",X"3A",X"FF",X"3C",X"FF",X"3F",X"FF",X"42",X"FF",X"44",X"FF",X"47",X"FF",
		X"4A",X"FF",X"4C",X"FF",X"4F",X"FF",X"52",X"FF",X"55",X"FF",X"57",X"FF",X"5A",X"FF",X"5D",X"FF",
		X"5F",X"FF",X"62",X"FF",X"66",X"FF",X"68",X"FF",X"6B",X"FF",X"6F",X"FF",X"72",X"FF",X"76",X"FF",
		X"79",X"FF",X"7C",X"FF",X"82",X"FF",X"86",X"FF",X"8B",X"FF",X"91",X"FF",X"94",X"FF",X"99",X"FF",
		X"9E",X"FF",X"A4",X"FF",X"A9",X"FF",X"AF",X"FF",X"B5",X"FF",X"BB",X"FF",X"C1",X"FF",X"C8",X"FF",
		X"CF",X"FF",X"D5",X"FF",X"DC",X"FF",X"E3",X"FF",X"EA",X"FF",X"F1",X"FF",X"F8",X"FF",X"00",X"00",
		X"00",X"00",X"08",X"00",X"0F",X"00",X"16",X"00",X"1D",X"00",X"24",X"00",X"2B",X"00",X"31",X"00",
		X"38",X"00",X"3F",X"00",X"45",X"00",X"4B",X"00",X"51",X"00",X"57",X"00",X"5C",X"00",X"62",X"00",
		X"67",X"00",X"6C",X"00",X"6F",X"00",X"6F",X"00",X"7A",X"00",X"7E",X"00",X"84",X"00",X"87",X"00",
		X"8A",X"00",X"8E",X"00",X"91",X"00",X"95",X"00",X"98",X"00",X"9A",X"00",X"9E",X"00",X"A1",X"00",
		X"A3",X"00",X"A6",X"00",X"A9",X"00",X"A6",X"00",X"AE",X"00",X"B1",X"00",X"B4",X"00",X"B6",X"00",
		X"B9",X"00",X"BC",X"00",X"BE",X"00",X"C1",X"00",X"C4",X"00",X"C6",X"00",X"C9",X"00",X"CC",X"00",
		X"CF",X"00",X"D1",X"00",X"D3",X"00",X"CF",X"00",X"D8",X"00",X"DA",X"00",X"DC",X"00",X"DE",X"00",
		X"E0",X"00",X"E1",X"00",X"E2",X"00",X"E3",X"00",X"E4",X"00",X"E5",X"00",X"E6",X"00",X"E7",X"00",
		X"00",X"01",X"FF",X"00",X"FE",X"00",X"FD",X"00",X"FC",X"00",X"FB",X"00",X"FA",X"00",X"F8",X"00",
		X"F6",X"00",X"F4",X"00",X"F2",X"00",X"F0",X"00",X"ED",X"00",X"EA",X"00",X"E8",X"00",X"E5",X"00",
		X"E2",X"00",X"DF",X"00",X"DC",X"00",X"D9",X"00",X"D6",X"00",X"D3",X"00",X"D0",X"00",X"CD",X"00",
		X"CA",X"00",X"C7",X"00",X"C4",X"00",X"C1",X"00",X"BE",X"00",X"BB",X"00",X"B8",X"00",X"B5",X"00",
		X"B2",X"00",X"AF",X"00",X"AB",X"00",X"A8",X"00",X"A5",X"00",X"A1",X"00",X"9D",X"00",X"99",X"00",
		X"96",X"00",X"92",X"00",X"8C",X"00",X"87",X"00",X"82",X"00",X"7B",X"00",X"78",X"00",X"72",X"00",
		X"6C",X"00",X"66",X"00",X"60",X"00",X"59",X"00",X"53",X"00",X"4C",X"00",X"45",X"00",X"3E",X"00",
		X"36",X"00",X"2F",X"00",X"28",X"00",X"20",X"00",X"18",X"00",X"10",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"FF",X"F0",X"FF",X"00",X"00",X"E0",X"FF",X"D8",X"FF",X"D1",X"FF",X"CA",X"FF",
		X"C2",X"FF",X"BB",X"FF",X"B4",X"FF",X"AD",X"FF",X"A7",X"FF",X"A0",X"FF",X"9A",X"FF",X"94",X"FF",
		X"8E",X"FF",X"88",X"FF",X"85",X"FF",X"88",X"FF",X"79",X"FF",X"74",X"FF",X"6E",X"FF",X"6A",X"FF",
		X"67",X"FF",X"63",X"FF",X"5F",X"FF",X"5B",X"FF",X"58",X"FF",X"55",X"FF",X"51",X"FF",X"4E",X"FF",
		X"4B",X"FF",X"48",X"FF",X"45",X"FF",X"45",X"FF",X"3F",X"FF",X"3C",X"FF",X"39",X"FF",X"36",X"FF",
		X"33",X"FF",X"30",X"FF",X"2D",X"FF",X"2A",X"FF",X"27",X"FF",X"24",X"FF",X"21",X"FF",X"1E",X"FF",
		X"1B",X"FF",X"18",X"FF",X"16",X"FF",X"13",X"FF",X"10",X"FF",X"0E",X"FF",X"0C",X"FF",X"0A",X"FF",
		X"08",X"FF",X"06",X"FF",X"05",X"FF",X"04",X"FF",X"03",X"FF",X"02",X"FF",X"01",X"FF",X"00",X"FF",
		X"00",X"FF",X"01",X"FF",X"02",X"FF",X"03",X"FF",X"04",X"FF",X"05",X"FF",X"06",X"FF",X"08",X"FF",
		X"0A",X"FF",X"0C",X"FF",X"0E",X"FF",X"10",X"FF",X"13",X"FF",X"16",X"FF",X"18",X"FF",X"1B",X"FF",
		X"1E",X"FF",X"21",X"FF",X"24",X"FF",X"27",X"FF",X"2A",X"FF",X"2D",X"FF",X"30",X"FF",X"33",X"FF",
		X"36",X"FF",X"39",X"FF",X"3C",X"FF",X"3F",X"FF",X"42",X"FF",X"45",X"FF",X"48",X"FF",X"4B",X"FF",
		X"4E",X"FF",X"51",X"FF",X"55",X"FF",X"58",X"FF",X"5B",X"FF",X"5F",X"FF",X"63",X"FF",X"67",X"FF",
		X"6A",X"FF",X"6E",X"FF",X"74",X"FF",X"79",X"FF",X"7E",X"FF",X"85",X"FF",X"88",X"FF",X"8E",X"FF",
		X"94",X"FF",X"9A",X"FF",X"A0",X"FF",X"A7",X"FF",X"AD",X"FF",X"B4",X"FF",X"BB",X"FF",X"C2",X"FF",
		X"CA",X"FF",X"D1",X"FF",X"D8",X"FF",X"E0",X"FF",X"E8",X"FF",X"F0",X"FF",X"F8",X"FF",X"00",X"00",
		X"00",X"00",X"08",X"00",X"10",X"00",X"18",X"00",X"20",X"00",X"28",X"00",X"2F",X"00",X"36",X"00",
		X"3E",X"00",X"45",X"00",X"4C",X"00",X"53",X"00",X"59",X"00",X"60",X"00",X"66",X"00",X"6C",X"00",
		X"72",X"00",X"78",X"00",X"7B",X"00",X"7B",X"00",X"87",X"00",X"8C",X"00",X"92",X"00",X"96",X"00",
		X"99",X"00",X"9D",X"00",X"A1",X"00",X"A5",X"00",X"A8",X"00",X"AB",X"00",X"AF",X"00",X"B2",X"00",
		X"B5",X"00",X"B8",X"00",X"BB",X"00",X"B8",X"00",X"C1",X"00",X"C4",X"00",X"C7",X"00",X"CA",X"00",
		X"CD",X"00",X"D0",X"00",X"D3",X"00",X"D6",X"00",X"D9",X"00",X"DC",X"00",X"DF",X"00",X"E2",X"00",
		X"E5",X"00",X"E8",X"00",X"EA",X"00",X"E5",X"00",X"F0",X"00",X"F2",X"00",X"F4",X"00",X"F6",X"00",
		X"F8",X"00",X"FA",X"00",X"FB",X"00",X"FC",X"00",X"FD",X"00",X"FE",X"00",X"FF",X"00",X"00",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
