`define BUILD_DATE "190320"
`define BUILD_TIME "164646"
