library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"11",X"33",X"22",X"00",X"00",X"55",X"55",X"55",X"55",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"66",X"66",X"00",
		X"66",X"77",X"DD",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"77",X"33",X"00",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"FF",X"FF",X"44",X"44",X"44",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"66",X"33",X"11",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"77",X"00",
		X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"33",X"11",X"11",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"44",X"77",X"77",X"00",
		X"11",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"44",X"44",X"44",X"44",X"77",X"77",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"FF",X"FF",X"00",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"EE",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"77",X"33",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"FF",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",
		X"BB",X"BB",X"BB",X"BB",X"FF",X"FF",X"00",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"11",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",X"00",X"00",X"77",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"77",X"FF",X"CC",X"CC",X"FF",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"EE",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"77",
		X"33",X"33",X"33",X"33",X"FF",X"EE",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"FF",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"88",X"22",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"33",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"EE",X"22",X"22",X"00",X"11",X"22",X"22",X"22",X"33",
		X"AA",X"AA",X"AA",X"22",X"00",X"00",X"00",X"EE",X"22",X"22",X"22",X"11",X"00",X"22",X"22",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",
		X"33",X"33",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"77",X"77",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",
		X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"EE",X"EE",X"EE",X"66",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"CC",X"00",X"22",X"EE",X"22",X"00",X"00",X"88",X"77",X"00",X"00",X"FF",X"44",X"00",X"00",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"22",X"44",X"88",X"77",X"00",X"88",X"DD",X"AA",X"88",X"88",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"22",X"44",X"88",X"77",X"00",X"99",X"AA",X"AA",X"AA",X"EE",
		X"22",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"88",X"77",X"00",X"CC",X"BB",X"88",X"88",X"CC",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"CC",X"22",X"22",X"CC",X"00",X"22",X"EE",X"22",X"77",X"88",X"88",X"77",X"00",X"00",X"FF",X"44",
		X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"22",X"22",X"AA",X"77",X"88",X"88",X"77",X"00",X"66",X"99",X"88",
		X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"77",X"88",X"88",X"77",X"00",X"88",X"DD",X"AA",
		X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"77",X"88",X"88",X"77",X"00",X"99",X"AA",X"AA",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"CC",X"00",X"88",X"77",X"00",X"77",X"88",X"88",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"20",X"90",X"80",X"00",X"00",X"30",X"30",X"10",X"10",X"00",X"00",
		X"41",X"21",X"12",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"0C",X"8C",X"0C",X"00",X"00",X"00",X"07",X"0F",X"0F",X"C3",X"1F",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"0F",X"2F",X"4F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"07",X"4F",X"0F",X"A7",X"87",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"D3",X"87",X"97",X"0F",X"2F",X"07",X"00",X"00",X"33",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"0E",X"8E",X"1F",X"0F",
		X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"4F",X"1F",X"0F",X"4F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"01",X"03",X"87",X"87",X"87",X"47",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"10",
		X"EF",X"47",X"07",X"07",X"03",X"01",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",
		X"0F",X"0B",X"0C",X"0F",X"01",X"00",X"00",X"00",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"68",X"68",X"68",X"6E",X"6E",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"68",X"68",X"68",X"68",X"68",X"0C",X"00",X"00",X"0F",X"0F",X"07",X"0C",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"20",
		X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"10",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"0C",X"0F",X"CF",X"2F",X"0F",X"0F",
		X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"30",X"52",X"61",X"F1",X"BC",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",
		X"D2",X"63",X"52",X"30",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"48",X"84",X"C2",X"E0",X"00",X"00",X"E0",X"B4",X"7C",X"E1",X"5B",X"A5",
		X"68",X"84",X"C0",X"80",X"00",X"00",X"00",X"00",X"F5",X"E1",X"5A",X"BE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"33",X"31",X"71",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F3",X"71",X"31",X"33",X"0F",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"8E",X"CF",X"88",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"CF",X"8E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F1",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",
		X"E0",X"F1",X"E0",X"E0",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"DD",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"EF",X"67",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"23",X"67",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"79",X"69",X"0F",X"1F",X"FF",X"FF",X"33",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"33",X"79",X"69",X"0F",X"1F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"88",X"00",X"88",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"88",X"00",X"88",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"00",X"33",X"74",X"74",X"F8",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"FF",X"F9",X"F9",X"F9",X"F8",X"74",X"74",X"33",X"00",
		X"FF",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"FF",
		X"00",X"CC",X"E2",X"E2",X"F1",X"F9",X"F9",X"F9",X"FF",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"F1",X"E2",X"E2",X"CC",X"00",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FF",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"E2",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"E2",X"E2",X"CC",X"00",
		X"00",X"33",X"74",X"74",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"74",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F8",X"F8",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"F1",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F1",X"F1",X"FF",X"00",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"F0",X"F9",X"F9",X"F9",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F0",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"0C",X"8C",X"0C",X"00",X"00",X"30",X"30",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"20",X"90",X"80",X"00",X"00",X"00",X"07",X"0F",X"0F",X"C3",X"1F",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"21",X"12",X"03",X"03",X"01",X"00",X"00",X"07",X"08",X"0F",X"2F",X"4F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"07",X"4F",X"0F",X"A7",X"87",X"00",X"00",X"00",X"08",X"0E",X"8E",X"1F",X"0F",
		X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"33",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"D3",X"87",X"97",X"0F",X"2F",X"07",X"00",X"00",X"4F",X"1F",X"0F",X"4F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"10",
		X"00",X"00",X"01",X"03",X"87",X"87",X"87",X"47",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"47",X"07",X"07",X"03",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"0C",X"68",X"68",X"68",X"6E",X"6E",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",
		X"00",X"00",X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"68",X"68",X"68",X"68",X"68",X"0C",X"00",X"00",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0B",X"0C",X"0F",X"01",X"00",X"00",X"00",X"0F",X"0F",X"07",X"0C",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"20",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0C",X"0F",X"CF",X"2F",X"0F",X"0F",
		X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"80",X"48",X"84",X"C2",X"E0",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",
		X"00",X"00",X"00",X"30",X"52",X"61",X"F1",X"BC",X"00",X"00",X"E0",X"B4",X"7C",X"E1",X"5B",X"A5",
		X"68",X"84",X"C0",X"80",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"D2",X"63",X"52",X"30",X"00",X"00",X"00",X"00",X"F5",X"E1",X"5A",X"BE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"33",X"31",X"71",X"F3",X"00",X"00",X"00",X"08",X"0C",X"8E",X"CF",X"88",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F3",X"71",X"31",X"33",X"0F",X"00",X"00",X"FF",X"88",X"CF",X"8E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"DD",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",
		X"E0",X"F1",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"CC",X"88",X"8C",X"4E",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"00",X"7F",X"BF",X"7F",X"AF",X"5F",X"7F",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"11",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"8C",X"08",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"00",X"7F",X"BF",X"7F",X"AF",X"5F",X"7F",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"11",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"EE",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"69",X"0F",X"71",X"69",X"0F",X"17",X"00",X"00",X"00",X"88",X"EE",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"77",X"33",X"00",X"00",X"00",
		X"00",X"EE",X"EE",X"EE",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"69",X"0F",X"71",X"69",X"0F",X"17",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",
		X"EE",X"66",X"66",X"EE",X"EE",X"EE",X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"EE",X"EE",X"EE",X"EE",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"EE",X"EE",X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0C",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0E",X"0E",
		X"00",X"00",X"00",X"08",X"08",X"08",X"0C",X"0C",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0C",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"0C",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"0C",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"10",X"F0",X"F0",X"F0",X"F3",X"F3",X"F0",X"00",X"F0",X"F1",X"F2",X"F2",X"F1",X"F1",X"F2",
		X"80",X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"00",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F0",X"F3",X"F3",X"F0",X"F0",X"F0",X"10",X"00",X"F2",X"F1",X"F1",X"F2",X"F2",X"F1",X"F0",X"00",
		X"00",X"C0",X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"10",X"F0",X"F0",X"F0",X"F3",X"F3",X"F0",X"00",X"F0",X"F1",X"F2",X"F2",X"F1",X"F1",X"F2",
		X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"C0",X"00",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F0",X"F3",X"F3",X"F0",X"F0",X"F0",X"10",X"00",X"F2",X"F1",X"F1",X"F2",X"F2",X"F1",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"00",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"11",X"00",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"00",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"11",X"00",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"00",X"FF",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"11",X"00",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"00",X"FF",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"11",X"00",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",X"FF",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"11",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"11",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"01",X"30",X"30",X"67",X"77",
		X"00",X"11",X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"67",X"30",X"30",X"01",X"00",X"00",X"00",
		X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"01",X"30",X"30",X"67",X"77",
		X"00",X"11",X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"67",X"30",X"30",X"01",X"00",X"00",X"00",
		X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"06",X"02",X"0C",X"00",X"02",X"02",X"0A",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"0F",X"04",X"02",X"01",X"02",X"0C",X"00",X"08",X"0E",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"02",X"0C",X"00",X"0C",X"02",X"02",X"02",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"09",X"09",X"09",X"07",X"00",X"0F",X"0C",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"77",X"00",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"CC",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"33",X"33",X"77",X"77",X"77",
		X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"01",X"02",X"04",X"0C",X"08",X"84",X"84",X"08",X"01",X"00",X"00",X"00",X"09",X"05",X"03",X"00",
		X"00",X"08",X"07",X"78",X"FA",X"F5",X"EA",X"7B",X"00",X"00",X"00",X"0B",X"B5",X"EA",X"77",X"32",
		X"08",X"84",X"84",X"08",X"0C",X"04",X"02",X"01",X"00",X"01",X"01",X"01",X"03",X"04",X"08",X"00",
		X"26",X"5D",X"B2",X"7C",X"07",X"00",X"00",X"00",X"72",X"E6",X"CC",X"FC",X"E3",X"0E",X"00",X"00",
		X"00",X"60",X"60",X"E0",X"E0",X"E8",X"CC",X"88",X"00",X"00",X"00",X"01",X"00",X"00",X"67",X"77",
		X"00",X"11",X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"00",X"00",X"F0",X"F8",X"FD",X"FF",X"FF",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"67",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"60",X"60",X"E0",X"E0",X"E8",X"CC",X"88",X"00",X"00",X"00",X"11",X"23",X"23",X"77",X"77",
		X"00",X"11",X"FF",X"1D",X"0C",X"0F",X"1F",X"FF",X"00",X"00",X"F0",X"F8",X"FD",X"FF",X"FF",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"23",X"23",X"11",X"00",X"00",X"00",
		X"FF",X"1D",X"0C",X"0F",X"1F",X"FF",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"33",X"77",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"77",X"77",X"33",X"11",X"11",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"33",X"77",X"77",X"FF",X"77",X"EE",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"33",X"33",X"11",X"11",X"11",X"00",X"00",X"88",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",X"EE",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",X"77",X"77",X"FF",X"FF",X"FF",
		X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"66",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"77",X"77",X"FF",
		X"00",X"88",X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"77",X"33",X"33",X"33",X"11",
		X"00",X"00",X"CC",X"EE",X"EE",X"EE",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",
		X"88",X"CC",X"EE",X"EE",X"EE",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",
		X"CC",X"EE",X"EE",X"EE",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"CC",X"EE",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"44",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"00",X"00",X"11",X"99",X"44",X"00",X"00",
		X"00",X"22",X"11",X"88",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"22",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
