library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu4_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu4_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"33",X"3A",X"33",X"74",X"93",X"3A",X"33",X"43",X"93",X"33",X"33",X"74",X"33",X"33",X"33",X"43",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"08",X"08",X"17",X"51",X"51",X"3B",X"41",X"3D",X"08",X"08",X"17",X"51",X"51",X"13",X"51",
		X"13",X"08",X"08",X"27",X"0A",X"51",X"13",X"51",X"13",X"08",X"08",X"08",X"17",X"51",X"5B",X"41",
		X"5D",X"08",X"07",X"08",X"17",X"51",X"3B",X"41",X"3D",X"08",X"08",X"18",X"1A",X"51",X"13",X"51",
		X"13",X"08",X"08",X"17",X"51",X"51",X"13",X"51",X"13",X"08",X"08",X"17",X"51",X"51",X"5B",X"41",
		X"5D",X"10",X"44",X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"44",X"44",X"33",X"33",X"44",X"44",
		X"33",X"33",X"47",X"44",X"33",X"33",X"44",X"44",X"33",X"33",X"44",X"43",X"33",X"33",X"44",X"43",
		X"33",X"33",X"08",X"08",X"17",X"51",X"3B",X"41",X"41",X"3D",X"19",X"19",X"1A",X"51",X"13",X"51",
		X"51",X"13",X"51",X"51",X"51",X"51",X"5B",X"41",X"41",X"5D",X"51",X"3E",X"3F",X"51",X"00",X"01",
		X"01",X"02",X"51",X"4E",X"4F",X"51",X"10",X"21",X"21",X"12",X"51",X"51",X"51",X"51",X"3B",X"41",
		X"41",X"3D",X"28",X"28",X"0A",X"51",X"13",X"51",X"51",X"13",X"08",X"08",X"17",X"51",X"5B",X"41",
		X"41",X"5D",X"10",X"44",X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"36",X"63",X"33",X"33",X"33",X"33",X"44",X"43",X"33",X"33",X"44",
		X"43",X"33",X"33",X"07",X"08",X"17",X"51",X"00",X"01",X"01",X"02",X"19",X"19",X"1A",X"51",X"10",
		X"21",X"21",X"12",X"28",X"28",X"0A",X"51",X"3B",X"41",X"41",X"3D",X"08",X"08",X"17",X"51",X"13",
		X"0E",X"0F",X"13",X"07",X"08",X"17",X"51",X"13",X"1E",X"1F",X"13",X"08",X"08",X"17",X"51",X"5B",
		X"41",X"41",X"5D",X"08",X"08",X"17",X"51",X"00",X"01",X"01",X"02",X"08",X"08",X"17",X"51",X"10",
		X"21",X"21",X"12",X"10",X"74",X"43",X"33",X"33",X"44",X"43",X"36",X"63",X"44",X"43",X"33",X"33",
		X"44",X"43",X"35",X"53",X"74",X"43",X"35",X"53",X"44",X"43",X"33",X"33",X"44",X"43",X"33",X"33",
		X"44",X"43",X"36",X"63",X"07",X"08",X"17",X"51",X"51",X"3B",X"3C",X"3D",X"08",X"08",X"17",X"51",
		X"51",X"4B",X"4C",X"4D",X"08",X"08",X"17",X"51",X"51",X"5B",X"5C",X"5D",X"08",X"18",X"1A",X"51",
		X"51",X"00",X"01",X"02",X"19",X"1A",X"51",X"51",X"51",X"10",X"21",X"12",X"51",X"51",X"51",X"51",
		X"51",X"3B",X"41",X"3D",X"28",X"28",X"0A",X"51",X"51",X"13",X"51",X"13",X"08",X"08",X"17",X"51",
		X"51",X"5B",X"41",X"5D",X"10",X"74",X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"44",X"43",X"33",
		X"33",X"44",X"43",X"33",X"33",X"44",X"33",X"33",X"63",X"33",X"33",X"33",X"33",X"44",X"43",X"33",
		X"33",X"44",X"43",X"33",X"33",X"51",X"51",X"51",X"51",X"51",X"3B",X"41",X"3D",X"28",X"28",X"0A",
		X"51",X"51",X"13",X"50",X"13",X"08",X"08",X"17",X"51",X"51",X"5B",X"41",X"5D",X"08",X"08",X"17",
		X"51",X"51",X"00",X"01",X"02",X"08",X"07",X"17",X"51",X"51",X"10",X"21",X"12",X"08",X"08",X"17",
		X"51",X"51",X"34",X"35",X"36",X"08",X"08",X"17",X"51",X"51",X"44",X"51",X"46",X"08",X"08",X"17",
		X"51",X"51",X"54",X"55",X"56",X"10",X"33",X"33",X"33",X"33",X"44",X"43",X"33",X"93",X"44",X"43",
		X"33",X"33",X"44",X"43",X"33",X"33",X"47",X"43",X"33",X"63",X"44",X"43",X"33",X"33",X"44",X"43",
		X"33",X"33",X"44",X"43",X"33",X"33",X"08",X"08",X"17",X"51",X"34",X"35",X"35",X"36",X"08",X"08",
		X"17",X"51",X"44",X"51",X"51",X"46",X"08",X"08",X"17",X"51",X"54",X"55",X"55",X"56",X"08",X"08",
		X"17",X"51",X"3B",X"41",X"41",X"3D",X"19",X"19",X"1A",X"51",X"13",X"51",X"51",X"13",X"51",X"51",
		X"51",X"51",X"5B",X"41",X"41",X"5D",X"51",X"00",X"01",X"01",X"01",X"01",X"01",X"02",X"51",X"10",
		X"21",X"21",X"21",X"21",X"21",X"12",X"10",X"44",X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"44",
		X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"66",X"66",X"66",X"08",X"07",X"17",X"51",X"51",X"3B",X"41",X"3D",X"08",
		X"08",X"17",X"51",X"51",X"13",X"50",X"13",X"08",X"08",X"17",X"51",X"51",X"5B",X"41",X"5D",X"18",
		X"19",X"1A",X"51",X"51",X"00",X"01",X"02",X"27",X"0A",X"51",X"51",X"51",X"10",X"21",X"12",X"08",
		X"27",X"0A",X"51",X"51",X"3B",X"41",X"3D",X"08",X"08",X"17",X"51",X"51",X"13",X"50",X"13",X"08",
		X"08",X"17",X"51",X"51",X"5B",X"41",X"5D",X"10",X"47",X"43",X"33",X"33",X"44",X"43",X"33",X"93",
		X"44",X"43",X"33",X"33",X"44",X"43",X"33",X"33",X"44",X"33",X"33",X"63",X"44",X"43",X"33",X"33",
		X"44",X"43",X"33",X"93",X"44",X"43",X"33",X"33",X"3B",X"41",X"3D",X"85",X"86",X"16",X"51",X"51",
		X"13",X"51",X"13",X"85",X"86",X"16",X"51",X"51",X"13",X"51",X"13",X"85",X"86",X"16",X"51",X"51",
		X"5B",X"41",X"5D",X"85",X"86",X"16",X"51",X"51",X"3B",X"41",X"3D",X"85",X"86",X"D1",X"D2",X"51",
		X"13",X"51",X"13",X"85",X"96",X"97",X"98",X"D3",X"13",X"51",X"13",X"A5",X"A6",X"A7",X"86",X"16",
		X"5B",X"41",X"5D",X"51",X"50",X"85",X"86",X"16",X"10",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",
		X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",X"33",
		X"3E",X"33",X"33",X"33",X"3E",X"33",X"33",X"93",X"3E",X"60",X"65",X"61",X"51",X"51",X"85",X"86",
		X"16",X"3B",X"41",X"3D",X"51",X"50",X"85",X"86",X"16",X"13",X"51",X"13",X"51",X"B5",X"B7",X"86",
		X"16",X"5B",X"41",X"5D",X"51",X"85",X"C6",X"C8",X"D4",X"3B",X"3C",X"3D",X"51",X"85",X"86",X"D5",
		X"51",X"4B",X"4C",X"4D",X"51",X"85",X"96",X"98",X"D3",X"5B",X"5C",X"5D",X"51",X"A5",X"A7",X"86",
		X"16",X"60",X"65",X"61",X"51",X"50",X"85",X"86",X"16",X"10",X"44",X"43",X"33",X"3E",X"33",X"33",
		X"93",X"3E",X"33",X"33",X"33",X"3E",X"33",X"33",X"33",X"3E",X"33",X"33",X"33",X"EE",X"33",X"33",
		X"33",X"3E",X"33",X"33",X"33",X"3E",X"44",X"43",X"93",X"3E",X"40",X"41",X"42",X"51",X"B5",X"B7",
		X"86",X"16",X"34",X"35",X"36",X"51",X"85",X"C6",X"C8",X"D4",X"44",X"51",X"46",X"51",X"85",X"86",
		X"D5",X"51",X"54",X"55",X"56",X"51",X"85",X"96",X"98",X"D3",X"60",X"65",X"61",X"50",X"A5",X"A7",
		X"86",X"16",X"3B",X"3C",X"3D",X"B5",X"B6",X"B7",X"86",X"16",X"4B",X"4C",X"4D",X"85",X"C6",X"C7",
		X"C8",X"D4",X"5B",X"5C",X"5D",X"85",X"86",X"E1",X"E0",X"51",X"10",X"33",X"33",X"33",X"3E",X"33",
		X"33",X"33",X"3E",X"33",X"33",X"33",X"EE",X"33",X"33",X"33",X"3E",X"44",X"49",X"33",X"3E",X"33",
		X"33",X"33",X"3E",X"33",X"33",X"33",X"3E",X"33",X"33",X"3E",X"EE",X"3B",X"41",X"3D",X"85",X"86",
		X"16",X"51",X"51",X"13",X"51",X"13",X"85",X"86",X"16",X"51",X"51",X"13",X"51",X"13",X"85",X"86",
		X"E4",X"51",X"51",X"5B",X"41",X"5D",X"85",X"96",X"98",X"D3",X"51",X"60",X"61",X"50",X"A5",X"A7",
		X"86",X"16",X"51",X"34",X"35",X"36",X"B5",X"B7",X"86",X"16",X"51",X"44",X"51",X"46",X"85",X"C6",
		X"C8",X"D4",X"51",X"54",X"55",X"56",X"85",X"86",X"F0",X"51",X"51",X"10",X"33",X"33",X"3E",X"EE",
		X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",X"33",X"EE",X"44",X"93",X"33",X"EE",
		X"33",X"33",X"33",X"EE",X"33",X"33",X"33",X"EE",X"33",X"33",X"3E",X"EE",X"51",X"51",X"50",X"85",
		X"86",X"16",X"51",X"51",X"51",X"51",X"B5",X"B7",X"86",X"16",X"51",X"51",X"51",X"51",X"85",X"C6",
		X"C8",X"D4",X"51",X"51",X"51",X"50",X"85",X"86",X"F0",X"51",X"51",X"51",X"B6",X"B6",X"B7",X"86",
		X"16",X"51",X"51",X"51",X"C7",X"C7",X"C7",X"C8",X"D4",X"51",X"51",X"51",X"25",X"25",X"25",X"E0",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"10",X"33",X"93",X"3E",
		X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"39",X"33",X"EE",X"EE",X"33",X"33",X"EE",
		X"EE",X"33",X"33",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"3B",X"41",X"41",
		X"3D",X"00",X"01",X"01",X"02",X"13",X"0E",X"0F",X"13",X"30",X"51",X"51",X"32",X"13",X"1E",X"1F",
		X"13",X"10",X"11",X"11",X"12",X"5B",X"41",X"41",X"5D",X"50",X"51",X"51",X"51",X"34",X"35",X"35",
		X"36",X"51",X"B5",X"B6",X"B6",X"44",X"51",X"51",X"46",X"51",X"85",X"C6",X"C7",X"44",X"51",X"51",
		X"46",X"51",X"85",X"86",X"E1",X"54",X"55",X"55",X"56",X"51",X"85",X"86",X"16",X"10",X"33",X"33",
		X"33",X"33",X"35",X"53",X"33",X"33",X"35",X"53",X"33",X"33",X"33",X"33",X"93",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"3E",X"33",X"33",X"33",X"3E",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"E3",X"E3",X"D2",X"51",X"51",X"51",X"51",X"51",X"97",X"97",
		X"98",X"D3",X"51",X"51",X"51",X"51",X"A6",X"A7",X"86",X"D1",X"D2",X"51",X"51",X"51",X"50",X"85",
		X"96",X"97",X"98",X"D3",X"51",X"51",X"51",X"A5",X"A6",X"A7",X"86",X"16",X"51",X"51",X"51",X"51",
		X"50",X"85",X"86",X"16",X"51",X"51",X"51",X"51",X"51",X"85",X"86",X"16",X"51",X"51",X"10",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"3E",X"EE",X"EE",X"33",X"3E",X"EE",X"EE",X"93",
		X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"33",X"93",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"3B",
		X"41",X"41",X"3D",X"51",X"85",X"86",X"16",X"13",X"51",X"51",X"13",X"51",X"85",X"86",X"D1",X"5B",
		X"41",X"41",X"5D",X"51",X"85",X"96",X"97",X"00",X"01",X"01",X"02",X"51",X"A5",X"A6",X"A6",X"10",
		X"11",X"11",X"12",X"50",X"51",X"51",X"51",X"3B",X"41",X"41",X"3D",X"51",X"51",X"51",X"51",X"13",
		X"51",X"51",X"13",X"51",X"3E",X"3F",X"51",X"5B",X"41",X"41",X"5D",X"51",X"4E",X"4F",X"51",X"10",
		X"33",X"33",X"33",X"3E",X"33",X"33",X"33",X"3E",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"51",X"50",X"51",X"51",X"51",X"50",X"51",X"51",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"30",X"51",X"51",X"51",X"51",X"51",X"51",X"32",X"10",X"22",X"22",X"22",X"22",X"22",X"22",X"12",
		X"10",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"39",X"33",X"39",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"36",X"66",X"66",
		X"63",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"30",X"51",X"51",X"51",X"51",X"51",X"51",
		X"32",X"10",X"11",X"11",X"11",X"11",X"11",X"11",X"12",X"51",X"51",X"50",X"51",X"51",X"51",X"50",
		X"51",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"25",X"25",X"25",X"25",X"25",X"25",X"25",X"25",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"93",
		X"33",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"B6",X"B6",X"B6",X"B7",X"86",X"16",X"51",X"51",X"C7",X"C7",X"C7",X"C7",X"C8",X"D4",
		X"51",X"51",X"25",X"25",X"25",X"25",X"E0",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"E3",X"E3",X"E3",X"E3",X"D2",X"51",
		X"51",X"51",X"97",X"97",X"97",X"97",X"98",X"D3",X"51",X"51",X"A6",X"A6",X"A6",X"A7",X"86",X"16",
		X"51",X"51",X"10",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"33",X"3E",X"EE",X"33",
		X"33",X"3E",X"EE",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"25",X"25",X"25",X"25",X"25",X"25",X"25",X"25",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"E3",X"E3",X"E3",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"50",X"B5",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B7",X"C6",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C8",X"07",X"F1",X"25",X"25",X"25",X"25",X"25",X"25",X"E0",
		X"51",X"51",X"51",X"51",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"D2",X"51",X"97",X"97",X"97",X"97",
		X"97",X"98",X"07",X"F2",X"A6",X"A6",X"A6",X"A6",X"A7",X"96",X"97",X"97",X"51",X"51",X"51",X"50",
		X"A5",X"A6",X"A6",X"A6",X"10",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"37",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"33",X"33",X"7E",X"33",X"33",X"33",
		X"33",X"33",X"39",X"33",X"33",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"B5",
		X"B6",X"B6",X"B6",X"B6",X"B6",X"51",X"50",X"85",X"C6",X"C7",X"C7",X"C7",X"C7",X"51",X"51",X"85",
		X"86",X"E1",X"25",X"25",X"25",X"51",X"51",X"85",X"86",X"D1",X"E3",X"E3",X"E3",X"51",X"50",X"85",
		X"96",X"97",X"97",X"97",X"97",X"51",X"51",X"A5",X"A6",X"A6",X"A6",X"A6",X"A6",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"39",X"33",
		X"33",X"33",X"33",X"33",X"EE",X"EE",X"33",X"33",X"EE",X"EE",X"39",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"01",X"02",X"0B",X"0B",X"03",X"04",X"10",X"11",
		X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"4E",X"4E",
		X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"14",X"14",
		X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",X"22",X"20",X"20",X"21",X"30",X"31",
		X"24",X"24",X"32",X"33",X"23",X"23",X"30",X"33",X"33",X"33",X"33",X"37",X"73",X"37",X"73",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"B4",
		X"4B",X"B4",X"4B",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",
		X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"4E",
		X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"14",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",X"22",X"20",X"20",X"21",X"23",
		X"23",X"23",X"23",X"23",X"23",X"23",X"30",X"30",X"33",X"33",X"33",X"33",X"37",X"73",X"37",X"73",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"B4",X"4B",X"B4",X"4B",X"44",X"44",X"44",X"44",X"60",X"0B",X"0B",X"61",X"04",X"00",X"00",X"00",
		X"10",X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",X"22",X"20",X"20",X"21",
		X"70",X"71",X"71",X"72",X"33",X"23",X"23",X"23",X"30",X"33",X"33",X"33",X"33",X"37",X"73",X"37",
		X"73",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"B4",X"4B",X"B4",X"4B",X"44",X"45",X"44",X"44",X"40",X"41",X"4E",X"4E",X"4E",X"03",X"42",
		X"00",X"10",X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"4E",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",X"22",X"20",X"20",
		X"21",X"50",X"51",X"24",X"24",X"24",X"32",X"52",X"23",X"30",X"34",X"DD",X"DD",X"33",X"37",X"73",
		X"37",X"73",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"B4",X"4B",X"B4",X"4B",X"44",X"44",X"44",X"54",X"00",X"00",X"05",X"02",X"0B",X"0B",
		X"03",X"04",X"10",X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"4E",X"4E",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",X"22",X"20",
		X"20",X"21",X"06",X"07",X"08",X"71",X"09",X"0A",X"23",X"23",X"30",X"33",X"33",X"33",X"33",X"37",
		X"73",X"37",X"73",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"B4",X"4B",X"B4",X"4B",X"55",X"54",X"55",X"44",X"00",X"00",X"15",X"16",X"17",
		X"18",X"19",X"1A",X"10",X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"4E",X"4E",X"4E",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",X"22",
		X"20",X"20",X"21",X"25",X"26",X"27",X"28",X"29",X"2A",X"23",X"23",X"30",X"33",X"88",X"00",X"88",
		X"37",X"73",X"37",X"73",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"B4",X"4B",X"B4",X"4B",X"88",X"00",X"88",X"44",X"0B",X"0B",X"0B",X"5C",
		X"5D",X"1A",X"00",X"00",X"10",X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"4E",X"4E",X"4E",X"4E",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",X"21",
		X"22",X"20",X"20",X"21",X"5E",X"5E",X"5E",X"5F",X"29",X"2A",X"23",X"23",X"30",X"EE",X"E2",X"88",
		X"33",X"37",X"73",X"37",X"73",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"B4",X"4B",X"B4",X"4B",X"EE",X"EE",X"88",X"44",X"00",X"00",X"00",
		X"6C",X"6D",X"6E",X"0B",X"0B",X"10",X"11",X"12",X"10",X"10",X"11",X"12",X"10",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"4E",X"4E",X"4E",X"4E",X"4E",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"20",X"20",
		X"21",X"22",X"20",X"20",X"21",X"23",X"23",X"23",X"7C",X"7D",X"7E",X"5E",X"5E",X"30",X"33",X"33",
		X"3E",X"EE",X"37",X"73",X"37",X"73",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"B4",X"4B",X"B4",X"4B",X"44",X"44",X"5E",X"EE",X"34",X"35",
		X"36",X"37",X"38",X"39",X"3A",X"3B",X"5B",X"6B",X"75",X"4E",X"76",X"5B",X"6B",X"4E",X"5B",X"6B",
		X"75",X"4E",X"76",X"5B",X"6B",X"4E",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"54",X"55",
		X"56",X"56",X"56",X"56",X"5A",X"4E",X"64",X"65",X"57",X"58",X"59",X"4E",X"6A",X"4E",X"64",X"65",
		X"67",X"68",X"69",X"4E",X"6A",X"4E",X"64",X"65",X"77",X"78",X"79",X"4E",X"6A",X"4E",X"30",X"34",
		X"44",X"44",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"34",X"44",X"44",X"33",X"35",
		X"55",X"55",X"33",X"35",X"DD",X"DD",X"33",X"35",X"D7",X"DD",X"33",X"35",X"DD",X"DD",X"33",X"64",
		X"65",X"4E",X"4E",X"4E",X"4E",X"6A",X"4E",X"64",X"65",X"57",X"58",X"59",X"4E",X"6A",X"4E",X"64",
		X"65",X"67",X"68",X"69",X"4E",X"6A",X"4E",X"64",X"65",X"77",X"78",X"79",X"4E",X"6A",X"4E",X"64",
		X"65",X"4E",X"4E",X"4E",X"4E",X"6A",X"4E",X"64",X"65",X"57",X"58",X"59",X"4E",X"6A",X"4E",X"64",
		X"65",X"67",X"68",X"69",X"4E",X"6A",X"4E",X"64",X"65",X"77",X"78",X"79",X"4E",X"6A",X"4E",X"30",
		X"35",X"DD",X"DD",X"33",X"35",X"DD",X"DD",X"33",X"35",X"D7",X"DD",X"33",X"35",X"DD",X"DD",X"33",
		X"35",X"DD",X"DD",X"33",X"35",X"DD",X"DD",X"33",X"35",X"D7",X"DD",X"33",X"35",X"DD",X"DD",X"33",
		X"7A",X"0B",X"63",X"63",X"63",X"63",X"0B",X"7A",X"0B",X"0C",X"0D",X"0E",X"0D",X"0E",X"0F",X"0B",
		X"63",X"1B",X"1C",X"1D",X"1C",X"1D",X"1E",X"63",X"63",X"1B",X"1C",X"1D",X"1F",X"1D",X"1E",X"63",
		X"63",X"2B",X"1C",X"2C",X"2D",X"2C",X"2E",X"63",X"63",X"2F",X"1C",X"3C",X"2D",X"3D",X"2E",X"63",
		X"0B",X"3E",X"3F",X"4C",X"3F",X"4D",X"53",X"0B",X"7A",X"0B",X"63",X"63",X"63",X"63",X"0B",X"7A",
		X"30",X"73",X"33",X"33",X"37",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"73",X"33",X"33",
		X"37",X"7A",X"0B",X"63",X"63",X"63",X"63",X"0B",X"7A",X"0B",X"0C",X"0E",X"0D",X"0D",X"66",X"0F",
		X"0B",X"63",X"2B",X"3D",X"2D",X"2D",X"62",X"7B",X"63",X"63",X"1B",X"1D",X"1C",X"1F",X"1D",X"1E",
		X"63",X"63",X"1B",X"1D",X"1F",X"1F",X"1D",X"1E",X"63",X"63",X"2F",X"3C",X"1C",X"1C",X"2C",X"2E",
		X"63",X"0B",X"3E",X"4C",X"3F",X"3F",X"4D",X"53",X"0B",X"7A",X"0B",X"63",X"63",X"63",X"63",X"0B",
		X"7A",X"30",X"73",X"33",X"33",X"37",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"73",X"33",
		X"33",X"37",X"7A",X"0B",X"63",X"63",X"63",X"63",X"0B",X"7A",X"0B",X"0C",X"0E",X"0D",X"66",X"0D",
		X"0F",X"0B",X"63",X"2F",X"74",X"1C",X"23",X"1C",X"7B",X"63",X"63",X"1B",X"1D",X"1C",X"1F",X"1F",
		X"1E",X"63",X"63",X"1B",X"1D",X"1F",X"1F",X"1F",X"1E",X"63",X"63",X"2F",X"3C",X"2D",X"62",X"1C",
		X"7B",X"63",X"0B",X"2B",X"62",X"1C",X"74",X"1C",X"7B",X"0B",X"0B",X"1B",X"1D",X"1C",X"1D",X"1F",
		X"1E",X"0B",X"30",X"73",X"33",X"33",X"37",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"0B",X"2F",X"3C",X"2D",X"3D",X"2D",X"2E",X"0B",X"0B",X"2F",X"23",X"1C",X"74",
		X"1C",X"7B",X"0B",X"63",X"2B",X"62",X"1C",X"74",X"1C",X"7B",X"63",X"63",X"1B",X"1D",X"1C",X"1D",
		X"1F",X"1E",X"63",X"63",X"1B",X"1D",X"1C",X"1D",X"1C",X"1E",X"63",X"63",X"1B",X"1D",X"1C",X"1D",
		X"1F",X"1E",X"63",X"0B",X"3E",X"4D",X"3F",X"4D",X"3F",X"53",X"0B",X"7A",X"0B",X"63",X"63",X"63",
		X"63",X"0B",X"7A",X"30",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"73",X"33",X"33",X"37",X"00",X"01",X"02",X"00",X"02",X"00",X"01",X"02",X"25",X"25",X"25",X"CB",
		X"CC",X"CD",X"CE",X"32",X"11",X"11",X"11",X"FE",X"30",X"DF",X"DE",X"32",X"AD",X"AE",X"AF",X"13",
		X"30",X"DF",X"DE",X"32",X"BD",X"BE",X"BF",X"13",X"30",X"DF",X"DE",X"32",X"01",X"01",X"01",X"FF",
		X"30",X"DF",X"DE",X"32",X"DA",X"DA",X"DA",X"DB",X"DC",X"DD",X"DE",X"32",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EB",X"12",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"34",X"33",X"33",X"33",X"34",
		X"33",X"00",X"03",X"34",X"33",X"00",X"03",X"34",X"33",X"33",X"33",X"34",X"33",X"44",X"44",X"44",
		X"33",X"33",X"33",X"33",X"33",X"00",X"01",X"02",X"00",X"02",X"00",X"01",X"02",X"30",X"51",X"C9",
		X"CB",X"CC",X"CB",X"CC",X"25",X"30",X"51",X"16",X"32",X"D7",X"D8",X"F9",X"11",X"30",X"51",X"16",
		X"32",X"30",X"32",X"13",X"AC",X"30",X"51",X"16",X"32",X"E7",X"E8",X"13",X"BC",X"30",X"51",X"16",
		X"32",X"F7",X"F8",X"EF",X"01",X"30",X"51",X"D9",X"DB",X"DC",X"DB",X"DC",X"DA",X"10",X"11",X"E9",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"CC",X"33",X"33",X"33",
		X"CC",X"33",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"33",X"33",X"44",
		X"44",X"44",X"33",X"33",X"33",X"33",X"01",X"01",X"02",X"00",X"01",X"01",X"01",X"02",X"CB",X"CC",
		X"25",X"25",X"25",X"CD",X"CE",X"32",X"12",X"10",X"11",X"11",X"FC",X"DF",X"DE",X"32",X"88",X"89",
		X"8A",X"8B",X"30",X"DF",X"DE",X"32",X"87",X"99",X"9A",X"9B",X"30",X"DF",X"DE",X"32",X"02",X"00",
		X"01",X"01",X"FD",X"DF",X"DE",X"32",X"DB",X"DC",X"DA",X"DA",X"DA",X"DD",X"DE",X"32",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EB",X"12",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"34",X"33",X"33",
		X"33",X"34",X"33",X"00",X"00",X"34",X"33",X"00",X"00",X"34",X"33",X"33",X"33",X"34",X"33",X"44",
		X"44",X"44",X"33",X"33",X"33",X"33",X"33",X"00",X"01",X"02",X"00",X"01",X"02",X"00",X"01",X"30",
		X"51",X"C9",X"25",X"CB",X"CC",X"CB",X"CC",X"30",X"51",X"16",X"51",X"32",X"D7",X"D8",X"F9",X"30",
		X"51",X"16",X"FA",X"12",X"10",X"12",X"13",X"30",X"51",X"16",X"32",X"8D",X"8E",X"8F",X"13",X"30",
		X"51",X"16",X"FB",X"01",X"01",X"02",X"EF",X"30",X"51",X"D9",X"DA",X"DA",X"DA",X"DB",X"DC",X"10",
		X"11",X"E9",X"EA",X"EA",X"EA",X"EA",X"EA",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"3C",X"C3",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"03",X"33",X"33",X"33",X"33",
		X"33",X"44",X"44",X"44",X"33",X"33",X"33",X"33",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"30",X"FA",X"11",X"11",X"11",X"11",X"FC",X"ED",X"30",X"32",X"88",X"89",X"8A",X"8B",X"30",X"ED",
		X"30",X"32",X"87",X"99",X"9A",X"9B",X"30",X"ED",X"E7",X"E8",X"8C",X"8D",X"8E",X"8F",X"30",X"ED",
		X"F7",X"F8",X"9C",X"9D",X"9E",X"9F",X"30",X"ED",X"30",X"FB",X"01",X"01",X"01",X"01",X"FD",X"ED",
		X"10",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"12",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"3C",X"33",X"00",X"00",X"3C",X"33",X"00",X"00",X"3C",X"33",X"00",X"00",X"3C",X"33",X"00",X"00",
		X"3C",X"33",X"33",X"33",X"3C",X"3C",X"CC",X"CC",X"C3",X"00",X"01",X"01",X"01",X"01",X"01",X"02",
		X"51",X"30",X"51",X"51",X"51",X"51",X"51",X"32",X"51",X"10",X"21",X"21",X"21",X"21",X"21",X"12",
		X"51",X"47",X"04",X"05",X"05",X"05",X"05",X"05",X"06",X"57",X"14",X"15",X"15",X"15",X"15",X"15",
		X"16",X"57",X"14",X"15",X"15",X"15",X"15",X"15",X"16",X"67",X"14",X"15",X"15",X"15",X"15",X"15",
		X"16",X"51",X"24",X"25",X"25",X"25",X"25",X"25",X"26",X"10",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"36",X"66",X"66",X"33",X"C5",X"55",X"55",X"53",X"C5",X"55",X"55",X"53",X"C5",X"55",
		X"55",X"53",X"C5",X"55",X"55",X"53",X"33",X"33",X"33",X"33",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"00",X"01",X"01",X"02",X"00",X"01",X"02",X"51",X"30",X"51",X"51",X"32",X"30",
		X"51",X"32",X"51",X"30",X"51",X"51",X"32",X"30",X"51",X"32",X"51",X"10",X"11",X"11",X"12",X"10",
		X"11",X"12",X"51",X"00",X"01",X"01",X"01",X"01",X"01",X"02",X"51",X"10",X"11",X"11",X"11",X"11",
		X"11",X"12",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"10",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"01",X"02",X"34",X"35",
		X"35",X"35",X"36",X"30",X"51",X"32",X"44",X"51",X"51",X"51",X"46",X"30",X"51",X"32",X"44",X"51",
		X"51",X"51",X"46",X"30",X"51",X"32",X"44",X"51",X"51",X"51",X"46",X"10",X"11",X"12",X"54",X"55",
		X"55",X"55",X"56",X"51",X"51",X"50",X"51",X"51",X"50",X"3E",X"3F",X"51",X"51",X"51",X"51",X"51",
		X"51",X"4E",X"4F",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"10",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"93",X"39",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"47",X"00",X"01",X"01",
		X"01",X"01",X"01",X"02",X"57",X"30",X"51",X"51",X"51",X"51",X"51",X"32",X"57",X"30",X"51",X"51",
		X"51",X"51",X"51",X"32",X"67",X"10",X"11",X"11",X"11",X"11",X"11",X"12",X"00",X"01",X"01",X"02",
		X"47",X"37",X"38",X"39",X"30",X"51",X"51",X"32",X"57",X"0E",X"0F",X"30",X"30",X"51",X"51",X"32",
		X"57",X"1E",X"1F",X"30",X"10",X"11",X"11",X"12",X"67",X"01",X"01",X"FD",X"10",X"C3",X"33",X"33",
		X"33",X"C3",X"33",X"33",X"33",X"C3",X"33",X"33",X"33",X"C3",X"33",X"33",X"33",X"33",X"33",X"CC",
		X"CC",X"33",X"33",X"C5",X"53",X"33",X"33",X"C5",X"53",X"33",X"33",X"C3",X"33",X"00",X"01",X"01",
		X"01",X"02",X"00",X"01",X"02",X"30",X"51",X"51",X"51",X"43",X"30",X"51",X"43",X"10",X"11",X"11",
		X"11",X"12",X"10",X"11",X"12",X"00",X"01",X"01",X"02",X"00",X"01",X"01",X"02",X"30",X"51",X"51",
		X"33",X"30",X"51",X"51",X"32",X"30",X"51",X"51",X"32",X"30",X"51",X"51",X"32",X"30",X"51",X"51",
		X"33",X"30",X"51",X"51",X"32",X"10",X"11",X"11",X"12",X"10",X"21",X"21",X"12",X"10",X"33",X"33",
		X"33",X"33",X"33",X"33",X"63",X"36",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"36",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"36",X"33",X"33",X"33",X"33",X"36",X"63",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"6A",X"6B",X"6B",X"6B",X"6C",X"25",X"CD",X"CE",X"6D",X"A8",
		X"A9",X"AA",X"30",X"EC",X"DF",X"DE",X"6D",X"B8",X"B9",X"BA",X"30",X"EC",X"DF",X"DE",X"6D",X"AB",
		X"B4",X"95",X"30",X"EC",X"DF",X"DE",X"6E",X"01",X"01",X"01",X"FD",X"EC",X"DF",X"DE",X"D9",X"DA",
		X"DA",X"DA",X"DA",X"DA",X"DD",X"DE",X"90",X"83",X"83",X"83",X"83",X"83",X"83",X"B0",X"10",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"43",X"3E",X"EE",X"3C",X"43",X"3E",X"EE",X"3C",X"43",X"3E",
		X"EE",X"3C",X"43",X"33",X"33",X"3C",X"43",X"44",X"44",X"44",X"43",X"33",X"33",X"33",X"33",X"FA",
		X"11",X"11",X"11",X"FC",X"51",X"00",X"02",X"32",X"A8",X"A9",X"AA",X"30",X"51",X"E7",X"E8",X"32",
		X"B8",X"B9",X"BA",X"30",X"51",X"F7",X"F8",X"32",X"AB",X"B4",X"95",X"30",X"51",X"10",X"12",X"7A",
		X"41",X"41",X"7B",X"7C",X"11",X"FC",X"51",X"32",X"A8",X"AA",X"13",X"A8",X"AA",X"30",X"EC",X"32",
		X"AB",X"95",X"13",X"AB",X"95",X"30",X"EC",X"FB",X"01",X"01",X"7D",X"01",X"01",X"FD",X"51",X"10",
		X"33",X"33",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",X"3E",X"EE",X"33",X"33",
		X"33",X"33",X"33",X"33",X"3E",X"E3",X"EE",X"3C",X"3E",X"E3",X"EE",X"3C",X"33",X"33",X"33",X"33",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"30",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"09",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"1B",X"25",X"25",X"25",X"25",X"25",X"25",X"25",X"25",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"E3",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"3A",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"5A",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"0B",X"11",X"11",X"0C",X"0D",X"B6",X"B6",X"B6",X"1C",X"01",X"01",X"1D",X"75",X"C7",
		X"C7",X"C7",X"29",X"11",X"11",X"2A",X"2B",X"25",X"25",X"25",X"1C",X"01",X"01",X"1D",X"B9",X"51",
		X"51",X"51",X"29",X"11",X"11",X"2A",X"B9",X"51",X"51",X"51",X"1C",X"01",X"01",X"1D",X"74",X"E3",
		X"E3",X"E3",X"29",X"11",X"11",X"2A",X"4A",X"97",X"97",X"97",X"5E",X"01",X"01",X"5F",X"66",X"A6",
		X"A6",X"A6",X"10",X"33",X"33",X"33",X"33",X"43",X"34",X"33",X"33",X"43",X"34",X"EE",X"EE",X"43",
		X"34",X"EE",X"EE",X"43",X"34",X"EE",X"EE",X"43",X"34",X"EE",X"EE",X"43",X"34",X"33",X"33",X"33",
		X"33",X"33",X"33",X"7A",X"8D",X"8E",X"8F",X"99",X"9D",X"9E",X"7A",X"9C",X"9D",X"9E",X"9F",X"8C",
		X"8D",X"8E",X"8F",X"9E",X"9F",X"AC",X"AD",X"AD",X"AE",X"8B",X"9D",X"8E",X"8F",X"AF",X"BC",X"BD",
		X"AF",X"9B",X"8D",X"8C",X"98",X"AF",X"BE",X"BF",X"AF",X"AB",X"9F",X"9C",X"9D",X"CC",X"AD",X"AD",
		X"CD",X"BB",X"9A",X"9E",X"9F",X"CF",X"DD",X"DE",X"DF",X"CE",X"9D",X"7A",X"8F",X"9C",X"9D",X"9E",
		X"9F",X"8C",X"7A",X"30",X"70",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",
		X"00",X"4C",X"C4",X"00",X"00",X"4C",X"C4",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"07",X"40",X"40",X"50",X"80",X"38",X"70",X"02",X"58",X"62",X"3C",X"3C",X"54",
		X"7C",X"38",X"6C",X"02",X"56",X"5E",X"3C",X"3C",X"58",X"78",X"3C",X"68",X"02",X"54",X"5E",X"38",
		X"38",X"5C",X"74",X"3C",X"64",X"02",X"54",X"5A",X"38",X"38",X"60",X"70",X"40",X"60",X"02",X"52",
		X"5A",X"34",X"34",X"64",X"6C",X"40",X"5C",X"02",X"52",X"56",X"38",X"32",X"68",X"68",X"44",X"58",
		X"02",X"52",X"56",X"40",X"3A",X"6C",X"60",X"44",X"4E",X"03",X"50",X"52",X"3C",X"38",X"70",X"58",
		X"48",X"48",X"03",X"4E",X"52",X"38",X"36",X"74",X"50",X"48",X"42",X"03",X"4E",X"50",X"34",X"34",
		X"78",X"48",X"4C",X"3C",X"03",X"4C",X"4E",X"30",X"32",X"7C",X"40",X"4C",X"36",X"03",X"4C",X"4E",
		X"28",X"30",X"80",X"40",X"50",X"30",X"03",X"4A",X"4C",X"30",X"38",X"84",X"38",X"50",X"2C",X"04",
		X"48",X"4A",X"2E",X"36",X"88",X"30",X"54",X"28",X"04",X"46",X"48",X"2C",X"34",X"8C",X"2C",X"54",
		X"24",X"04",X"44",X"46",X"2A",X"32",X"90",X"28",X"58",X"20",X"04",X"42",X"44",X"28",X"30",X"94",
		X"24",X"58",X"1C",X"04",X"40",X"42",X"26",X"30",X"98",X"20",X"5C",X"18",X"04",X"40",X"40",X"38",
		X"2C",X"9C",X"1E",X"5C",X"14",X"05",X"3E",X"3E",X"34",X"26",X"A0",X"1C",X"60",X"10",X"05",X"3C",
		X"3C",X"30",X"20",X"A4",X"18",X"60",X"0C",X"05",X"3A",X"3A",X"2C",X"18",X"A8",X"14",X"64",X"08",
		X"05",X"38",X"38",X"28",X"08",X"C0",X"08",X"FF",X"04",X"06",X"30",X"30",X"14",X"0F",X"76",X"1D",
		X"19",X"18",X"17",X"1B",X"1F",X"76",X"67",X"6F",X"6E",X"62",X"45",X"80",X"46",X"80",X"47",X"80",
		X"48",X"80",X"49",X"00",X"48",X"00",X"47",X"00",X"46",X"00",X"45",X"40",X"46",X"40",X"47",X"40",
		X"48",X"40",X"49",X"C0",X"48",X"C0",X"47",X"C0",X"46",X"C0",X"5F",X"06",X"43",X"44",X"45",X"40",
		X"40",X"45",X"44",X"43",X"59",X"5A",X"FF",X"59",X"57",X"D9",X"57",X"D7",X"00",X"00",X"57",X"DA",
		X"57",X"D8",X"9E",X"AF",X"9F",X"92",X"00",X"00",X"9E",X"CB",X"A0",X"14",X"9B",X"B2",X"9B",X"FD",
		X"9C",X"9D",X"9C",X"58",X"9C",X"DC",X"9D",X"2E",X"E0",X"01",X"04",X"60",X"60",X"EF",X"FC",X"90",
		X"04",X"30",X"E0",X"EF",X"40",X"01",X"04",X"A0",X"FC",X"20",X"30",X"EF",X"F5",X"14",X"F5",X"1F",
		X"F5",X"2A",X"F5",X"35",X"05",X"00",X"01",X"08",X"01",X"F8",X"01",X"10",X"01",X"F0",X"01",X"05",
		X"00",X"11",X"FA",X"01",X"06",X"01",X"0C",X"11",X"F4",X"11",X"05",X"00",X"01",X"FA",X"11",X"06",
		X"11",X"F4",X"21",X"0C",X"21",X"05",X"00",X"11",X"F8",X"01",X"08",X"01",X"F8",X"21",X"08",X"21",
		X"01",X"01",X"00",X"00",X"01",X"08",X"00",X"00",X"01",X"10",X"00",X"00",X"01",X"08",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"08",X"00",X"00",X"01",X"10",
		X"00",X"00",X"01",X"08",X"00",X"00",X"01",X"01",X"FE",X"FF",X"00",X"00",X"FE",X"F8",X"00",X"00",
		X"FE",X"F0",X"00",X"00",X"FE",X"F8",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"FE",X"F8",X"00",X"00",X"FE",X"F0",X"00",X"00",X"FE",X"F8",X"00",X"00",X"FE",X"FF",
		X"80",X"FF",X"FF",X"80",X"00",X"FF",X"FF",X"00",X"A2",X"A4",X"A3",X"22",X"A3",X"A7",X"A4",X"24",
		X"A4",X"C2",X"A5",X"45",X"A1",X"E3",X"A5",X"19",X"A5",X"55",X"A5",X"2F",X"A5",X"35",X"01",X"01",
		X"01",X"01",X"01",X"01",X"00",X"FF",X"FE",X"01",X"01",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",
		X"0D",X"44",X"43",X"43",X"42",X"42",X"41",X"41",X"40",X"40",X"A3",X"7C",X"A3",X"8F",X"A3",X"7C",
		X"A3",X"9B",X"25",X"26",X"27",X"24",X"27",X"26",X"25",X"24",X"F5",X"EE",X"F5",X"FE",X"F6",X"0E",
		X"F6",X"1E",X"F6",X"2E",X"F6",X"3E",X"F6",X"2E",X"F6",X"1E",X"F6",X"0E",X"F5",X"FE",X"60",X"61",
		X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"69",X"6A",
		X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"72",X"73",
		X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"7B",X"7C",
		X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"84",X"85",
		X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"8D",X"8E",
		X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"94",X"93",X"92",X"91",X"90",X"8F",X"8E",X"96",X"97",
		X"98",X"97",X"4F",X"40",X"54",X"40",X"50",X"40",X"54",X"40",X"51",X"40",X"54",X"40",X"52",X"40",
		X"54",X"40",X"53",X"40",X"54",X"40",X"00",X"C0",X"40",X"80",X"3D",X"39",X"34",X"30",X"2C",X"28",
		X"25",X"22",X"20",X"1E",X"1C",X"1A",X"18",X"17",X"15",X"14",X"3E",X"39",X"35",X"31",X"2E",X"2A",
		X"27",X"25",X"22",X"20",X"1E",X"1C",X"1A",X"19",X"17",X"16",X"3E",X"3A",X"36",X"33",X"2F",X"2C",
		X"29",X"27",X"24",X"22",X"20",X"1E",X"1C",X"1B",X"19",X"18",X"3E",X"3B",X"37",X"34",X"31",X"2E",
		X"2B",X"28",X"26",X"24",X"22",X"20",X"1E",X"1D",X"1B",X"1A",X"3E",X"3B",X"38",X"35",X"32",X"2F",
		X"2C",X"2A",X"28",X"25",X"23",X"22",X"20",X"1E",X"1D",X"1C",X"3E",X"3B",X"38",X"36",X"33",X"30",
		X"2E",X"2B",X"29",X"27",X"25",X"23",X"21",X"20",X"1E",X"1D",X"3E",X"3C",X"39",X"36",X"34",X"31",
		X"2F",X"2C",X"2A",X"28",X"26",X"25",X"23",X"21",X"20",X"1E",X"3F",X"3C",X"39",X"37",X"34",X"32",
		X"30",X"2D",X"2B",X"29",X"28",X"26",X"24",X"23",X"21",X"20",X"20",X"0D",X"08",X"06",X"04",X"04",
		X"03",X"03",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"33",X"20",X"16",X"10",X"0D",X"0B",
		X"09",X"08",X"07",X"06",X"06",X"05",X"05",X"04",X"04",X"04",X"38",X"2A",X"20",X"19",X"15",X"11",
		X"0F",X"0D",X"0C",X"0A",X"09",X"09",X"08",X"07",X"07",X"06",X"3A",X"2F",X"27",X"20",X"1B",X"17",
		X"14",X"12",X"10",X"0E",X"0D",X"0C",X"0B",X"0A",X"0A",X"09",X"3B",X"33",X"2B",X"25",X"20",X"1C",
		X"19",X"16",X"14",X"12",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"3C",X"35",X"2E",X"29",X"24",X"20",
		X"1C",X"1A",X"17",X"15",X"14",X"12",X"11",X"10",X"0F",X"0E",X"3D",X"37",X"31",X"2C",X"27",X"23",
		X"20",X"1D",X"1A",X"18",X"16",X"15",X"13",X"12",X"11",X"10",X"3D",X"38",X"33",X"2E",X"2A",X"26",
		X"23",X"20",X"1D",X"1B",X"19",X"17",X"16",X"15",X"13",X"12",X"00",X"06",X"0C",X"12",X"19",X"1F",
		X"25",X"2B",X"31",X"38",X"3E",X"44",X"4A",X"50",X"56",X"5C",X"61",X"67",X"6D",X"73",X"78",X"7E",
		X"83",X"88",X"8E",X"93",X"98",X"9D",X"A2",X"A7",X"AB",X"B0",X"B5",X"B9",X"BD",X"C1",X"C5",X"C9",
		X"CD",X"D1",X"D4",X"D8",X"DB",X"DE",X"E1",X"E4",X"E7",X"EA",X"EC",X"EE",X"F1",X"F3",X"F4",X"F6",
		X"F8",X"F9",X"FB",X"FC",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"01",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FD",X"FC",X"FB",X"F9",X"F8",X"F6",X"F4",X"F3",X"F1",X"EE",X"EC",X"EA",X"E7",X"E4",X"E1",X"DE",
		X"DB",X"D8",X"D4",X"D1",X"CD",X"C9",X"C5",X"C1",X"BD",X"B9",X"B5",X"B0",X"AB",X"A7",X"A2",X"9D",
		X"98",X"93",X"8E",X"88",X"83",X"7E",X"78",X"73",X"6D",X"67",X"61",X"5C",X"56",X"50",X"4A",X"44",
		X"3E",X"38",X"31",X"2B",X"25",X"1F",X"19",X"12",X"0C",X"06",X"00",X"01",X"00",X"FF",X"00",X"A0",
		X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"99",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"03",
		X"28",X"01",X"58",X"04",X"70",X"02",X"D8",X"05",X"25",X"01",X"55",X"02",X"87",X"05",X"30",X"07",
		X"E0",X"02",X"6C",X"02",X"63",X"06",X"BE",X"07",X"88",X"06",X"C8",X"03",X"91",X"00",X"00",X"5A",
		X"59",X"58",X"57",X"56",X"3B",X"3C",X"3D",X"3C",X"38",X"39",X"3A",X"39",X"43",X"44",X"45",X"40",
		X"5A",X"59",X"58",X"57",X"56",X"05",X"1F",X"01",X"2F",X"1D",X"01",X"00",X"05",X"3F",X"01",X"2F",
		X"1D",X"00",X"00",X"02",X"67",X"05",X"30",X"1E",X"0A",X"00",X"06",X"7F",X"02",X"48",X"1F",X"00",
		X"00",X"01",X"8F",X"02",X"48",X"20",X"00",X"00",X"01",X"6F",X"02",X"48",X"20",X"01",X"00",X"03",
		X"4F",X"02",X"88",X"21",X"00",X"00",X"03",X"27",X"02",X"88",X"21",X"01",X"00",X"02",X"CF",X"03",
		X"18",X"22",X"00",X"00",X"02",X"CF",X"03",X"38",X"22",X"00",X"00",X"02",X"CF",X"03",X"58",X"22",
		X"00",X"00",X"02",X"BF",X"05",X"60",X"23",X"00",X"00",X"02",X"9F",X"05",X"60",X"23",X"00",X"00",
		X"07",X"17",X"05",X"50",X"23",X"0C",X"00",X"07",X"37",X"05",X"50",X"23",X"0C",X"00",X"02",X"CF",
		X"05",X"80",X"24",X"00",X"00",X"01",X"3F",X"06",X"08",X"25",X"00",X"00",X"02",X"67",X"01",X"28",
		X"26",X"00",X"00",X"02",X"67",X"01",X"48",X"26",X"00",X"00",X"02",X"CF",X"01",X"08",X"27",X"00",
		X"00",X"02",X"CF",X"01",X"38",X"27",X"01",X"00",X"01",X"FF",X"01",X"08",X"28",X"00",X"00",X"01",
		X"DF",X"01",X"08",X"28",X"00",X"00",X"01",X"BF",X"01",X"08",X"28",X"00",X"00",X"F9",X"29",X"F9",
		X"61",X"F9",X"99",X"F9",X"D1",X"FA",X"09",X"F8",X"F1",X"FA",X"09",X"F9",X"D1",X"F9",X"99",X"F9",
		X"61",X"03",X"C0",X"05",X"58",X"00",X"00",X"01",X"03",X"E0",X"05",X"58",X"00",X"00",X"01",X"04",
		X"00",X"05",X"58",X"00",X"00",X"01",X"04",X"20",X"05",X"58",X"00",X"00",X"01",X"03",X"D0",X"05",
		X"58",X"01",X"00",X"01",X"03",X"F0",X"05",X"58",X"01",X"00",X"01",X"04",X"10",X"05",X"58",X"01",
		X"00",X"01",X"04",X"30",X"05",X"58",X"01",X"00",X"01",X"06",X"FF",X"07",X"88",X"0A",X"00",X"01",
		X"07",X"1F",X"07",X"88",X"03",X"15",X"01",X"07",X"3F",X"07",X"88",X"04",X"15",X"01",X"07",X"5F",
		X"07",X"88",X"05",X"15",X"01",X"07",X"7F",X"07",X"88",X"06",X"15",X"01",X"07",X"9F",X"07",X"88",
		X"07",X"15",X"01",X"07",X"BF",X"07",X"88",X"08",X"15",X"01",X"07",X"DF",X"07",X"88",X"09",X"15",
		X"01",X"01",X"4F",X"03",X"C8",X"12",X"00",X"01",X"01",X"6F",X"03",X"E8",X"12",X"02",X"01",X"01",
		X"6F",X"04",X"48",X"12",X"03",X"01",X"01",X"4F",X"04",X"68",X"12",X"05",X"01",X"00",X"EF",X"04",
		X"68",X"12",X"06",X"01",X"00",X"CF",X"04",X"48",X"12",X"08",X"01",X"00",X"CF",X"03",X"E8",X"12",
		X"09",X"01",X"00",X"EF",X"03",X"C8",X"12",X"0B",X"01",X"00",X"27",X"07",X"00",X"13",X"03",X"01",
		X"00",X"47",X"07",X"20",X"14",X"03",X"01",X"00",X"67",X"07",X"40",X"15",X"03",X"01",X"00",X"87",
		X"07",X"60",X"16",X"04",X"01",X"00",X"37",X"07",X"10",X"17",X"04",X"01",X"00",X"57",X"07",X"30",
		X"18",X"03",X"01",X"00",X"77",X"07",X"50",X"19",X"03",X"01",X"00",X"97",X"07",X"70",X"1A",X"03",
		X"01",X"04",X"77",X"03",X"F8",X"1B",X"00",X"01",X"04",X"67",X"03",X"D8",X"1B",X"02",X"01",X"04",
		X"67",X"03",X"B8",X"1B",X"03",X"01",X"04",X"67",X"03",X"98",X"1B",X"04",X"01",X"04",X"47",X"03",
		X"78",X"1B",X"05",X"01",X"04",X"27",X"03",X"70",X"1B",X"07",X"01",X"04",X"07",X"03",X"88",X"1B",
		X"09",X"01",X"03",X"FF",X"03",X"A8",X"1B",X"0B",X"01",X"05",X"6F",X"04",X"C0",X"1C",X"08",X"01",
		X"05",X"4F",X"04",X"C8",X"1C",X"07",X"01",X"05",X"2F",X"04",X"D0",X"1C",X"06",X"01",X"05",X"0F",
		X"04",X"D8",X"1C",X"05",X"01",X"04",X"EF",X"04",X"E0",X"1C",X"04",X"01",X"04",X"CF",X"04",X"E8",
		X"1C",X"03",X"01",X"04",X"AF",X"04",X"F0",X"1C",X"02",X"01",X"04",X"8F",X"04",X"F8",X"1C",X"01",
		X"01",X"FA",X"93",X"FA",X"9D",X"FA",X"AE",X"FA",X"AD",X"FA",X"AC",X"FA",X"AB",X"FA",X"AA",X"FA",
		X"A9",X"FA",X"A8",X"FA",X"A7",X"FA",X"C4",X"FA",X"C5",X"FA",X"C6",X"FA",X"C7",X"FA",X"C8",X"FA",
		X"C9",X"FA",X"CA",X"FA",X"CB",X"FA",X"DB",X"FA",X"E8",X"FA",X"EC",X"FA",X"F0",X"FA",X"F4",X"FA",
		X"F9",X"FA",X"FE",X"FB",X"02",X"FB",X"06",X"FB",X"0A",X"FB",X"1F",X"FB",X"2F",X"FB",X"39",X"FB",
		X"44",X"FB",X"4F",X"FB",X"58",X"FB",X"3B",X"FB",X"68",X"FB",X"75",X"FB",X"82",X"FB",X"3E",X"FB",
		X"8B",X"FB",X"6C",X"41",X"1D",X"32",X"1D",X"42",X"1D",X"32",X"1D",X"41",X"FE",X"31",X"1D",X"42",
		X"1D",X"32",X"1D",X"42",X"1D",X"31",X"FE",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"2C",
		X"2C",X"24",X"0E",X"2C",X"2C",X"2A",X"0E",X"2C",X"2C",X"26",X"0E",X"28",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"FD",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"1C",X"1C",X"14",X"0E",
		X"1C",X"1C",X"1A",X"0E",X"1C",X"1C",X"16",X"0E",X"1C",X"1A",X"FC",X"14",X"44",X"4C",X"44",X"24",
		X"2C",X"24",X"34",X"3C",X"34",X"14",X"1C",X"FF",X"0D",X"14",X"01",X"FE",X"09",X"18",X"01",X"FE",
		X"05",X"1C",X"01",X"FE",X"01",X"1F",X"11",X"01",X"FE",X"01",X"2F",X"21",X"01",X"FE",X"05",X"2C",
		X"01",X"FE",X"09",X"28",X"01",X"FE",X"0D",X"24",X"01",X"FE",X"62",X"32",X"34",X"34",X"64",X"61",
		X"23",X"21",X"83",X"81",X"43",X"41",X"74",X"1F",X"13",X"74",X"43",X"83",X"23",X"65",X"FF",X"01",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"74",X"58",X"74",X"57",X"72",X"01",X"FE",X"24",
		X"24",X"81",X"47",X"72",X"17",X"51",X"38",X"61",X"FF",X"01",X"46",X"01",X"47",X"4F",X"01",X"47",
		X"4F",X"4F",X"01",X"FE",X"02",X"1F",X"1F",X"14",X"02",X"48",X"02",X"1F",X"1F",X"02",X"FE",X"24",
		X"2F",X"2D",X"48",X"1F",X"1F",X"12",X"38",X"FF",X"25",X"2A",X"2F",X"2A",X"01",X"4F",X"41",X"01",
		X"1F",X"1F",X"1A",X"01",X"3F",X"31",X"01",X"FF",X"01",X"23",X"2F",X"2F",X"01",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"25",X"01",X"FE",X"01",X"4F",X"42",X"02",X"2F",X"2F",X"2F",X"23",X"02",X"3F",X"32",
		X"01",X"FE",X"01",X"2F",X"2F",X"2F",X"29",X"02",X"44",X"01",X"FE",X"46",X"4E",X"1F",X"15",X"3F",
		X"35",X"2F",X"25",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"FF",X"80",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"00",X"00",X"00",X"80",X"00",X"80",X"FF",X"80",X"FF",X"80",X"FF",X"80",
		X"00",X"80",X"00",X"80",X"FF",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"FF",X"80",X"FF",X"80",X"00",X"80",
		X"00",X"80",X"00",X"80",X"FF",X"80",X"FF",X"80",X"00",X"80",X"FF",X"80",X"00",X"01",X"02",X"03",
		X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"0F",X"0E",X"0D",
		X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"80",X"00",X"00",
		X"C0",X"A0",X"E0",X"00",X"40",X"60",X"20",X"FC",X"51",X"FC",X"4D",X"FC",X"49",X"FC",X"45",X"FC",
		X"41",X"FC",X"3D",X"FC",X"39",X"FC",X"35",X"FC",X"31",X"FC",X"2D",X"FC",X"29",X"FC",X"25",X"FC",
		X"21",X"E1",X"E2",X"E3",X"E4",X"DD",X"DE",X"DF",X"E0",X"D9",X"DA",X"DB",X"DC",X"D5",X"D6",X"D7",
		X"D8",X"D1",X"D2",X"D3",X"D4",X"CD",X"CE",X"CF",X"D0",X"C9",X"CA",X"CB",X"CC",X"C5",X"C6",X"C7",
		X"C8",X"C1",X"C2",X"C3",X"C4",X"BD",X"BE",X"BF",X"C0",X"B9",X"BA",X"BB",X"BC",X"B5",X"B6",X"B7",
		X"B8",X"FF",X"FF",X"FF",X"FF",X"13",X"C5",X"12",X"C5",X"11",X"C5",X"13",X"C4",X"12",X"C4",X"11",
		X"C4",X"13",X"C3",X"12",X"C3",X"11",X"83",X"12",X"83",X"13",X"83",X"11",X"84",X"12",X"84",X"13",
		X"84",X"11",X"85",X"12",X"85",X"13",X"05",X"12",X"05",X"11",X"05",X"13",X"04",X"12",X"04",X"11",
		X"04",X"13",X"03",X"12",X"03",X"11",X"43",X"12",X"43",X"13",X"43",X"11",X"44",X"12",X"44",X"13",
		X"44",X"11",X"45",X"12",X"45",X"01",X"01",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"00",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"14",X"80",X"15",X"80",X"16",X"80",X"17",X"80",X"18",X"00",X"17",
		X"00",X"16",X"00",X"15",X"00",X"14",X"40",X"15",X"40",X"16",X"40",X"17",X"40",X"18",X"C0",X"17",
		X"C0",X"16",X"C0",X"15",X"C0",X"19",X"80",X"1A",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"00",X"1C",
		X"00",X"1B",X"00",X"1A",X"00",X"19",X"40",X"1A",X"40",X"1B",X"40",X"1C",X"40",X"1D",X"C0",X"1C",
		X"C0",X"1B",X"C0",X"1A",X"C0",X"04",X"0C",X"04",X"0A",X"06",X"0A",X"06",X"08",X"08",X"08",X"08",
		X"06",X"0A",X"06",X"0A",X"04",X"0C",X"04",X"0A",X"04",X"0A",X"06",X"08",X"06",X"08",X"08",X"06",
		X"08",X"06",X"0A",X"04",X"0A",X"91",X"F2",X"92",X"32",X"92",X"26",X"91",X"FA",X"91",X"FE",X"92",
		X"02",X"92",X"06",X"92",X"0E",X"92",X"16",X"92",X"1A",X"92",X"1E",X"92",X"22",X"92",X"3E",X"92",
		X"42",X"92",X"46",X"92",X"4A",X"92",X"58",X"92",X"5D",X"92",X"67",X"92",X"6C",X"92",X"71",X"92",
		X"12",X"92",X"7B",X"92",X"0A",X"92",X"80",X"92",X"8A",X"92",X"8F",X"92",X"94",X"B3",X"02",X"B3",
		X"1F",X"B3",X"28",X"B3",X"49",X"B3",X"58",X"B3",X"F2",X"B4",X"2A",X"B4",X"69",X"B5",X"55",X"B3",
		X"57",X"B3",X"F1",X"B3",X"FE",X"B4",X"38",X"B4",X"80",X"B5",X"80",X"0F",X"00",X"0A",X"0B",X"0C",
		X"0D",X"0E",X"0F",X"00",X"01",X"02",X"06",X"0A",X"0E",X"0C",X"0D",X"5D",X"A0",X"00",X"2D",X"C3",
		X"51",X"E5",X"00",X"70",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"9E",X"81",X"9E",X"81",X"9E",X"81",X"9E",X"81",X"9E",X"81",X"9E",X"81",X"9E",X"B6",X"6A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
