library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_1 is
	type rom is array(0 to  7167) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",
		X"00",X"00",X"40",X"42",X"7F",X"7F",X"40",X"40",X"00",X"62",X"73",X"79",X"59",X"5D",X"4F",X"46",
		X"00",X"20",X"61",X"49",X"4D",X"4F",X"7B",X"31",X"00",X"18",X"1C",X"16",X"13",X"7F",X"7F",X"10",
		X"00",X"27",X"67",X"45",X"45",X"45",X"7D",X"38",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",
		X"00",X"03",X"03",X"71",X"79",X"0D",X"07",X"03",X"00",X"36",X"4F",X"4D",X"59",X"59",X"76",X"30",
		X"00",X"06",X"4F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"7C",X"7E",X"13",X"11",X"13",X"7E",X"7C",
		X"00",X"7F",X"7F",X"49",X"49",X"49",X"7F",X"36",X"00",X"1C",X"3E",X"63",X"41",X"41",X"63",X"22",
		X"00",X"7F",X"7F",X"41",X"41",X"63",X"3E",X"1C",X"00",X"00",X"7F",X"7F",X"49",X"49",X"49",X"41",
		X"00",X"7F",X"7F",X"09",X"09",X"09",X"09",X"01",X"00",X"1C",X"3E",X"63",X"41",X"49",X"79",X"79",
		X"00",X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"41",X"7F",X"7F",X"41",X"41",
		X"00",X"20",X"60",X"40",X"40",X"40",X"7F",X"3F",X"00",X"7F",X"7F",X"18",X"3C",X"76",X"63",X"41",
		X"00",X"00",X"7F",X"7F",X"40",X"40",X"40",X"40",X"00",X"7F",X"7F",X"0E",X"1C",X"0E",X"7F",X"7F",
		X"00",X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",
		X"00",X"7F",X"7F",X"11",X"11",X"11",X"1F",X"0E",X"00",X"3E",X"7F",X"41",X"51",X"71",X"3F",X"5E",
		X"00",X"7F",X"7F",X"11",X"31",X"79",X"6F",X"4E",X"00",X"26",X"6F",X"49",X"49",X"4B",X"7A",X"30",
		X"00",X"00",X"01",X"01",X"7F",X"7F",X"01",X"01",X"00",X"3F",X"7F",X"40",X"40",X"40",X"7F",X"3F",
		X"00",X"0F",X"1F",X"38",X"70",X"38",X"1F",X"0F",X"00",X"1F",X"7F",X"38",X"1C",X"38",X"7F",X"1F",
		X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"00",X"03",X"0F",X"78",X"78",X"0F",X"03",
		X"00",X"61",X"71",X"79",X"5D",X"4F",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"12",X"1E",X"00",X"7E",X"5A",X"5A",X"00",
		X"7E",X"12",X"1E",X"00",X"7E",X"12",X"1E",X"00",X"7E",X"5A",X"5A",X"00",X"7E",X"12",X"2E",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"7F",X"40",X"40",X"40",X"40",X"40",X"40",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"10",X"00",X"22",X"00",X"10",X"04",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"10",X"00",X"48",X"00",X"00",X"20",X"00",X"08",X"40",X"00",X"10",X"04",
		X"00",X"00",X"00",X"01",X"00",X"10",X"00",X"00",X"02",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"02",X"00",X"24",X"00",X"08",X"41",X"04",X"00",X"09",X"01",X"04",X"90",X"04",X"20",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"10",X"80",X"00",X"00",X"20",X"00",X"80",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"80",X"04",X"00",X"20",X"05",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"41",X"08",X"00",X"20",X"81",X"00",X"10",X"00",X"00",X"82",X"00",X"04",X"00",X"20",
		X"00",X"00",X"24",X"00",X"04",X"01",X"10",X"00",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"04",X"40",X"08",X"20",X"02",X"00",X"20",X"04",X"80",X"01",X"08",X"20",X"02",X"00",X"04",X"01",
		X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"10",X"00",X"04",X"00",X"01",X"00",X"04",X"00",X"00",X"09",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C6",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"92",X"F6",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DE",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DE",X"92",X"F2",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"DE",X"92",X"F2",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"50",X"60",X"F0",X"D4",X"5A",X"88",X"A8",X"50",X"A0",X"CC",X"70",X"78",X"40",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"04",X"06",X"04",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"6E",X"76",X"7F",X"5D",X"7F",X"77",X"7F",X"5E",X"76",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"CC",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"CC",X"F8",X"20",X"10",X"10",X"E0",
		X"30",X"79",X"77",X"EF",X"EF",X"DF",X"DF",X"DF",X"EF",X"EF",X"77",X"79",X"31",X"02",X"01",X"00",
		X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"10",X"5C",X"54",X"74",X"10",X"00",
		X"00",X"00",X"7C",X"20",X"7C",X"64",X"7C",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"00",X"03",X"1F",X"11",X"1B",X"11",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"80",X"70",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"80",X"60",X"60",X"00",X"00",X"00",
		X"00",X"0C",X"02",X"A2",X"12",X"12",X"0C",X"00",X"00",X"00",X"BE",X"00",X"00",X"BE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E6",X"B2",X"9E",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C6",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"9E",X"92",X"F2",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E6",X"B2",X"9E",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"24",X"FE",X"20",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"FE",X"92",X"F6",X"00",X"FE",X"82",X"FE",X"82",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"08",X"1D",X"1F",X"3F",X"3E",X"3E",X"0E",X"04",X"00",X"00",X"00",
		X"00",X"04",X"8C",X"9E",X"9C",X"9E",X"1F",X"1F",X"1F",X"1F",X"1B",X"97",X"86",X"46",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"08",X"1D",X"1F",X"3F",X"3E",X"3E",X"0E",X"04",X"00",X"00",X"00",
		X"00",X"00",X"10",X"0C",X"1C",X"9E",X"9F",X"9F",X"99",X"87",X"07",X"16",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"08",X"1A",X"1F",X"3F",X"3E",X"3E",X"0E",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"56",X"56",X"17",X"1B",X"1F",X"1F",X"1F",X"9F",X"86",X"46",X"00",X"00",
		X"00",X"00",X"00",X"03",X"3F",X"1F",X"11",X"1B",X"1B",X"11",X"1F",X"3F",X"01",X"00",X"00",X"00",
		X"00",X"06",X"03",X"13",X"9F",X"9E",X"94",X"1E",X"1E",X"24",X"2E",X"3F",X"0E",X"07",X"0E",X"0C",
		X"00",X"00",X"00",X"01",X"3F",X"1F",X"11",X"1B",X"1B",X"11",X"1F",X"3F",X"03",X"00",X"00",X"00",
		X"0C",X"0E",X"07",X"0B",X"3F",X"2E",X"24",X"1E",X"1E",X"94",X"9E",X"9F",X"13",X"03",X"06",X"00",
		X"00",X"00",X"00",X"01",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"03",X"00",X"00",X"00",
		X"0C",X"0E",X"07",X"2B",X"2F",X"2F",X"1F",X"1F",X"1F",X"9F",X"9F",X"9F",X"1B",X"07",X"0E",X"00",
		X"00",X"00",X"00",X"03",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"01",X"00",X"00",X"00",
		X"00",X"0E",X"07",X"1B",X"9F",X"9F",X"9F",X"1F",X"1F",X"1F",X"2F",X"2F",X"2B",X"07",X"0E",X"0C",
		X"00",X"00",X"00",X"03",X"3F",X"1F",X"11",X"1B",X"1B",X"11",X"1F",X"3F",X"03",X"00",X"00",X"00",
		X"0C",X"0E",X"07",X"1B",X"9F",X"9E",X"94",X"1E",X"1E",X"94",X"9E",X"9F",X"1B",X"07",X"0E",X"0C",
		X"00",X"00",X"00",X"03",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"03",X"00",X"00",X"00",
		X"0C",X"0E",X"07",X"1B",X"9F",X"9F",X"9F",X"1F",X"1F",X"9F",X"9F",X"9F",X"1B",X"07",X"0E",X"0C",
		X"00",X"00",X"80",X"80",X"10",X"08",X"1D",X"1F",X"3F",X"3E",X"3E",X"0E",X"04",X"00",X"00",X"00",
		X"00",X"00",X"11",X"0F",X"1C",X"9E",X"9F",X"9F",X"99",X"87",X"47",X"76",X"18",X"00",X"00",X"00",
		X"00",X"00",X"80",X"03",X"3F",X"1F",X"11",X"1B",X"1B",X"11",X"1F",X"3F",X"03",X"00",X"00",X"00",
		X"00",X"01",X"03",X"1F",X"9F",X"9E",X"94",X"1E",X"1E",X"14",X"5E",X"7F",X"1B",X"07",X"0E",X"0C",
		X"00",X"80",X"C0",X"83",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"03",X"00",X"00",X"00",
		X"00",X"00",X"03",X"1F",X"9F",X"9F",X"9F",X"1F",X"1F",X"1F",X"DF",X"DF",X"1B",X"07",X"0E",X"0C",
		X"C0",X"C0",X"80",X"83",X"3F",X"1F",X"11",X"1B",X"1B",X"11",X"1F",X"3F",X"83",X"80",X"C0",X"C0",
		X"00",X"01",X"03",X"0F",X"8F",X"8F",X"8A",X"0F",X"0F",X"8A",X"8F",X"8F",X"0F",X"03",X"01",X"00",
		X"C0",X"C0",X"80",X"83",X"3F",X"1F",X"11",X"1B",X"1B",X"11",X"1F",X"3F",X"83",X"80",X"C0",X"C0",
		X"00",X"01",X"03",X"0F",X"8F",X"8F",X"8A",X"0F",X"0F",X"8A",X"8F",X"8F",X"0F",X"03",X"01",X"00",
		X"00",X"F0",X"E0",X"80",X"01",X"02",X"00",X"03",X"00",X"00",X"02",X"01",X"80",X"E0",X"F0",X"00",
		X"00",X"01",X"03",X"0F",X"8F",X"8F",X"8A",X"0F",X"0F",X"8A",X"8F",X"8F",X"0F",X"03",X"01",X"00",
		X"60",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"80",X"80",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"60",
		X"00",X"00",X"01",X"01",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"01",X"01",X"00",X"00",
		X"80",X"C0",X"0C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0C",X"C0",X"C0",X"80",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"00",X"30",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"30",X"00",X"00",X"00",
		X"04",X"0C",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"0C",X"04",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",
		X"08",X"0C",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"10",X"10",X"10",X"08",X"04",X"00",X"00",X"40",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"84",X"88",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"40",X"00",X"01",X"04",X"08",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"04",X"10",X"10",X"00",X"00",X"00",X"00",X"40",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"04",X"01",X"00",X"40",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"40",X"50",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"80",
		X"00",X"00",X"00",X"80",X"80",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"01",X"02",X"20",X"40",X"40",X"00",X"00",X"00",X"01",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"90",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"28",X"00",X"14",X"40",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"80",X"80",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",
		X"00",X"00",X"48",X"00",X"08",X"20",X"0B",X"10",X"49",X"02",X"14",X"80",X"00",X"12",X"00",X"40",
		X"82",X"80",X"80",X"80",X"02",X"00",X"03",X"00",X"00",X"01",X"00",X"00",X"80",X"80",X"80",X"80",
		X"E0",X"F0",X"FC",X"FE",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",
		X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",
		X"C0",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"E0",X"F8",X"FC",X"FE",X"FE",X"F3",X"FF",X"FF",X"FF",X"FF",X"F3",X"FE",X"FE",X"FC",X"F8",X"E0",
		X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",
		X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",
		X"07",X"1F",X"3F",X"7E",X"7E",X"FA",X"FC",X"FF",X"FF",X"FC",X"FA",X"7E",X"7E",X"3F",X"1F",X"07",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"18",X"3E",X"7F",X"7B",X"FB",X"FB",X"F7",X"FF",X"FF",X"F7",X"FB",X"FB",X"7B",X"7F",X"3E",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"70",X"70",X"D8",X"D8",X"E8",X"E8",X"F8",X"F8",X"E8",X"E8",X"D8",X"D8",X"70",X"70",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"88",X"00",X"A0",X"80",X"A0",X"00",X"88",X"80",X"A0",X"A0",X"88",X"00",X"A0",X"48",
		X"00",X"80",X"E0",X"F0",X"F0",X"78",X"F8",X"F8",X"F8",X"F8",X"78",X"F0",X"F0",X"E0",X"80",X"00",
		X"00",X"07",X"1F",X"3F",X"3E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3E",X"3F",X"1F",X"07",X"00",
		X"25",X"E0",X"FC",X"FD",X"AC",X"1E",X"BE",X"FE",X"FE",X"BE",X"1E",X"AC",X"FD",X"F8",X"E2",X"01",
		X"10",X"01",X"07",X"2F",X"0E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0E",X"0F",X"07",X"09",X"00",
		X"C0",X"F0",X"7C",X"3E",X"3F",X"3F",X"7F",X"FF",X"FF",X"FE",X"FC",X"F0",X"E0",X"C0",X"80",X"80",
		X"07",X"18",X"10",X"20",X"28",X"A8",X"B6",X"F8",X"FF",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"03",
		X"C0",X"60",X"20",X"10",X"18",X"1C",X"3E",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"C0",
		X"03",X"84",X"98",X"B0",X"70",X"34",X"3B",X"3C",X"3F",X"3F",X"7F",X"5F",X"DF",X"1F",X"0F",X"03",
		X"80",X"C0",X"F0",X"FC",X"FE",X"7F",X"BF",X"BF",X"3F",X"3F",X"7F",X"FE",X"F0",X"E0",X"C0",X"00",
		X"03",X"07",X"1F",X"1F",X"38",X"F3",X"60",X"20",X"20",X"20",X"70",X"38",X"3F",X"1F",X"0F",X"07",
		X"C0",X"E0",X"F8",X"FC",X"7E",X"BE",X"5F",X"5F",X"1E",X"1E",X"3C",X"7C",X"F8",X"E0",X"C0",X"80",
		X"03",X"0F",X"0F",X"1F",X"3C",X"79",X"30",X"30",X"30",X"70",X"F8",X"3C",X"1F",X"07",X"03",X"01",
		X"80",X"C0",X"F0",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"FA",X"F9",X"FC",X"F0",X"E0",X"C0",X"00",
		X"03",X"07",X"1F",X"1F",X"3F",X"FF",X"7F",X"3F",X"3F",X"3F",X"7F",X"3F",X"3F",X"1F",X"0F",X"07",
		X"C0",X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"E0",X"C0",X"80",
		X"03",X"0F",X"0F",X"1F",X"3F",X"7F",X"3F",X"3F",X"3F",X"7F",X"FF",X"3F",X"1F",X"07",X"03",X"01",
		X"00",X"80",X"E0",X"F0",X"F0",X"78",X"38",X"38",X"38",X"38",X"78",X"F0",X"E0",X"C0",X"00",X"00",
		X"8E",X"9F",X"7F",X"7F",X"F8",X"F0",X"E0",X"E8",X"E8",X"E4",X"F0",X"F8",X"FF",X"7F",X"BF",X"9C",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"8C",X"9E",X"7F",X"7F",X"F8",X"F0",X"E0",X"E8",X"E8",X"E4",X"F0",X"F8",X"7F",X"7E",X"9C",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"88",X"80",X"80",X"92",X"80",X"08",X"40",X"84",X"88",X"80",X"20",X"84",X"80",X"40",X"40",
		X"00",X"00",X"C0",X"A0",X"F8",X"E8",X"7C",X"F8",X"FC",X"E8",X"F8",X"F0",X"40",X"80",X"00",X"00",
		X"8E",X"9F",X"7F",X"7F",X"E3",X"C1",X"91",X"90",X"BC",X"90",X"C1",X"E3",X"FF",X"7F",X"BF",X"9C",
		X"89",X"C0",X"64",X"DA",X"7C",X"3C",X"96",X"1E",X"9F",X"1B",X"3E",X"7A",X"DE",X"F8",X"60",X"CA",
		X"05",X"23",X"07",X"9F",X"FC",X"38",X"32",X"31",X"32",X"30",X"38",X"FC",X"9B",X"0F",X"2F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"C0",X"C0",X"E4",X"C0",X"C8",X"E2",X"C0",X"C8",X"E2",X"C0",X"C0",X"EA",X"C0",
		X"C0",X"EA",X"C0",X"C0",X"E2",X"C8",X"C0",X"E2",X"C8",X"C0",X"E4",X"C0",X"C0",X"E0",X"C0",X"00",
		X"80",X"80",X"C0",X"80",X"80",X"C8",X"80",X"90",X"C4",X"80",X"90",X"C4",X"80",X"80",X"D4",X"80",
		X"80",X"D4",X"80",X"80",X"C4",X"90",X"80",X"C4",X"90",X"80",X"C8",X"80",X"80",X"C0",X"80",X"00",
		X"00",X"00",X"80",X"00",X"00",X"90",X"00",X"20",X"88",X"00",X"20",X"88",X"00",X"00",X"A8",X"00",
		X"00",X"A8",X"00",X"00",X"88",X"20",X"00",X"88",X"20",X"00",X"90",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"40",X"10",X"00",X"40",X"10",X"00",X"00",X"50",X"00",
		X"00",X"50",X"00",X"00",X"10",X"40",X"00",X"10",X"40",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"20",X"00",X"80",X"20",X"00",X"00",X"A0",X"00",
		X"00",X"A0",X"00",X"00",X"20",X"80",X"00",X"20",X"80",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"40",X"00",
		X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"80",X"00",
		X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"06",X"06",X"07",X"06",X"06",X"07",X"06",X"06",X"07",X"06",X"06",X"07",X"06",X"06",X"07",X"06",
		X"06",X"07",X"06",X"06",X"07",X"06",X"06",X"07",X"06",X"06",X"07",X"06",X"06",X"07",X"06",X"00",
		X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",
		X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"0C",X"0E",X"0C",X"00",
		X"18",X"18",X"1C",X"18",X"18",X"1C",X"18",X"19",X"1C",X"18",X"19",X"1C",X"18",X"18",X"1D",X"18",
		X"18",X"1D",X"18",X"18",X"1C",X"19",X"18",X"1C",X"19",X"18",X"1C",X"18",X"18",X"1C",X"18",X"00",
		X"30",X"30",X"38",X"30",X"30",X"39",X"30",X"32",X"38",X"30",X"32",X"38",X"30",X"30",X"3A",X"30",
		X"30",X"3A",X"30",X"30",X"38",X"32",X"30",X"38",X"32",X"30",X"39",X"30",X"30",X"38",X"30",X"00",
		X"60",X"60",X"70",X"60",X"60",X"72",X"60",X"64",X"71",X"60",X"64",X"71",X"60",X"60",X"75",X"60",
		X"60",X"75",X"60",X"60",X"71",X"64",X"60",X"71",X"64",X"60",X"72",X"60",X"60",X"70",X"60",X"00",
		X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",
		X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"0E",X"06",X"00",
		X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",
		X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"1C",X"0C",X"00",
		X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",
		X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"38",X"18",X"00",
		X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",
		X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"70",X"30",X"00",
		X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",
		X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"E0",X"60",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",
		X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",
		X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"00",
		X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",
		X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",X"00",
		X"00",X"00",X"78",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"78",X"00",X"00",
		X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",
		X"00",X"00",X"1E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1E",X"00",X"00",
		X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"62",X"40",X"42",X"02",X"42",X"06",X"02",X"02",X"06",X"06",X"02",X"06",
		X"06",X"06",X"06",X"02",X"06",X"02",X"02",X"02",X"06",X"00",X"02",X"40",X"02",X"38",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C4",X"80",X"84",X"04",X"84",X"0C",X"04",X"04",X"0C",X"0C",X"04",X"0C",
		X"0C",X"0C",X"0C",X"04",X"0C",X"04",X"04",X"04",X"0C",X"00",X"04",X"80",X"04",X"70",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"88",X"00",X"08",X"08",X"08",X"18",X"08",X"08",X"18",X"18",X"08",X"18",
		X"18",X"18",X"18",X"08",X"18",X"08",X"08",X"08",X"18",X"00",X"08",X"00",X"08",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"80",X"10",X"00",X"10",X"10",X"10",X"30",X"10",X"10",X"30",X"30",X"10",X"30",
		X"30",X"30",X"30",X"10",X"30",X"10",X"10",X"10",X"30",X"00",X"10",X"00",X"10",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"20",X"20",X"60",X"20",X"20",X"60",X"60",X"20",X"60",
		X"60",X"60",X"60",X"20",X"60",X"20",X"20",X"20",X"60",X"00",X"20",X"00",X"20",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"40",X"40",X"C0",X"40",X"40",X"C0",X"C0",X"40",X"C0",
		X"C0",X"C0",X"C0",X"40",X"C0",X"40",X"40",X"40",X"C0",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"07",X"06",X"04",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"0C",X"08",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"18",X"10",X"10",X"00",X"10",X"01",X"00",X"00",X"01",X"01",X"00",X"01",
		X"01",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"10",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"38",X"31",X"20",X"21",X"01",X"21",X"03",X"01",X"01",X"03",X"03",X"01",X"03",
		X"03",X"03",X"03",X"01",X"03",X"01",X"01",X"01",X"03",X"00",X"01",X"20",X"01",X"1C",X"00",X"00",
		X"D0",X"78",X"BC",X"FE",X"74",X"7A",X"FC",X"F8",X"7C",X"FA",X"FE",X"7C",X"3A",X"7C",X"F4",X"FE",
		X"FE",X"F4",X"7C",X"3A",X"7C",X"FE",X"FA",X"7C",X"F8",X"FC",X"7A",X"74",X"FE",X"BC",X"78",X"00",
		X"A0",X"F0",X"78",X"FC",X"E8",X"F4",X"F8",X"F0",X"F8",X"F4",X"FC",X"F8",X"74",X"F8",X"E8",X"FC",
		X"FC",X"E8",X"F8",X"74",X"F8",X"FC",X"F4",X"F8",X"F0",X"F8",X"F4",X"E8",X"FC",X"78",X"F0",X"00",
		X"40",X"E0",X"F0",X"F8",X"D0",X"E8",X"F0",X"E0",X"F0",X"E8",X"F8",X"F0",X"E8",X"F0",X"D0",X"F8",
		X"F8",X"D0",X"F0",X"E8",X"F0",X"F8",X"E8",X"F0",X"E0",X"F0",X"E8",X"D0",X"F8",X"F0",X"E0",X"00",
		X"80",X"C0",X"E0",X"F0",X"A0",X"D0",X"E0",X"C0",X"E0",X"D0",X"F0",X"E0",X"D0",X"E0",X"A0",X"F0",
		X"F0",X"A0",X"E0",X"D0",X"E0",X"F0",X"D0",X"E0",X"C0",X"E0",X"D0",X"A0",X"F0",X"E0",X"C0",X"00",
		X"00",X"80",X"C0",X"E0",X"40",X"A0",X"C0",X"80",X"C0",X"A0",X"E0",X"C0",X"A0",X"C0",X"40",X"E0",
		X"E0",X"40",X"C0",X"A0",X"C0",X"E0",X"A0",X"C0",X"80",X"C0",X"A0",X"40",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"80",X"C0",X"80",X"40",X"80",X"00",X"80",X"40",X"C0",X"80",X"40",X"80",X"80",X"C0",
		X"C0",X"80",X"80",X"40",X"80",X"C0",X"40",X"80",X"00",X"80",X"40",X"80",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"80",X"00",X"00",X"80",
		X"80",X"00",X"00",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"03",X"01",X"02",X"03",X"01",X"01",X"03",X"03",X"01",X"03",X"03",X"01",X"00",X"01",X"03",X"03",
		X"03",X"03",X"01",X"00",X"01",X"03",X"03",X"01",X"03",X"03",X"01",X"01",X"03",X"02",X"01",X"00",
		X"06",X"03",X"05",X"07",X"03",X"03",X"07",X"07",X"03",X"07",X"07",X"03",X"01",X"03",X"07",X"07",
		X"07",X"07",X"03",X"01",X"03",X"07",X"07",X"03",X"07",X"07",X"03",X"03",X"07",X"05",X"03",X"00",
		X"0D",X"07",X"0B",X"0F",X"07",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",
		X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"07",X"07",X"0F",X"0B",X"07",X"00",
		X"1A",X"0F",X"17",X"1F",X"0E",X"0F",X"1F",X"1F",X"0F",X"1F",X"1F",X"0F",X"07",X"0F",X"1E",X"1F",
		X"1F",X"1E",X"0F",X"07",X"0F",X"1F",X"1F",X"0F",X"1F",X"1F",X"0F",X"0E",X"1F",X"17",X"0F",X"00",
		X"34",X"1E",X"2F",X"3F",X"1D",X"1E",X"3F",X"3E",X"1F",X"3E",X"3F",X"1F",X"0E",X"1F",X"3D",X"3F",
		X"3F",X"3D",X"1F",X"0E",X"1F",X"3F",X"3E",X"1F",X"3E",X"3F",X"1E",X"1D",X"3F",X"2F",X"1E",X"00",
		X"68",X"3C",X"5E",X"7F",X"3A",X"3D",X"7E",X"7C",X"3E",X"7D",X"7F",X"3E",X"1D",X"3E",X"7A",X"7F",
		X"7F",X"7A",X"3E",X"1D",X"3E",X"7F",X"7D",X"3E",X"7C",X"7E",X"3D",X"3A",X"7F",X"5E",X"3C",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
