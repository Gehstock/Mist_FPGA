library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity satans_hollow_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of satans_hollow_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"FE",X"01",X"7F",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"5F",X"05",X"7F",X"05",X"FF",X"57",X"FE",
		X"A3",X"FF",X"F3",X"FC",X"C0",X"03",X"07",X"FF",X"17",X"FF",X"05",X"7D",X"00",X"5F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"F3",X"FF",X"F3",X"AB",X"A3",X"AB",
		X"FC",X"17",X"F1",X"7F",X"FC",X"17",X"FF",X"F1",X"FE",X"AC",X"7F",X"FF",X"D5",X"55",X"3F",X"FF",
		X"00",X"03",X"03",X"FF",X"FF",X"FF",X"00",X"0F",X"EA",X"FF",X"EA",X"FF",X"FF",X"FC",X"FF",X"FD",
		X"3F",X"FA",X"0F",X"FE",X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"03",X"FF",X"3F",X"00",X"05",X"FF",X"17",X"AF",X"57",X"FF",X"05",X"7F",X"00",X"00",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"3F",X"FA",
		X"00",X"0F",X"FF",X"FA",X"FF",X"AA",X"FF",X"AA",X"55",X"AA",X"00",X"AA",X"FF",X"EA",X"FF",X"EA",
		X"F0",X"00",X"0F",X"FF",X"7E",X"FF",X"1F",X"FF",X"C5",X"55",X"30",X"00",X"0F",X"CF",X"FF",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"01",X"00",X"FC",X"FF",X"FC",
		X"FF",X"F3",X"FF",X"F0",X"FF",X"FC",X"FF",X"F0",X"00",X"F3",X"FF",X"F0",X"55",X"54",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"F3",X"FF",X"4F",X"FF",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FA",X"AA",X"EA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"00",X"FF",X"03",X"F0",X"0F",X"F0",X"0F",X"00",X"3F",X"00",X"FF",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"03",X"FF",X"00",X"FC",X"0F",X"00",
		X"00",X"3F",X"03",X"FC",X"0F",X"C0",X"0F",X"00",X"30",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",
		X"3F",X"FF",X"FF",X"FF",X"00",X"FF",X"03",X"FF",X"00",X"FF",X"F0",X"15",X"FD",X"55",X"F0",X"15",
		X"03",X"FF",X"00",X"15",X"C0",X"01",X"FC",X"00",X"FF",X"03",X"00",X"0F",X"00",X"FF",X"0F",X"FF",
		X"FF",X"D5",X"0F",X"D5",X"00",X"05",X"00",X"00",X"00",X"0F",X"00",X"05",X"00",X"15",X"00",X"FF",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"30",X"3F",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"03",X"00",X"FF",X"00",X"0C",
		X"55",X"4F",X"55",X"F0",X"FD",X"5C",X"FF",X"FF",X"0F",X"F0",X"0F",X"05",X"00",X"FF",X"01",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"50",X"FF",X"54",X"0F",
		X"FF",X"55",X"55",X"55",X"55",X"55",X"3F",X"F5",X"FF",X"57",X"FF",X"15",X"FF",X"C5",X"FF",X"F3",
		X"55",X"54",X"05",X"40",X"15",X"00",X"55",X"53",X"FF",X"FD",X"55",X"55",X"55",X"55",X"FF",X"D5",
		X"05",X"D5",X"F5",X"F5",X"F5",X"FD",X"F5",X"FD",X"F5",X"FF",X"D5",X"FF",X"55",X"7F",X"55",X"7D",
		X"00",X"13",X"00",X"4F",X"01",X"5F",X"55",X"5F",X"45",X"4F",X"15",X"3F",X"14",X"FD",X"11",X"F5",
		X"01",X"D5",X"00",X"75",X"00",X"5D",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",
		X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"55",X"00",X"57",X"00",X"1F",X"15",X"7F",X"05",X"FF",
		X"FC",X"55",X"3C",X"55",X"3C",X"55",X"3C",X"55",X"0D",X"55",X"05",X"55",X"05",X"55",X"15",X"55",
		X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FC",X"55",X"FC",X"55",X"FC",X"55",X"FC",X"55",X"FC",X"55",
		X"F1",X"55",X"F1",X"55",X"F1",X"55",X"F1",X"55",X"51",X"55",X"7C",X"55",X"7C",X"55",X"FC",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"3D",X"55",X"3D",X"55",X"3D",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"02",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"02",X"0A",X"AA",X"0A",X"AA",X"08",X"02",X"08",X"02",X"00",X"00",
		X"00",X"00",X"0A",X"82",X"0A",X"82",X"08",X"82",X"08",X"82",X"08",X"AA",X"08",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"82",X"08",X"82",X"08",X"82",X"08",X"82",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"00",X"20",X"00",X"20",X"02",X"A0",X"02",X"A0",X"00",X"00",
		X"00",X"00",X"08",X"AA",X"08",X"AA",X"08",X"82",X"08",X"82",X"08",X"82",X"0A",X"82",X"00",X"00",
		X"00",X"00",X"08",X"2A",X"08",X"2A",X"08",X"22",X"08",X"22",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"00",X"08",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"82",X"08",X"82",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"22",X"08",X"22",X"0A",X"A2",X"0A",X"A2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"20",X"08",X"20",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"0A",X"AA",X"0A",X"22",X"0A",X"22",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"08",X"02",X"08",X"02",X"08",X"02",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"02",X"A8",X"0A",X"AA",X"0A",X"0A",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"08",X"02",X"08",X"82",X"08",X"82",X"08",X"82",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"20",X"08",X"20",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"08",X"2A",X"08",X"2A",X"08",X"02",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"00",X"20",X"00",X"20",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"08",X"02",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"08",X"02",X"08",X"02",X"00",X"00",
		X"08",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"02",X"08",X"02",X"00",X"2A",X"00",X"2A",X"00",X"00",
		X"00",X"00",X"08",X"02",X"08",X"0A",X"0A",X"28",X"02",X"A0",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"08",X"00",X"0A",X"AA",X"08",X"00",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"00",X"A8",X"02",X"80",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"02",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"A0",X"0A",X"A0",X"08",X"20",X"08",X"20",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"08",X"0A",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"8A",X"0A",X"AA",X"08",X"A0",X"08",X"80",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"AA",X"08",X"AA",X"08",X"82",X"08",X"82",X"0A",X"82",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"08",X"02",X"0A",X"AA",X"0A",X"AA",X"08",X"02",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"00",X"02",X"00",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"08",X"00",X"0A",X"A0",X"00",X"2A",X"0A",X"AA",X"0A",X"A0",X"08",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"00",X"02",X"0A",X"AA",X"00",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"08",X"02",X"0A",X"2A",X"00",X"A0",X"0A",X"80",X"0A",X"20",X"08",X"0A",X"00",X"00",
		X"00",X"00",X"08",X"00",X"0A",X"00",X"00",X"AA",X"02",X"AA",X"0A",X"80",X"08",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"0A",X"02",X"0A",X"82",X"08",X"A2",X"08",X"2A",X"08",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3D",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"3D",X"55",X"3D",X"55",X"3D",X"55",X"3D",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",
		X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"01",
		X"00",X"00",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"2A",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"AF",X"FF",X"AF",X"FE",X"BF",X"FF",X"AF",X"F5",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"BF",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9A",X"4A",X"96",X"52",X"55",X"52",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"5A",X"AA",X"5A",X"AA",X"55",X"FF",X"55",X"AA",
		X"9A",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"95",X"AA",X"55",X"AA",X"55",X"AA",X"A5",X"AA",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"55",X"02",X"55",X"56",X"55",X"56",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"5A",X"AA",X"50",X"AA",X"55",X"2A",X"55",X"6A",X"55",X"40",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"99",X"69",X"AA",X"A9",X"95",X"9A",X"A9",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"56",X"AA",X"A6",
		X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"80",X"55",X"4A",X"55",X"4A",X"55",X"4A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"42",X"A9",X"50",X"A5",X"94",X"95",X"A4",X"95",X"A4",X"15",X"A5",X"05",X"A5",X"45",X"A9",X"45",
		X"A5",X"09",X"A9",X"45",X"A9",X"45",X"A9",X"41",X"A9",X"41",X"A9",X"51",X"AA",X"51",X"AA",X"51",
		X"AA",X"95",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",
		X"15",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"2A",X"14",X"2A",X"50",X"AA",
		X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"2A",
		X"55",X"10",X"55",X"04",X"55",X"05",X"55",X"45",X"55",X"41",X"55",X"49",X"55",X"49",X"55",X"49",
		X"54",X"AA",X"A5",X"0A",X"A5",X"4A",X"F5",X"4A",X"A5",X"4A",X"65",X"42",X"69",X"50",X"69",X"54",
		X"FF",X"D4",X"FF",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"FD",X"55",X"55",X"55",X"55",
		X"94",X"94",X"94",X"94",X"94",X"94",X"F5",X"14",X"A9",X"52",X"A9",X"52",X"A9",X"52",X"BD",X"0A",
		X"4A",X"A5",X"4A",X"A5",X"52",X"A5",X"52",X"95",X"52",X"95",X"52",X"94",X"52",X"92",X"52",X"92",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"95",X"25",X"95",X"29",X"55",X"2A",X"54",X"2A",X"50",X"AA",X"52",X"AA",X"52",X"AA",X"52",X"AA",
		X"A9",X"52",X"A9",X"42",X"A9",X"4A",X"A9",X"4A",X"A5",X"0A",X"A5",X"2A",X"95",X"2A",X"95",X"29",
		X"AA",X"52",X"AA",X"52",X"A9",X"50",X"A9",X"44",X"A9",X"44",X"A9",X"45",X"A9",X"45",X"A9",X"41",
		X"52",X"AA",X"54",X"AA",X"54",X"2A",X"55",X"2A",X"55",X"0A",X"55",X"4A",X"55",X"42",X"55",X"52",
		X"55",X"52",X"55",X"54",X"95",X"54",X"95",X"55",X"95",X"55",X"95",X"55",X"A5",X"55",X"A5",X"55",
		X"52",X"A9",X"52",X"A6",X"52",X"A6",X"52",X"99",X"50",X"A6",X"54",X"99",X"54",X"66",X"54",X"99",
		X"94",X"A6",X"94",X"29",X"95",X"26",X"95",X"09",X"95",X"4A",X"95",X"49",X"A5",X"42",X"A5",X"52",
		X"95",X"0A",X"A5",X"4A",X"A5",X"4A",X"A5",X"4A",X"A5",X"42",X"A9",X"52",X"A9",X"52",X"A9",X"52",
		X"AD",X"51",X"FD",X"51",X"FD",X"51",X"FD",X"54",X"FD",X"54",X"BD",X"50",X"FF",X"51",X"AB",X"45",
		X"A9",X"54",X"A5",X"54",X"A5",X"50",X"A5",X"52",X"A5",X"42",X"A5",X"49",X"95",X"05",X"55",X"2A",
		X"66",X"66",X"99",X"99",X"66",X"66",X"99",X"99",X"66",X"66",X"99",X"99",X"66",X"66",X"99",X"99",
		X"6E",X"54",X"9B",X"54",X"6E",X"54",X"99",X"54",X"ED",X"54",X"B9",X"54",X"AD",X"54",X"A9",X"54",
		X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"54",X"AA",X"54",X"AA",X"54",X"AA",X"54",X"AA",X"54",X"A9",X"50",X"A9",X"52",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"65",X"55",X"69",X"55",X"A9",X"55",X"A9",X"55",X"96",X"55",X"96",X"55",X"A9",X"55",X"95",X"A5",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"95",
		X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"95",X"A5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"9A",X"A9",X"5A",X"AA",X"AA",X"A6",X"AA",X"A6",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"AA",X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",X"6A",X"95",X"AA",X"6A",X"AA",X"AA",X"AA",
		X"A9",X"5A",X"AA",X"56",X"AA",X"95",X"AA",X"A5",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"56",X"55",X"5A",X"55",X"6A",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",
		X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"54",X"55",X"52",X"55",X"4A",X"55",X"0A",X"54",X"2A",X"54",X"AA",X"52",X"AA",X"42",X"AA",
		X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"D5",
		X"AA",X"82",X"A8",X"08",X"80",X"A0",X"2A",X"82",X"AA",X"28",X"80",X"AA",X"AA",X"AA",X"AA",X"0A",
		X"AA",X"8B",X"02",X"8F",X"22",X"8C",X"22",X"80",X"20",X"02",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"2A",X"A8",X"2A",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",
		X"AA",X"8A",X"AA",X"8A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",
		X"AF",X"FC",X"FF",X"02",X"F0",X"0A",X"00",X"AA",X"0A",X"AB",X"AA",X"AE",X"AA",X"FA",X"AB",X"AA",
		X"AA",X"FC",X"FF",X"02",X"C0",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"B0",
		X"54",X"00",X"14",X"2A",X"10",X"FF",X"13",X"FF",X"0F",X"C0",X"3C",X"00",X"00",X"AA",X"82",X"AA",
		X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"0A",
		X"55",X"55",X"55",X"54",X"55",X"40",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",X"55",X"4A",
		X"00",X"0F",X"FF",X"FA",X"FE",X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"00",X"00",X"2A",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"52",X"AA",X"52",X"AA",X"4A",X"AA",X"4A",X"AA",X"4A",X"AA",X"4A",X"AA",X"4A",X"AA",X"6A",X"AA",
		X"55",X"40",X"55",X"42",X"55",X"2A",X"55",X"2A",X"54",X"AA",X"54",X"AA",X"54",X"AA",X"54",X"FF",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"EA",X"AA",X"AA",
		X"2A",X"AF",X"2B",X"FF",X"3F",X"FF",X"3F",X"FC",X"3F",X"F0",X"30",X"00",X"00",X"00",X"80",X"2A",
		X"54",X"3F",X"54",X"00",X"54",X"00",X"54",X"2A",X"54",X"2A",X"54",X"2A",X"54",X"2A",X"50",X"AA",
		X"55",X"52",X"55",X"52",X"55",X"4A",X"55",X"4A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"03",X"C0",X"0F",X"C0",X"3F",X"C0",X"FF",X"C0",X"FF",X"FF",
		X"00",X"08",X"00",X"28",X"00",X"A8",X"02",X"A8",X"0A",X"A0",X"2A",X"A0",X"AA",X"80",X"FF",X"FF",
		X"FF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",
		X"FD",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D5",
		X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",
		X"55",X"55",X"55",X"55",X"59",X"AA",X"59",X"AA",X"59",X"96",X"59",X"96",X"5A",X"96",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"55",X"65",X"55",X"65",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"5A",X"55",X"6A",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",
		X"55",X"55",X"55",X"5A",X"55",X"5A",X"55",X"56",X"55",X"56",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"C0",X"00",X"00",X"03",
		X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"55",X"AA",X"55",X"A5",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"2A",X"82",X"8A",X"A0",X"82",X"A8",X"A0",X"2A",X"82",X"AA",X"8A",X"A8",X"2A",X"A0",X"AA",X"A8",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A8",X"AA",X"A2",X"AA",X"0A",X"80",X"A8",X"2A",X"A2",X"AA",X"A8",X"02",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"03",X"00",X"02",X"C0",X"02",X"C0",X"00",X"B0",X"00",X"2C",X"00",X"2C",X"00",X"0B",X"00",X"02",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"AA",X"A2",X"A0",X"2A",X"8A",X"A8",X"2A",X"A2",X"AA",X"8A",X"AA",X"2A",X"0A",X"AA",
		X"55",X"5F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"0A",X"B0",X"AB",X"00",X"C0",X"00",
		X"FC",X"3F",X"FC",X"F3",X"F3",X"C3",X"F3",X"03",X"F3",X"C3",X"F0",X"F3",X"F0",X"3F",X"F0",X"0F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F0",X"0F",X"F0",X"3F",X"F0",X"F3",X"F0",X"C3",X"F3",X"03",X"F3",X"C3",X"FC",X"33",X"FC",X"3F",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"59",X"56",X"59",X"56",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"56",X"5A",X"AA",X"5A",X"AA",X"59",X"56",X"59",X"56",X"55",X"55",
		X"55",X"55",X"5A",X"96",X"5A",X"96",X"59",X"96",X"59",X"96",X"59",X"AA",X"59",X"AA",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"59",X"96",X"59",X"96",X"59",X"96",X"59",X"96",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"55",X"65",X"55",X"65",X"56",X"A5",X"56",X"A5",X"55",X"55",
		X"55",X"55",X"59",X"AA",X"59",X"AA",X"59",X"96",X"59",X"96",X"59",X"96",X"5A",X"96",X"55",X"55",
		X"55",X"55",X"59",X"6A",X"59",X"6A",X"59",X"66",X"59",X"66",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"59",X"55",X"59",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"59",X"96",X"59",X"96",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"5A",X"AA",X"5A",X"AA",X"59",X"66",X"59",X"66",X"5A",X"A6",X"5A",X"A6",X"55",X"55",
		X"00",X"A0",X"02",X"A0",X"0A",X"E0",X"2B",X"E0",X"AF",X"E0",X"BF",X"E0",X"FF",X"EA",X"FF",X"FF",
		X"55",X"55",X"59",X"56",X"59",X"96",X"59",X"96",X"59",X"96",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"2A",X"A8",X"80",X"02",X"88",X"22",X"88",X"22",X"88",X"22",X"82",X"82",X"80",X"02",X"2A",X"A8",
		X"55",X"55",X"55",X"56",X"59",X"56",X"59",X"56",X"59",X"56",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"5A",X"9A",X"5A",X"AA",X"59",X"A5",X"59",X"95",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"56",X"A9",X"5A",X"AA",X"5A",X"5A",X"59",X"56",X"5A",X"AA",X"5A",X"AA",X"55",X"55",
		X"55",X"55",X"59",X"56",X"59",X"56",X"5A",X"AA",X"5A",X"AA",X"59",X"56",X"59",X"56",X"55",X"55",
		X"55",X"55",X"5A",X"55",X"59",X"56",X"5A",X"AA",X"5A",X"AA",X"59",X"56",X"5A",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
