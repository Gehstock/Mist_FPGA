library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"51",X"32",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"02",X"44",X"88",
		X"32",X"65",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"48",X"6E",X"44",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"8E",X"76",X"9F",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"66",X"FD",X"55",X"8A",
		X"7C",X"BD",X"27",X"0A",X"AA",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"22",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"8C",X"E2",X"77",X"11",X"00",X"22",X"00",X"00",
		X"00",X"00",X"C8",X"CC",X"E6",X"15",X"AA",X"33",X"00",X"00",X"00",X"11",X"44",X"45",X"22",X"10",
		X"00",X"00",X"88",X"44",X"22",X"88",X"91",X"33",X"00",X"00",X"CC",X"02",X"B3",X"55",X"EC",X"EF",
		X"7D",X"8A",X"33",X"48",X"22",X"99",X"00",X"00",X"44",X"00",X"10",X"22",X"11",X"00",X"00",X"00",
		X"DD",X"88",X"00",X"E6",X"44",X"00",X"00",X"00",X"C8",X"2A",X"55",X"2A",X"22",X"66",X"00",X"00",
		X"07",X"78",X"F7",X"FC",X"FC",X"F7",X"F0",X"FF",X"00",X"01",X"03",X"16",X"34",X"3C",X"3C",X"3C",
		X"00",X"08",X"0C",X"86",X"C2",X"C3",X"C3",X"C3",X"0E",X"E1",X"FE",X"F2",X"F3",X"FF",X"F0",X"FE",
		X"FF",X"F0",X"FF",X"FC",X"FC",X"F6",X"78",X"07",X"3C",X"3C",X"3C",X"34",X"16",X"03",X"01",X"00",
		X"C3",X"C3",X"C3",X"C2",X"86",X"0C",X"08",X"00",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",X"E1",X"0E",
		X"44",X"22",X"77",X"1F",X"7F",X"0F",X"FF",X"0F",X"88",X"44",X"22",X"11",X"99",X"77",X"33",X"33",
		X"11",X"22",X"44",X"88",X"99",X"EE",X"CC",X"CC",X"22",X"44",X"EE",X"0F",X"6F",X"6F",X"FF",X"0F",
		X"7F",X"0F",X"FF",X"0F",X"7F",X"0F",X"77",X"88",X"33",X"33",X"77",X"BB",X"11",X"22",X"44",X"88",
		X"CC",X"CC",X"EE",X"DD",X"88",X"44",X"22",X"11",X"EF",X"0F",X"FF",X"0F",X"EF",X"0F",X"EE",X"11",
		X"00",X"C0",X"E0",X"E0",X"C0",X"8B",X"1E",X"3C",X"00",X"10",X"31",X"31",X"10",X"00",X"03",X"0F",
		X"E0",X"F8",X"F8",X"E0",X"44",X"0C",X"CE",X"0F",X"00",X"10",X"10",X"00",X"00",X"0F",X"C7",X"C7",
		X"3C",X"1E",X"8B",X"C0",X"E0",X"E0",X"C0",X"00",X"0F",X"03",X"00",X"10",X"31",X"31",X"10",X"00",
		X"0F",X"CE",X"0C",X"44",X"E0",X"F8",X"F8",X"E0",X"C7",X"C7",X"0F",X"00",X"00",X"10",X"10",X"00",
		X"01",X"01",X"03",X"83",X"C7",X"83",X"16",X"34",X"00",X"00",X"30",X"73",X"70",X"70",X"30",X"00",
		X"00",X"00",X"C0",X"EC",X"E0",X"E0",X"C0",X"00",X"08",X"08",X"0C",X"1C",X"3E",X"1C",X"86",X"C2",
		X"34",X"37",X"07",X"07",X"27",X"AF",X"03",X"01",X"00",X"00",X"00",X"60",X"F6",X"F0",X"F0",X"60",
		X"00",X"00",X"00",X"60",X"F6",X"F0",X"F0",X"60",X"C2",X"CE",X"0E",X"0E",X"4E",X"5F",X"0C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",
		X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"CC",X"F8",X"F8",X"F8",X"E1",X"E1",X"E1",X"E1",
		X"7F",X"3F",X"3F",X"33",X"00",X"00",X"00",X"00",X"09",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"C3",X"C3",X"C3",X"87",X"87",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"38",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"00",X"00",X"0C",X"7F",X"7F",X"7F",X"FE",X"FE",
		X"87",X"87",X"87",X"C3",X"C3",X"03",X"00",X"00",X"34",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"FE",X"FE",X"7F",X"7F",X"7F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"C0",X"87",X"87",X"87",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"30",X"37",X"33",X"33",X"33",X"11",X"11",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"87",X"87",X"87",X"C0",
		X"0C",X"06",X"06",X"07",X"07",X"06",X"06",X"0C",X"03",X"66",X"EE",X"FA",X"FA",X"EE",X"66",X"03",
		X"00",X"00",X"00",X"03",X"95",X"2A",X"55",X"AA",X"CC",X"C8",X"20",X"10",X"00",X"00",X"11",X"11",
		X"33",X"31",X"40",X"80",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"0C",X"56",X"AB",X"55",X"AA",
		X"00",X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",
		X"00",X"00",X"00",X"22",X"FF",X"FF",X"00",X"00",X"00",X"00",X"44",X"44",X"77",X"77",X"44",X"44",
		X"00",X"22",X"33",X"99",X"99",X"DD",X"FF",X"66",X"00",X"66",X"77",X"77",X"55",X"55",X"44",X"44",
		X"00",X"00",X"11",X"99",X"DD",X"FF",X"BB",X"11",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",
		X"00",X"88",X"CC",X"66",X"33",X"FF",X"FF",X"00",X"00",X"11",X"11",X"11",X"11",X"77",X"77",X"11",
		X"00",X"77",X"77",X"55",X"55",X"55",X"DD",X"88",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",
		X"00",X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"33",X"33",X"11",X"99",X"DD",X"77",X"33",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"00",
		X"00",X"66",X"FF",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"55",X"77",X"33",
		X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"88",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CC",X"66",X"33",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"66",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"00",
		X"00",X"00",X"33",X"66",X"CC",X"88",X"00",X"00",X"00",X"00",X"66",X"33",X"11",X"00",X"00",X"00",
		X"55",X"AA",X"5D",X"A6",X"03",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"10",X"20",X"C8",X"CC",
		X"EE",X"33",X"11",X"99",X"DD",X"99",X"BB",X"EE",X"77",X"CC",X"88",X"99",X"BB",X"99",X"DD",X"77",
		X"00",X"CC",X"EE",X"33",X"11",X"33",X"EE",X"CC",X"00",X"77",X"77",X"11",X"11",X"11",X"77",X"77",
		X"00",X"FF",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",X"77",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"CC",X"EE",X"33",X"11",X"11",X"33",X"22",X"00",X"11",X"33",X"66",X"44",X"44",X"66",X"22",
		X"00",X"FF",X"FF",X"11",X"11",X"33",X"EE",X"CC",X"00",X"77",X"77",X"44",X"44",X"66",X"33",X"11",
		X"00",X"00",X"FF",X"FF",X"99",X"99",X"99",X"11",X"00",X"00",X"77",X"77",X"44",X"44",X"44",X"44",
		X"00",X"FF",X"FF",X"99",X"99",X"99",X"99",X"11",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"EE",X"33",X"11",X"99",X"99",X"99",X"00",X"11",X"33",X"66",X"44",X"44",X"77",X"77",
		X"00",X"FF",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",X"77",X"77",X"00",X"00",X"00",X"77",X"77",
		X"00",X"00",X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"44",X"44",X"77",X"77",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"22",X"66",X"44",X"44",X"66",X"77",X"33",
		X"00",X"FF",X"FF",X"88",X"CC",X"66",X"33",X"11",X"00",X"77",X"77",X"11",X"33",X"77",X"66",X"44",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"44",X"44",X"44",X"44",
		X"00",X"FF",X"FF",X"EE",X"CC",X"EE",X"FF",X"FF",X"00",X"77",X"77",X"00",X"11",X"00",X"77",X"77",
		X"00",X"FF",X"FF",X"EE",X"CC",X"88",X"FF",X"FF",X"00",X"77",X"77",X"00",X"11",X"33",X"77",X"77",
		X"00",X"EE",X"FF",X"11",X"11",X"11",X"FF",X"EE",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"EE",X"00",X"77",X"77",X"11",X"11",X"11",X"11",X"00",
		X"08",X"08",X"00",X"00",X"80",X"40",X"31",X"33",X"55",X"AA",X"45",X"9A",X"0C",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"11",X"11",X"99",X"FF",X"EE",X"00",X"77",X"77",X"11",X"33",X"77",X"66",X"44",
		X"00",X"66",X"FF",X"99",X"99",X"BB",X"AA",X"00",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",
		X"00",X"00",X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"FF",X"FF",X"88",X"00",X"88",X"FF",X"FF",X"00",X"00",X"11",X"33",X"77",X"33",X"11",X"00",
		X"00",X"FF",X"FF",X"88",X"CC",X"88",X"FF",X"FF",X"00",X"11",X"77",X"33",X"11",X"33",X"77",X"11",
		X"00",X"33",X"77",X"EE",X"CC",X"EE",X"77",X"33",X"00",X"66",X"77",X"33",X"11",X"33",X"77",X"66",
		X"00",X"00",X"33",X"FF",X"88",X"88",X"FF",X"33",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"00",
		X"00",X"11",X"11",X"99",X"DD",X"FF",X"77",X"33",X"00",X"66",X"77",X"77",X"55",X"44",X"44",X"44",
		X"00",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"00",X"00",X"00",
		X"00",X"22",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"44",X"00",
		X"00",X"00",X"00",X"22",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"00",X"00",
		X"00",X"00",X"03",X"0E",X"5D",X"AA",X"55",X"AA",X"CC",X"C8",X"20",X"10",X"01",X"01",X"03",X"02",
		X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E1",X"C3",X"86",X"84",X"84",X"84",X"84",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"84",X"84",X"84",X"84",X"86",X"C3",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"F0",X"78",X"3C",X"16",X"12",X"12",X"12",X"12",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"12",X"12",X"12",X"12",X"16",X"3C",X"78",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"0C",
		X"E1",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"12",X"12",X"12",X"16",X"3C",X"79",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"84",X"84",X"84",X"84",X"86",X"C3",X"E9",X"FC",
		X"F3",X"79",X"3C",X"16",X"12",X"12",X"12",X"12",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"E9",X"C3",X"86",X"84",X"84",X"84",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FC",
		X"F3",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"12",X"12",X"12",X"12",X"12",X"13",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"84",X"84",X"84",X"8C",X"CC",
		X"33",X"13",X"12",X"12",X"12",X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"8C",X"84",X"84",X"84",X"84",X"84",X"84",
		X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",
		X"12",X"12",X"12",X"12",X"33",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"84",X"84",X"84",X"84",X"CC",X"EE",X"FF",X"FF",
		X"FF",X"EF",X"77",X"33",X"12",X"12",X"12",X"12",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"EE",X"CC",X"84",X"84",X"84",X"84",
		X"00",X"00",X"00",X"00",X"33",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",
		X"FF",X"EF",X"77",X"33",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"EE",X"CC",X"00",X"00",X"00",X"00",
		X"12",X"12",X"12",X"12",X"33",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"84",X"CC",X"EE",X"FF",X"FF",
		X"FF",X"EF",X"77",X"33",X"12",X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"EE",X"CC",X"84",X"84",X"84",X"84",
		X"FF",X"EF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"EE",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",
		X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"11",X"33",X"33",X"3F",X"F3",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CF",X"FC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"EF",X"FF",X"33",X"12",X"12",X"12",X"12",X"F1",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"FF",X"CC",X"84",X"84",X"84",X"84",
		X"9F",X"EF",X"FF",X"33",X"00",X"00",X"00",X"00",X"F1",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"FF",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"11",X"33",X"33",X"33",X"73",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"EF",X"FF",X"33",X"12",X"12",X"12",X"12",X"91",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"FF",X"CC",X"84",X"84",X"84",X"84",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"FF",X"CC",X"00",X"00",X"00",X"00",
		X"9F",X"EF",X"FF",X"33",X"00",X"00",X"00",X"00",X"91",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"12",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"3F",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CF",X"FC",X"84",X"84",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"12",X"12",X"F3",X"3F",X"11",X"11",X"00",X"00",X"00",X"00",
		X"FC",X"CF",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",X"84",X"84",
		X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"3F",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CF",X"FC",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"00",X"00",X"F3",X"3F",X"11",X"11",X"00",X"00",X"00",X"00",
		X"FC",X"CF",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",X"00",X"00",
		X"12",X"02",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"B3",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"84",X"84",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"12",X"12",X"73",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",X"04",X"84",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"B3",
		X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"00",X"00",X"73",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"12",X"12",X"12",X"12",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"F8",X"84",X"84",X"84",X"84",X"CC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"F3",X"3F",X"33",X"33",X"11",X"11",X"00",X"00",
		X"FC",X"CF",X"CC",X"CC",X"88",X"88",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"F8",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",
		X"12",X"12",X"12",X"12",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"84",X"84",X"84",X"80",X"CC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"73",X"33",X"33",X"33",X"11",X"11",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"91",
		X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"B3",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"9F",X"EF",X"FF",X"33",X"00",X"00",X"73",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"FF",X"CC",X"00",X"00",
		X"66",X"FF",X"FF",X"FE",X"FD",X"97",X"C2",X"1F",X"00",X"00",X"00",X"19",X"59",X"3C",X"1E",X"3C",
		X"00",X"88",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",
		X"3C",X"0F",X"1F",X"FF",X"FF",X"FF",X"77",X"00",X"0F",X"07",X"0C",X"08",X"11",X"11",X"00",X"00",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"CC",X"00",X"00",X"1F",X"3F",X"9F",X"FF",X"FF",X"FF",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"66",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"07",X"1D",X"AA",X"55",X"AA",X"55",X"AA",X"CC",X"C8",X"21",X"03",X"13",X"06",X"15",X"26",
		X"33",X"31",X"48",X"0C",X"04",X"8E",X"46",X"8A",X"00",X"0E",X"47",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"2E",X"07",X"00",X"15",X"26",X"17",X"02",X"03",X"21",X"C8",X"CC",
		X"46",X"8A",X"06",X"8C",X"0C",X"48",X"31",X"33",X"55",X"AA",X"55",X"AA",X"55",X"8B",X"0E",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"00",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"11",X"FF",X"00",X"FF",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",
		X"33",X"FF",X"FF",X"8F",X"0F",X"0F",X"6F",X"6F",X"00",X"00",X"11",X"11",X"33",X"33",X"33",X"73",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"1F",X"0F",X"0F",X"6F",X"6F",
		X"6F",X"FF",X"FF",X"33",X"00",X"00",X"00",X"00",X"91",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"FF",X"FF",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"B3",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"73",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"91",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"1F",
		X"0F",X"0F",X"6F",X"6F",X"6F",X"FF",X"FF",X"33",X"73",X"33",X"33",X"33",X"11",X"11",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"0F",X"0F",X"6F",X"6F",X"6F",X"FF",X"FF",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"43",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"10",X"08",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"87",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"F0",X"10",
		X"0F",X"0F",X"0F",X"0F",X"87",X"61",X"10",X"00",X"87",X"43",X"21",X"21",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"87",X"43",
		X"08",X"0F",X"0F",X"87",X"43",X"21",X"21",X"21",X"21",X"21",X"21",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"87",X"00",X"00",X"0C",X"0F",X"0F",X"4B",X"38",X"08",
		X"21",X"21",X"21",X"29",X"0F",X"0F",X"C3",X"30",X"00",X"86",X"87",X"87",X"43",X"21",X"10",X"00",
		X"43",X"43",X"87",X"0E",X"0E",X"0C",X"08",X"00",X"08",X"08",X"08",X"18",X"69",X"0F",X"0F",X"0E",
		X"00",X"0F",X"F0",X"F0",X"F0",X"80",X"12",X"34",X"06",X"69",X"78",X"78",X"70",X"30",X"00",X"00",
		X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"16",X"78",X"F0",X"F0",X"F0",X"78",X"F0",X"C0",
		X"78",X"F0",X"E0",X"E1",X"F0",X"F0",X"F0",X"F0",X"00",X"01",X"16",X"78",X"78",X"78",X"70",X"30",
		X"24",X"78",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"80",X"00",X"07",X"78",X"F0",X"F0",X"F0",X"C0",
		X"3C",X"F0",X"F0",X"87",X"80",X"00",X"00",X"00",X"00",X"03",X"34",X"78",X"78",X"78",X"68",X"68",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"78",X"80",X"E0",X"F0",X"F0",X"3C",X"12",X"01",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"68",X"78",X"34",X"34",X"12",X"01",X"00",X"00",
		X"78",X"78",X"78",X"F0",X"E0",X"C0",X"08",X"00",X"00",X"00",X"00",X"07",X"78",X"78",X"07",X"00",
		X"10",X"61",X"87",X"0F",X"0F",X"29",X"21",X"43",X"00",X"00",X"30",X"C3",X"87",X"87",X"86",X"00",
		X"08",X"0C",X"0C",X"0E",X"86",X"87",X"43",X"43",X"C3",X"0F",X"0F",X"1C",X"0C",X"08",X"08",X"0C",
		X"43",X"87",X"0F",X"0E",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"10",X"21",X"43",X"43",X"43",X"43",
		X"87",X"86",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"04",X"06",X"16",X"87",X"43",X"43",X"21",X"00",
		X"33",X"31",X"40",X"80",X"08",X"08",X"0C",X"8C",X"00",X"00",X"0C",X"8F",X"45",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"2A",X"1F",X"03",X"00",X"00",X"13",X"03",X"01",X"01",X"10",X"20",X"C8",X"CC",
		X"04",X"0C",X"08",X"08",X"80",X"40",X"31",X"33",X"55",X"AA",X"55",X"AB",X"07",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"87",X"0F",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"71",X"F1",X"E1",X"07",X"03",X"03",X"06",X"06",
		X"88",X"66",X"00",X"08",X"0E",X"0F",X"87",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"61",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"03",X"03",X"07",X"E1",X"F1",X"71",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"01",X"00",X"00",X"30",X"30",X"10",
		X"68",X"78",X"78",X"3C",X"06",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"01",X"0F",X"03",
		X"02",X"02",X"02",X"06",X"3C",X"78",X"78",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"87",X"0F",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"F0",X"E1",X"07",X"03",X"03",X"06",X"06",
		X"88",X"66",X"00",X"08",X"0E",X"0F",X"87",X"87",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"03",X"03",X"07",X"E1",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"01",X"00",X"00",X"30",X"30",X"10",
		X"68",X"7A",X"7A",X"3C",X"06",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"01",X"0F",X"03",
		X"02",X"02",X"02",X"06",X"3C",X"7A",X"7A",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"60",X"78",X"78",X"3F",X"3C",X"0F",X"0F",X"07",X"60",X"E1",X"E1",X"CF",X"C3",X"0F",X"0F",X"0E",
		X"00",X"03",X"0F",X"0C",X"19",X"22",X"22",X"00",X"00",X"0C",X"0F",X"03",X"01",X"00",X"00",X"00",
		X"02",X"02",X"03",X"07",X"0F",X"78",X"F0",X"E0",X"04",X"04",X"0C",X"0E",X"0F",X"E1",X"F0",X"70",
		X"00",X"00",X"60",X"70",X"00",X"08",X"0F",X"00",X"00",X"00",X"60",X"E0",X"00",X"01",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"60",X"78",X"78",X"3C",X"3C",X"0F",X"0F",X"07",X"60",X"E1",X"E1",X"C3",X"C3",X"0F",X"0F",X"0E",
		X"00",X"03",X"0F",X"0C",X"19",X"22",X"22",X"00",X"00",X"0C",X"0F",X"03",X"01",X"00",X"00",X"00",
		X"02",X"02",X"03",X"07",X"0F",X"78",X"F6",X"E0",X"04",X"04",X"0C",X"0E",X"0F",X"E1",X"F6",X"70",
		X"00",X"00",X"60",X"70",X"00",X"08",X"0F",X"00",X"00",X"00",X"60",X"E0",X"00",X"01",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"0E",X"06",X"02",X"03",X"03",X"C0",X"A4",X"00",X"01",X"03",X"06",X"86",X"86",
		X"30",X"07",X"0F",X"08",X"00",X"88",X"44",X"00",X"E0",X"C3",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"12",X"12",X"06",X"06",X"0C",X"08",X"00",X"00",X"C2",X"C2",X"87",X"07",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"03",X"30",X"30",X"E0",X"C0",X"00",X"03",X"0F",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"0E",X"0F",X"01",X"22",X"44",X"00",X"00",
		X"30",X"12",X"00",X"08",X"0C",X"06",X"16",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"0C",
		X"34",X"34",X"1E",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"3C",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"04",X"0C",X"0C",
		X"C0",X"C0",X"70",X"30",X"00",X"0C",X"0F",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"06",X"06",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F4",
		X"00",X"00",X"02",X"02",X"03",X"03",X"07",X"87",X"00",X"00",X"00",X"00",X"00",X"38",X"78",X"0F",
		X"E0",X"48",X"0C",X"04",X"00",X"80",X"80",X"80",X"F4",X"70",X"03",X"07",X"03",X"03",X"07",X"07",
		X"87",X"0F",X"0F",X"0C",X"08",X"08",X"00",X"00",X"0F",X"09",X"00",X"00",X"00",X"10",X"10",X"00",
		X"80",X"80",X"80",X"00",X"04",X"0C",X"48",X"E0",X"07",X"07",X"03",X"03",X"07",X"03",X"70",X"F4",
		X"44",X"33",X"08",X"08",X"0C",X"0F",X"0F",X"87",X"00",X"10",X"10",X"00",X"00",X"00",X"09",X"0F",
		X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"F4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"07",X"03",X"03",X"02",X"02",X"00",X"00",X"0F",X"78",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C8",X"C8",X"C8",X"80",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",
		X"03",X"03",X"03",X"03",X"07",X"87",X"87",X"07",X"00",X"00",X"08",X"78",X"F8",X"3C",X"3C",X"1E",
		X"08",X"0C",X"0C",X"04",X"00",X"C0",X"C0",X"40",X"00",X"01",X"03",X"01",X"01",X"03",X"03",X"03",
		X"0F",X"0F",X"0F",X"0C",X"08",X"00",X"00",X"00",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"C0",X"00",X"04",X"0C",X"0C",X"08",X"03",X"03",X"03",X"01",X"01",X"03",X"01",X"00",
		X"22",X"11",X"00",X"08",X"0C",X"0F",X"0F",X"0F",X"00",X"88",X"00",X"00",X"00",X"00",X"09",X"0F",
		X"80",X"C8",X"C8",X"C8",X"80",X"00",X"00",X"00",X"70",X"F0",X"F0",X"70",X"00",X"00",X"00",X"00",
		X"07",X"87",X"87",X"07",X"03",X"03",X"03",X"03",X"1E",X"3C",X"3C",X"F8",X"78",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"0F",X"0F",X"03",X"00",X"00",X"00",
		X"10",X"39",X"3C",X"3C",X"1E",X"0F",X"07",X"07",X"80",X"C8",X"C0",X"C0",X"80",X"0C",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"00",X"00",X"00",
		X"03",X"01",X"01",X"03",X"16",X"3C",X"10",X"00",X"0E",X"48",X"68",X"68",X"E0",X"E0",X"C0",X"00",
		X"00",X"03",X"0F",X"0F",X"0C",X"11",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"10",X"31",X"30",X"30",X"10",X"03",X"0F",X"0F",X"80",X"C9",X"C3",X"C3",X"87",X"0F",X"0E",X"0E",
		X"00",X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"21",X"61",X"61",X"70",X"70",X"30",X"00",X"0C",X"08",X"08",X"0C",X"86",X"C3",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0E",X"0F",X"01",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0E",X"0F",X"0F",X"07",X"07",X"60",X"F0",X"F0",X"F0",X"60",X"0F",X"0F",X"0F",
		X"0C",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"00",X"00",
		X"03",X"01",X"01",X"03",X"07",X"0E",X"00",X"00",X"0F",X"1E",X"78",X"F0",X"F7",X"70",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"08",X"00",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"60",X"F0",X"F0",X"F0",X"60",X"0F",X"0F",X"0F",X"00",X"00",X"02",X"07",X"0F",X"0F",X"0E",X"0E",
		X"22",X"00",X"00",X"00",X"60",X"70",X"00",X"00",X"03",X"10",X"10",X"10",X"10",X"00",X"00",X"00",
		X"0F",X"87",X"E1",X"F0",X"FE",X"E0",X"00",X"00",X"0C",X"08",X"08",X"0C",X"0E",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",
		X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"11",X"11",X"33",X"33",X"77",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"CC",X"CC",X"88",X"88",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"BF",X"CF",X"33",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"77",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"EE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"88",X"00",X"00",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"00",X"00",X"11",X"77",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"00",X"00",X"33",X"77",X"DF",X"BF",X"7F",X"7F",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"77",X"33",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"04",X"0C",X"09",X"09",
		X"00",X"00",X"00",X"10",X"16",X"0F",X"0F",X"0F",X"00",X"00",X"E0",X"F0",X"C3",X"C4",X"C4",X"E6",
		X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"09",X"09",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"07",X"09",X"0F",X"16",X"10",X"00",X"00",X"00",X"E6",X"C4",X"C4",X"C3",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"07",X"0C",X"00",X"03",X"06",X"0D",X"0D",X"87",X"0E",X"03",X"00",X"0C",X"0E",X"0F",X"0F",X"1E",
		X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F7",X"19",X"08",X"0F",X"07",X"00",X"00",X"F0",X"FE",X"89",X"01",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"80",X"0C",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"04",X"0C",X"08",X"08",
		X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"00",X"60",X"F0",X"F0",X"69",X"6A",X"6A",X"7B",
		X"06",X"06",X"06",X"0C",X"80",X"00",X"00",X"00",X"08",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"0B",X"0C",X"07",X"07",X"03",X"00",X"00",X"00",X"7B",X"6A",X"6A",X"69",X"F0",X"F0",X"60",X"00",
		X"00",X"00",X"00",X"80",X"0E",X"03",X"03",X"8B",X"02",X"02",X"00",X"06",X"0E",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"00",X"60",X"F0",X"F0",X"78",X"3D",X"3D",X"3D",
		X"8B",X"03",X"03",X"0E",X"80",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0E",X"06",X"00",X"02",X"02",
		X"0D",X"0E",X"0F",X"07",X"03",X"00",X"00",X"00",X"3D",X"35",X"3D",X"78",X"F0",X"F0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"07",X"0C",X"00",X"00",X"03",X"0E",X"0D",X"0D",X"0E",X"03",X"00",X"00",X"0C",X"0F",X"0F",X"0F",
		X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"00",
		X"0F",X"F0",X"F7",X"19",X"08",X"0F",X"07",X"00",X"0F",X"F0",X"FF",X"88",X"00",X"0F",X"0F",X"00",
		X"00",X"08",X"0B",X"00",X"00",X"00",X"08",X"08",X"00",X"01",X"0D",X"00",X"00",X"00",X"01",X"01",
		X"0F",X"0F",X"08",X"00",X"07",X"0F",X"0E",X"0D",X"0F",X"0F",X"01",X"00",X"0E",X"0F",X"0F",X"0F",
		X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"00",
		X"0D",X"F7",X"F0",X"97",X"09",X"08",X"0F",X"07",X"0F",X"FE",X"F0",X"9E",X"09",X"01",X"0F",X"0E",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"48",X"00",X"01",X"03",X"06",X"04",X"01",X"01",X"01",
		X"00",X"08",X"00",X"07",X"0F",X"07",X"0B",X"1E",X"00",X"00",X"00",X"0C",X"78",X"78",X"F0",X"F7",
		X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"F1",X"F1",X"F1",X"E1",X"70",X"00",X"00",X"CC",X"CC",X"01",X"03",X"0F",X"0C",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"02",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"21",
		X"00",X"00",X"00",X"03",X"E1",X"E1",X"F0",X"FE",X"00",X"01",X"00",X"0E",X"0D",X"0B",X"0F",X"87",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"33",X"33",X"08",X"0C",X"0F",X"03",X"00",X"00",X"C3",X"F8",X"F8",X"F8",X"78",X"E0",X"00",X"00",
		X"00",X"88",X"00",X"00",X"88",X"88",X"88",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"FF",X"00",X"00",X"FF",X"88",X"FF",X"00",X"33",X"FF",X"00",X"00",X"FF",X"11",X"FF",X"00",
		X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"11",X"FF",X"00",X"FF",X"11",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"12",X"21",X"73",X"73",X"73",X"51",X"88",X"88",X"48",X"84",X"EC",X"EC",X"EC",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"11",X"11",X"12",X"21",X"73",X"73",X"00",X"00",X"88",X"88",X"48",X"84",X"EC",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"73",X"51",X"00",X"00",X"02",X"00",X"01",X"20",X"EC",X"A8",X"00",X"08",X"80",X"04",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"11",X"11",X"21",X"12",X"73",X"73",X"00",X"00",X"88",X"88",X"84",X"48",X"EC",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"73",X"51",X"00",X"02",X"10",X"00",X"20",X"01",X"EC",X"A8",X"00",X"00",X"40",X"08",X"00",X"40",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"4B",X"0F",X"03",X"07",X"1E",X"2D",X"4B",X"5A",X"34",X"34",
		X"08",X"0C",X"86",X"0F",X"0F",X"4B",X"87",X"1E",X"03",X"07",X"0F",X"3C",X"4B",X"A5",X"C3",X"F0",
		X"0E",X"86",X"0C",X"86",X"87",X"0F",X"0E",X"08",X"12",X"07",X"1E",X"2D",X"3C",X"16",X"12",X"01",
		X"D2",X"B4",X"4B",X"E1",X"78",X"E1",X"0F",X"69",X"A5",X"0F",X"87",X"A5",X"D2",X"B4",X"87",X"0D",
		X"E0",X"F2",X"F2",X"E0",X"44",X"0C",X"CE",X"0F",X"00",X"10",X"30",X"30",X"10",X"00",X"03",X"0F",
		X"00",X"C4",X"E4",X"E0",X"C0",X"8B",X"1E",X"3C",X"00",X"10",X"10",X"00",X"00",X"0F",X"C7",X"C7",
		X"0F",X"CE",X"0C",X"44",X"E0",X"F2",X"F2",X"E0",X"0F",X"03",X"00",X"10",X"30",X"30",X"10",X"00",
		X"3C",X"1E",X"8B",X"C0",X"E0",X"E4",X"C4",X"00",X"C7",X"C7",X"0F",X"00",X"00",X"10",X"10",X"00",
		X"E0",X"F8",X"F8",X"E0",X"44",X"0C",X"CE",X"0F",X"00",X"10",X"31",X"31",X"10",X"00",X"03",X"0F",
		X"00",X"C0",X"E0",X"E0",X"C0",X"8B",X"1E",X"3C",X"00",X"10",X"10",X"00",X"00",X"0F",X"C7",X"C7",
		X"0F",X"CE",X"0C",X"44",X"E0",X"F8",X"F8",X"E0",X"0F",X"03",X"00",X"10",X"31",X"31",X"10",X"00",
		X"3C",X"1E",X"8B",X"C0",X"E0",X"E0",X"C0",X"00",X"C7",X"C7",X"0F",X"00",X"00",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"F2",X"F0",X"00",X"06",X"07",X"03",X"03",X"01",X"01",X"F1",
		X"10",X"10",X"18",X"1F",X"0F",X"0F",X"3C",X"3C",X"C0",X"E4",X"F0",X"E0",X"40",X"08",X"0C",X"C2",
		X"F8",X"2C",X"8C",X"4E",X"0E",X"0E",X"0C",X"00",X"F0",X"F0",X"74",X"20",X"00",X"00",X"00",X"00",
		X"16",X"96",X"03",X"01",X"30",X"70",X"72",X"30",X"C7",X"CF",X"0F",X"0F",X"AF",X"97",X"C1",X"80",
		X"00",X"00",X"C0",X"E0",X"E0",X"EC",X"C0",X"00",X"00",X"00",X"30",X"70",X"70",X"73",X"30",X"00",
		X"01",X"01",X"03",X"83",X"C7",X"83",X"16",X"34",X"08",X"08",X"0C",X"1C",X"3E",X"1C",X"86",X"C2",
		X"00",X"00",X"00",X"60",X"F0",X"F0",X"F6",X"60",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F6",X"60",
		X"34",X"37",X"07",X"07",X"27",X"AF",X"03",X"01",X"C2",X"CE",X"0E",X"0E",X"4E",X"5F",X"0C",X"08",
		X"00",X"00",X"C0",X"EC",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"30",X"73",X"70",X"70",X"30",X"00",
		X"01",X"01",X"03",X"83",X"C7",X"83",X"16",X"34",X"08",X"08",X"0C",X"1C",X"3E",X"1C",X"86",X"C2",
		X"00",X"00",X"00",X"60",X"F6",X"F0",X"F0",X"60",X"00",X"00",X"00",X"60",X"F6",X"F0",X"F0",X"60",
		X"34",X"37",X"07",X"07",X"27",X"AF",X"03",X"01",X"C2",X"CE",X"0E",X"0E",X"4E",X"5F",X"0C",X"08",
		X"0C",X"0E",X"0F",X"0F",X"87",X"C2",X"0E",X"0C",X"00",X"06",X"07",X"07",X"1E",X"3C",X"1E",X"16",
		X"03",X"07",X"0F",X"87",X"2D",X"5A",X"D2",X"3C",X"01",X"0B",X"0F",X"96",X"96",X"4B",X"E1",X"A5",
		X"84",X"0E",X"0F",X"87",X"87",X"0F",X"0A",X"00",X"03",X"01",X"03",X"16",X"16",X"03",X"03",X"01",
		X"B4",X"78",X"E1",X"2D",X"96",X"C3",X"83",X"08",X"5A",X"C3",X"A5",X"C3",X"5A",X"3C",X"07",X"03",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0E",X"0E",X"0C",X"00",X"03",X"03",X"16",X"25",X"3C",X"3C",X"1E",
		X"0F",X"0F",X"69",X"87",X"0F",X"A5",X"2D",X"D2",X"00",X"0C",X"0F",X"0F",X"69",X"96",X"C3",X"B4",
		X"0E",X"4A",X"87",X"C3",X"0F",X"0E",X"0C",X"00",X"5A",X"69",X"1E",X"2D",X"34",X"16",X"03",X"00",
		X"3C",X"96",X"A5",X"D2",X"69",X"C3",X"0F",X"0C",X"87",X"0F",X"C3",X"96",X"78",X"2D",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"DE",
		X"FF",X"EE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ED",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"30",X"B7",X"7B",X"00",X"00",X"00",X"00",X"00",X"C0",X"88",X"CD",
		X"02",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B7",X"7B",X"30",X"00",X"00",X"00",X"00",X"00",X"CC",X"88",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"30",X"7B",X"B7",X"00",X"00",X"00",X"00",X"00",X"C0",X"88",X"CC",
		X"81",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7B",X"B7",X"30",X"00",X"00",X"00",X"00",X"00",X"CC",X"89",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"0E",X"0E",X"0C",X"00",X"08",X"0C",X"06",X"07",X"07",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"06",X"4B",X"BD",X"78",X"F0",X"00",X"01",X"05",X"1E",X"AD",X"C3",X"97",X"E3",
		X"0C",X"08",X"08",X"00",X"86",X"4B",X"0F",X"06",X"02",X"03",X"01",X"00",X"04",X"07",X"03",X"03",
		X"BC",X"7D",X"29",X"56",X"83",X"09",X"08",X"00",X"FB",X"E5",X"B4",X"0F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"0C",X"0E",X"0E",X"0F",X"0F",X"06",X"03",X"07",X"07",X"07",X"03",X"01",X"00",X"00",
		X"08",X"0C",X"0E",X"0E",X"0D",X"09",X"01",X"03",X"00",X"0C",X"0E",X"05",X"01",X"0B",X"0F",X"0F",
		X"00",X"00",X"08",X"0C",X"0C",X"0C",X"08",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"07",X"03",X"00",
		X"07",X"07",X"0E",X"0C",X"08",X"08",X"00",X"00",X"0E",X"0F",X"07",X"07",X"0F",X"0F",X"07",X"03",
		X"00",X"08",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"0E",X"0C",X"00",X"00",X"00",X"00",X"04",X"0C",X"0E",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"80",X"00",X"00",X"60",X"80",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"D0",X"70",X"B0",X"63",X"00",X"00",X"00",X"40",X"F0",X"E4",X"F8",X"6C",
		X"00",X"40",X"00",X"80",X"80",X"40",X"00",X"00",X"20",X"10",X"00",X"00",X"10",X"20",X"00",X"00",
		X"C3",X"73",X"E1",X"B2",X"20",X"10",X"00",X"00",X"B4",X"6C",X"F1",X"D0",X"A0",X"40",X"00",X"00",
		X"00",X"00",X"40",X"80",X"80",X"00",X"80",X"C8",X"00",X"00",X"20",X"10",X"00",X"00",X"20",X"10",
		X"00",X"00",X"20",X"90",X"F1",X"73",X"F4",X"ED",X"00",X"00",X"80",X"D8",X"FE",X"F4",X"7B",X"79",
		X"C8",X"A0",X"00",X"80",X"80",X"40",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"20",X"00",X"00",
		X"FE",X"F4",X"F3",X"F3",X"90",X"20",X"00",X"00",X"3C",X"7B",X"F5",X"FE",X"D8",X"80",X"40",X"00",
		X"00",X"20",X"40",X"80",X"80",X"D8",X"EC",X"E8",X"00",X"40",X"20",X"10",X"11",X"B1",X"73",X"71",
		X"90",X"71",X"77",X"FF",X"E3",X"C3",X"AD",X"1E",X"90",X"EC",X"E6",X"FE",X"7E",X"3F",X"97",X"C3",
		X"E8",X"EC",X"D8",X"88",X"80",X"40",X"20",X"00",X"75",X"77",X"B1",X"10",X"10",X"20",X"40",X"00",
		X"3C",X"9E",X"CF",X"E7",X"F7",X"76",X"71",X"90",X"87",X"5B",X"3C",X"7C",X"FF",X"EE",X"E8",X"90",
		X"C0",X"16",X"40",X"1C",X"20",X"00",X"00",X"00",X"10",X"60",X"50",X"82",X"60",X"02",X"00",X"00",
		X"40",X"0C",X"08",X"80",X"00",X"80",X"00",X"00",X"00",X"80",X"C1",X"00",X"02",X"00",X"20",X"00",
		X"60",X"90",X"02",X"08",X"86",X"50",X"68",X"80",X"10",X"00",X"00",X"00",X"60",X"10",X"42",X"30",
		X"00",X"00",X"04",X"1C",X"00",X"08",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"C0",X"E4",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"E4",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"31",X"10",X"00",X"00",X"00",X"00",X"00",X"E0",X"EC",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CC",X"CC",X"88",X"88",X"88",X"66",X"FF",X"FF",X"FF",X"FE",X"76",X"32",X"32",
		X"11",X"BB",X"FF",X"F0",X"F0",X"F0",X"FE",X"FC",X"CC",X"FF",X"FF",X"F1",X"F0",X"F0",X"FE",X"F6",
		X"CC",X"CC",X"AA",X"FF",X"FF",X"F7",X"E6",X"C4",X"76",X"77",X"33",X"11",X"00",X"11",X"11",X"33",
		X"F1",X"F1",X"FF",X"FE",X"FC",X"F8",X"F9",X"FB",X"F0",X"F1",X"FF",X"F1",X"F0",X"F0",X"FC",X"FE",
		X"80",X"E6",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"33",X"33",X"11",X"00",X"00",X"11",X"11",X"11",
		X"FB",X"F9",X"FC",X"FE",X"FF",X"F8",X"F0",X"F0",X"FE",X"FC",X"F0",X"F1",X"FF",X"F1",X"F0",X"F8",
		X"00",X"88",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"33",X"33",X"77",X"77",X"76",X"32",X"31",X"11",
		X"FF",X"FF",X"FF",X"F1",X"F0",X"F0",X"FF",X"DD",X"F9",X"F3",X"F1",X"F8",X"F1",X"F3",X"FF",X"CC");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
