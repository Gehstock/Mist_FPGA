library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity satans_hollow_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of satans_hollow_sp_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"DD",X"D7",X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"77",X"DD",X"DD",X"70",X"67",X"7D",X"67",X"70",
		X"67",X"7D",X"67",X"70",X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"66",X"D7",
		X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"DD",X"D7",X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"DD",X"DD",X"70",X"60",X"7D",X"67",X"70",
		X"60",X"7D",X"67",X"70",X"00",X"77",X"77",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"66",X"D7",
		X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"0D",X"77",X"00",
		X"00",X"ED",X"DD",X"D7",X"00",X"D7",X"66",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"77",X"0D",X"DD",X"70",X"67",X"DD",X"67",X"70",
		X"67",X"7D",X"67",X"70",X"77",X"07",X"77",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"66",X"D7",
		X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"DF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"DD",X"0D",X"77",X"00",
		X"07",X"DD",X"DD",X"D7",X"07",X"77",X"66",X"00",X"77",X"07",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"0D",X"DD",X"70",X"60",X"DD",X"67",X"70",
		X"60",X"7D",X"67",X"70",X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"66",X"D7",
		X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"0D",X"77",X"00",
		X"00",X"ED",X"DD",X"D7",X"00",X"D7",X"66",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"77",X"0D",X"DD",X"70",X"67",X"7D",X"67",X"70",
		X"67",X"7D",X"67",X"70",X"77",X"07",X"77",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"77",X"00",X"00",X"ED",X"DD",X"00",X"00",X"D7",X"66",X"D7",
		X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"DD",X"0D",X"77",X"00",
		X"07",X"DD",X"DD",X"D7",X"07",X"77",X"66",X"00",X"77",X"07",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"0D",X"DD",X"70",X"60",X"7D",X"67",X"70",
		X"60",X"7D",X"67",X"70",X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"DD",X"0D",X"77",X"00",X"07",X"DD",X"DD",X"00",X"07",X"77",X"66",X"D7",
		X"77",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"43",X"00",X"00",X"01",X"41",X"00",X"00",X"14",X"43",X"00",X"00",X"32",X"41",X"10",
		X"10",X"32",X"43",X"21",X"41",X"11",X"11",X"42",X"14",X"01",X"00",X"24",X"01",X"01",X"01",X"22",
		X"01",X"19",X"13",X"31",X"00",X"99",X"13",X"10",X"00",X"CC",X"33",X"00",X"00",X"99",X"33",X"00",
		X"01",X"19",X"13",X"00",X"01",X"01",X"01",X"01",X"14",X"11",X"11",X"14",X"41",X"33",X"22",X"14",
		X"10",X"22",X"44",X"44",X"00",X"32",X"11",X"14",X"00",X"14",X"00",X"14",X"10",X"42",X"00",X"01",
		X"31",X"22",X"00",X"00",X"C1",X"23",X"00",X"00",X"C3",X"11",X"00",X"00",X"41",X"00",X"00",X"00",
		X"31",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"0C",X"C9",X"00",X"00",X"0C",X"C9",
		X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"C9",X"00",X"0F",X"00",X"C9",X"00",X"FC",X"00",X"99",
		X"00",X"FC",X"00",X"99",X"00",X"FF",X"09",X"09",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"9F",X"90",X"00",X"00",X"9F",X"99",X"00",X"00",X"F0",X"F9",
		X"00",X"00",X"F0",X"F9",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"F9",X"0C",
		X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"9C",X"00",X"00",X"9C",X"9C",X"00",X"00",X"9C",X"0F",
		X"00",X"00",X"CC",X"F0",X"00",X"0F",X"C0",X"F0",X"00",X"9C",X"00",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"FF",X"00",X"99",X"00",X"0F",X"00",X"B9",X"00",
		X"09",X"09",X"BB",X"00",X"09",X"99",X"9B",X"99",X"09",X"99",X"9B",X"99",X"09",X"99",X"9B",X"00",
		X"09",X"99",X"9B",X"00",X"09",X"99",X"9B",X"99",X"FF",X"09",X"9B",X"99",X"00",X"00",X"9B",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"05",X"09",X"00",X"00",X"55",X"66",X"00",
		X"00",X"55",X"6C",X"00",X"00",X"05",X"CC",X"00",X"00",X"FF",X"CC",X"60",X"00",X"5F",X"CC",X"60",
		X"00",X"F5",X"CC",X"60",X"00",X"55",X"6C",X"60",X"99",X"90",X"66",X"60",X"90",X"06",X"96",X"60",
		X"90",X"06",X"96",X"60",X"00",X"06",X"06",X"60",X"00",X"06",X"66",X"00",X"00",X"06",X"66",X"00",
		X"00",X"06",X"C6",X"00",X"00",X"06",X"CC",X"00",X"00",X"06",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"BB",X"C0",X"00",X"00",X"BB",X"CC",X"00",X"BB",X"BB",X"CC",X"00",X"00",X"BB",X"CC",X"00",
		X"00",X"BB",X"C0",X"00",X"00",X"B0",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"99",X"00",X"00",X"DD",X"9C",X"00",X"00",X"0D",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"90",X"00",X"00",X"DD",X"C9",X"00",X"00",X"0D",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"90",
		X"00",X"00",X"02",X"99",X"33",X"00",X"92",X"99",X"93",X"99",X"92",X"22",X"33",X"92",X"99",X"90",
		X"00",X"00",X"29",X"90",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"02",X"99",
		X"00",X"00",X"02",X"90",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"09",X"00",X"00",X"BB",X"B9",X"00",X"00",X"9B",X"BB",X"1B",X"00",X"00",X"BB",X"B1",X"00",
		X"00",X"B9",X"BB",X"00",X"00",X"1B",X"1B",X"00",X"09",X"C1",X"11",X"00",X"A1",X"C1",X"B1",X"00",
		X"BA",X"AA",X"B1",X"00",X"BB",X"1C",X"BB",X"10",X"9B",X"1C",X"BB",X"19",X"BB",X"11",X"11",X"11",
		X"BB",X"11",X"19",X"11",X"BB",X"91",X"91",X"1B",X"BB",X"B9",X"99",X"1B",X"BB",X"BB",X"B9",X"1B",
		X"BB",X"BB",X"91",X"1B",X"BB",X"11",X"19",X"11",X"BB",X"11",X"11",X"11",X"9B",X"1C",X"BB",X"19",
		X"BB",X"1C",X"BB",X"00",X"99",X"AA",X"9B",X"00",X"9A",X"C1",X"11",X"00",X"A1",X"C1",X"1B",X"00",
		X"09",X"1B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"1B",X"B9",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"BB",X"0F",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"09",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",
		X"CC",X"00",X"99",X"00",X"C9",X"77",X"99",X"70",X"99",X"FF",X"99",X"FA",X"C9",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"19",X"00",X"00",X"BB",X"11",X"00",X"00",X"BB",X"11",X"00",X"00",X"BB",X"11",
		X"00",X"00",X"BA",X"1C",X"00",X"00",X"BA",X"AC",X"00",X"00",X"AA",X"AA",X"00",X"00",X"A1",X"CC",
		X"00",X"00",X"11",X"C1",X"00",X"00",X"0B",X"C1",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"B9",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"11",X"BB",X"00",X"00",X"1B",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"1B",X"00",X"00",X"91",X"1B",X"00",X"00",X"99",X"1B",X"00",X"00",X"19",X"11",X"00",X"00",
		X"BB",X"11",X"00",X"00",X"BB",X"1B",X"00",X"00",X"9B",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",
		X"B1",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"97",X"88",X"88",X"88",X"99",
		X"88",X"88",X"88",X"79",X"88",X"88",X"88",X"79",X"88",X"88",X"88",X"97",X"88",X"88",X"88",X"99",
		X"88",X"88",X"8F",X"99",X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"99",X"88",X"88",X"89",X"99",
		X"88",X"88",X"99",X"99",X"88",X"88",X"99",X"9C",X"88",X"88",X"99",X"9A",X"88",X"88",X"FF",X"99",
		X"88",X"88",X"F8",X"99",X"88",X"88",X"88",X"99",X"88",X"88",X"F8",X"99",X"88",X"88",X"89",X"9C",
		X"88",X"88",X"8F",X"99",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"79",X"88",X"88",X"88",X"99",
		X"88",X"88",X"88",X"97",X"88",X"88",X"8F",X"77",X"88",X"88",X"89",X"99",X"88",X"88",X"F8",X"99",
		X"88",X"88",X"99",X"9F",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"9B",X"B9",X"19",X"00",X"9B",X"B9",X"11",X"00",X"9B",X"B9",X"11",X"00",X"9B",X"B9",X"1C",
		X"00",X"99",X"9B",X"CC",X"00",X"99",X"BB",X"CC",X"00",X"99",X"BB",X"CC",X"00",X"09",X"BB",X"AA",
		X"00",X"09",X"BB",X"C1",X"00",X"09",X"BB",X"CB",X"00",X"00",X"BB",X"1B",X"00",X"00",X"99",X"BB",
		X"00",X"0A",X"91",X"BB",X"00",X"AA",X"B1",X"BB",X"00",X"A0",X"BC",X"BB",X"00",X"00",X"BB",X"9B",
		X"00",X"00",X"BB",X"B9",X"00",X"00",X"B0",X"99",X"00",X"09",X"9B",X"99",X"00",X"91",X"99",X"99",
		X"00",X"11",X"09",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"11",X"9B",X"00",X"99",X"CC",X"9B",X"00",X"19",X"11",X"91",X"00",X"19",X"CC",X"91",X"00",
		X"11",X"11",X"91",X"00",X"BB",X"9C",X"11",X"00",X"BB",X"91",X"1B",X"00",X"BB",X"B9",X"B0",X"00",
		X"B1",X"11",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B1",X"11",X"00",X"00",X"B9",X"11",X"00",X"00",
		X"9B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"1B",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"DF",X"DE",X"00",X"00",X"FF",X"DE",X"00",X"00",X"FD",X"DE",X"00",
		X"00",X"FD",X"E0",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"EE",X"00",X"00",X"0D",X"ED",X"00",
		X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"30",X"00",X"03",X"00",X"33",X"00",X"34",X"00",X"33",
		X"00",X"02",X"00",X"33",X"00",X"00",X"33",X"22",X"00",X"00",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"22",X"33",X"22",X"00",X"00",X"22",X"33",X"00",X"00",X"23",X"30",X"00",X"00",X"23",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"C5",X"00",X"00",X"50",X"CC",X"00",
		X"00",X"5C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"5C",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"C5",X"CC",X"00",X"00",X"CC",X"5C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"99",X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"CC",X"00",X"55",X"00",X"CC",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"CC",X"00",
		X"99",X"55",X"99",X"CC",X"99",X"55",X"99",X"CC",X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",X"99",
		X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",X"99",X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"CC",X"55",X"CC",X"CC",X"CC",X"55",X"CC",X"CC",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"55",
		X"CC",X"99",X"55",X"55",X"CC",X"99",X"55",X"55",X"55",X"99",X"99",X"55",X"55",X"99",X"99",X"95",
		X"59",X"99",X"99",X"CC",X"99",X"99",X"99",X"CC",X"55",X"99",X"F9",X"55",X"55",X"99",X"FF",X"55",
		X"CC",X"99",X"9F",X"99",X"CC",X"99",X"FF",X"95",X"CC",X"99",X"9F",X"55",X"CC",X"99",X"99",X"55",
		X"55",X"55",X"99",X"CC",X"55",X"55",X"99",X"CC",X"55",X"99",X"99",X"55",X"55",X"99",X"99",X"55",
		X"CC",X"99",X"55",X"99",X"CC",X"99",X"55",X"99",X"00",X"95",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"CC",X"55",X"CC",X"00",X"CC",X"55",X"CC",X"CC",X"00",X"55",X"00",X"CC",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"FF",X"09",
		X"00",X"09",X"FC",X"09",X"00",X"00",X"FC",X"99",X"09",X"00",X"FC",X"99",X"09",X"99",X"CC",X"99",
		X"9C",X"99",X"FF",X"90",X"99",X"99",X"FF",X"CC",X"CC",X"CC",X"CC",X"99",X"FC",X"99",X"CC",X"99",
		X"FF",X"FC",X"CC",X"99",X"99",X"CF",X"FF",X"90",X"99",X"CF",X"F9",X"99",X"99",X"99",X"CC",X"99",
		X"09",X"C9",X"C9",X"99",X"09",X"CC",X"99",X"99",X"00",X"FF",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"FF",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"90",X"99",
		X"00",X"99",X"99",X"00",X"00",X"FF",X"99",X"00",X"09",X"CC",X"99",X"99",X"09",X"C9",X"99",X"99",
		X"99",X"99",X"CC",X"99",X"99",X"CF",X"F9",X"99",X"99",X"CF",X"FF",X"90",X"FF",X"FC",X"CC",X"99",
		X"99",X"99",X"99",X"99",X"CC",X"CC",X"CC",X"99",X"99",X"99",X"9F",X"CC",X"9C",X"99",X"9F",X"90",
		X"09",X"99",X"99",X"99",X"09",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"09",X"9C",X"09",
		X"00",X"99",X"9F",X"09",X"00",X"99",X"9F",X"09",X"00",X"99",X"99",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"FC",X"00",X"C9",X"99",X"F9",X"09",X"C9",X"00",X"99",X"9C",X"90",X"99",
		X"C9",X"99",X"00",X"99",X"C9",X"0C",X"99",X"99",X"CC",X"00",X"09",X"09",X"00",X"00",X"00",X"09",
		X"00",X"90",X"00",X"C9",X"00",X"C9",X"00",X"C9",X"00",X"CC",X"00",X"C9",X"00",X"CC",X"00",X"C9",
		X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"CC",X"09",X"00",X"00",X"99",
		X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"99",
		X"00",X"00",X"0C",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"30",
		X"00",X"00",X"02",X"33",X"33",X"00",X"32",X"33",X"93",X"33",X"32",X"22",X"33",X"32",X"33",X"30",
		X"00",X"00",X"23",X"30",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"23",X"00",X"00",X"02",X"33",
		X"00",X"00",X"02",X"30",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"22",X"00",X"00",X"04",X"22",X"00",X"00",X"24",X"02",X"00",X"00",X"44",X"02",X"00",
		X"00",X"34",X"02",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"22",X"02",X"00",X"00",X"33",X"02",X"00",X"00",X"03",X"22",X"00",X"00",X"00",X"22",X"30",
		X"00",X"00",X"33",X"30",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"23",X"33",
		X"00",X"22",X"22",X"33",X"00",X"33",X"22",X"33",X"02",X"33",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"33",X"32",X"00",X"00",X"33",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"03",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",
		X"00",X"20",X"33",X"00",X"00",X"22",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"23",X"00",
		X"00",X"33",X"23",X"30",X"00",X"33",X"22",X"30",X"00",X"03",X"23",X"30",X"00",X"00",X"33",X"30",
		X"00",X"00",X"33",X"30",X"00",X"00",X"23",X"04",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"13",X"33",X"00",X"00",X"13",X"39",
		X"00",X"00",X"03",X"33",X"00",X"00",X"23",X"00",X"00",X"20",X"23",X"00",X"00",X"32",X"23",X"00",
		X"00",X"33",X"23",X"00",X"00",X"33",X"23",X"00",X"00",X"03",X"23",X"00",X"00",X"03",X"23",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"60",X"22",X"00",X"00",X"66",X"32",X"00",
		X"00",X"66",X"32",X"00",X"00",X"66",X"32",X"00",X"00",X"66",X"32",X"00",X"00",X"06",X"32",X"00",
		X"00",X"66",X"32",X"00",X"00",X"06",X"33",X"00",X"00",X"66",X"33",X"00",X"00",X"66",X"33",X"00",
		X"00",X"06",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"34",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"24",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"02",X"20",X"00",
		X"00",X"02",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"02",X"00",X"00",X"03",X"23",X"00",X"00",X"03",X"23",X"00",X"00",X"03",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"30",X"00",X"00",X"33",X"30",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"32",X"66",X"00",X"00",X"32",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"20",X"66",X"00",
		X"00",X"20",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"40",X"00",X"20",X"00",X"93",X"00",X"20",X"00",X"13",X"00",X"22",X"00",X"93",
		X"00",X"32",X"03",X"40",X"00",X"32",X"30",X"00",X"00",X"32",X"20",X"00",X"00",X"32",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"22",
		X"00",X"22",X"00",X"30",X"00",X"23",X"22",X"00",X"00",X"23",X"23",X"00",X"00",X"23",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"32",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"30",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"39",
		X"00",X"32",X"00",X"33",X"00",X"32",X"03",X"00",X"00",X"32",X"32",X"00",X"00",X"32",X"20",X"00",
		X"00",X"33",X"20",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"03",X"33",X"22",X"00",
		X"03",X"33",X"32",X"00",X"03",X"32",X"33",X"00",X"40",X"33",X"23",X"22",X"00",X"33",X"22",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"0C",X"99",
		X"00",X"00",X"C9",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"99",X"00",X"99",X"CC",
		X"09",X"00",X"00",X"C9",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"CC",X"00",X"99",X"00",X"C9",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"90",X"00",X"99",
		X"00",X"00",X"00",X"99",X"9C",X"00",X"09",X"99",X"C9",X"0C",X"99",X"00",X"C9",X"09",X"99",X"00",
		X"99",X"99",X"00",X"00",X"F9",X"99",X"09",X"00",X"FC",X"00",X"C9",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"80",X"00",
		X"00",X"88",X"88",X"00",X"08",X"88",X"88",X"00",X"08",X"88",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"88",X"88",X"00",X"88",X"85",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"C8",X"88",X"80",
		X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"CC",X"C8",X"88",X"88",X"99",X"88",X"88",
		X"88",X"5C",X"CC",X"88",X"88",X"88",X"89",X"88",X"88",X"58",X"88",X"88",X"88",X"98",X"88",X"88",
		X"88",X"C5",X"88",X"80",X"88",X"5C",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"88",X"88",X"00",X"08",X"88",X"88",X"00",X"08",X"88",X"88",X"00",X"00",X"88",X"88",X"00",
		X"00",X"88",X"80",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"FF",X"00",X"99",X"00",X"0F",X"00",X"B9",X"00",
		X"09",X"09",X"BB",X"00",X"09",X"99",X"9B",X"99",X"09",X"99",X"9B",X"99",X"09",X"99",X"9B",X"00",
		X"09",X"99",X"9B",X"00",X"09",X"99",X"9B",X"99",X"FF",X"09",X"9B",X"99",X"00",X"00",X"9B",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"DD",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"09",X"CC",X"00",X"00",X"90",X"9C",X"00",
		X"00",X"00",X"9C",X"00",X"00",X"00",X"F9",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"F0",X"00",
		X"00",X"09",X"00",X"00",X"00",X"90",X"C0",X"00",X"00",X"90",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"09",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"9C",X"00",
		X"00",X"00",X"9C",X"00",X"00",X"09",X"F9",X"00",X"00",X"99",X"90",X"00",X"00",X"90",X"F0",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"50",X"00",X"00",
		X"55",X"55",X"00",X"00",X"05",X"F5",X"00",X"00",X"05",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"22",X"00",X"00",X"04",X"22",X"00",X"00",X"94",X"02",X"00",X"00",X"44",X"02",X"00",
		X"00",X"94",X"02",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"22",X"02",X"00",X"00",X"99",X"02",X"00",X"00",X"09",X"22",X"00",X"00",X"00",X"22",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"29",X"99",
		X"00",X"22",X"22",X"99",X"00",X"99",X"22",X"99",X"02",X"99",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",
		X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",
		X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",X"99",X"99",X"99",X"EE",X"00",X"00",X"FF",X"EE",
		X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",
		X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",
		X"00",X"20",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"29",X"90",X"00",X"99",X"22",X"90",X"00",X"09",X"29",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"29",X"04",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"19",X"33",X"00",X"00",X"19",X"39",
		X"00",X"00",X"09",X"33",X"00",X"00",X"29",X"00",X"00",X"20",X"29",X"00",X"00",X"92",X"29",X"00",
		X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"29",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"60",X"22",X"00",X"00",X"66",X"92",X"00",
		X"00",X"66",X"92",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"92",X"00",X"00",X"06",X"92",X"00",
		X"00",X"66",X"92",X"00",X"00",X"06",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",
		X"00",X"06",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"94",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"02",X"20",X"00",
		X"00",X"02",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"02",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"20",X"66",X"00",
		X"00",X"20",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"40",X"00",X"20",X"00",X"93",X"00",X"20",X"00",X"13",X"00",X"22",X"00",X"93",
		X"00",X"92",X"09",X"40",X"00",X"92",X"90",X"00",X"00",X"92",X"20",X"00",X"00",X"92",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"22",
		X"00",X"22",X"00",X"90",X"00",X"29",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"33",X"00",X"99",X"00",X"39",
		X"00",X"92",X"00",X"33",X"00",X"92",X"09",X"00",X"00",X"92",X"92",X"00",X"00",X"92",X"20",X"00",
		X"00",X"99",X"20",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"22",X"00",
		X"09",X"99",X"92",X"00",X"09",X"92",X"99",X"00",X"40",X"99",X"29",X"22",X"00",X"99",X"22",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
