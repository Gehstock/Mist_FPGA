library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr2_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr2_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"C0",X"30",X"00",X"00",X"C0",X"70",X"00",X"00",X"C0",X"78",X"00",X"00",X"C4",X"3C",X"01",
		X"00",X"CC",X"3C",X"01",X"00",X"CC",X"79",X"00",X"00",X"C8",X"73",X"00",X"00",X"C0",X"77",X"00",
		X"00",X"80",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"53",X"00",X"00",X"88",X"21",X"00",X"00",X"88",X"21",X"00",X"00",X"88",X"21",X"00",X"00",
		X"88",X"21",X"00",X"00",X"88",X"21",X"00",X"00",X"88",X"21",X"00",X"00",X"00",X"53",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FD",X"10",X"00",X"CC",X"C4",X"30",X"00",
		X"66",X"E6",X"70",X"00",X"E6",X"F2",X"10",X"00",X"E2",X"F3",X"00",X"00",X"22",X"F3",X"00",X"00",
		X"22",X"F3",X"00",X"00",X"E2",X"F3",X"00",X"00",X"E6",X"F2",X"10",X"00",X"66",X"E6",X"70",X"00",
		X"CC",X"C4",X"30",X"00",X"88",X"FD",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"70",X"00",
		X"00",X"F0",X"30",X"00",X"00",X"F0",X"10",X"00",X"00",X"F0",X"00",X"00",X"00",X"70",X"00",X"10",
		X"00",X"30",X"80",X"10",X"00",X"10",X"C0",X"10",X"00",X"00",X"E0",X"10",X"00",X"00",X"F0",X"10",
		X"00",X"80",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2C",X"C3",X"00",X"00",X"E0",X"D2",X"30",X"00",X"2C",X"E1",X"70",X"01",
		X"E0",X"D2",X"10",X"01",X"2C",X"E1",X"30",X"01",X"E0",X"F0",X"70",X"01",X"2C",X"4B",X"10",X"01",
		X"E0",X"F0",X"10",X"01",X"2C",X"0F",X"70",X"01",X"E0",X"F0",X"10",X"01",X"2C",X"0F",X"30",X"01",
		X"68",X"E1",X"70",X"01",X"A4",X"D2",X"20",X"00",X"A4",X"D2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"70",X"00",
		X"10",X"FC",X"73",X"00",X"90",X"BE",X"73",X"00",X"F0",X"1F",X"73",X"00",X"90",X"BE",X"73",X"00",
		X"10",X"FC",X"FB",X"00",X"00",X"E0",X"F8",X"11",X"00",X"00",X"EE",X"11",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"FF",X"1F",X"01",X"CC",X"FF",X"13",X"01",X"EE",X"FF",X"13",X"01",X"EE",X"FF",X"3E",X"17",
		X"CC",X"F7",X"FE",X"0F",X"88",X"F7",X"FF",X"09",X"CC",X"F7",X"FF",X"09",X"EE",X"F7",X"FF",X"9F",
		X"EE",X"F7",X"FF",X"FF",X"CC",X"F7",X"FE",X"FF",X"88",X"FF",X"FE",X"FF",X"CC",X"FF",X"FE",X"77",
		X"EE",X"FF",X"FE",X"77",X"EE",X"FF",X"FE",X"33",X"CC",X"FF",X"FE",X"11",X"88",X"77",X"FC",X"00",
		X"CC",X"FF",X"77",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"F3",X"FF",X"17",X"CC",X"FB",X"FF",X"0F",
		X"88",X"FB",X"FF",X"09",X"88",X"F3",X"FF",X"09",X"CC",X"F7",X"FF",X"17",X"EE",X"F7",X"FF",X"33",
		X"EE",X"F7",X"FF",X"33",X"CC",X"F7",X"FF",X"17",X"88",X"F3",X"FF",X"09",X"88",X"FB",X"FF",X"09",
		X"CC",X"FB",X"FF",X"0F",X"EE",X"F3",X"FF",X"17",X"EE",X"FF",X"FF",X"00",X"CC",X"FF",X"77",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"11",X"EE",X"00",X"EE",X"FF",X"FF",X"17",X"EE",X"FF",X"FF",X"0F",
		X"CC",X"FB",X"FF",X"0D",X"88",X"F1",X"FF",X"0D",X"CC",X"B1",X"FE",X"17",X"EE",X"31",X"FE",X"33",
		X"EE",X"31",X"FE",X"33",X"CC",X"B1",X"FE",X"17",X"88",X"F1",X"FF",X"0D",X"CC",X"FB",X"FF",X"0D",
		X"EE",X"FF",X"FF",X"0F",X"EE",X"FF",X"FF",X"17",X"CC",X"11",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"33",X"00",X"00",X"CC",X"77",X"00",X"00",X"88",X"3E",X"00",X"00",X"CC",X"3E",X"00",X"00",
		X"CC",X"3A",X"00",X"00",X"88",X"3A",X"00",X"01",X"CC",X"3A",X"00",X"00",X"CC",X"3E",X"00",X"00",
		X"CC",X"76",X"00",X"00",X"CC",X"3E",X"00",X"00",X"88",X"3E",X"00",X"00",X"CC",X"3A",X"00",X"00",
		X"CC",X"3A",X"00",X"00",X"88",X"3A",X"00",X"01",X"CC",X"3E",X"00",X"00",X"CC",X"32",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"0F",X"07",X"00",X"2A",X"E1",X"3C",X"01",X"2E",X"F0",X"78",X"03",
		X"A6",X"F0",X"F8",X"13",X"A6",X"00",X"40",X"13",X"84",X"60",X"50",X"13",X"84",X"60",X"58",X"03",
		X"84",X"60",X"58",X"03",X"84",X"60",X"50",X"13",X"A6",X"E0",X"50",X"13",X"A6",X"E0",X"D8",X"13",
		X"2E",X"F0",X"78",X"03",X"2A",X"E1",X"3C",X"01",X"22",X"0F",X"07",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"0E",X"0F",X"00",X"44",X"C3",X"78",X"03",X"4C",X"E1",X"F0",X"07",
		X"4C",X"F0",X"F0",X"37",X"4C",X"FE",X"F7",X"26",X"4C",X"F2",X"F5",X"26",X"08",X"F2",X"F5",X"07",
		X"88",X"F2",X"F5",X"07",X"CC",X"F2",X"F5",X"26",X"6E",X"F2",X"F4",X"26",X"3B",X"F2",X"F4",X"37",
		X"19",X"E1",X"F0",X"07",X"11",X"C3",X"78",X"03",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"00",X"11",X"C3",X"78",X"03",X"19",X"E1",X"F0",X"07",
		X"3B",X"F0",X"F0",X"37",X"6E",X"FE",X"F7",X"04",X"CC",X"F2",X"F5",X"04",X"88",X"F2",X"F5",X"07",
		X"08",X"F2",X"F5",X"07",X"4C",X"F2",X"F5",X"04",X"4C",X"F2",X"F4",X"04",X"4C",X"F2",X"F4",X"37",
		X"4C",X"E1",X"F0",X"07",X"44",X"C3",X"78",X"03",X"44",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"0F",X"07",X"00",X"2A",X"E1",X"3C",X"01",X"2E",X"F0",X"78",X"03",
		X"A6",X"F0",X"F8",X"13",X"A6",X"E0",X"50",X"13",X"84",X"C0",X"40",X"13",X"84",X"90",X"68",X"03",
		X"84",X"30",X"78",X"03",X"84",X"50",X"60",X"13",X"A6",X"C0",X"40",X"13",X"A6",X"E0",X"D8",X"13",
		X"2E",X"F0",X"78",X"03",X"2A",X"E1",X"3C",X"01",X"22",X"0F",X"07",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"0E",X"0F",X"00",X"44",X"C3",X"78",X"03",X"4C",X"E1",X"F0",X"07",
		X"4C",X"F0",X"F0",X"37",X"4C",X"F2",X"F4",X"26",X"4C",X"F6",X"F6",X"26",X"08",X"FC",X"F2",X"07",
		X"88",X"F8",X"F1",X"07",X"CC",X"F4",X"F3",X"26",X"6E",X"F6",X"F6",X"26",X"3B",X"F2",X"F4",X"37",
		X"19",X"E1",X"F0",X"07",X"11",X"C3",X"78",X"03",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"00",X"11",X"C3",X"78",X"03",X"19",X"E1",X"F0",X"07",
		X"3B",X"F0",X"F0",X"37",X"6E",X"F2",X"F4",X"04",X"CC",X"F6",X"F6",X"04",X"88",X"FC",X"F2",X"07",
		X"08",X"F8",X"F1",X"07",X"4C",X"F4",X"F3",X"04",X"4C",X"F6",X"F6",X"04",X"4C",X"F2",X"F4",X"37",
		X"4C",X"E1",X"F0",X"07",X"44",X"C3",X"78",X"03",X"44",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"0F",X"07",X"00",X"2A",X"E1",X"3C",X"01",X"2E",X"F0",X"78",X"03",
		X"A6",X"F0",X"F8",X"13",X"A6",X"F0",X"50",X"13",X"84",X"F0",X"50",X"13",X"84",X"F0",X"58",X"03",
		X"84",X"00",X"48",X"03",X"84",X"F0",X"50",X"13",X"A6",X"F0",X"50",X"13",X"A6",X"F0",X"D8",X"13",
		X"2E",X"F0",X"78",X"03",X"2A",X"E1",X"3C",X"01",X"22",X"0F",X"07",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"0E",X"0F",X"00",X"44",X"C3",X"78",X"03",X"4C",X"E1",X"F0",X"07",
		X"4C",X"F0",X"F0",X"37",X"4C",X"F0",X"F4",X"26",X"4C",X"F0",X"F4",X"26",X"08",X"F0",X"F4",X"07",
		X"88",X"FE",X"F7",X"07",X"CC",X"F0",X"F4",X"26",X"6E",X"F0",X"F4",X"26",X"3B",X"F0",X"F4",X"37",
		X"19",X"E1",X"F0",X"07",X"11",X"C3",X"78",X"03",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"00",X"11",X"C3",X"78",X"03",X"19",X"E1",X"F0",X"07",
		X"3B",X"F0",X"F0",X"37",X"6E",X"F0",X"F4",X"04",X"CC",X"F0",X"F4",X"04",X"88",X"F0",X"F4",X"07",
		X"08",X"FE",X"F7",X"07",X"4C",X"F0",X"F4",X"04",X"4C",X"F0",X"F4",X"04",X"4C",X"F0",X"F4",X"37",
		X"4C",X"E1",X"F0",X"07",X"44",X"C3",X"78",X"03",X"44",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"0F",X"07",X"00",X"2A",X"E1",X"3C",X"01",X"2E",X"F0",X"78",X"03",
		X"A6",X"F0",X"F8",X"13",X"A6",X"00",X"40",X"13",X"84",X"B0",X"50",X"13",X"84",X"B0",X"58",X"03",
		X"84",X"B0",X"58",X"03",X"84",X"80",X"50",X"13",X"A6",X"20",X"40",X"13",X"A6",X"60",X"E8",X"13",
		X"2E",X"F0",X"78",X"03",X"2A",X"E1",X"3C",X"01",X"22",X"FF",X"07",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"0E",X"0F",X"00",X"44",X"C3",X"78",X"03",X"4C",X"E1",X"F0",X"07",
		X"4C",X"F0",X"F0",X"37",X"4C",X"FE",X"F7",X"26",X"4C",X"F8",X"F4",X"26",X"08",X"F8",X"F4",X"07",
		X"88",X"F8",X"F4",X"07",X"CC",X"FE",X"F4",X"26",X"6E",X"FA",X"F7",X"26",X"3B",X"F2",X"F3",X"37",
		X"19",X"E1",X"F0",X"07",X"11",X"C3",X"78",X"03",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"00",X"11",X"C3",X"78",X"03",X"19",X"E1",X"F0",X"07",
		X"3B",X"F0",X"F0",X"37",X"6E",X"FE",X"F7",X"04",X"CC",X"F8",X"F4",X"04",X"88",X"F8",X"F4",X"07",
		X"08",X"F8",X"F4",X"07",X"4C",X"FE",X"F4",X"04",X"4C",X"FA",X"F7",X"04",X"4C",X"F2",X"F3",X"37",
		X"4C",X"E1",X"F0",X"07",X"44",X"C3",X"78",X"03",X"44",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"0F",X"07",X"00",X"2A",X"E1",X"3C",X"01",X"2E",X"F0",X"78",X"03",
		X"A6",X"F0",X"F8",X"13",X"A6",X"00",X"70",X"13",X"84",X"50",X"60",X"13",X"84",X"D0",X"48",X"03",
		X"84",X"D0",X"58",X"03",X"84",X"D0",X"40",X"13",X"A6",X"50",X"60",X"13",X"A6",X"00",X"F8",X"13",
		X"2E",X"F0",X"78",X"03",X"2A",X"E1",X"3C",X"01",X"22",X"0F",X"07",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"0E",X"0F",X"00",X"44",X"C3",X"78",X"03",X"4C",X"E1",X"F0",X"07",
		X"4C",X"F0",X"F0",X"37",X"4C",X"FE",X"F1",X"26",X"4C",X"F4",X"F3",X"26",X"08",X"F4",X"F6",X"07",
		X"88",X"F4",X"F4",X"07",X"CC",X"F4",X"F6",X"26",X"6E",X"F4",X"F3",X"26",X"3B",X"FE",X"F1",X"37",
		X"19",X"E1",X"F0",X"07",X"11",X"C3",X"78",X"03",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"00",X"11",X"C3",X"78",X"03",X"19",X"E1",X"F0",X"07",
		X"3B",X"F0",X"F0",X"37",X"6E",X"FE",X"F1",X"04",X"CC",X"F4",X"F3",X"04",X"88",X"F4",X"F6",X"37",
		X"08",X"F4",X"F4",X"37",X"4C",X"F4",X"F6",X"04",X"4C",X"F4",X"F3",X"04",X"4C",X"FE",X"F1",X"37",
		X"4C",X"E1",X"F0",X"07",X"44",X"C3",X"78",X"03",X"44",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"4C",X"3C",X"00",X"00",X"4C",X"7C",X"00",X"00",X"4C",X"7C",X"00",X"00",
		X"4C",X"7C",X"00",X"00",X"4C",X"38",X"00",X"00",X"4C",X"38",X"00",X"00",X"08",X"3C",X"00",X"00",
		X"08",X"3C",X"00",X"00",X"4C",X"38",X"00",X"00",X"4C",X"38",X"00",X"00",X"4C",X"7C",X"00",X"00",
		X"4C",X"7C",X"00",X"00",X"4C",X"7C",X"00",X"00",X"4C",X"3C",X"00",X"00",X"08",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"10",X"00",X"00",X"F3",X"F0",X"10",X"88",X"F1",X"F0",X"30",
		X"CC",X"F1",X"F0",X"70",X"CC",X"F0",X"F0",X"70",X"CC",X"F3",X"F0",X"52",X"CC",X"F1",X"78",X"61",
		X"C4",X"F0",X"78",X"77",X"EE",X"96",X"78",X"FC",X"EE",X"96",X"4B",X"B8",X"E6",X"B4",X"87",X"21",
		X"CC",X"F0",X"87",X"30",X"88",X"F1",X"D2",X"10",X"00",X"F0",X"F0",X"10",X"00",X"C0",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",X"88",X"F1",X"F0",X"10",X"CC",X"F0",X"F0",X"30",
		X"EE",X"F0",X"F0",X"30",X"E6",X"F0",X"F0",X"21",X"EE",X"F1",X"78",X"30",X"EE",X"F0",X"78",X"FF",
		X"E6",X"F0",X"78",X"B8",X"EE",X"96",X"4B",X"30",X"EE",X"96",X"87",X"21",X"E6",X"B4",X"87",X"30",
		X"CC",X"F0",X"D2",X"30",X"88",X"F1",X"F0",X"10",X"00",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"70",X"00",X"00",X"F0",X"F0",X"10",X"CC",X"F0",X"F0",X"10",X"C4",X"F0",X"F0",X"21",
		X"EE",X"F0",X"78",X"30",X"E6",X"F0",X"78",X"FF",X"EE",X"F1",X"78",X"B9",X"CC",X"F0",X"78",X"30",
		X"C4",X"F0",X"C3",X"61",X"CC",X"3C",X"1E",X"70",X"CC",X"3D",X"1E",X"70",X"CC",X"78",X"B4",X"30",
		X"88",X"F1",X"F0",X"30",X"00",X"F3",X"F0",X"10",X"00",X"C0",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",
		X"88",X"F1",X"F0",X"10",X"CC",X"F0",X"F0",X"30",X"EE",X"F0",X"F0",X"30",X"E6",X"F0",X"F0",X"21",
		X"EE",X"F1",X"78",X"30",X"EE",X"F0",X"78",X"33",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"F0",X"78",X"30",X"EE",X"96",X"4B",X"30",
		X"EE",X"96",X"87",X"21",X"E6",X"B4",X"87",X"30",X"CC",X"F0",X"D2",X"30",X"88",X"F1",X"F0",X"10",
		X"00",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"C0",X"F0",X"30",X"00",X"E0",X"F0",X"30",X"88",X"F1",X"F0",X"52",X"88",X"F0",X"F0",X"61",
		X"CC",X"F1",X"F0",X"61",X"CC",X"F1",X"F0",X"01",X"CC",X"F7",X"78",X"00",X"88",X"F3",X"0F",X"33",
		X"88",X"11",X"00",X"EE",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"11",X"00",X"00",
		X"88",X"71",X"00",X"00",X"CC",X"F3",X"10",X"00",X"CC",X"3D",X"61",X"00",X"CC",X"3C",X"96",X"01",
		X"88",X"78",X"96",X"61",X"88",X"F1",X"87",X"61",X"00",X"F0",X"96",X"21",X"00",X"E0",X"F0",X"30",
		X"00",X"80",X"F0",X"10",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"96",X"01",X"00",X"C0",X"9E",X"01",X"00",X"E0",X"9E",X"01",X"00",X"E0",X"9E",X"01",X"00",
		X"E0",X"DE",X"11",X"00",X"E0",X"9E",X"01",X"00",X"E0",X"1E",X"01",X"00",X"E0",X"1E",X"01",X"00",
		X"E0",X"1E",X"01",X"00",X"C4",X"1E",X"01",X"00",X"CC",X"1E",X"01",X"00",X"88",X"3F",X"01",X"00",
		X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",
		X"88",X"3F",X"01",X"00",X"CC",X"1E",X"01",X"00",X"C4",X"1E",X"01",X"00",X"E0",X"1E",X"01",X"00",
		X"E0",X"1E",X"01",X"00",X"E0",X"1E",X"01",X"00",X"E0",X"9E",X"01",X"00",X"E0",X"DE",X"11",X"00",
		X"E0",X"9E",X"01",X"00",X"E0",X"9E",X"01",X"00",X"C0",X"9E",X"01",X"00",X"80",X"96",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8C",X"01",X"00",X"00",X"CE",X"33",X"00",X"00",X"EE",X"37",X"00",
		X"00",X"CE",X"77",X"00",X"00",X"CC",X"37",X"00",X"00",X"08",X"13",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8C",X"01",X"00",X"00",X"CE",X"13",X"00",X"00",X"EE",X"33",X"00",
		X"00",X"EE",X"33",X"00",X"00",X"EE",X"33",X"00",X"00",X"CE",X"13",X"00",X"00",X"8C",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CE",X"13",X"00",X"00",X"EF",X"37",X"00",X"00",X"FF",X"77",X"00",
		X"00",X"EF",X"37",X"00",X"00",X"CE",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"08",X"02",X"00",
		X"00",X"8C",X"72",X"00",X"00",X"CE",X"C6",X"00",X"00",X"E3",X"B9",X"00",X"88",X"F1",X"4E",X"00",
		X"80",X"FE",X"51",X"00",X"00",X"ED",X"B2",X"00",X"00",X"C2",X"8D",X"00",X"00",X"84",X"35",X"00",
		X"00",X"08",X"22",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"08",X"13",X"00",
		X"00",X"8C",X"24",X"00",X"00",X"CE",X"59",X"00",X"00",X"E3",X"D6",X"00",X"88",X"F1",X"51",X"00",
		X"80",X"FE",X"BE",X"00",X"00",X"ED",X"6D",X"00",X"00",X"C2",X"A2",X"00",X"00",X"84",X"12",X"00",
		X"00",X"08",X"31",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"88",X"21",X"00",
		X"00",X"C4",X"55",X"00",X"00",X"E2",X"A9",X"00",X"00",X"3D",X"26",X"00",X"80",X"1E",X"A5",X"00",
		X"08",X"E1",X"4E",X"00",X"00",X"D3",X"9D",X"00",X"00",X"2E",X"52",X"00",X"00",X"4C",X"62",X"00",
		X"00",X"88",X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"C2",X"90",X"F0",X"00",X"42",X"F0",X"80",X"10",
		X"42",X"00",X"00",X"10",X"42",X"EE",X"00",X"10",X"42",X"EE",X"03",X"10",X"40",X"6E",X"04",X"10",
		X"42",X"6E",X"04",X"10",X"42",X"66",X"03",X"10",X"C2",X"66",X"00",X"10",X"82",X"70",X"80",X"10",
		X"02",X"C0",X"C0",X"00",X"00",X"80",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"07",X"00",X"08",X"03",X"0C",X"01",X"0C",X"00",X"00",X"03",
		X"04",X"00",X"66",X"02",X"06",X"54",X"FF",X"06",X"02",X"FE",X"FF",X"04",X"02",X"EE",X"99",X"15",
		X"02",X"EE",X"FF",X"15",X"02",X"FE",X"99",X"04",X"06",X"54",X"FF",X"06",X"04",X"00",X"66",X"02",
		X"0C",X"00",X"00",X"03",X"08",X"03",X"0C",X"01",X"00",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"06",X"10",X"00",X"00",X"00",X"20",X"00",
		X"00",X"06",X"40",X"00",X"00",X"0F",X"80",X"00",X"00",X"0F",X"10",X"10",X"00",X"06",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"10",X"00",X"00",X"3C",X"30",X"00",X"00",X"1E",X"21",X"00",X"00",X"1E",X"21",X"00",X"00",
		X"3C",X"30",X"00",X"00",X"E0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"88",X"BF",X"8F",X"11",X"88",X"DF",X"AF",X"11",X"88",X"DF",X"AF",X"11",
		X"88",X"3F",X"FF",X"11",X"88",X"FF",X"FF",X"11",X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",
		X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",X"88",X"FF",X"FF",X"11",X"88",X"3F",X"CF",X"11",
		X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",X"00",X"FF",X"FF",X"00",
		X"88",X"FF",X"FF",X"11",X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",
		X"88",X"3F",X"CF",X"11",X"88",X"FF",X"FF",X"11",X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",
		X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",X"88",X"FF",X"FF",X"11",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"88",X"FF",X"FF",X"11",X"88",X"FF",X"FF",X"11",X"88",X"DF",X"DF",X"11",
		X"88",X"1F",X"8F",X"11",X"88",X"DF",X"FF",X"11",X"88",X"FF",X"FF",X"11",X"88",X"FF",X"FF",X"11",
		X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"88",X"FF",X"FF",X"11",X"88",X"9F",X"DF",X"11",X"88",X"5F",X"BF",X"11",
		X"88",X"5F",X"BF",X"11",X"88",X"5F",X"BF",X"11",X"88",X"DF",X"CF",X"11",X"88",X"FF",X"FF",X"11",
		X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"88",X"FF",X"FF",X"11",X"88",X"3F",X"FF",X"11",X"88",X"BF",X"EF",X"11",
		X"88",X"BF",X"DF",X"11",X"88",X"1F",X"8F",X"11",X"88",X"BF",X"FF",X"11",X"88",X"FF",X"FF",X"11",
		X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"88",X"FF",X"FF",X"11",X"88",X"3F",X"CF",X"11",X"88",X"DF",X"AF",X"11",
		X"88",X"DF",X"AF",X"11",X"88",X"DF",X"AF",X"11",X"88",X"3F",X"FF",X"11",X"88",X"FF",X"FF",X"11",
		X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"88",X"FF",X"FF",X"11",X"88",X"3F",X"DF",X"11",X"88",X"DF",X"AF",X"11",
		X"88",X"DF",X"AF",X"11",X"88",X"DF",X"AF",X"11",X"88",X"3F",X"DF",X"11",X"88",X"FF",X"FF",X"11",
		X"88",X"3F",X"CF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"DF",X"BF",X"11",X"88",X"3F",X"CF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"00",X"F0",X"F0",X"00",
		X"80",X"F0",X"F0",X"10",X"80",X"F0",X"F0",X"10",X"C0",X"F0",X"F0",X"30",X"C0",X"F0",X"F0",X"30",
		X"C0",X"F0",X"F0",X"30",X"C0",X"F0",X"F0",X"30",X"80",X"F0",X"F0",X"10",X"80",X"F0",X"F0",X"10",
		X"00",X"F0",X"F0",X"00",X"00",X"C0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"33",X"00",X"00",X"6E",X"67",X"00",X"00",X"3F",X"CF",X"00",X"00",X"1F",X"8F",X"00",X"00",
		X"1F",X"8F",X"00",X"00",X"3F",X"CF",X"00",X"00",X"6E",X"67",X"00",X"00",X"CC",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"82",X"13",X"6D",X"10",X"86",X"DB",X"6D",X"32",
		X"82",X"DB",X"6D",X"32",X"82",X"DB",X"6D",X"32",X"82",X"DB",X"2D",X"32",X"80",X"DB",X"0F",X"32",
		X"82",X"DB",X"09",X"32",X"86",X"DB",X"09",X"32",X"82",X"DB",X"0F",X"32",X"02",X"9B",X"6D",X"32",
		X"02",X"88",X"6D",X"10",X"00",X"00",X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"8A",X"21",X"B6",X"11",X"8E",X"6D",X"B6",X"13",
		X"8A",X"6D",X"B6",X"13",X"8A",X"6D",X"3E",X"13",X"8A",X"6D",X"3E",X"13",X"88",X"6D",X"E1",X"13",
		X"8A",X"6D",X"18",X"13",X"8E",X"6D",X"18",X"13",X"8A",X"6D",X"96",X"13",X"02",X"29",X"B6",X"13",
		X"02",X"08",X"B6",X"11",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"0A",X"23",X"DB",X"01",X"0E",X"B6",X"DB",X"21",
		X"0A",X"B6",X"DB",X"21",X"0A",X"B6",X"5B",X"21",X"0A",X"B6",X"1F",X"21",X"08",X"B6",X"1F",X"21",
		X"0A",X"B6",X"19",X"21",X"0E",X"B6",X"19",X"21",X"0A",X"B6",X"9F",X"21",X"02",X"B2",X"DB",X"21",
		X"02",X"80",X"DB",X"01",X"00",X"00",X"DB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"00",X"C0",X"F0",X"F0",X"10",
		X"0C",X"0F",X"0F",X"03",X"CC",X"3F",X"8C",X"33",X"C0",X"78",X"84",X"30",X"0C",X"0F",X"0F",X"03",
		X"88",X"FF",X"FF",X"11",X"80",X"F0",X"70",X"00",X"0C",X"0F",X"0F",X"00",X"EE",X"FF",X"FF",X"00",
		X"C0",X"F0",X"70",X"00",X"08",X"00",X"02",X"00",X"0C",X"07",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"00",X"CC",X"FF",X"FF",X"11",
		X"C0",X"1E",X"C3",X"30",X"0C",X"0F",X"0C",X"03",X"CC",X"7F",X"8C",X"33",X"C0",X"F0",X"F0",X"30",
		X"08",X"0F",X"0F",X"01",X"88",X"FF",X"77",X"00",X"C0",X"F0",X"F0",X"00",X"0E",X"0F",X"0F",X"00",
		X"CC",X"FF",X"77",X"00",X"08",X"00",X"02",X"00",X"0C",X"07",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F0",X"00",X"0C",X"0F",X"0F",X"01",
		X"CC",X"1F",X"CF",X"33",X"C0",X"3C",X"84",X"30",X"0C",X"0F",X"0C",X"03",X"CC",X"FF",X"FF",X"33",
		X"80",X"F0",X"F0",X"10",X"08",X"0F",X"07",X"00",X"CC",X"FF",X"FF",X"00",X"E0",X"F0",X"F0",X"00",
		X"0C",X"0F",X"07",X"00",X"08",X"00",X"02",X"00",X"0C",X"07",X"0F",X"01",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
