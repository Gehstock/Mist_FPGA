library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gravitar_pgm_rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gravitar_pgm_rom1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"A9",X"16",X"85",X"00",X"85",X"01",X"A9",X"08",X"85",X"EB",X"85",X"EC",X"A9",X"00",X"85",X"D0",
		X"85",X"4F",X"20",X"2D",X"DE",X"20",X"9E",X"CB",X"20",X"C2",X"E1",X"20",X"A6",X"CA",X"A9",X"00",
		X"85",X"F2",X"20",X"36",X"90",X"20",X"97",X"90",X"20",X"72",X"CD",X"AD",X"00",X"78",X"29",X"10",
		X"D0",X"EC",X"4C",X"8B",X"ED",X"A9",X"A6",X"CF",X"B5",X"00",X"AA",X"A5",X"FA",X"10",X"0B",X"BD",
		X"7A",X"90",X"48",X"BD",X"79",X"90",X"48",X"4C",X"52",X"90",X"BD",X"54",X"90",X"48",X"BD",X"53",
		X"90",X"48",X"60",X"51",X"50",X"FF",X"4F",X"91",X"53",X"BD",X"57",X"D3",X"93",X"ED",X"50",X"58",
		X"51",X"06",X"52",X"A2",X"92",X"B4",X"92",X"7B",X"93",X"5A",X"55",X"F2",X"91",X"0B",X"93",X"4A",
		X"92",X"13",X"CB",X"34",X"94",X"A8",X"94",X"01",X"95",X"51",X"50",X"FF",X"4F",X"91",X"53",X"BD",
		X"57",X"21",X"91",X"ED",X"50",X"58",X"51",X"06",X"52",X"A2",X"92",X"B4",X"92",X"7B",X"93",X"5A",
		X"55",X"75",X"91",X"0B",X"93",X"B5",X"91",X"A6",X"CF",X"E6",X"4F",X"A5",X"D0",X"D0",X"3B",X"A5",
		X"F1",X"29",X"03",X"D0",X"04",X"A9",X"02",X"85",X"D6",X"A0",X"FF",X"A5",X"D6",X"F0",X"17",X"C9",
		X"02",X"A5",X"1D",X"90",X"09",X"29",X"40",X"F0",X"05",X"A0",X"02",X"4C",X"C6",X"90",X"A5",X"1D",
		X"29",X"20",X"F0",X"02",X"A0",X"00",X"98",X"30",X"0E",X"95",X"00",X"24",X"F9",X"30",X"08",X"A9",
		X"FF",X"85",X"F9",X"A9",X"04",X"85",X"FC",X"4C",X"E0",X"90",X"24",X"F9",X"30",X"02",X"C6",X"F9",
		X"60",X"A9",X"FF",X"85",X"FA",X"A9",X"01",X"8D",X"00",X"20",X"A9",X"E2",X"8D",X"01",X"20",X"A9",
		X"20",X"8D",X"03",X"20",X"8D",X"03",X"24",X"A9",X"00",X"85",X"00",X"A9",X"00",X"85",X"EB",X"20",
		X"C2",X"E1",X"E6",X"4F",X"A5",X"42",X"C9",X"01",X"B0",X"04",X"A9",X"01",X"85",X"42",X"A9",X"00",
		X"85",X"F2",X"20",X"36",X"90",X"20",X"72",X"CD",X"AD",X"00",X"78",X"29",X"10",X"F0",X"E3",X"4C",
		X"3A",X"E8",X"20",X"07",X"C7",X"20",X"D1",X"98",X"20",X"60",X"9F",X"A5",X"88",X"F0",X"1B",X"20",
		X"98",X"95",X"20",X"64",X"97",X"20",X"7E",X"98",X"20",X"11",X"97",X"20",X"3D",X"C4",X"20",X"E8",
		X"A0",X"20",X"D2",X"BE",X"20",X"B2",X"BD",X"20",X"30",X"BE",X"20",X"EE",X"C4",X"20",X"D9",X"9D",
		X"20",X"05",X"9E",X"20",X"7E",X"9C",X"20",X"B1",X"9C",X"20",X"A6",X"BF",X"20",X"BE",X"BC",X"20",
		X"2F",X"BC",X"20",X"D5",X"C3",X"20",X"6F",X"C8",X"20",X"85",X"C0",X"20",X"72",X"C9",X"20",X"12",
		X"9C",X"A9",X"02",X"85",X"EB",X"60",X"A9",X"01",X"85",X"CE",X"A5",X"88",X"F0",X"18",X"20",X"D1",
		X"98",X"20",X"98",X"95",X"20",X"A7",X"97",X"20",X"11",X"97",X"20",X"3D",X"C4",X"20",X"E5",X"C1",
		X"20",X"9F",X"BB",X"20",X"B3",X"C0",X"20",X"63",X"9C",X"20",X"33",X"9B",X"20",X"8E",X"C5",X"20",
		X"D5",X"C3",X"20",X"30",X"BE",X"20",X"07",X"C7",X"20",X"6F",X"C8",X"20",X"85",X"C0",X"20",X"3E",
		X"9C",X"A9",X"0A",X"85",X"EB",X"60",X"A9",X"01",X"85",X"CE",X"A9",X"60",X"85",X"30",X"A5",X"88",
		X"F0",X"0F",X"20",X"98",X"95",X"20",X"7E",X"98",X"20",X"11",X"97",X"20",X"D1",X"98",X"20",X"3D",
		X"C4",X"A6",X"86",X"20",X"3C",X"9B",X"20",X"04",X"9D",X"20",X"9E",X"C5",X"20",X"F3",X"BB",X"20",
		X"07",X"C7",X"20",X"7B",X"BF",X"20",X"6F",X"C8",X"20",X"85",X"C0",X"20",X"3E",X"9C",X"A9",X"0A",
		X"85",X"EB",X"60",X"A9",X"01",X"85",X"CE",X"A6",X"CF",X"B5",X"88",X"F0",X"1B",X"20",X"D1",X"98",
		X"20",X"98",X"95",X"20",X"A7",X"97",X"20",X"11",X"97",X"20",X"3D",X"C4",X"20",X"E5",X"C1",X"20",
		X"62",X"BC",X"20",X"76",X"96",X"20",X"B3",X"C0",X"20",X"9F",X"BB",X"20",X"63",X"9C",X"20",X"33",
		X"9B",X"20",X"8E",X"C5",X"20",X"D5",X"C3",X"20",X"30",X"BE",X"20",X"07",X"C7",X"20",X"6F",X"C8",
		X"20",X"85",X"C0",X"20",X"3E",X"9C",X"A5",X"F0",X"29",X"C0",X"C9",X"C0",X"F0",X"06",X"A9",X"02",
		X"05",X"F5",X"85",X"F5",X"A6",X"CF",X"A9",X"0A",X"95",X"EB",X"60",X"A9",X"01",X"85",X"CE",X"A9",
		X"60",X"85",X"30",X"A6",X"CF",X"B5",X"88",X"F0",X"0F",X"20",X"98",X"95",X"20",X"7E",X"98",X"20",
		X"11",X"97",X"20",X"D1",X"98",X"20",X"3D",X"C4",X"A6",X"86",X"20",X"3C",X"9B",X"20",X"04",X"9D",
		X"20",X"9E",X"C5",X"20",X"F3",X"BB",X"20",X"62",X"BB",X"20",X"07",X"C7",X"20",X"62",X"BC",X"20",
		X"76",X"96",X"20",X"7B",X"BF",X"20",X"6F",X"C8",X"20",X"85",X"C0",X"20",X"3E",X"9C",X"A5",X"F0",
		X"29",X"C0",X"C9",X"C0",X"F0",X"06",X"A9",X"02",X"05",X"F5",X"85",X"F5",X"A6",X"CF",X"A9",X"0A",
		X"95",X"EB",X"60",X"20",X"C8",X"C9",X"20",X"CC",X"92",X"20",X"E6",X"E4",X"A9",X"00",X"85",X"D0",
		X"85",X"FC",X"85",X"F9",X"60",X"AD",X"6D",X"04",X"10",X"11",X"A0",X"FF",X"84",X"30",X"A6",X"CF",
		X"AC",X"6C",X"04",X"B9",X"6F",X"04",X"95",X"00",X"20",X"D7",X"51",X"60",X"A5",X"D0",X"F8",X"A2",
		X"02",X"BD",X"63",X"01",X"18",X"6D",X"57",X"04",X"8D",X"57",X"04",X"BD",X"65",X"01",X"6D",X"58",
		X"04",X"8D",X"58",X"04",X"AD",X"59",X"04",X"69",X"00",X"8D",X"59",X"04",X"CA",X"D0",X"E2",X"D8",
		X"AD",X"4E",X"04",X"18",X"6D",X"54",X"04",X"8D",X"54",X"04",X"AD",X"4F",X"04",X"6D",X"55",X"04",
		X"8D",X"55",X"04",X"AD",X"56",X"04",X"69",X"00",X"8D",X"56",X"04",X"60",X"A5",X"30",X"48",X"C9",
		X"FF",X"D0",X"03",X"20",X"0B",X"E1",X"68",X"C9",X"80",X"90",X"1B",X"20",X"6F",X"C8",X"C6",X"30",
		X"A9",X"00",X"85",X"F5",X"A6",X"CF",X"BD",X"7A",X"01",X"C9",X"01",X"D0",X"06",X"A9",X"01",X"05",
		X"F5",X"85",X"F5",X"4C",X"6B",X"93",X"A6",X"CF",X"B5",X"F6",X"29",X"01",X"D0",X"06",X"20",X"F3",
		X"53",X"4C",X"47",X"93",X"20",X"04",X"54",X"A9",X"07",X"8D",X"38",X"01",X"A9",X"F9",X"8D",X"39",
		X"01",X"A9",X"01",X"85",X"28",X"85",X"29",X"A9",X"18",X"95",X"00",X"BD",X"7A",X"01",X"C9",X"01",
		X"D0",X"09",X"A9",X"FE",X"25",X"F5",X"85",X"F5",X"FE",X"7A",X"01",X"A6",X"CF",X"A9",X"0C",X"95",
		X"EB",X"60",X"A9",X"00",X"A2",X"05",X"95",X"12",X"CA",X"10",X"FB",X"60",X"A5",X"30",X"A0",X"01",
		X"A6",X"CF",X"B5",X"4D",X"AA",X"A5",X"30",X"DD",X"B6",X"93",X"90",X"05",X"C6",X"30",X"4C",X"A0",
		X"93",X"A5",X"D0",X"D0",X"05",X"A9",X"24",X"4C",X"9C",X"93",X"A9",X"08",X"A6",X"CF",X"95",X"00",
		X"88",X"10",X"DD",X"A9",X"EB",X"25",X"F4",X"85",X"F4",X"A9",X"FD",X"25",X"F5",X"85",X"F5",X"A6",
		X"CF",X"A9",X"06",X"95",X"EB",X"60",X"81",X"81",X"81",X"64",X"60",X"81",X"81",X"81",X"50",X"60",
		X"81",X"81",X"70",X"81",X"60",X"02",X"02",X"02",X"03",X"03",X"02",X"02",X"02",X"03",X"03",X"02",
		X"02",X"03",X"02",X"03",X"20",X"07",X"C7",X"20",X"D1",X"98",X"20",X"60",X"9F",X"A6",X"CF",X"B5",
		X"88",X"F0",X"21",X"20",X"98",X"95",X"20",X"64",X"97",X"20",X"7E",X"98",X"20",X"11",X"97",X"20",
		X"3D",X"C4",X"20",X"E8",X"A0",X"20",X"D2",X"BE",X"20",X"62",X"BC",X"20",X"B2",X"BD",X"20",X"94",
		X"BB",X"20",X"30",X"BE",X"20",X"EE",X"C4",X"20",X"D9",X"9D",X"20",X"05",X"9E",X"20",X"7E",X"9C",
		X"20",X"B1",X"9C",X"20",X"A6",X"BF",X"20",X"BE",X"BC",X"20",X"2F",X"BC",X"20",X"D5",X"C3",X"20",
		X"76",X"96",X"20",X"6F",X"C8",X"20",X"85",X"C0",X"20",X"72",X"C9",X"20",X"12",X"9C",X"A6",X"CF",
		X"A9",X"02",X"95",X"EB",X"60",X"A9",X"38",X"85",X"0F",X"A2",X"FF",X"86",X"10",X"E8",X"8E",X"36",
		X"01",X"8D",X"37",X"01",X"86",X"0D",X"86",X"0E",X"86",X"1E",X"86",X"4B",X"8E",X"44",X"01",X"8E",
		X"6E",X"04",X"8E",X"7D",X"01",X"8E",X"7E",X"01",X"86",X"F5",X"A9",X"A0",X"8D",X"7C",X"01",X"A9",
		X"04",X"85",X"27",X"85",X"11",X"85",X"4C",X"86",X"EE",X"86",X"CF",X"86",X"F6",X"8E",X"3C",X"01",
		X"85",X"28",X"85",X"29",X"A9",X"06",X"8D",X"38",X"01",X"A9",X"FA",X"8D",X"39",X"01",X"A9",X"02",
		X"85",X"49",X"85",X"E3",X"20",X"1D",X"DE",X"20",X"19",X"54",X"20",X"72",X"93",X"20",X"67",X"54",
		X"20",X"A9",X"50",X"A9",X"80",X"85",X"30",X"A9",X"01",X"85",X"CE",X"AD",X"BE",X"59",X"85",X"18",
		X"A9",X"22",X"85",X"00",X"A9",X"10",X"95",X"EB",X"60",X"20",X"E7",X"98",X"20",X"B1",X"95",X"20",
		X"07",X"C7",X"20",X"64",X"97",X"20",X"B3",X"C0",X"20",X"63",X"9C",X"20",X"8E",X"C5",X"20",X"33",
		X"9B",X"20",X"D5",X"C3",X"20",X"82",X"95",X"A9",X"14",X"20",X"63",X"95",X"85",X"F4",X"A9",X"80",
		X"05",X"F2",X"85",X"F2",X"A9",X"10",X"85",X"EB",X"60",X"CE",X"7C",X"01",X"D0",X"13",X"AC",X"7E",
		X"01",X"C8",X"B9",X"F1",X"94",X"8D",X"7D",X"01",X"B9",X"F9",X"94",X"8D",X"7C",X"01",X"8C",X"7E",
		X"01",X"60",X"08",X"01",X"04",X"00",X"02",X"08",X"01",X"00",X"04",X"02",X"20",X"20",X"36",X"0E",
		X"01",X"FF",X"20",X"07",X"C7",X"A5",X"88",X"F0",X"3C",X"20",X"D9",X"94",X"20",X"E7",X"98",X"20",
		X"60",X"9F",X"20",X"65",X"96",X"20",X"64",X"97",X"20",X"7E",X"98",X"20",X"6F",X"95",X"20",X"3A",
		X"97",X"20",X"E8",X"A0",X"20",X"E3",X"C4",X"20",X"25",X"BF",X"20",X"62",X"BC",X"20",X"EE",X"C4",
		X"20",X"D9",X"9D",X"20",X"05",X"9E",X"20",X"D5",X"C3",X"20",X"7E",X"9C",X"20",X"B1",X"9C",X"20",
		X"A6",X"BF",X"20",X"BE",X"BC",X"20",X"6F",X"C8",X"20",X"85",X"C0",X"A9",X"7F",X"25",X"F2",X"85",
		X"F2",X"A9",X"60",X"20",X"63",X"95",X"85",X"F4",X"20",X"72",X"C9",X"20",X"82",X"95",X"A9",X"12",
		X"85",X"EB",X"60",X"A6",X"D6",X"F0",X"05",X"09",X"08",X"4C",X"6E",X"95",X"29",X"F7",X"60",X"AD",
		X"7D",X"01",X"29",X"04",X"F0",X"02",X"C6",X"11",X"AD",X"7D",X"01",X"29",X"08",X"F0",X"02",X"E6",
		X"11",X"60",X"A5",X"00",X"A8",X"C9",X"08",X"D0",X"02",X"A0",X"24",X"C9",X"0A",X"D0",X"02",X"A0",
		X"16",X"84",X"00",X"A9",X"FF",X"85",X"3F",X"60",X"A9",X"00",X"85",X"4C",X"A5",X"1D",X"29",X"10",
		X"D0",X"01",X"60",X"18",X"F8",X"A5",X"48",X"69",X"06",X"85",X"48",X"D8",X"85",X"4C",X"20",X"EF",
		X"E0",X"A5",X"11",X"29",X"0F",X"A8",X"A5",X"1E",X"4A",X"4A",X"B0",X"06",X"B9",X"54",X"97",X"4C",
		X"C5",X"95",X"B9",X"44",X"97",X"85",X"1A",X"A5",X"28",X"85",X"19",X"20",X"6E",X"DE",X"A4",X"1E",
		X"46",X"1C",X"66",X"1B",X"46",X"1C",X"66",X"1B",X"46",X"1C",X"66",X"1B",X"A5",X"1B",X"59",X"55",
		X"96",X"85",X"1B",X"A5",X"1C",X"59",X"55",X"96",X"85",X"1C",X"A5",X"17",X"18",X"65",X"1B",X"85",
		X"17",X"A5",X"16",X"65",X"1C",X"85",X"16",X"10",X"05",X"A9",X"FF",X"4C",X"00",X"96",X"A9",X"00",
		X"85",X"15",X"98",X"4A",X"4A",X"A5",X"11",X"29",X"0F",X"A8",X"B0",X"06",X"B9",X"44",X"97",X"4C",
		X"15",X"96",X"B9",X"54",X"97",X"85",X"1A",X"A5",X"29",X"85",X"19",X"20",X"6E",X"DE",X"A4",X"1E",
		X"46",X"1C",X"66",X"1B",X"46",X"1C",X"66",X"1B",X"46",X"1C",X"66",X"1B",X"A5",X"1B",X"59",X"5D",
		X"96",X"85",X"1B",X"A5",X"1C",X"59",X"5D",X"96",X"85",X"1C",X"A5",X"14",X"18",X"65",X"1B",X"85",
		X"14",X"A5",X"13",X"65",X"1C",X"85",X"13",X"10",X"05",X"A9",X"FF",X"4C",X"50",X"96",X"A9",X"00",
		X"85",X"12",X"4C",X"D3",X"96",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"A9",X"00",X"85",X"4C",X"AD",X"7D",X"01",X"29",X"02",X"F0",X"05",
		X"85",X"4C",X"4C",X"B1",X"95",X"60",X"A6",X"CF",X"BD",X"68",X"01",X"1D",X"6A",X"01",X"1D",X"6C",
		X"01",X"F0",X"41",X"A5",X"48",X"F0",X"3A",X"F8",X"BD",X"68",X"01",X"38",X"E5",X"48",X"9D",X"68",
		X"01",X"B0",X"16",X"BD",X"6A",X"01",X"E9",X"00",X"9D",X"6A",X"01",X"08",X"C9",X"21",X"B0",X"08",
		X"BD",X"6C",X"01",X"D0",X"03",X"20",X"D3",X"E0",X"28",X"B0",X"15",X"BD",X"6C",X"01",X"E9",X"00",
		X"9D",X"6C",X"01",X"B0",X"0B",X"A9",X"00",X"9D",X"68",X"01",X"9D",X"6A",X"01",X"9D",X"6C",X"01",
		X"D8",X"4C",X"CE",X"96",X"A9",X"FF",X"85",X"30",X"95",X"42",X"A9",X"0A",X"95",X"00",X"A9",X"00",
		X"85",X"48",X"60",X"A0",X"00",X"AE",X"38",X"01",X"A5",X"16",X"10",X"0F",X"CD",X"39",X"01",X"B0",
		X"07",X"AD",X"39",X"01",X"85",X"16",X"84",X"17",X"4C",X"F4",X"96",X"CD",X"38",X"01",X"90",X"04",
		X"84",X"17",X"86",X"16",X"A5",X"13",X"10",X"0F",X"CD",X"39",X"01",X"B0",X"07",X"AD",X"39",X"01",
		X"85",X"13",X"84",X"14",X"4C",X"10",X"97",X"CD",X"38",X"01",X"90",X"04",X"86",X"13",X"84",X"14",
		X"60",X"A6",X"CF",X"BD",X"68",X"01",X"1D",X"6A",X"01",X"1D",X"6C",X"01",X"F0",X"25",X"A5",X"1D",
		X"29",X"04",X"F0",X"08",X"E6",X"27",X"A5",X"27",X"29",X"3F",X"85",X"11",X"A5",X"1D",X"29",X"08",
		X"F0",X"08",X"C6",X"27",X"A5",X"27",X"29",X"3F",X"85",X"11",X"A5",X"11",X"4A",X"4A",X"4A",X"29",
		X"06",X"85",X"1E",X"60",X"00",X"19",X"32",X"4A",X"62",X"79",X"8E",X"A2",X"B5",X"C6",X"D5",X"E2",
		X"ED",X"F5",X"FB",X"FF",X"FF",X"FB",X"F5",X"ED",X"E2",X"D5",X"C6",X"B5",X"A2",X"8E",X"79",X"62",
		X"4A",X"32",X"19",X"00",X"A6",X"CF",X"B5",X"4D",X"AA",X"BD",X"31",X"C1",X"29",X"10",X"D0",X"37",
		X"BD",X"31",X"C1",X"29",X"20",X"D0",X"1B",X"A6",X"CF",X"B5",X"F6",X"29",X"04",X"D0",X"14",X"A5",
		X"17",X"38",X"E5",X"18",X"85",X"17",X"A5",X"16",X"E9",X"00",X"85",X"16",X"A5",X"15",X"E9",X"00",
		X"85",X"15",X"60",X"A5",X"17",X"18",X"65",X"18",X"85",X"17",X"A5",X"16",X"69",X"00",X"85",X"16",
		X"A5",X"15",X"69",X"00",X"85",X"15",X"60",X"A5",X"0F",X"38",X"E5",X"52",X"85",X"38",X"A5",X"10",
		X"E5",X"51",X"85",X"7B",X"85",X"39",X"A5",X"0D",X"38",X"E5",X"54",X"85",X"3A",X"A5",X"0E",X"E5",
		X"53",X"85",X"3B",X"85",X"7C",X"20",X"49",X"98",X"A4",X"CF",X"B9",X"00",X"00",X"C9",X"08",X"D0",
		X"0D",X"B9",X"F6",X"00",X"29",X"04",X"F0",X"06",X"A5",X"7B",X"49",X"80",X"85",X"7B",X"A5",X"17",
		X"A6",X"7B",X"30",X"14",X"38",X"E5",X"38",X"85",X"17",X"A5",X"16",X"E9",X"00",X"85",X"16",X"A5",
		X"15",X"E9",X"00",X"85",X"15",X"4C",X"09",X"98",X"18",X"65",X"38",X"85",X"17",X"A5",X"16",X"69",
		X"00",X"85",X"16",X"A5",X"15",X"69",X"00",X"85",X"15",X"B9",X"00",X"00",X"C9",X"08",X"D0",X"0D",
		X"B9",X"F6",X"00",X"29",X"04",X"F0",X"06",X"A5",X"7C",X"49",X"80",X"85",X"7C",X"A5",X"14",X"A6",
		X"7C",X"30",X"14",X"38",X"E5",X"3A",X"85",X"14",X"A5",X"13",X"E9",X"00",X"85",X"13",X"A5",X"12",
		X"E9",X"00",X"85",X"12",X"4C",X"48",X"98",X"18",X"65",X"3A",X"85",X"14",X"A5",X"13",X"69",X"00",
		X"85",X"13",X"A5",X"12",X"69",X"00",X"85",X"12",X"60",X"A2",X"02",X"A0",X"00",X"B5",X"39",X"10",
		X"0B",X"98",X"38",X"F5",X"38",X"95",X"38",X"98",X"F5",X"39",X"95",X"39",X"CA",X"CA",X"10",X"ED",
		X"A2",X"02",X"A0",X"03",X"56",X"39",X"76",X"38",X"88",X"10",X"F9",X"56",X"38",X"56",X"38",X"B5",
		X"38",X"4A",X"18",X"75",X"38",X"09",X"03",X"95",X"38",X"CA",X"CA",X"10",X"E5",X"60",X"A6",X"CF",
		X"B5",X"4D",X"AA",X"BD",X"31",X"C1",X"29",X"20",X"D0",X"3C",X"A2",X"03",X"A4",X"49",X"B5",X"14",
		X"F0",X"2F",X"B5",X"12",X"30",X"17",X"B5",X"14",X"38",X"F9",X"C7",X"98",X"95",X"14",X"B5",X"13",
		X"E9",X"00",X"95",X"13",X"B5",X"12",X"E9",X"00",X"95",X"12",X"4C",X"C1",X"98",X"B5",X"14",X"18",
		X"79",X"C7",X"98",X"95",X"14",X"B5",X"13",X"69",X"00",X"95",X"13",X"B5",X"12",X"69",X"00",X"95",
		X"12",X"CA",X"CA",X"CA",X"10",X"C8",X"60",X"03",X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"02",
		X"02",X"A6",X"CF",X"B5",X"88",X"D0",X"01",X"60",X"A5",X"1D",X"29",X"01",X"F0",X"09",X"F8",X"A9",
		X"20",X"18",X"65",X"48",X"85",X"48",X"D8",X"A5",X"0B",X"18",X"65",X"17",X"85",X"0B",X"A5",X"0F",
		X"65",X"16",X"85",X"0F",X"A5",X"10",X"65",X"15",X"30",X"0A",X"C9",X"05",X"90",X"06",X"A0",X"00",
		X"84",X"0F",X"A9",X"05",X"85",X"10",X"A6",X"CF",X"B5",X"00",X"C9",X"24",X"F0",X"04",X"C9",X"08",
		X"D0",X"09",X"20",X"7E",X"9A",X"20",X"8E",X"99",X"4C",X"45",X"99",X"C9",X"1C",X"D0",X"13",X"A9",
		X"FE",X"85",X"21",X"A9",X"02",X"85",X"22",X"A9",X"02",X"85",X"23",X"A9",X"FE",X"85",X"24",X"4C",
		X"42",X"99",X"A9",X"FD",X"85",X"21",X"A9",X"02",X"85",X"22",X"A9",X"03",X"85",X"23",X"A9",X"FD",
		X"85",X"24",X"20",X"37",X"9A",X"A5",X"0C",X"18",X"65",X"14",X"85",X"0C",X"A5",X"0D",X"65",X"13",
		X"85",X"0D",X"A5",X"0E",X"65",X"12",X"85",X"0E",X"A5",X"7A",X"F0",X"03",X"20",X"60",X"99",X"60",
		X"24",X"7A",X"10",X"16",X"A9",X"00",X"38",X"E5",X"14",X"85",X"14",X"A9",X"00",X"E5",X"13",X"85",
		X"13",X"A9",X"00",X"E5",X"12",X"85",X"12",X"4C",X"8D",X"99",X"A9",X"00",X"38",X"E5",X"17",X"85",
		X"17",X"A9",X"00",X"E5",X"16",X"85",X"16",X"A9",X"00",X"E5",X"15",X"85",X"15",X"60",X"A6",X"CF",
		X"B5",X"4D",X"AA",X"BD",X"31",X"C1",X"29",X"F0",X"F0",X"17",X"BD",X"FA",X"99",X"85",X"21",X"BD",
		X"0A",X"9A",X"85",X"22",X"BD",X"19",X"9A",X"85",X"23",X"BD",X"28",X"9A",X"85",X"24",X"4C",X"37",
		X"9A",X"A5",X"12",X"25",X"0E",X"A6",X"30",X"E0",X"50",X"B0",X"05",X"C9",X"FF",X"4C",X"C2",X"99",
		X"C9",X"FD",X"B0",X"0F",X"C9",X"10",X"90",X"0B",X"20",X"C8",X"9A",X"20",X"A5",X"9A",X"68",X"68",
		X"4C",X"5F",X"99",X"A5",X"12",X"30",X"22",X"A5",X"0E",X"A6",X"30",X"E0",X"50",X"B0",X"05",X"C9",
		X"01",X"4C",X"E6",X"99",X"C9",X"02",X"90",X"11",X"F0",X"0F",X"C9",X"10",X"B0",X"0B",X"20",X"C8",
		X"9A",X"20",X"A5",X"9A",X"68",X"68",X"4C",X"5F",X"99",X"60",X"00",X"00",X"00",X"FA",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"FA",X"00",X"F8",X"00",X"00",X"00",X"06",X"03",X"00",
		X"00",X"00",X"04",X"03",X"00",X"00",X"06",X"00",X"08",X"00",X"00",X"00",X"06",X"08",X"00",X"00",
		X"00",X"08",X"08",X"00",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"FA",X"F8",X"00",X"00",X"00",
		X"00",X"F8",X"00",X"00",X"F8",X"00",X"F8",X"A9",X"00",X"85",X"7A",X"A5",X"0E",X"10",X"11",X"C5",
		X"24",X"B0",X"0A",X"A9",X"80",X"85",X"7A",X"A9",X"08",X"85",X"0D",X"E6",X"0E",X"4C",X"5E",X"9A",
		X"C5",X"23",X"90",X"0A",X"A9",X"80",X"85",X"7A",X"A9",X"F7",X"85",X"0D",X"C6",X"0E",X"A5",X"10",
		X"10",X"0F",X"C5",X"21",X"B0",X"08",X"A9",X"40",X"85",X"7A",X"A9",X"FF",X"85",X"0F",X"4C",X"7D",
		X"9A",X"C5",X"22",X"90",X"08",X"A9",X"40",X"85",X"7A",X"A9",X"00",X"85",X"0F",X"60",X"A5",X"7A",
		X"D0",X"22",X"18",X"A5",X"2E",X"65",X"14",X"85",X"2E",X"A5",X"2F",X"65",X"13",X"85",X"2F",X"24",
		X"12",X"30",X"07",X"90",X"02",X"E6",X"2A",X"4C",X"9E",X"9A",X"B0",X"02",X"C6",X"2A",X"A5",X"2A",
		X"29",X"0F",X"85",X"2A",X"60",X"A5",X"2C",X"18",X"65",X"14",X"85",X"2C",X"A5",X"2D",X"65",X"13",
		X"85",X"2D",X"24",X"12",X"30",X"07",X"90",X"02",X"E6",X"2B",X"4C",X"C1",X"9A",X"B0",X"02",X"C6",
		X"2B",X"A5",X"2B",X"29",X"0F",X"85",X"2B",X"60",X"A2",X"16",X"BD",X"73",X"02",X"38",X"E5",X"14",
		X"9D",X"73",X"02",X"BD",X"5C",X"02",X"E5",X"13",X"9D",X"5C",X"02",X"BD",X"45",X"02",X"E5",X"12",
		X"9D",X"45",X"02",X"20",X"0A",X"9B",X"E0",X"02",X"B0",X"1C",X"BD",X"12",X"01",X"38",X"E5",X"14",
		X"9D",X"12",X"01",X"BD",X"16",X"01",X"E5",X"13",X"9D",X"16",X"01",X"BD",X"1A",X"01",X"E5",X"12",
		X"9D",X"1A",X"01",X"20",X"0A",X"9B",X"CA",X"10",X"C1",X"60",X"BD",X"45",X"02",X"10",X"0A",X"C9",
		X"F8",X"B0",X"03",X"4C",X"21",X"9B",X"4C",X"20",X"9B",X"C9",X"08",X"90",X"03",X"4C",X"21",X"9B",
		X"60",X"BD",X"45",X"02",X"30",X"06",X"38",X"E9",X"10",X"4C",X"2F",X"9B",X"18",X"69",X"10",X"9D",
		X"45",X"02",X"60",X"A2",X"01",X"20",X"3C",X"9B",X"CA",X"10",X"FA",X"60",X"A9",X"03",X"8D",X"3F",
		X"01",X"A9",X"FB",X"8D",X"40",X"01",X"8D",X"42",X"01",X"A9",X"04",X"8D",X"41",X"01",X"A4",X"CF",
		X"B9",X"E3",X"00",X"85",X"7B",X"B9",X"3C",X"01",X"F0",X"01",X"60",X"BD",X"34",X"01",X"F0",X"01",
		X"60",X"BD",X"0C",X"01",X"10",X"2C",X"2C",X"40",X"01",X"10",X"1B",X"CD",X"40",X"01",X"D0",X"1F",
		X"C5",X"10",X"B0",X"18",X"E0",X"02",X"90",X"0E",X"A9",X"00",X"9D",X"24",X"01",X"9D",X"20",X"01",
		X"9D",X"1C",X"01",X"4C",X"89",X"9B",X"20",X"9B",X"9D",X"4C",X"8F",X"9B",X"20",X"9B",X"9D",X"4C",
		X"C1",X"9B",X"CD",X"40",X"01",X"D0",X"22",X"C5",X"10",X"90",X"18",X"E0",X"02",X"90",X"0E",X"A9",
		X"00",X"9D",X"24",X"01",X"9D",X"20",X"01",X"9D",X"1C",X"01",X"4C",X"B0",X"9B",X"20",X"9B",X"9D",
		X"4C",X"B6",X"9B",X"20",X"9B",X"9D",X"4C",X"C1",X"9B",X"CD",X"3F",X"01",X"90",X"03",X"20",X"B1",
		X"9D",X"BD",X"04",X"01",X"18",X"7D",X"1C",X"01",X"9D",X"04",X"01",X"BD",X"08",X"01",X"7D",X"20",
		X"01",X"9D",X"08",X"01",X"BD",X"0C",X"01",X"7D",X"24",X"01",X"9D",X"0C",X"01",X"BD",X"18",X"01",
		X"10",X"0B",X"CD",X"42",X"01",X"D0",X"03",X"20",X"6C",X"9D",X"4C",X"F5",X"9B",X"CD",X"41",X"01",
		X"90",X"03",X"20",X"82",X"9D",X"BD",X"10",X"01",X"18",X"7D",X"28",X"01",X"9D",X"10",X"01",X"BD",
		X"14",X"01",X"7D",X"2C",X"01",X"9D",X"14",X"01",X"BD",X"18",X"01",X"7D",X"30",X"01",X"9D",X"18",
		X"01",X"60",X"A5",X"4F",X"29",X"FF",X"D0",X"25",X"AD",X"4E",X"04",X"29",X"01",X"D0",X"1E",X"A6",
		X"CF",X"18",X"B5",X"E5",X"69",X"01",X"C9",X"10",X"90",X"02",X"A9",X"10",X"95",X"E5",X"B5",X"49",
		X"A8",X"B9",X"5B",X"9C",X"18",X"75",X"E7",X"10",X"02",X"A9",X"80",X"95",X"E7",X"60",X"A5",X"4F",
		X"29",X"FF",X"D0",X"16",X"AD",X"4E",X"04",X"29",X"03",X"D0",X"0F",X"A6",X"CF",X"B5",X"E3",X"18",
		X"69",X"01",X"C9",X"07",X"90",X"02",X"A9",X"07",X"95",X"E3",X"60",X"01",X"02",X"03",X"04",X"05",
		X"06",X"07",X"08",X"A2",X"01",X"20",X"04",X"9D",X"CA",X"10",X"FA",X"60",X"BD",X"00",X"01",X"D0",
		X"09",X"20",X"CA",X"9D",X"20",X"D1",X"9D",X"4C",X"7D",X"9C",X"DE",X"00",X"01",X"60",X"A9",X"01",
		X"85",X"21",X"A6",X"CF",X"B5",X"E5",X"85",X"7B",X"A2",X"03",X"20",X"10",X"9D",X"CA",X"C6",X"21",
		X"10",X"F8",X"60",X"03",X"03",X"03",X"00",X"00",X"04",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"01",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"A5",X"37",X"D0",X"4E",X"A6",X"CF",X"B5",X"E5",X"85",X"7B",X"B5",X"4D",X"AA",X"BD",X"31",
		X"C1",X"29",X"08",X"D0",X"3E",X"BD",X"93",X"9C",X"8D",X"3F",X"01",X"BD",X"A2",X"9C",X"8D",X"40",
		X"01",X"A9",X"F7",X"8D",X"42",X"01",X"A9",X"09",X"8D",X"41",X"01",X"A9",X"01",X"85",X"21",X"A2",
		X"03",X"20",X"5B",X"9B",X"BD",X"18",X"01",X"10",X"0C",X"C9",X"F8",X"B0",X"05",X"A9",X"07",X"9D",
		X"18",X"01",X"4C",X"FE",X"9C",X"C9",X"08",X"90",X"05",X"A9",X"F9",X"9D",X"18",X"01",X"CA",X"C6",
		X"21",X"10",X"DE",X"60",X"A4",X"CF",X"B9",X"E3",X"00",X"85",X"7B",X"B9",X"3C",X"01",X"D0",X"5B",
		X"BD",X"00",X"01",X"D0",X"53",X"BD",X"08",X"01",X"85",X"38",X"BD",X"0C",X"01",X"85",X"39",X"BD",
		X"14",X"01",X"85",X"3A",X"BD",X"18",X"01",X"85",X"3B",X"20",X"6F",X"A5",X"86",X"24",X"20",X"99",
		X"A4",X"A6",X"24",X"E0",X"03",X"D0",X"06",X"20",X"6C",X"9D",X"4C",X"56",X"9D",X"E0",X"02",X"D0",
		X"06",X"20",X"82",X"9D",X"4C",X"56",X"9D",X"A5",X"55",X"29",X"02",X"D0",X"06",X"20",X"82",X"9D",
		X"4C",X"56",X"9D",X"20",X"6C",X"9D",X"A5",X"55",X"29",X"01",X"D0",X"06",X"20",X"B1",X"9D",X"4C",
		X"65",X"9D",X"20",X"9B",X"9D",X"4C",X"6B",X"9D",X"DE",X"00",X"01",X"60",X"A9",X"00",X"9D",X"30",
		X"01",X"AD",X"0A",X"60",X"9D",X"28",X"01",X"29",X"0F",X"9D",X"00",X"01",X"A5",X"7B",X"9D",X"2C",
		X"01",X"60",X"A9",X"00",X"38",X"E5",X"7B",X"9D",X"2C",X"01",X"AD",X"0A",X"60",X"9D",X"28",X"01",
		X"29",X"0F",X"9D",X"00",X"01",X"A9",X"FF",X"9D",X"30",X"01",X"60",X"A9",X"00",X"9D",X"24",X"01",
		X"AD",X"0A",X"60",X"9D",X"1C",X"01",X"29",X"07",X"9D",X"00",X"01",X"A5",X"7B",X"9D",X"20",X"01",
		X"60",X"A9",X"00",X"38",X"E5",X"7B",X"9D",X"20",X"01",X"AD",X"0A",X"60",X"9D",X"1C",X"01",X"29",
		X"07",X"9D",X"00",X"01",X"A9",X"FF",X"9D",X"24",X"01",X"60",X"AD",X"0A",X"60",X"30",X"E2",X"10",
		X"CA",X"AD",X"0A",X"60",X"30",X"AC",X"4C",X"6C",X"9D",X"A6",X"CF",X"B5",X"4D",X"AA",X"BD",X"31",
		X"C1",X"30",X"21",X"A5",X"37",X"D0",X"1D",X"A5",X"10",X"D0",X"0B",X"A5",X"30",X"F0",X"04",X"A9",
		X"80",X"85",X"37",X"4C",X"04",X"9E",X"30",X"0C",X"C9",X"03",X"90",X"08",X"A5",X"30",X"30",X"04",
		X"A9",X"40",X"85",X"37",X"60",X"24",X"37",X"10",X"26",X"A5",X"30",X"F0",X"20",X"38",X"E9",X"04",
		X"85",X"30",X"20",X"5C",X"9E",X"A5",X"0E",X"10",X"0A",X"C9",X"FF",X"B0",X"03",X"20",X"AD",X"9E",
		X"4C",X"2A",X"9E",X"C9",X"01",X"90",X"03",X"20",X"8E",X"9E",X"4C",X"2F",X"9E",X"85",X"37",X"24",
		X"37",X"50",X"28",X"A5",X"30",X"30",X"20",X"18",X"69",X"04",X"85",X"30",X"20",X"75",X"9E",X"A5",
		X"0E",X"10",X"0A",X"C9",X"FF",X"B0",X"03",X"20",X"8E",X"9E",X"4C",X"54",X"9E",X"C9",X"01",X"90",
		X"03",X"20",X"AD",X"9E",X"4C",X"5B",X"9E",X"A9",X"00",X"85",X"37",X"60",X"A5",X"0F",X"18",X"69",
		X"10",X"85",X"0F",X"90",X"02",X"E6",X"10",X"A5",X"66",X"18",X"69",X"10",X"85",X"66",X"90",X"02",
		X"E6",X"67",X"4C",X"CC",X"9E",X"A5",X"0F",X"38",X"E9",X"10",X"85",X"0F",X"B0",X"02",X"C6",X"10",
		X"A5",X"66",X"38",X"E9",X"10",X"85",X"66",X"B0",X"02",X"C6",X"67",X"4C",X"F1",X"9E",X"A5",X"0D",
		X"38",X"E9",X"09",X"85",X"0D",X"B0",X"02",X"C6",X"0E",X"A5",X"2D",X"18",X"69",X"09",X"85",X"2D",
		X"90",X"08",X"A5",X"2B",X"69",X"00",X"29",X"0F",X"85",X"2B",X"4C",X"3B",X"9F",X"A5",X"0D",X"18",
		X"69",X"09",X"85",X"0D",X"90",X"02",X"E6",X"0E",X"A5",X"2D",X"38",X"E9",X"09",X"85",X"2D",X"B0",
		X"08",X"A5",X"2B",X"E9",X"00",X"29",X"0F",X"85",X"2B",X"4C",X"16",X"9F",X"A2",X"16",X"BD",X"17",
		X"02",X"18",X"69",X"10",X"9D",X"17",X"02",X"90",X"03",X"FE",X"00",X"02",X"E0",X"02",X"B0",X"0D",
		X"BD",X"0A",X"01",X"69",X"10",X"9D",X"0A",X"01",X"90",X"03",X"FE",X"0E",X"01",X"CA",X"10",X"DE",
		X"60",X"A2",X"16",X"BD",X"17",X"02",X"38",X"E9",X"10",X"9D",X"17",X"02",X"B0",X"03",X"DE",X"00",
		X"02",X"E0",X"02",X"B0",X"0D",X"BD",X"0A",X"01",X"E9",X"0F",X"9D",X"0A",X"01",X"B0",X"03",X"DE",
		X"0E",X"01",X"CA",X"10",X"DE",X"60",X"A2",X"16",X"BD",X"5C",X"02",X"18",X"69",X"09",X"9D",X"5C",
		X"02",X"90",X"03",X"FE",X"45",X"02",X"E0",X"02",X"B0",X"0D",X"BD",X"16",X"01",X"69",X"09",X"9D",
		X"16",X"01",X"90",X"03",X"FE",X"1A",X"01",X"CA",X"10",X"DE",X"60",X"A2",X"16",X"BD",X"5C",X"02",
		X"38",X"E9",X"09",X"9D",X"5C",X"02",X"B0",X"03",X"DE",X"45",X"02",X"E0",X"02",X"B0",X"0D",X"BD",
		X"16",X"01",X"E9",X"08",X"9D",X"16",X"01",X"B0",X"03",X"DE",X"1A",X"01",X"CA",X"10",X"DE",X"60",
		X"A9",X"00",X"38",X"E5",X"2D",X"85",X"44",X"A9",X"F8",X"E9",X"00",X"85",X"45",X"A5",X"2B",X"0A",
		X"A8",X"A5",X"66",X"18",X"71",X"62",X"85",X"46",X"A5",X"67",X"C8",X"71",X"62",X"88",X"85",X"47",
		X"A2",X"03",X"86",X"21",X"A6",X"21",X"BD",X"EC",X"02",X"D0",X"03",X"4C",X"5A",X"A0",X"BD",X"64",
		X"02",X"38",X"E5",X"44",X"85",X"38",X"BD",X"4D",X"02",X"E5",X"45",X"85",X"39",X"18",X"65",X"2B",
		X"29",X"0F",X"85",X"22",X"A5",X"2B",X"85",X"23",X"A0",X"03",X"B9",X"44",X"00",X"99",X"31",X"00",
		X"88",X"10",X"F7",X"A5",X"23",X"0A",X"A8",X"E6",X"32",X"A5",X"33",X"18",X"71",X"5C",X"85",X"33",
		X"A5",X"34",X"C8",X"71",X"5C",X"88",X"85",X"34",X"E6",X"23",X"A5",X"23",X"29",X"0F",X"85",X"23",
		X"C5",X"22",X"D0",X"DF",X"A8",X"B1",X"5E",X"D0",X"03",X"4C",X"5A",X"A0",X"85",X"23",X"B1",X"60",
		X"A8",X"20",X"B7",X"A0",X"90",X"6D",X"B1",X"56",X"F0",X"69",X"B1",X"5A",X"85",X"19",X"BD",X"64",
		X"02",X"38",X"E5",X"31",X"85",X"24",X"BD",X"4D",X"02",X"E5",X"32",X"10",X"07",X"A9",X"00",X"38");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
