library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg2_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg2_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"3C",X"66",X"42",X"42",X"42",X"66",X"3C",X"00",X"00",X"00",X"22",X"7E",X"02",X"00",X"00",
		X"00",X"26",X"6E",X"4A",X"4A",X"4A",X"7A",X"32",X"00",X"44",X"46",X"52",X"52",X"52",X"7E",X"6C",
		X"00",X"0C",X"1C",X"34",X"64",X"44",X"7E",X"04",X"00",X"74",X"56",X"52",X"52",X"52",X"5E",X"0C",
		X"00",X"3C",X"76",X"52",X"52",X"52",X"5E",X"0C",X"00",X"40",X"42",X"46",X"4C",X"58",X"70",X"60",
		X"00",X"2C",X"7E",X"52",X"52",X"52",X"7E",X"2C",X"00",X"30",X"7A",X"4A",X"4A",X"4A",X"6E",X"3C",
		X"00",X"1E",X"34",X"64",X"44",X"64",X"34",X"1E",X"00",X"7E",X"52",X"52",X"52",X"52",X"7E",X"2C",
		X"00",X"3C",X"66",X"42",X"42",X"42",X"42",X"42",X"00",X"7E",X"42",X"42",X"42",X"42",X"66",X"3C",
		X"00",X"7E",X"52",X"52",X"52",X"52",X"42",X"42",X"00",X"7E",X"50",X"50",X"50",X"50",X"40",X"40",
		X"00",X"3C",X"66",X"42",X"42",X"4A",X"6A",X"2E",X"00",X"7E",X"10",X"10",X"10",X"10",X"10",X"7E",
		X"00",X"00",X"00",X"42",X"7E",X"42",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",X"02",X"06",X"7C",
		X"00",X"7E",X"06",X"0C",X"18",X"34",X"66",X"42",X"00",X"7E",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"7E",X"30",X"18",X"0C",X"18",X"30",X"7E",X"00",X"7E",X"60",X"30",X"18",X"0C",X"06",X"7E",
		X"00",X"3C",X"66",X"42",X"42",X"42",X"66",X"3C",X"00",X"7E",X"48",X"48",X"48",X"48",X"78",X"30",
		X"00",X"3C",X"66",X"42",X"4A",X"4C",X"66",X"3A",X"00",X"7E",X"48",X"48",X"48",X"4E",X"7A",X"32",
		X"00",X"24",X"76",X"52",X"5A",X"4A",X"6E",X"24",X"00",X"40",X"40",X"40",X"7E",X"40",X"40",X"40",
		X"00",X"7C",X"06",X"02",X"02",X"02",X"06",X"7C",X"00",X"70",X"1C",X"06",X"02",X"06",X"1C",X"70",
		X"00",X"7C",X"06",X"0C",X"18",X"0C",X"06",X"7C",X"00",X"42",X"66",X"2C",X"18",X"34",X"66",X"42",
		X"00",X"60",X"30",X"18",X"0E",X"18",X"30",X"60",X"00",X"42",X"46",X"4E",X"5A",X"72",X"62",X"42",
		X"00",X"20",X"60",X"40",X"5A",X"50",X"70",X"20",X"00",X"00",X"00",X"00",X"7A",X"60",X"00",X"00",
		X"00",X"6C",X"7E",X"52",X"42",X"16",X"1C",X"10",X"00",X"30",X"78",X"7C",X"3E",X"7C",X"78",X"30",
		X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7C",X"82",X"BA",X"AA",X"AA",X"82",X"7C",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"68",X"70",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"D8",X"D8",X"F8",X"78",X"FC",X"00",X"00",X"04",X"0C",X"1C",X"3C",X"7C",X"7A",
		X"FE",X"FE",X"74",X"34",X"30",X"30",X"00",X"00",X"7F",X"79",X"3F",X"06",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"38",X"0C",X"04",X"46",X"E2",X"E2",X"00",X"07",X"1C",X"30",X"26",X"6F",X"4F",X"59",
		X"E2",X"E2",X"46",X"04",X"0C",X"38",X"E0",X"00",X"5F",X"49",X"6F",X"26",X"30",X"1C",X"07",X"00",
		X"00",X"FE",X"0F",X"0F",X"0F",X"0F",X"FE",X"00",X"F0",X"FF",X"F0",X"00",X"00",X"F0",X"FF",X"F0",
		X"00",X"00",X"0F",X"FF",X"0F",X"C0",X"F0",X"3C",X"00",X"00",X"F0",X"FF",X"3C",X"0F",X"03",X"F0",
		X"FF",X"0F",X"00",X"00",X"0F",X"FF",X"0F",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"EF",X"3F",X"3F",X"EF",X"00",X"00",X"F0",X"FF",X"F1",X"00",X"00",X"F1",X"FF",
		X"00",X"00",X"00",X"0F",X"FF",X"8F",X"8F",X"8F",X"F0",X"00",X"00",X"F0",X"FF",X"F1",X"F1",X"F1",
		X"CF",X"CF",X"1F",X"00",X"00",X"0F",X"FF",X"0F",X"F3",X"F3",X"F8",X"00",X"00",X"F0",X"FF",X"F1",
		X"C0",X"F8",X"3E",X"0F",X"0F",X"00",X"00",X"1F",X"F1",X"F1",X"F9",X"7F",X"3E",X"00",X"00",X"7E",
		X"1F",X"0E",X"8F",X"CF",X"CF",X"FF",X"7E",X"00",X"FF",X"F3",X"F3",X"F1",X"70",X"F8",X"F8",X"00",
		X"00",X"0F",X"7F",X"CF",X"40",X"40",X"CF",X"7F",X"00",X"00",X"00",X"F3",X"FE",X"FE",X"F3",X"00",
		X"0F",X"00",X"00",X"0F",X"FF",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"FF",X"F0",X"00",X"00",
		X"0F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"60",X"30",X"18",X"30",X"60",X"FF",X"00",X"3F",X"08",X"18",X"10",X"10",X"18",X"08",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"81",X"81",X"81",X"81",X"C3",X"7E",
		X"00",X"1E",X"33",X"21",X"21",X"21",X"33",X"1E",X"00",X"03",X"03",X"00",X"3C",X"F8",X"F0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"98",X"08",X"08",X"98",X"F0",X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"0F",
		X"98",X"08",X"08",X"98",X"F0",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"07",X"1F",X"1F",X"3F",X"3F",X"3F",X"00",X"00",X"E0",X"F8",X"F8",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"E0",X"00",X"00",X"3F",X"3F",X"3F",X"1F",X"1F",X"07",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"1F",X"3F",X"3F",X"3F",X"00",X"00",X"E0",X"F9",X"F9",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"98",X"08",X"08",X"98",X"F0",X"9F",X"0F",X"0F",X"9F",X"FF",X"07",X"00",X"00",
		X"00",X"00",X"F7",X"9F",X"0F",X"0F",X"9F",X"FF",X"98",X"08",X"08",X"98",X"F8",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"00",X"3F",X"3F",X"3F",X"1F",X"1F",X"07",X"07",X"0F",
		X"3F",X"7F",X"3F",X"3F",X"7F",X"7F",X"3F",X"7F",X"00",X"B2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"FE",X"FE",X"FC",X"FC",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4D",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",
		X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3F",X"1F",X"1F",X"1F",X"9F",X"FF",X"FF",X"FF",X"FB",X"F8",X"F4",X"FA",X"F1",
		X"5F",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"E1",X"F6",X"F8",X"F0",X"F6",X"FF",X"FF",X"FF",
		X"1F",X"3F",X"3F",X"3F",X"1F",X"00",X"07",X"1F",X"00",X"00",X"00",X"81",X"81",X"C7",X"C7",X"CF",
		X"F8",X"E0",X"F0",X"98",X"08",X"08",X"98",X"F0",X"9B",X"0B",X"0B",X"99",X"F1",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"99",X"09",X"0B",X"9B",X"F3",X"98",X"08",X"08",X"98",X"F0",X"00",X"E0",X"F8",
		X"DF",X"FF",X"FF",X"BF",X"9F",X"00",X"00",X"00",X"1F",X"07",X"00",X"01",X"01",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",
		X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"3F",X"7F",X"3F",X"7F",X"3F",X"3F",X"7F",X"7F",X"3F",X"1F",
		X"00",X"B0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"32",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"FC",X"FE",X"FE",X"FC",X"FC",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0D",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"4C",X"00",
		X"F8",X"E0",X"07",X"1F",X"1F",X"3F",X"3F",X"3F",X"FC",X"FC",X"FC",X"F9",X"F9",X"E3",X"03",X"03",
		X"3F",X"3F",X"3F",X"9F",X"9F",X"C7",X"C0",X"C0",X"1F",X"07",X"E0",X"F8",X"F8",X"FC",X"FC",X"FC",
		X"03",X"03",X"E3",X"F9",X"F9",X"FC",X"FC",X"FC",X"3F",X"3F",X"3F",X"1F",X"1F",X"07",X"E0",X"F8",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"E0",X"07",X"1F",X"C0",X"C0",X"C7",X"9F",X"9F",X"3F",X"3F",X"3F",
		X"F8",X"E0",X"F7",X"9F",X"0F",X"0F",X"9F",X"FF",X"FC",X"FC",X"FC",X"99",X"09",X"0B",X"9B",X"F3",
		X"3F",X"3F",X"3F",X"9F",X"9F",X"C7",X"C7",X"CF",X"1F",X"07",X"E0",X"F9",X"F9",X"FF",X"FF",X"FF",
		X"9B",X"0B",X"0B",X"99",X"F9",X"FC",X"FC",X"FC",X"9F",X"0F",X"0F",X"9F",X"FF",X"07",X"E0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"07",X"1F",X"DF",X"FF",X"FF",X"BF",X"9F",X"3F",X"3F",X"3F",
		X"03",X"03",X"07",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"03",
		X"00",X"00",X"E0",X"F8",X"F8",X"FC",X"FF",X"FF",X"00",X"00",X"07",X"1F",X"1F",X"3F",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F8",X"F8",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"3F",X"1F",X"1F",X"07",X"00",X"00",X"FF",X"FF",X"FC",X"F8",X"F8",X"E0",X"00",X"00",
		X"3F",X"7F",X"3F",X"1F",X"1F",X"07",X"07",X"1F",X"1F",X"07",X"07",X"1F",X"1F",X"3F",X"3F",X"7F",
		X"00",X"02",X"07",X"9F",X"9F",X"FF",X"FF",X"FF",X"00",X"80",X"E0",X"F9",X"F9",X"FF",X"FF",X"FF",
		X"F8",X"E0",X"E0",X"F8",X"F8",X"FC",X"FE",X"FC",X"FE",X"FC",X"FC",X"F8",X"F8",X"E0",X"E0",X"F8",
		X"FF",X"FF",X"FF",X"F9",X"F9",X"E0",X"40",X"00",X"FF",X"FF",X"FF",X"9F",X"9F",X"07",X"01",X"00",
		X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F8",
		X"3F",X"7F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"3F",X"7F",
		X"F8",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"FE",X"FC",X"FE",X"FC",X"FC",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"1F",X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"0F",
		X"00",X"00",X"F0",X"98",X"08",X"08",X"98",X"F0",X"00",X"00",X"F0",X"98",X"08",X"08",X"98",X"F8",
		X"98",X"08",X"08",X"98",X"F0",X"00",X"00",X"00",X"98",X"08",X"08",X"98",X"F0",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"3F",X"7F",X"3F",X"7F",X"3F",X"3F",X"7F",X"7F",X"3F",X"1F",
		X"00",X"B0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"32",X"FF",X"9F",X"0F",X"0F",X"9F",X"FF",
		X"FE",X"FC",X"FE",X"9E",X"0C",X"0C",X"9C",X"F8",X"98",X"0C",X"0E",X"9E",X"FC",X"FC",X"FE",X"FC",
		X"9F",X"0F",X"0F",X"9F",X"FF",X"7F",X"0D",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"4C",X"00",
		X"1F",X"3F",X"3F",X"3F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"07",X"07",X"0F",
		X"00",X"00",X"E0",X"F9",X"F9",X"FF",X"FF",X"FF",X"00",X"00",X"F7",X"9F",X"0F",X"0F",X"9F",X"FF",
		X"FC",X"FC",X"FC",X"98",X"08",X"08",X"98",X"F0",X"98",X"08",X"08",X"98",X"F8",X"FC",X"FC",X"FC",
		X"9F",X"0F",X"0F",X"9F",X"FF",X"07",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"00",
		X"3F",X"7F",X"3F",X"1F",X"1F",X"07",X"07",X"1F",X"1F",X"3F",X"3F",X"3F",X"1F",X"3F",X"3F",X"7F",
		X"00",X"02",X"F7",X"9F",X"0F",X"0F",X"9F",X"FF",X"00",X"80",X"E0",X"F9",X"F9",X"FF",X"FF",X"FF",
		X"98",X"08",X"08",X"98",X"F8",X"FC",X"FE",X"FC",X"FE",X"FC",X"FC",X"98",X"08",X"08",X"98",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"40",X"00",X"9F",X"0F",X"0F",X"9F",X"FF",X"07",X"01",X"00",
		X"FF",X"FF",X"FF",X"9F",X"0F",X"0F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"0F",X"0F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"1F",X"08",X"08",X"08",X"04",X"00",X"0E",X"11",X"11",X"1A",X"0F",X"00",X"1F",X"10",X"10",
		X"18",X"0F",X"00",X"7F",X"04",X"0A",X"0B",X"09",X"00",X"09",X"15",X"15",X"15",X"12",X"00",X"0E",
		X"11",X"11",X"11",X"11",X"00",X"0E",X"11",X"11",X"11",X"0E",X"00",X"1F",X"08",X"08",X"08",X"04",
		X"00",X"1F",X"10",X"10",X"18",X"0F",X"00",X"0E",X"11",X"11",X"1A",X"0F",X"00",X"1F",X"10",X"0F",
		X"10",X"0F",X"00",X"0E",X"15",X"15",X"15",X"0C",X"00",X"09",X"15",X"15",X"15",X"12",X"00",X"0E",
		X"11",X"11",X"11",X"11",X"00",X"0E",X"15",X"15",X"15",X"0C",X"00",X"1F",X"10",X"10",X"18",X"0F",
		X"00",X"0E",X"15",X"15",X"15",X"0C",X"00",X"00",X"00",X"10",X"7F",X"11",X"00",X"00",X"2F",X"00",
		X"00",X"1F",X"10",X"0F",X"10",X"0F",X"00",X"0E",X"15",X"15",X"15",X"0C",X"00",X"00",X"00",X"00",
		X"78",X"FC",X"FE",X"FF",X"FF",X"FF",X"DF",X"1F",X"00",X"03",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"1F",X"1F",X"1F",X"7F",X"FF",X"FF",X"FE",X"FC",X"F8",X"E0",X"00",X"00",X"01",X"07",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FC",X"E0",X"80",X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"FE",X"FF",X"FF",X"7F",X"1F",X"1F",X"1F",X"1F",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"F0",X"FC",X"FE",X"FC",X"F8",X"F8",X"FC",X"FF",X"FF",X"7F",X"3F",X"7F",
		X"1F",X"7F",X"FF",X"FF",X"FE",X"FC",X"FE",X"FF",X"00",X"00",X"01",X"07",X"1F",X"3F",X"1F",X"07",
		X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FC",X"F8",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"7F",X"1F",X"1F",X"1F",X"1F",X"DF",X"FF",X"01",X"00",X"00",X"E0",X"F8",X"FF",X"FF",X"FF",
		X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"F8",X"F9",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"3F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"C0",
		X"80",X"80",X"C3",X"C7",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"C3",X"81",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F3",X"E3",X"C3",X"C1",X"80",X"80",X"80",
		X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C1",X"E3",X"FF",X"FF",X"FF",X"FF",X"0F",X"03",X"0F",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FC",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"3F",X"7F",X"7F",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FF",X"7F",X"7F",X"3F",
		X"F8",X"F0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"0F",X"1F",X"3F",X"1F",X"0F",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"C0",X"80",X"00",
		X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FE",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",X"00",
		X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"FC",X"7E",X"7E",X"3E",X"3F",X"3F",X"1F",X"1F",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"3F",X"7E",X"7E",X"7C",X"FC",X"FC",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3E",X"7E",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"00",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"7C",X"7E",X"7E",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",
		X"00",X"00",X"00",X"80",X"C0",X"F0",X"FC",X"FF",X"7E",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",
		X"F0",X"F0",X"F0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FD",X"FB",X"73",X"07",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"7F",X"3F",X"1F",X"FF",X"FF",X"3F",X"0F",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"7F",X"FE",X"FE",X"FC",X"FC",X"F8",
		X"87",X"01",X"00",X"C7",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"03",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"00",X"01",X"3F",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FE",X"7C",X"00",X"00",X"00",
		X"FD",X"F9",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FE",X"F8",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"7F",X"7F",X"FE",X"FC",X"F8",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FE",X"FC",X"F0",X"C0",X"00",
		X"00",X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FE",X"7F",X"7F",X"3F",X"1F",X"0F",X"03",
		X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F4",X"E0",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",
		X"1C",X"78",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"FF",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"C3",
		X"E0",X"E0",X"C7",X"C3",X"FF",X"FF",X"FF",X"DF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"80",X"20",X"00",X"00",X"00",X"00",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"3F",X"3F",X"3F",X"DF",X"EE",X"EE",X"C0",X"C0",X"C0",X"80",X"0F",X"3F",X"7F",X"7F",
		X"8F",X"03",X"8F",X"DF",X"FF",X"7E",X"1C",X"00",X"7F",X"7E",X"3F",X"3F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"EF",X"CF",X"07",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"A0",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",
		X"F0",X"E0",X"C4",X"00",X"00",X"00",X"00",X"00",X"BF",X"8F",X"C3",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F3",X"E0",X"C3",X"C3",X"C3",X"83",X"03",X"03",X"01",X"00",
		X"F0",X"FC",X"FC",X"F0",X"B8",X"38",X"00",X"00",X"E0",X"E1",X"F9",X"FD",X"FD",X"E8",X"60",X"00",
		X"00",X"00",X"01",X"03",X"03",X"02",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"01",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"3F",X"3F",X"1F",X"1F",
		X"F0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"40",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"00",X"00",X"10",X"38",X"3C",X"7E",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",
		X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"03",X"01",
		X"0F",X"1B",X"10",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"08",X"08",X"08",X"08",
		X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"01",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"C0",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",
		X"00",X"80",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"3F",X"FF",X"FF",X"FF",X"00",X"00",
		X"3F",X"03",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"1F",X"00",X"1F",X"FF",X"FF",X"E0",X"00",
		X"03",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FC",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"F0",X"F0",
		X"FF",X"03",X"03",X"03",X"03",X"03",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"F8",X"FF",X"FF",X"80",X"80",X"F0",X"FE",X"FF",X"9F",
		X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"83",X"80",X"00",X"00",X"00",X"00",X"03",X"03",
		X"87",X"FF",X"FF",X"FE",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"3F",X"7F",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"FE",X"8F",X"07",X"03",X"03",X"01",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"FF",X"E0",X"71",X"7F",X"3F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"FF",X"7F",X"3F",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"3F",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"07",X"FF",X"FF",X"F9",X"01",X"F9",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"15",X"15",X"15",X"0C",X"00",X"00",X"0F",X"1E",X"3C",X"78",X"F0",X"E1",X"C3",X"87");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
