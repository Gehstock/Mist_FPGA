library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity popeye_ch_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of popeye_ch_bits is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"32",X"63",X"63",X"63",X"26",X"1C",X"00",X"18",X"1C",X"18",X"18",X"18",X"18",X"7E",
		X"00",X"3E",X"63",X"70",X"3C",X"1E",X"07",X"7F",X"00",X"7E",X"30",X"18",X"3C",X"60",X"63",X"3E",
		X"00",X"38",X"3C",X"36",X"33",X"7F",X"30",X"30",X"00",X"3F",X"03",X"3F",X"60",X"60",X"63",X"3E",
		X"00",X"3C",X"06",X"03",X"3F",X"63",X"63",X"3E",X"00",X"7F",X"63",X"30",X"18",X"0C",X"0C",X"0C",
		X"00",X"1E",X"23",X"27",X"1C",X"7B",X"61",X"3E",X"00",X"3E",X"63",X"63",X"7E",X"60",X"30",X"1E",
		X"00",X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"3F",X"63",X"63",X"3F",X"63",X"63",X"3F",
		X"00",X"3C",X"66",X"03",X"03",X"03",X"66",X"3C",X"00",X"1F",X"33",X"63",X"63",X"63",X"33",X"1F",
		X"00",X"7E",X"06",X"06",X"3E",X"06",X"06",X"7E",X"00",X"7F",X"03",X"03",X"3F",X"03",X"03",X"03",
		X"00",X"7C",X"06",X"03",X"73",X"63",X"66",X"7C",X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",
		X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"7E",X"00",X"60",X"60",X"60",X"60",X"60",X"63",X"3E",
		X"00",X"63",X"33",X"1B",X"0F",X"1F",X"3B",X"73",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"7E",
		X"00",X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"63",X"67",X"6F",X"7F",X"7B",X"73",X"63",
		X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"3F",X"63",X"63",X"63",X"3F",X"03",X"03",
		X"00",X"3E",X"63",X"63",X"63",X"7B",X"33",X"5E",X"00",X"3F",X"63",X"63",X"73",X"1F",X"3B",X"73",
		X"00",X"1E",X"33",X"03",X"3E",X"60",X"63",X"3E",X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"18",
		X"00",X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",
		X"00",X"63",X"63",X"6B",X"7F",X"7F",X"36",X"22",X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",
		X"00",X"66",X"66",X"24",X"3C",X"18",X"18",X"18",X"00",X"7F",X"70",X"38",X"1C",X"0E",X"07",X"7F",
		X"00",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"18",X"18",X"10",X"10",X"08",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"08",X"49",X"2A",X"1C",X"2A",X"49",X"08",
		X"00",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3C",X"00",X"3C",X"00",X"00",X"00",X"36",X"36",X"7F",X"36",X"36",X"7F",X"36",
		X"00",X"1C",X"22",X"22",X"18",X"08",X"00",X"08",X"00",X"00",X"18",X"18",X"00",X"00",X"18",X"18",
		X"00",X"60",X"70",X"38",X"18",X"04",X"01",X"03",X"00",X"08",X"18",X"08",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"24",X"12",X"36",X"36",X"00",X"00",X"00",
		X"00",X"6C",X"6C",X"48",X"24",X"00",X"00",X"00",X"00",X"00",X"4C",X"4C",X"4C",X"4C",X"7C",X"38",
		X"00",X"00",X"0F",X"1B",X"1B",X"1B",X"0F",X"03",X"00",X"00",X"00",X"DE",X"96",X"9E",X"86",X"86",
		X"00",X"00",X"00",X"3B",X"09",X"39",X"21",X"B9",X"00",X"3C",X"42",X"99",X"85",X"99",X"42",X"3C",
		X"00",X"00",X"DB",X"A8",X"88",X"00",X"00",X"00",X"00",X"00",X"E0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"78",X"08",X"38",X"60",X"60",X"38",X"00",X"00",X"0C",X"1A",X"1A",X"1A",X"1A",X"0C",
		X"00",X"00",X"8C",X"4E",X"4C",X"4C",X"4C",X"9E",X"00",X"00",X"31",X"6B",X"6B",X"6B",X"6B",X"31",
		X"00",X"00",X"8C",X"5A",X"58",X"4C",X"46",X"9E",X"00",X"00",X"9E",X"48",X"4C",X"58",X"58",X"8E",
		X"00",X"00",X"9E",X"42",X"4E",X"58",X"58",X"8E",X"00",X"00",X"9C",X"42",X"4E",X"5A",X"5A",X"8C",
		X"00",X"00",X"19",X"B5",X"B5",X"B5",X"B5",X"19",X"00",X"00",X"63",X"D6",X"D6",X"D6",X"D6",X"63",
		X"FE",X"FF",X"A8",X"AD",X"8D",X"AD",X"FF",X"FE",X"7F",X"FF",X"A8",X"AA",X"AC",X"8A",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"1C",X"3C",X"3C",X"1C",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3B",X"7D",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"F7",
		X"FF",X"FF",X"FF",X"5F",X"3F",X"0F",X"00",X"00",X"FB",X"FF",X"FF",X"FF",X"BD",X"7D",X"FB",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DF",X"FF",X"FF",X"FF",X"BE",X"DC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"BF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FF",X"BF",X"FB",X"FF",
		X"00",X"00",X"00",X"00",X"20",X"30",X"38",X"3C",X"3C",X"38",X"30",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"E6",X"80",X"E0",X"F8",X"E6",X"67",X"1F",X"07",X"01",
		X"67",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E7",X"E7",X"FF",
		X"FF",X"E7",X"E7",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"67",
		X"E6",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"67",X"E6",X"F8",X"E0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"36",X"36",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"10",X"00",X"E0",X"60",X"60",X"E0",X"00",X"FF",X"00",X"00",X"DC",X"D5",X"D5",X"D4",
		X"00",X"FF",X"00",X"00",X"B9",X"9A",X"BA",X"19",X"00",X"7F",X"80",X"00",X"75",X"35",X"75",X"33",
		X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"73",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"B6",X"9A",X"92",X"12",X"9E",X"0C",X"00",X"01",X"02",X"12",X"82",X"D1",X"B2",X"8C",
		X"00",X"00",X"00",X"30",X"4A",X"3E",X"09",X"70",X"00",X"00",X"00",X"90",X"88",X"DC",X"FE",X"25",
		X"00",X"10",X"18",X"4C",X"EE",X"FF",X"FF",X"C9",X"5A",X"32",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5B",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"40",X"40",X"20",X"20",X"00",X"00",X"00",X"03",X"04",X"04",X"08",X"08",
		X"10",X"10",X"08",X"08",X"04",X"84",X"82",X"42",X"10",X"10",X"20",X"20",X"41",X"42",X"82",X"84",
		X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",X"41",X"21",X"20",X"10",X"10",X"08",X"08",X"04",
		X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"00",X"01",X"01",X"02",X"02",X"00",X"00",X"00",X"00",
		X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"03",X"00",X"00",X"00",X"80",X"F0",X"FC",X"FE",X"FF",
		X"00",X"80",X"C0",X"EF",X"9F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"C1",X"0F",
		X"01",X"07",X"F7",X"CF",X"3F",X"FF",X"07",X"F0",X"00",X"00",X"3F",X"FF",X"FF",X"F2",X"FC",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"03",X"FF",X"01",X"01",X"02",X"02",X"04",X"08",X"08",
		X"FF",X"00",X"00",X"00",X"00",X"FC",X"04",X"08",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FD",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",
		X"F8",X"00",X"00",X"00",X"00",X"FF",X"80",X"40",X"FF",X"80",X"80",X"40",X"40",X"20",X"10",X"10",
		X"10",X"20",X"20",X"40",X"80",X"80",X"00",X"00",X"08",X"10",X"20",X"20",X"00",X"00",X"01",X"02",
		X"40",X"20",X"10",X"10",X"08",X"04",X"84",X"42",X"08",X"04",X"04",X"02",X"01",X"01",X"00",X"00",
		X"02",X"04",X"08",X"08",X"10",X"20",X"20",X"40",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"E0",X"F0",X"E0",X"D0",X"D0",X"D0",X"C9",X"CF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"F9",X"F9",X"F9",X"FB",X"FB",X"FB",X"FF",X"FF",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"20",X"10",X"10",X"08",X"04",X"04",X"00",
		X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"F0",X"F0",X"F7",X"EF",X"EF",X"EF",X"CF",X"DF",
		X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"9F",X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F9",X"E3",X"0F",X"FF",X"1F",X"EF",X"FF",X"FF",X"FF",X"7F",X"80",
		X"FF",X"FE",X"F8",X"03",X"83",X"FD",X"FE",X"FF",X"FF",X"FF",X"01",X"FC",X"FF",X"FF",X"CF",X"83",
		X"FF",X"FF",X"FC",X"F8",X"F9",X"F9",X"FD",X"FF",X"0F",X"E7",X"FB",X"FD",X"3F",X"CF",X"E7",X"F3",
		X"00",X"03",X"07",X"0F",X"0E",X"0F",X"0F",X"0F",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"F7",X"FB",X"FB",X"FB",X"FB",X"FB",X"F8",X"F8",X"E3",X"87",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"07",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"80",X"C0",X"C0",X"E0",X"F8",X"FF",X"7F",X"BF",
		X"FF",X"FF",X"DF",X"BF",X"7F",X"7F",X"FF",X"FF",X"F3",X"F3",X"E3",X"E7",X"FF",X"FF",X"7E",X"1C",
		X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"37",X"8F",X"77",X"FB",X"FF",X"FF",X"7F",X"1F",X"80",
		X"FF",X"7F",X"1E",X"CE",X"E6",X"E6",X"F3",X"F2",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F1",X"F3",X"F3",X"E3",X"E3",X"E7",X"C7",X"CF",X"8F",X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"B8",X"C3",X"FF",X"FF",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"08",X"04",X"04",X"84",X"84",X"84",X"84",X"42",
		X"01",X"01",X"01",X"00",X"00",X"00",X"C0",X"30",X"FF",X"FE",X"FC",X"F8",X"E0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"FF",X"FF",X"3F",X"0F",X"87",X"E3",X"F8",X"FE",X"33",X"38",X"3C",X"1E",X"1F",X"0F",X"07",X"01",
		X"10",X"21",X"21",X"21",X"21",X"21",X"22",X"42",X"42",X"42",X"C2",X"02",X"02",X"01",X"01",X"01",
		X"0C",X"03",X"00",X"00",X"80",X"60",X"18",X"06",X"00",X"60",X"18",X"06",X"01",X"00",X"00",X"00",
		X"00",X"00",X"18",X"60",X"80",X"00",X"00",X"00",X"30",X"C0",X"00",X"00",X"01",X"06",X"18",X"60",
		X"42",X"42",X"43",X"40",X"40",X"80",X"80",X"80",X"81",X"61",X"19",X"06",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"86",X"98",X"60",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"BC",X"DC",X"BC",X"DC",
		X"03",X"07",X"1C",X"3F",X"3F",X"7F",X"FF",X"FD",X"B8",X"70",X"C0",X"E0",X"A0",X"A0",X"90",X"40",
		X"7D",X"BB",X"C7",X"FF",X"7D",X"1C",X"06",X"02",X"FF",X"9F",X"0F",X"07",X"07",X"07",X"0F",X"9F",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"03",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"07",X"0F",X"1F",X"3F",X"3F",X"FC",X"FC",X"FC",X"FC",X"FC",X"7C",X"3C",X"3C",
		X"FF",X"FF",X"FF",X"E1",X"C0",X"80",X"00",X"00",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"3E",X"3E",X"7E",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"0B",X"73",X"83",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"03",X"FC",X"00",X"00",X"00",X"00",X"40",X"38",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B8",X"8C",X"9C",X"A0",X"AC",X"BC",X"00",X"00",X"73",X"59",X"5B",X"79",X"7B",X"5B",
		X"00",X"00",X"01",X"07",X"FC",X"FF",X"FF",X"FF",X"23",X"77",X"DE",X"3E",X"FC",X"FF",X"FF",X"FF",
		X"14",X"BE",X"F7",X"73",X"39",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"E0",X"BF",X"FF",X"FF",X"FF",
		X"6E",X"FF",X"FF",X"5D",X"33",X"3E",X"77",X"77",X"E6",X"EE",X"CC",X"9C",X"3C",X"FF",X"FF",X"FF",
		X"76",X"FF",X"FF",X"6A",X"9C",X"FC",X"EE",X"F6",X"F3",X"7B",X"79",X"7C",X"37",X"FF",X"FF",X"FF",
		X"76",X"FF",X"FF",X"F7",X"6D",X"0E",X"0B",X"0B",X"1B",X"1B",X"1B",X"3B",X"37",X"37",X"77",X"77",
		X"7C",X"FE",X"FF",X"FF",X"AE",X"54",X"D0",X"70",X"F8",X"F8",X"E8",X"EC",X"EC",X"F4",X"F6",X"F6",
		X"00",X"00",X"09",X"0F",X"0F",X"1F",X"1B",X"1B",X"00",X"00",X"90",X"F0",X"F0",X"F8",X"E8",X"E8",
		X"00",X"00",X"09",X"0D",X"0F",X"1F",X"3F",X"77",X"00",X"00",X"10",X"10",X"B0",X"F8",X"FC",X"F6",
		X"00",X"00",X"00",X"08",X"1C",X"3F",X"FB",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"77",X"7F",X"7F",X"7F",X"3E",X"1C",X"08",X"00",X"00",X"78",X"20",X"30",X"60",X"60",X"38",
		X"00",X"00",X"2C",X"AC",X"BC",X"BC",X"AC",X"AC",X"00",X"00",X"E7",X"95",X"15",X"D7",X"97",X"F5",
		X"3F",X"FE",X"FC",X"F8",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"03",X"07",X"0F",X"0F",X"1F",X"3F",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3E",X"3E",X"3E",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"C0",X"FC",X"FF",X"F8",X"C0",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"3E",X"1E",X"0F",X"0F",X"07",X"03",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
