library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_program is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"C3",X"00",X"30",X"FF",X"FF",X"FF",X"FF",X"F1",X"C5",X"D5",X"DD",X"E5",X"FD",X"E5",X"E5",
		X"E5",X"21",X"44",X"11",X"E3",X"F5",X"C9",X"00",X"E7",X"CA",X"34",X"0F",X"C3",X"3A",X"0F",X"00",
		X"FD",X"21",X"40",X"0F",X"C3",X"28",X"0F",X"00",X"FD",X"21",X"58",X"0F",X"C3",X"28",X"0F",X"00",
		X"FD",X"21",X"70",X"0F",X"C3",X"28",X"0F",X"00",X"08",X"D9",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"00",X"A0",X"ED",X"57",X"DD",X"21",X"56",X"30",X"87",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"38",X"00",X"FF",X"FF",X"FF",X"FF",X"CD",X"73",X"00",
		X"C3",X"9A",X"01",X"CD",X"4C",X"11",X"3A",X"24",X"60",X"32",X"45",X"50",X"3A",X"25",X"60",X"32",
		X"4A",X"50",X"3A",X"26",X"60",X"32",X"4F",X"50",X"01",X"10",X"00",X"11",X"50",X"50",X"21",X"14",
		X"60",X"ED",X"B0",X"21",X"C3",X"60",X"11",X"00",X"6B",X"01",X"0A",X"00",X"C5",X"D5",X"3A",X"5F",
		X"66",X"B7",X"20",X"04",X"ED",X"B0",X"18",X"14",X"06",X"05",X"7E",X"ED",X"44",X"C6",X"0E",X"12",
		X"23",X"13",X"7E",X"ED",X"44",X"C6",X"10",X"12",X"23",X"13",X"10",X"EE",X"E1",X"C1",X"CD",X"00",
		X"31",X"00",X"00",X"2A",X"09",X"60",X"7C",X"B5",X"CA",X"17",X"11",X"2B",X"22",X"09",X"60",X"C3",
		X"17",X"11",X"CD",X"73",X"00",X"21",X"BF",X"60",X"34",X"7E",X"E6",X"0F",X"F5",X"CC",X"7F",X"03",
		X"F1",X"FE",X"01",X"20",X"0E",X"11",X"01",X"00",X"DD",X"21",X"B2",X"93",X"FD",X"21",X"FC",X"60",
		X"CD",X"6C",X"02",X"DD",X"21",X"27",X"60",X"DD",X"35",X"00",X"28",X"0A",X"DD",X"23",X"DD",X"23",
		X"DD",X"23",X"DD",X"23",X"18",X"F1",X"DD",X"7E",X"01",X"DD",X"77",X"00",X"21",X"19",X"01",X"DD",
		X"E5",X"E5",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"E9",X"DD",X"E1",X"18",X"DF",X"F1",X"F1",X"21",
		X"AE",X"60",X"7E",X"B7",X"28",X"0C",X"35",X"E6",X"07",X"C2",X"9A",X"01",X"CD",X"44",X"12",X"C3",
		X"9A",X"01",X"3A",X"00",X"60",X"4F",X"CB",X"11",X"06",X"02",X"FD",X"21",X"AF",X"60",X"CB",X"11",
		X"FD",X"7E",X"01",X"38",X"1C",X"FD",X"34",X"01",X"11",X"04",X"00",X"FD",X"19",X"10",X"EF",X"C3",
		X"9A",X"01",X"AF",X"32",X"B0",X"60",X"32",X"B4",X"60",X"3E",X"C8",X"32",X"AE",X"60",X"C3",X"9A",
		X"01",X"B7",X"28",X"E4",X"FE",X"01",X"38",X"EA",X"C5",X"FD",X"E5",X"AF",X"FD",X"77",X"01",X"FD",
		X"6E",X"00",X"26",X"00",X"CD",X"00",X"35",X"00",X"CD",X"C8",X"10",X"CD",X"65",X"12",X"FD",X"21",
		X"0B",X"60",X"DD",X"21",X"FC",X"60",X"CD",X"46",X"10",X"3A",X"CD",X"60",X"4F",X"87",X"E6",X"02",
		X"B1",X"32",X"CD",X"60",X"FD",X"E1",X"C1",X"C3",X"48",X"01",X"3A",X"00",X"B8",X"FD",X"E1",X"DD",
		X"E1",X"D9",X"3E",X"01",X"32",X"00",X"A0",X"00",X"08",X"C9",X"21",X"00",X"50",X"06",X"08",X"36",
		X"00",X"23",X"10",X"FB",X"AF",X"32",X"C0",X"50",X"18",X"33",X"DD",X"36",X"00",X"FF",X"DD",X"7E",
		X"00",X"FE",X"FF",X"00",X"00",X"DD",X"36",X"00",X"00",X"DD",X"7E",X"00",X"B7",X"00",X"00",X"DD",
		X"23",X"0B",X"78",X"B1",X"20",X"E4",X"E9",X"F5",X"C5",X"DD",X"E5",X"FD",X"E5",X"DD",X"2E",X"20",
		X"AF",X"06",X"08",X"0E",X"00",X"FD",X"60",X"FD",X"6F",X"FD",X"25",X"FD",X"7E",X"00",X"81",X"4F",
		X"FD",X"23",X"FD",X"7C",X"DD",X"BD",X"20",X"F3",X"DD",X"26",X"20",X"79",X"DD",X"BC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"E1",X"DD",X"E1",X"C1",X"F1",
		X"C9",X"21",X"00",X"68",X"21",X"1B",X"02",X"16",X"33",X"18",X"DB",X"3E",X"FF",X"32",X"32",X"60",
		X"32",X"00",X"A0",X"ED",X"56",X"AF",X"ED",X"47",X"00",X"06",X"0A",X"3A",X"32",X"60",X"B7",X"28",
		X"10",X"21",X"B8",X"0B",X"2B",X"7C",X"B5",X"20",X"FB",X"3A",X"00",X"B8",X"10",X"ED",X"C3",X"98",
		X"0C",X"3E",X"01",X"ED",X"47",X"21",X"05",X"00",X"CD",X"90",X"0F",X"DD",X"21",X"27",X"60",X"DD",
		X"36",X"00",X"01",X"DD",X"36",X"01",X"01",X"21",X"1D",X"01",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"3E",X"01",X"32",X"AF",X"60",X"32",X"B3",X"60",X"C3",X"E6",X"1A",X"CF",X"DD",X"E5",X"E1",X"CB",
		X"D4",X"06",X"03",X"FD",X"7E",X"02",X"1F",X"1F",X"1F",X"1F",X"CD",X"88",X"02",X"FD",X"7E",X"02",
		X"CD",X"88",X"02",X"FD",X"2B",X"10",X"EC",X"C9",X"E6",X"0F",X"28",X"02",X"16",X"FF",X"C6",X"30",
		X"CB",X"22",X"38",X"01",X"AF",X"DD",X"77",X"00",X"00",X"DD",X"23",X"2B",X"C9",X"CF",X"06",X"03",
		X"DD",X"E5",X"E1",X"CB",X"DC",X"FD",X"7E",X"02",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CD",X"C0",X"02",X"FD",X"7E",X"02",X"E6",X"0F",X"CD",X"C0",X"02",X"FD",X"2B",X"10",X"E6",X"C9",
		X"B7",X"28",X"02",X"16",X"FF",X"C6",X"30",X"CB",X"22",X"38",X"01",X"AF",X"DD",X"77",X"00",X"00",
		X"D5",X"11",X"E0",X"FF",X"19",X"DD",X"19",X"D1",X"C9",X"CF",X"21",X"4E",X"61",X"06",X"03",X"3A",
		X"71",X"61",X"E6",X"03",X"EE",X"03",X"3D",X"C5",X"06",X"0A",X"36",X"44",X"23",X"10",X"FB",X"C1",
		X"B8",X"30",X"16",X"F5",X"3A",X"71",X"61",X"E6",X"03",X"5F",X"FE",X"02",X"20",X"01",X"1C",X"78",
		X"EE",X"03",X"83",X"F6",X"80",X"77",X"F1",X"18",X"02",X"36",X"00",X"23",X"10",X"D9",X"CD",X"62",
		X"03",X"06",X"27",X"C5",X"01",X"00",X"04",X"FD",X"7E",X"00",X"E6",X"F0",X"CD",X"5C",X"03",X"FD",
		X"7E",X"00",X"E6",X"0F",X"CD",X"5C",X"03",X"FD",X"23",X"10",X"EC",X"71",X"23",X"C1",X"10",X"E3",
		X"06",X"27",X"1E",X"03",X"C5",X"01",X"00",X"04",X"FD",X"7E",X"F4",X"E6",X"F0",X"CD",X"5C",X"03",
		X"FD",X"7E",X"F4",X"E6",X"0F",X"CD",X"5C",X"03",X"FD",X"23",X"10",X"EC",X"71",X"23",X"C1",X"1D",
		X"20",X"07",X"11",X"E8",X"FF",X"FD",X"19",X"1E",X"03",X"10",X"D9",X"C9",X"28",X"01",X"37",X"CB",
		X"11",X"C9",X"21",X"00",X"61",X"3A",X"71",X"61",X"E6",X"03",X"FE",X"01",X"20",X"05",X"FD",X"21",
		X"C9",X"17",X"C9",X"38",X"05",X"FD",X"21",X"65",X"18",X"C9",X"FD",X"21",X"2D",X"17",X"C9",X"21",
		X"CD",X"60",X"CB",X"46",X"C0",X"21",X"02",X"60",X"CB",X"46",X"28",X"1B",X"11",X"01",X"00",X"DD",
		X"21",X"80",X"92",X"FD",X"21",X"72",X"61",X"CD",X"9E",X"02",X"16",X"00",X"DD",X"21",X"00",X"91",
		X"FD",X"21",X"5C",X"66",X"CD",X"9E",X"02",X"21",X"02",X"60",X"CB",X"4E",X"C8",X"2A",X"73",X"61",
		X"FD",X"21",X"BC",X"93",X"CD",X"BE",X"03",X"2A",X"5D",X"66",X"FD",X"21",X"5C",X"90",X"7C",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",X"4F",X"7C",X"E6",X"0F",X"67",X"06",X"04",X"CB",
		X"3C",X"CB",X"1D",X"10",X"FA",X"FD",X"E5",X"C5",X"22",X"0B",X"60",X"DD",X"21",X"0B",X"60",X"DD",
		X"36",X"02",X"00",X"CD",X"EC",X"10",X"C1",X"45",X"E1",X"78",X"B7",X"28",X"1B",X"05",X"78",X"D6",
		X"04",X"38",X"0B",X"47",X"00",X"00",X"CB",X"D4",X"71",X"CB",X"94",X"2B",X"18",X"F0",X"3E",X"FB",
		X"80",X"00",X"CB",X"D4",X"00",X"CB",X"94",X"2B",X"00",X"00",X"CB",X"D4",X"00",X"CB",X"94",X"2D",
		X"7D",X"E6",X"1F",X"20",X"F3",X"C9",X"FD",X"7E",X"0A",X"E6",X"07",X"FD",X"21",X"48",X"04",X"87",
		X"5F",X"16",X"00",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"11",X"E0",X"FF",X"06",X"04",
		X"C5",X"E5",X"06",X"04",X"DD",X"7E",X"00",X"77",X"CB",X"DC",X"71",X"CB",X"9C",X"19",X"DD",X"23",
		X"10",X"F2",X"E1",X"23",X"C1",X"10",X"E9",X"C9",X"24",X"92",X"06",X"93",X"46",X"91",X"05",X"93",
		X"45",X"91",X"2E",X"92",X"DD",X"21",X"A1",X"15",X"06",X"0A",X"FD",X"7E",X"00",X"CD",X"6F",X"04",
		X"FD",X"7E",X"00",X"1F",X"1F",X"1F",X"1F",X"CD",X"6F",X"04",X"FD",X"23",X"10",X"EC",X"C9",X"DD",
		X"5E",X"00",X"DD",X"56",X"01",X"19",X"E6",X"0F",X"5F",X"DD",X"7E",X"02",X"93",X"77",X"CB",X"DC",
		X"71",X"CB",X"9C",X"11",X"03",X"00",X"DD",X"19",X"C9",X"06",X"03",X"DD",X"21",X"C9",X"04",X"21",
		X"D8",X"60",X"7E",X"E5",X"FD",X"21",X"B9",X"04",X"87",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"6E",
		X"00",X"FD",X"66",X"01",X"DD",X"E5",X"C5",X"DD",X"22",X"FA",X"60",X"E9",X"C1",X"DD",X"E1",X"E1",
		X"23",X"11",X"06",X"00",X"DD",X"19",X"10",X"DA",X"C9",X"DB",X"04",X"89",X"05",X"DE",X"04",X"F8",
		X"05",X"F3",X"05",X"81",X"06",X"D3",X"06",X"97",X"07",X"4E",X"61",X"D5",X"60",X"DC",X"60",X"59",
		X"61",X"D6",X"60",X"DE",X"60",X"64",X"61",X"D7",X"60",X"E0",X"60",X"C3",X"AC",X"04",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"34",X"7E",X"FE",X"40",X"20",X"40",X"F5",X"E5",X"DD",X"E5",X"23",X"23",
		X"23",X"34",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"E5",X"FD",X"E1",X"3A",X"CB",X"60",X"FD",X"5E",
		X"06",X"CB",X"3F",X"53",X"CB",X"3A",X"92",X"6F",X"3A",X"CC",X"60",X"FD",X"56",X"07",X"92",X"67",
		X"FD",X"75",X"00",X"FD",X"74",X"01",X"FD",X"73",X"13",X"FD",X"72",X"19",X"AF",X"FD",X"77",X"12",
		X"FD",X"77",X"18",X"CD",X"AA",X"12",X"DD",X"E1",X"E1",X"F1",X"E6",X"07",X"C2",X"AC",X"04",X"7E",
		X"FE",X"48",X"38",X"03",X"3E",X"88",X"96",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"E5",X"FD",
		X"E1",X"DD",X"21",X"B1",X"14",X"F5",X"87",X"5F",X"16",X"00",X"DD",X"19",X"0E",X"17",X"CD",X"16",
		X"04",X"F1",X"FD",X"E1",X"CB",X"67",X"28",X"04",X"0E",X"18",X"18",X"02",X"0E",X"19",X"CD",X"54",
		X"04",X"CD",X"92",X"12",X"C3",X"AC",X"04",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"FD",X"E1",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"34",X"7E",X"FE",X"60",X"38",X"45",X"AF",X"77",X"F5",X"3A",
		X"CD",X"66",X"B7",X"CC",X"7B",X"12",X"F1",X"18",X"38",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",
		X"FD",X"E1",X"FD",X"CB",X"0A",X"7E",X"CA",X"AC",X"04",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"34",
		X"7E",X"FE",X"60",X"38",X"1C",X"AF",X"77",X"F5",X"E5",X"E5",X"3A",X"CD",X"66",X"B7",X"CC",X"7B",
		X"12",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"35",X"E1",X"20",X"04",X"23",X"23",X"23",X"34",X"E1",
		X"F1",X"E6",X"07",X"C2",X"AC",X"04",X"7E",X"FE",X"30",X"38",X"03",X"3E",X"58",X"96",X"F5",X"DD",
		X"21",X"41",X"15",X"87",X"5F",X"16",X"00",X"DD",X"19",X"FD",X"E5",X"0E",X"1D",X"CD",X"16",X"04",
		X"FD",X"E1",X"F1",X"CB",X"5F",X"28",X"04",X"0E",X"1A",X"18",X"02",X"0E",X"1B",X"CD",X"54",X"04",
		X"C3",X"AC",X"04",X"21",X"67",X"05",X"18",X"03",X"21",X"DE",X"04",X"E5",X"DD",X"E5",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"7E",X"FE",X"50",X"20",X"05",X"F5",X"CD",X"C4",X"12",X"F1",X"FE",X"80",
		X"20",X"04",X"23",X"23",X"23",X"34",X"3A",X"71",X"61",X"5F",X"16",X"00",X"FD",X"21",X"65",X"06",
		X"FD",X"19",X"FD",X"4E",X"00",X"CD",X"51",X"08",X"DD",X"7E",X"13",X"DD",X"77",X"E9",X"DD",X"7E",
		X"19",X"DD",X"77",X"EA",X"CD",X"20",X"32",X"DD",X"09",X"DD",X"36",X"01",X"02",X"F5",X"CD",X"A0",
		X"32",X"00",X"00",X"00",X"3E",X"04",X"DD",X"77",X"00",X"F1",X"FE",X"12",X"DD",X"E1",X"30",X"13",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"23",X"23",X"36",X"05",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"36",X"FF",X"E1",X"E9",X"03",X"03",X"03",X"00",X"04",X"04",X"04",X"00",X"05",X"05",X"05",
		X"00",X"06",X"06",X"06",X"00",X"07",X"07",X"07",X"00",X"08",X"08",X"08",X"00",X"09",X"09",X"09",
		X"00",X"DD",X"E5",X"CD",X"A9",X"12",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"E5",X"FD",X"E1",X"FD",
		X"34",X"00",X"FD",X"7E",X"00",X"FE",X"08",X"38",X"12",X"FD",X"E5",X"F5",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"E5",X"FD",X"E1",X"FD",X"34",X"03",X"F1",X"FD",X"E1",X"FD",X"E5",X"11",X"A8",X"37",
		X"FD",X"19",X"E6",X"07",X"C6",X"25",X"00",X"00",X"00",X"FD",X"E1",X"3A",X"CB",X"60",X"FD",X"96",
		X"E9",X"30",X"02",X"ED",X"44",X"FE",X"0A",X"30",X"05",X"3E",X"04",X"32",X"EC",X"60",X"DD",X"E1",
		X"C3",X"67",X"05",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"E5",X"FD",X"E1",X"34",X"CB",X"46",X"CA",
		X"67",X"05",X"FD",X"5E",X"E9",X"3A",X"CB",X"60",X"93",X"30",X"1B",X"ED",X"44",X"FE",X"0C",X"30",
		X"4A",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"23",X"23",X"34",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"36",X"00",X"C3",X"67",X"05",X"FE",X"0C",X"38",X"E7",X"7B",X"FE",X"16",X"1D",X"0E",X"80",
		X"30",X"31",X"3A",X"71",X"61",X"5F",X"16",X"00",X"21",X"70",X"07",X"19",X"7E",X"FD",X"77",X"00",
		X"CD",X"40",X"32",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"23",X"23",X"23",X"36",X"01",X"C3",X"67",X"05",X"7B",X"FE",X"F6",X"1C",X"0E",
		X"00",X"30",X"CF",X"FD",X"73",X"E9",X"FD",X"36",X"EA",X"10",X"7B",X"21",X"8F",X"07",X"E6",X"07",
		X"5F",X"16",X"00",X"19",X"7E",X"B1",X"CD",X"40",X"32",X"FD",X"19",X"FD",X"36",X"01",X"0E",X"21",
		X"5F",X"66",X"AE",X"FD",X"77",X"00",X"3A",X"1E",X"60",X"B7",X"CC",X"E1",X"12",X"C3",X"67",X"05",
		X"08",X"09",X"0A",X"00",X"06",X"07",X"08",X"00",X"04",X"05",X"06",X"03",X"04",X"05",X"00",X"02",
		X"03",X"04",X"00",X"01",X"02",X"03",X"00",X"01",X"01",X"02",X"00",X"01",X"01",X"01",X"00",X"28",
		X"29",X"2A",X"2B",X"2B",X"2A",X"29",X"28",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"7E",X"B7",X"20",
		X"2E",X"E5",X"DD",X"E5",X"F5",X"FD",X"21",X"0E",X"60",X"DD",X"21",X"0B",X"60",X"CD",X"96",X"10",
		X"21",X"C8",X"00",X"DD",X"21",X"0E",X"60",X"CD",X"C8",X"10",X"CD",X"C2",X"26",X"CD",X"60",X"35",
		X"FD",X"21",X"0B",X"60",X"DD",X"21",X"0E",X"60",X"CD",X"96",X"10",X"F1",X"DD",X"E1",X"E1",X"FE",
		X"0F",X"D2",X"E5",X"07",X"34",X"CD",X"60",X"32",X"19",X"3A",X"5F",X"66",X"EE",X"27",X"77",X"23",
		X"36",X"02",X"C3",X"67",X"05",X"E5",X"FD",X"E1",X"C3",X"12",X"07",X"DD",X"21",X"4E",X"61",X"FD",
		X"21",X"D8",X"60",X"06",X"03",X"16",X"00",X"21",X"E2",X"60",X"DD",X"CB",X"0A",X"7E",X"20",X"0B",
		X"36",X"00",X"23",X"36",X"00",X"FD",X"36",X"00",X"00",X"18",X"20",X"DD",X"7E",X"0A",X"E6",X"07",
		X"FD",X"E5",X"FD",X"21",X"45",X"08",X"87",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"77",
		X"FD",X"7E",X"01",X"23",X"77",X"FD",X"E1",X"FD",X"36",X"00",X"01",X"23",X"FD",X"23",X"1E",X"0B",
		X"DD",X"19",X"10",X"C6",X"DD",X"21",X"DC",X"60",X"DD",X"36",X"00",X"03",X"DD",X"36",X"02",X"07",
		X"DD",X"36",X"04",X"0C",X"C9",X"86",X"D8",X"BE",X"C8",X"4E",X"C8",X"BE",X"D0",X"4E",X"D0",X"86",
		X"88",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"E5",X"DD",X"E1",X"DD",X"5E",X"00",X"16",X"00",X"CB",
		X"7B",X"28",X"01",X"15",X"CB",X"23",X"CD",X"8C",X"08",X"DD",X"5E",X"12",X"DD",X"56",X"13",X"19",
		X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"5E",X"01",X"16",X"FF",X"CD",X"8C",X"08",X"DD",X"5E",
		X"18",X"DD",X"56",X"19",X"19",X"DD",X"75",X"18",X"DD",X"74",X"19",X"C9",X"06",X"08",X"21",X"00",
		X"00",X"79",X"29",X"87",X"30",X"01",X"19",X"10",X"F9",X"C9",X"DD",X"21",X"0E",X"60",X"CD",X"C0",
		X"10",X"20",X"06",X"21",X"EC",X"60",X"CB",X"C6",X"C9",X"DD",X"21",X"0E",X"60",X"CD",X"8E",X"10",
		X"3A",X"0E",X"60",X"FE",X"99",X"20",X"05",X"3E",X"60",X"32",X"0E",X"60",X"3A",X"BF",X"60",X"E6",
		X"0F",X"FE",X"06",X"20",X"26",X"06",X"02",X"DD",X"21",X"06",X"93",X"FD",X"21",X"0E",X"60",X"11",
		X"03",X"00",X"C5",X"D5",X"CD",X"A0",X"02",X"21",X"02",X"60",X"CB",X"46",X"D1",X"C1",X"28",X"0B",
		X"FD",X"21",X"10",X"60",X"DD",X"21",X"46",X"91",X"CD",X"A0",X"02",X"06",X"03",X"DD",X"21",X"06",
		X"09",X"DD",X"22",X"FA",X"60",X"C5",X"DD",X"E5",X"CD",X"12",X"09",X"DD",X"E1",X"C1",X"11",X"04",
		X"00",X"DD",X"19",X"10",X"EC",X"C9",X"D8",X"60",X"DC",X"60",X"D9",X"60",X"DE",X"60",X"DA",X"60",
		X"E0",X"60",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7E",X"E5",X"E6",X"07",X"FD",X"21",X"2D",X"09",
		X"87",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E9",X"37",X"09",X"78",
		X"09",X"D7",X"09",X"EA",X"09",X"13",X"0A",X"CD",X"EA",X"0A",X"E1",X"E5",X"11",X"FD",X"FF",X"19",
		X"35",X"E1",X"C0",X"34",X"21",X"D8",X"60",X"06",X"03",X"CB",X"A6",X"23",X"10",X"FB",X"3A",X"CB",
		X"60",X"CB",X"3F",X"D6",X"44",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"E5",X"FD",X"E1",X"FD",X"36",
		X"01",X"2A",X"FD",X"77",X"00",X"FD",X"36",X"13",X"86",X"FD",X"36",X"19",X"E8",X"FD",X"36",X"12",
		X"00",X"FD",X"36",X"18",X"00",X"C3",X"C5",X"12",X"21",X"EC",X"60",X"CB",X"4E",X"E1",X"C0",X"E5",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"0E",X"03",X"CD",X"57",X"08",X"DD",X"6E",X"13",X"DD",X"75",
		X"E9",X"DD",X"66",X"19",X"DD",X"74",X"EA",X"01",X"A8",X"37",X"DD",X"09",X"DD",X"36",X"01",X"02",
		X"E6",X"07",X"C6",X"8C",X"00",X"00",X"00",X"7C",X"FE",X"12",X"30",X"04",X"E1",X"36",X"03",X"C9",
		X"ED",X"5B",X"CB",X"60",X"7A",X"94",X"30",X"02",X"ED",X"44",X"FE",X"08",X"30",X"08",X"7B",X"95",
		X"30",X"02",X"ED",X"44",X"FE",X"08",X"E1",X"D0",X"36",X"02",X"2B",X"2B",X"2B",X"36",X"1E",X"21",
		X"EC",X"60",X"CB",X"CE",X"C3",X"4D",X"14",X"CD",X"EA",X"0A",X"E1",X"E5",X"2B",X"2B",X"2B",X"35",
		X"E1",X"C0",X"36",X"01",X"21",X"EC",X"60",X"CB",X"8E",X"C9",X"DD",X"6E",X"02",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"E5",X"FD",X"E1",X"FD",X"36",X"EA",X"12",X"FD",X"7E",X"E9",X"FE",X"86",X"E1",
		X"36",X"04",X"38",X"05",X"21",X"E5",X"12",X"18",X"03",X"21",X"28",X"12",X"FD",X"75",X"00",X"FD",
		X"74",X"01",X"C9",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"E5",X"FD",X"E1",X"FD",X"6E",X"E9",X"FD",
		X"66",X"EA",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"CD",X"03",X"10",X"28",X"40",X"7C",X"BA",X"28",
		X"07",X"38",X"03",X"25",X"18",X"02",X"24",X"24",X"7D",X"BB",X"0E",X"00",X"28",X"0B",X"38",X"05",
		X"2D",X"0E",X"02",X"18",X"01",X"2C",X"CD",X"6A",X"14",X"FD",X"75",X"E9",X"FD",X"74",X"EA",X"7D",
		X"21",X"8F",X"07",X"E6",X"07",X"5F",X"16",X"00",X"19",X"7E",X"B1",X"11",X"18",X"03",X"FD",X"19",
		X"CD",X"20",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"C9",X"01",X"00",X"0A",
		X"DD",X"21",X"B2",X"0A",X"CD",X"BE",X"2D",X"79",X"FE",X"09",X"E1",X"20",X"08",X"36",X"00",X"2B",
		X"2B",X"2B",X"36",X"14",X"C9",X"87",X"DD",X"21",X"C6",X"0A",X"87",X"5F",X"16",X"00",X"DD",X"19",
		X"DD",X"7E",X"02",X"A6",X"C0",X"06",X"03",X"21",X"D8",X"60",X"DD",X"7E",X"02",X"B6",X"DD",X"A6",
		X"03",X"77",X"23",X"10",X"F5",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"75",X"00",X"FD",X"74",
		X"01",X"C9",X"28",X"12",X"28",X"F8",X"40",X"F8",X"60",X"F8",X"86",X"F8",X"E5",X"12",X"E5",X"F8",
		X"CB",X"F8",X"B3",X"F8",X"86",X"E8",X"28",X"F8",X"00",X"FF",X"40",X"F8",X"00",X"FF",X"60",X"F8",
		X"20",X"FF",X"86",X"F8",X"10",X"DF",X"86",X"E8",X"00",X"EF",X"E5",X"F8",X"00",X"FF",X"CB",X"F8",
		X"00",X"FF",X"B3",X"F8",X"20",X"FF",X"86",X"F8",X"10",X"DF",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"11",X"A8",X"37",X"19",X"3A",X"BF",X"60",X"E6",X"07",X"C6",X"94",X"00",X"23",X"36",X"02",X"C9",
		X"CF",X"21",X"81",X"93",X"01",X"1A",X"1F",X"11",X"18",X"00",X"CD",X"FF",X"0B",X"CD",X"62",X"03",
		X"DD",X"21",X"81",X"93",X"01",X"03",X"27",X"C5",X"06",X"04",X"4E",X"CB",X"11",X"30",X"0A",X"FD",
		X"7E",X"00",X"1F",X"1F",X"1F",X"1F",X"CD",X"84",X"0B",X"DD",X"23",X"CB",X"11",X"30",X"06",X"FD",
		X"7E",X"00",X"CD",X"84",X"0B",X"DD",X"23",X"FD",X"23",X"10",X"E0",X"23",X"C1",X"0D",X"20",X"07",
		X"11",X"C8",X"FF",X"DD",X"19",X"0E",X"03",X"10",X"CE",X"01",X"03",X"27",X"C5",X"06",X"04",X"4E",
		X"CB",X"11",X"30",X"0A",X"FD",X"7E",X"F4",X"1F",X"1F",X"1F",X"1F",X"CD",X"84",X"0B",X"DD",X"23",
		X"CB",X"11",X"30",X"06",X"FD",X"7E",X"F4",X"CD",X"84",X"0B",X"DD",X"23",X"FD",X"23",X"10",X"E0",
		X"23",X"C1",X"0D",X"20",X"0C",X"0E",X"03",X"11",X"C8",X"FF",X"DD",X"19",X"11",X"E8",X"FF",X"FD",
		X"19",X"10",X"C9",X"C9",X"E6",X"0F",X"FD",X"E5",X"FD",X"21",X"A8",X"0B",X"87",X"5F",X"16",X"00",
		X"FD",X"19",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"DD",X"E5",X"11",X"00",X"08",X"DD",X"19",X"FD",
		X"7E",X"01",X"DD",X"77",X"00",X"DD",X"E1",X"FD",X"E1",X"C9",X"04",X"18",X"05",X"19",X"06",X"1A",
		X"07",X"1B",X"CF",X"21",X"00",X"90",X"36",X"00",X"23",X"7C",X"FE",X"48",X"20",X"F8",X"C9",X"CF",
		X"5E",X"23",X"56",X"23",X"D5",X"DD",X"E1",X"CD",X"38",X"10",X"10",X"F4",X"C9",X"CF",X"E5",X"0E",
		X"04",X"C5",X"21",X"48",X"93",X"CD",X"E0",X"0B",X"C1",X"E1",X"DD",X"21",X"A8",X"92",X"18",X"0C",
		X"C5",X"E5",X"CD",X"17",X"0C",X"E1",X"C1",X"13",X"23",X"10",X"F5",X"C9",X"5E",X"23",X"56",X"23",
		X"D5",X"FD",X"E1",X"16",X"00",X"59",X"CD",X"9D",X"02",X"DD",X"23",X"10",X"EF",X"C9",X"CF",X"C5",
		X"E5",X"41",X"72",X"CD",X"D0",X"32",X"00",X"00",X"D5",X"11",X"E0",X"FF",X"19",X"D1",X"10",X"F2",
		X"E1",X"C1",X"23",X"10",X"EA",X"C9",X"CF",X"1A",X"FE",X"24",X"C8",X"77",X"CD",X"D0",X"32",X"00",
		X"00",X"13",X"D5",X"11",X"E0",X"FF",X"19",X"D1",X"18",X"ED",X"CF",X"1A",X"FE",X"24",X"C8",X"77",
		X"00",X"00",X"00",X"00",X"00",X"2B",X"13",X"18",X"F2",X"CF",X"11",X"BA",X"1A",X"0E",X"17",X"21",
		X"1C",X"90",X"C3",X"2B",X"0C",X"32",X"C0",X"50",X"DD",X"21",X"00",X"90",X"01",X"00",X"08",X"DD",
		X"36",X"00",X"00",X"DD",X"23",X"0B",X"78",X"B1",X"20",X"F5",X"32",X"C0",X"50",X"21",X"01",X"19",
		X"01",X"E0",X"FF",X"DD",X"21",X"10",X"93",X"FD",X"21",X"10",X"47",X"7E",X"FE",X"24",X"28",X"0E",
		X"DD",X"77",X"00",X"FD",X"36",X"00",X"03",X"23",X"DD",X"09",X"FD",X"09",X"18",X"ED",X"7A",X"32",
		X"B0",X"92",X"7B",X"32",X"90",X"92",X"06",X"0A",X"21",X"20",X"66",X"32",X"C0",X"50",X"2B",X"7C",
		X"B5",X"20",X"F8",X"10",X"F3",X"C3",X"01",X"00",X"32",X"C0",X"50",X"F3",X"21",X"00",X"44",X"36",
		X"00",X"32",X"C0",X"50",X"23",X"7C",X"FE",X"48",X"20",X"F5",X"21",X"0B",X"19",X"11",X"00",X"00",
		X"18",X"AE",X"21",X"CD",X"60",X"CB",X"56",X"C0",X"CB",X"46",X"C2",X"34",X"0D",X"21",X"00",X"60",
		X"CB",X"7E",X"3E",X"02",X"20",X"02",X"3E",X"04",X"F5",X"21",X"00",X"60",X"CB",X"56",X"CA",X"E9",
		X"0C",X"21",X"00",X"60",X"CB",X"4E",X"CA",X"FD",X"0C",X"F1",X"CD",X"28",X"0D",X"C6",X"05",X"21",
		X"5F",X"66",X"00",X"32",X"80",X"98",X"C3",X"89",X"04",X"C1",X"3A",X"CB",X"60",X"90",X"FE",X"24",
		X"30",X"02",X"3E",X"24",X"32",X"CB",X"60",X"38",X"E1",X"1E",X"00",X"18",X"10",X"21",X"CB",X"60",
		X"F1",X"86",X"FE",X"EC",X"38",X"02",X"3E",X"EC",X"77",X"30",X"CF",X"1E",X"80",X"3A",X"80",X"98",
		X"CB",X"47",X"20",X"02",X"1C",X"00",X"CD",X"28",X"0D",X"C6",X"07",X"E6",X"7F",X"83",X"21",X"5F",
		X"66",X"00",X"32",X"80",X"98",X"C3",X"89",X"04",X"21",X"70",X"61",X"3E",X"08",X"96",X"00",X"00",
		X"4F",X"87",X"81",X"C9",X"3A",X"BF",X"60",X"E6",X"07",X"20",X"56",X"3A",X"CB",X"60",X"21",X"C3",
		X"60",X"BE",X"30",X"05",X"96",X"ED",X"44",X"18",X"01",X"96",X"FE",X"6F",X"7E",X"30",X"3F",X"3A",
		X"CE",X"60",X"D6",X"05",X"38",X"37",X"FE",X"07",X"30",X"33",X"4F",X"2A",X"C3",X"60",X"7C",X"FE",
		X"78",X"30",X"2A",X"79",X"DD",X"21",X"B6",X"0D",X"87",X"5F",X"16",X"00",X"DD",X"19",X"EB",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"7A",X"D6",X"15",X"E9",X"87",X"ED",X"44",X"18",X"0C",X"CB",X"3F",
		X"18",X"F8",X"AF",X"18",X"05",X"CB",X"3F",X"18",X"01",X"87",X"83",X"18",X"01",X"AF",X"32",X"60",
		X"66",X"3A",X"60",X"66",X"B7",X"CA",X"DA",X"0C",X"21",X"CB",X"60",X"96",X"30",X"0D",X"ED",X"44",
		X"FE",X"04",X"DA",X"DA",X"0C",X"3E",X"02",X"F5",X"C3",X"E9",X"0C",X"FE",X"04",X"DA",X"DA",X"0C",
		X"3E",X"02",X"F5",X"C3",X"FD",X"0C",X"79",X"0D",X"7A",X"0D",X"7E",X"0D",X"82",X"0D",X"85",X"0D",
		X"8A",X"0D",X"89",X"0D",X"CD",X"AA",X"12",X"11",X"D6",X"1A",X"21",X"F0",X"96",X"7E",X"FE",X"02",
		X"28",X"04",X"0E",X"02",X"18",X"02",X"0E",X"00",X"CB",X"94",X"C3",X"17",X"0C",X"11",X"A1",X"1A",
		X"21",X"5F",X"92",X"7E",X"FE",X"02",X"28",X"04",X"0E",X"02",X"18",X"02",X"0E",X"00",X"CB",X"94",
		X"C3",X"17",X"0C",X"F5",X"E5",X"FD",X"2E",X"FF",X"DD",X"2E",X"FF",X"DD",X"2C",X"DD",X"26",X"87",
		X"DD",X"24",X"DD",X"7E",X"00",X"FD",X"BD",X"00",X"20",X"10",X"DD",X"7D",X"57",X"FD",X"2C",X"FD",
		X"5D",X"EB",X"E9",X"DD",X"26",X"FF",X"FD",X"2E",X"FF",X"DD",X"E1",X"F1",X"C9",X"21",X"61",X"47",
		X"C5",X"11",X"03",X"00",X"FD",X"19",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"FD",X"46",X"02",X"DD",
		X"7E",X"03",X"77",X"DD",X"35",X"02",X"20",X"0F",X"DD",X"7E",X"04",X"DD",X"77",X"02",X"DD",X"7E",
		X"03",X"3D",X"E6",X"03",X"DD",X"77",X"03",X"19",X"10",X"E5",X"C1",X"10",X"D3",X"C9",X"6E",X"6D",
		X"71",X"6A",X"E0",X"FF",X"19",X"01",X"00",X"1E",X"20",X"00",X"19",X"FF",X"FF",X"1D",X"E0",X"FF",
		X"18",X"01",X"00",X"1C",X"20",X"00",X"17",X"FF",X"FF",X"1B",X"E0",X"FF",X"16",X"01",X"00",X"1A",
		X"20",X"00",X"15",X"FF",X"FF",X"19",X"E0",X"FF",X"14",X"01",X"00",X"18",X"20",X"00",X"13",X"FF",
		X"FF",X"18",X"CF",X"0E",X"01",X"11",X"9A",X"08",X"C3",X"9A",X"0F",X"CF",X"0E",X"01",X"11",X"B2",
		X"0C",X"C3",X"9A",X"0F",X"CF",X"11",X"18",X"72",X"21",X"81",X"93",X"01",X"1A",X"04",X"CD",X"FE",
		X"0B",X"21",X"9C",X"93",X"CD",X"FE",X"0B",X"21",X"85",X"93",X"01",X"04",X"17",X"CD",X"FE",X"0B",
		X"21",X"C5",X"90",X"CD",X"FF",X"0B",X"0E",X"07",X"CD",X"0C",X"10",X"3A",X"AD",X"60",X"4F",X"0C",
		X"3E",X"08",X"91",X"47",X"5F",X"AF",X"83",X"10",X"FD",X"DD",X"21",X"00",X"68",X"DD",X"36",X"00",
		X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"01",X"DD",X"36",X"03",X"00",X"DD",X"77",X"04",
		X"11",X"F3",X"0D",X"0E",X"07",X"C3",X"9A",X"0F",X"CF",X"11",X"DD",X"0D",X"0E",X"0F",X"C3",X"9A",
		X"0F",X"CF",X"11",X"C4",X"0D",X"0E",X"0A",X"C3",X"9A",X"0F",X"CF",X"11",X"9A",X"08",X"C3",X"BD",
		X"0F",X"CF",X"11",X"F3",X"0D",X"C3",X"BD",X"0F",X"CF",X"11",X"DD",X"0D",X"CD",X"BD",X"0F",X"06",
		X"10",X"21",X"13",X"90",X"36",X"00",X"2B",X"10",X"FB",X"C9",X"CF",X"11",X"C4",X"0D",X"C3",X"BD",
		X"0F",X"CF",X"11",X"B2",X"0C",X"C3",X"BD",X"0F",X"7C",X"87",X"84",X"5F",X"16",X"00",X"FD",X"19",
		X"26",X"60",X"FD",X"E9",X"1E",X"18",X"FD",X"19",X"FD",X"E9",X"1E",X"30",X"FD",X"19",X"FD",X"E9",
		X"CB",X"46",X"C9",X"CB",X"4E",X"C9",X"CB",X"56",X"C9",X"CB",X"5E",X"C9",X"CB",X"66",X"C9",X"CB",
		X"6E",X"C9",X"CB",X"76",X"C9",X"CB",X"7E",X"C9",X"CB",X"C6",X"C9",X"CB",X"CE",X"C9",X"CB",X"D6",
		X"C9",X"CB",X"DE",X"C9",X"CB",X"E6",X"C9",X"CB",X"EE",X"C9",X"CB",X"F6",X"C9",X"CB",X"FE",X"C9",
		X"CB",X"86",X"C9",X"CB",X"8E",X"C9",X"CB",X"96",X"C9",X"CB",X"9E",X"C9",X"CB",X"A6",X"C9",X"CB",
		X"AE",X"C9",X"CB",X"B6",X"C9",X"CB",X"BE",X"C9",X"00",X"2A",X"09",X"60",X"7C",X"B5",X"C9",X"CF",
		X"22",X"09",X"60",X"CD",X"88",X"0F",X"20",X"FB",X"C9",X"CF",X"C5",X"D5",X"11",X"4F",X"60",X"21",
		X"4B",X"60",X"01",X"25",X"00",X"F3",X"ED",X"B8",X"D1",X"C1",X"DD",X"21",X"27",X"60",X"DD",X"71",
		X"00",X"DD",X"71",X"01",X"DD",X"73",X"02",X"DD",X"72",X"03",X"FB",X"C9",X"CF",X"DD",X"21",X"27",
		X"60",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"7E",X"01",X"B7",X"C8",X"CD",X"03",X"10",X"28",
		X"0A",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"18",X"E6",X"F3",X"DD",X"7E",X"04",X"DD",
		X"77",X"00",X"DD",X"7E",X"06",X"DD",X"77",X"02",X"DD",X"7E",X"07",X"DD",X"77",X"03",X"DD",X"7E",
		X"05",X"DD",X"77",X"01",X"B7",X"28",X"0A",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"18",
		X"DB",X"FB",X"C9",X"00",X"E5",X"37",X"3F",X"ED",X"52",X"E1",X"C9",X"CF",X"2A",X"AB",X"60",X"ED",
		X"5F",X"8C",X"6F",X"3A",X"FC",X"60",X"8D",X"67",X"22",X"AB",X"60",X"1E",X"00",X"51",X"06",X"08",
		X"04",X"CB",X"22",X"30",X"FB",X"CB",X"1A",X"ED",X"52",X"30",X"01",X"19",X"CB",X"3A",X"CB",X"1B",
		X"10",X"F5",X"7D",X"32",X"AD",X"60",X"C9",X"00",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",
		X"DD",X"36",X"02",X"00",X"C9",X"00",X"DD",X"7E",X"00",X"FD",X"86",X"00",X"27",X"DD",X"77",X"00",
		X"DD",X"7E",X"01",X"FD",X"8E",X"01",X"27",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"FD",X"8E",X"02",
		X"27",X"DD",X"77",X"02",X"C9",X"00",X"DD",X"7E",X"00",X"FD",X"96",X"00",X"27",X"DD",X"77",X"00",
		X"DD",X"7E",X"01",X"FD",X"9E",X"01",X"27",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"FD",X"9E",X"02",
		X"27",X"DD",X"77",X"02",X"C9",X"CF",X"FD",X"21",X"12",X"11",X"C3",X"46",X"10",X"CF",X"FD",X"21",
		X"12",X"11",X"C3",X"66",X"10",X"00",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"FD",X"7E",X"01",X"DD",
		X"77",X"01",X"FD",X"7E",X"02",X"DD",X"77",X"02",X"C9",X"00",X"DD",X"7E",X"02",X"FD",X"BE",X"02",
		X"C0",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"C0",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"C9",X"00",
		X"FD",X"21",X"13",X"11",X"C3",X"AA",X"10",X"CF",X"01",X"10",X"27",X"CD",X"DA",X"10",X"01",X"64",
		X"00",X"CD",X"DA",X"10",X"0E",X"01",X"CD",X"DA",X"10",X"C9",X"AF",X"ED",X"42",X"38",X"05",X"C6",
		X"01",X"27",X"18",X"F7",X"09",X"DD",X"77",X"02",X"DD",X"2B",X"C9",X"00",X"21",X"00",X"00",X"01",
		X"01",X"00",X"CD",X"01",X"11",X"0E",X"64",X"CD",X"01",X"11",X"01",X"10",X"27",X"CD",X"01",X"11",
		X"C9",X"DD",X"7E",X"00",X"C6",X"01",X"27",X"D6",X"01",X"28",X"04",X"27",X"09",X"18",X"F8",X"DD",
		X"23",X"C9",X"01",X"00",X"00",X"00",X"CF",X"CD",X"00",X"34",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3A",X"00",X"B0",X"32",X"02",X"60",X"3A",X"5F",X"66",X"B7",X"C8",X"2A",X"00",
		X"60",X"7D",X"E6",X"70",X"6F",X"7C",X"E6",X"0F",X"B5",X"CB",X"64",X"28",X"02",X"CB",X"FF",X"32",
		X"00",X"60",X"C9",X"C9",X"E1",X"FD",X"E1",X"DD",X"E1",X"D1",X"C1",X"C9",X"06",X"03",X"DD",X"21",
		X"CC",X"66",X"C5",X"DD",X"E5",X"CD",X"63",X"11",X"DD",X"E1",X"C1",X"11",X"10",X"00",X"DD",X"19",
		X"10",X"F0",X"C9",X"DD",X"7E",X"01",X"B7",X"C8",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"E5",X"FD",
		X"E1",X"DD",X"35",X"01",X"20",X"05",X"FD",X"36",X"04",X"00",X"C9",X"DD",X"7E",X"00",X"E6",X"03",
		X"28",X"43",X"DD",X"35",X"03",X"20",X"3E",X"DD",X"7E",X"02",X"DD",X"77",X"03",X"DD",X"CB",X"00",
		X"66",X"20",X"1C",X"FD",X"34",X"04",X"FD",X"7E",X"04",X"FE",X"0B",X"38",X"28",X"DD",X"CB",X"00",
		X"4E",X"20",X"06",X"FD",X"36",X"04",X"00",X"18",X"1C",X"DD",X"CB",X"00",X"E6",X"18",X"16",X"FD",
		X"35",X"04",X"F2",X"C5",X"11",X"DD",X"CB",X"00",X"46",X"20",X"06",X"FD",X"36",X"04",X"0A",X"18",
		X"04",X"DD",X"CB",X"00",X"A6",X"DD",X"7E",X"00",X"E6",X"0C",X"C8",X"DD",X"35",X"05",X"C0",X"DD",
		X"7E",X"04",X"DD",X"77",X"05",X"DD",X"35",X"07",X"28",X"3F",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",
		X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"DD",X"CB",X"00",X"6E",X"20",X"03",X"19",X"18",X"03",X"AF",
		X"ED",X"52",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"7D",X"E6",X"0F",X"FD",X"77",X"00",X"7D",X"1F",
		X"1F",X"1F",X"1F",X"E6",X"0F",X"FD",X"77",X"01",X"7C",X"E6",X"0F",X"FD",X"77",X"02",X"7C",X"1F",
		X"1F",X"1F",X"1F",X"E6",X"0F",X"FD",X"77",X"03",X"C9",X"DD",X"7E",X"06",X"DD",X"77",X"07",X"DD",
		X"CB",X"00",X"6E",X"20",X"13",X"DD",X"CB",X"00",X"5E",X"28",X"05",X"DD",X"CB",X"00",X"EE",X"C9",
		X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"18",X"BA",X"DD",X"CB",X"00",X"56",X"28",X"F2",X"DD",X"CB",
		X"00",X"AE",X"C9",X"CF",X"3E",X"03",X"21",X"4F",X"12",X"32",X"24",X"60",X"C3",X"8E",X"14",X"00",
		X"00",X"01",X"00",X"0D",X"08",X"05",X"02",X"02",X"01",X"01",X"03",X"03",X"15",X"60",X"05",X"00",
		X"00",X"01",X"00",X"01",X"CF",X"3E",X"03",X"21",X"6C",X"12",X"18",X"DD",X"00",X"00",X"01",X"00",
		X"0D",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"60",X"CF",X"3E",X"0E",X"21",X"83",
		X"12",X"18",X"C6",X"04",X"02",X"00",X"00",X"0D",X"02",X"50",X"04",X"04",X"00",X"00",X"00",X"00",
		X"15",X"60",X"CF",X"3E",X"02",X"21",X"9A",X"12",X"18",X"AF",X"00",X"03",X"00",X"00",X"06",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"60",X"CF",X"3E",X"02",X"21",X"B5",X"12",X"32",
		X"25",X"60",X"C3",X"98",X"14",X"00",X"02",X"00",X"00",X"0D",X"12",X"08",X"01",X"01",X"00",X"00",
		X"00",X"00",X"1A",X"60",X"CF",X"3E",X"05",X"21",X"CC",X"12",X"18",X"E3",X"00",X"00",X"03",X"00",
		X"06",X"29",X"80",X"10",X"10",X"01",X"01",X"90",X"90",X"1A",X"60",X"02",X"00",X"00",X"01",X"00",
		X"01",X"CF",X"3E",X"02",X"21",X"E9",X"12",X"18",X"C6",X"08",X"02",X"00",X"00",X"06",X"12",X"14",
		X"04",X"04",X"00",X"00",X"00",X"00",X"1A",X"60",X"CF",X"3E",X"0E",X"21",X"00",X"13",X"18",X"AF",
		X"00",X"00",X"03",X"00",X"0D",X"2C",X"18",X"00",X"00",X"01",X"01",X"10",X"10",X"1A",X"60",X"20",
		X"00",X"00",X"02",X"00",X"02",X"CF",X"3E",X"00",X"21",X"21",X"13",X"32",X"26",X"60",X"C3",X"A2",
		X"14",X"00",X"04",X"02",X"00",X"0D",X"12",X"0A",X"01",X"01",X"00",X"00",X"00",X"00",X"1F",X"60",
		X"CF",X"3E",X"0A",X"21",X"38",X"13",X"18",X"E3",X"00",X"04",X"00",X"00",X"0D",X"16",X"1E",X"03",
		X"03",X"03",X"03",X"03",X"03",X"1F",X"60",X"07",X"00",X"50",X"00",X"50",X"00",X"CF",X"3E",X"00",
		X"21",X"55",X"13",X"18",X"C6",X"00",X"08",X"00",X"00",X"0D",X"1D",X"1E",X"03",X"03",X"01",X"01",
		X"06",X"06",X"1F",X"60",X"01",X"00",X"00",X"01",X"00",X"01",X"CF",X"3E",X"00",X"32",X"24",X"60",
		X"3E",X"01",X"32",X"25",X"60",X"3E",X"02",X"32",X"26",X"60",X"21",X"C7",X"13",X"E5",X"E5",X"CD",
		X"8E",X"14",X"E1",X"CD",X"98",X"14",X"E1",X"CD",X"A2",X"14",X"3E",X"15",X"32",X"D4",X"66",X"3E",
		X"1A",X"32",X"E4",X"66",X"3E",X"1F",X"32",X"F4",X"66",X"21",X"ED",X"60",X"34",X"7E",X"FE",X"06",
		X"38",X"02",X"AF",X"77",X"FD",X"21",X"D8",X"13",X"87",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"6E",
		X"00",X"FD",X"66",X"01",X"22",X"D8",X"66",X"22",X"DA",X"66",X"22",X"E8",X"66",X"22",X"EA",X"66",
		X"22",X"F8",X"66",X"22",X"FA",X"66",X"C9",X"00",X"00",X"00",X"00",X"08",X"1E",X"0A",X"03",X"03",
		X"01",X"01",X"03",X"03",X"15",X"60",X"02",X"00",X"80",X"00",X"00",X"01",X"C0",X"00",X"80",X"01",
		X"40",X"01",X"00",X"01",X"CF",X"21",X"04",X"00",X"CD",X"90",X"0F",X"3E",X"03",X"32",X"24",X"60",
		X"3E",X"07",X"32",X"25",X"60",X"3E",X"08",X"32",X"26",X"60",X"21",X"2B",X"14",X"E5",X"E5",X"CD",
		X"8E",X"14",X"E1",X"CD",X"98",X"14",X"E1",X"CD",X"A2",X"14",X"3E",X"15",X"32",X"D4",X"66",X"3E",
		X"1A",X"32",X"E4",X"66",X"3E",X"1F",X"32",X"F4",X"66",X"21",X"ED",X"60",X"34",X"7E",X"FE",X"08",
		X"38",X"02",X"AF",X"77",X"FD",X"21",X"3C",X"14",X"C3",X"A8",X"13",X"00",X"03",X"00",X"00",X"0D",
		X"0C",X"09",X"00",X"00",X"01",X"01",X"05",X"05",X"15",X"60",X"03",X"00",X"30",X"00",X"28",X"00",
		X"20",X"00",X"18",X"00",X"10",X"00",X"50",X"00",X"58",X"00",X"60",X"00",X"CF",X"3E",X"07",X"21",
		X"55",X"14",X"C3",X"AF",X"12",X"00",X"03",X"00",X"00",X"0D",X"2C",X"48",X"00",X"00",X"01",X"01",
		X"12",X"12",X"1A",X"60",X"24",X"00",X"C0",X"01",X"C0",X"01",X"CF",X"3A",X"BF",X"60",X"E6",X"1F",
		X"C0",X"3E",X"02",X"21",X"E9",X"12",X"CD",X"1B",X"13",X"3E",X"1F",X"32",X"F4",X"66",X"C9",X"CF",
		X"3E",X"00",X"21",X"00",X"13",X"CD",X"49",X"12",X"3E",X"15",X"32",X"D4",X"66",X"C9",X"DD",X"21",
		X"15",X"60",X"FD",X"21",X"CC",X"66",X"18",X"12",X"DD",X"21",X"1A",X"60",X"FD",X"21",X"DC",X"66",
		X"18",X"08",X"DD",X"21",X"1F",X"60",X"FD",X"21",X"EC",X"66",X"06",X"05",X"7E",X"DD",X"77",X"00",
		X"DD",X"23",X"23",X"10",X"F7",X"06",X"10",X"7E",X"FD",X"77",X"00",X"23",X"FD",X"23",X"10",X"F7",
		X"C9",X"08",X"0C",X"10",X"09",X"3C",X"5C",X"5D",X"14",X"27",X"5F",X"5E",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"CE",X"CF",X"14",X"27",X"D0",X"D1",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"D2",X"D3",X"14",X"27",X"D4",X"D5",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"D6",X"D7",X"14",X"27",X"D8",X"D9",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"DA",X"DB",X"14",X"27",X"DC",X"DD",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"DE",X"DF",X"14",X"27",X"E0",X"E1",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"E2",X"E3",X"14",X"27",X"E4",X"E5",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0C",X"10",X"09",X"3C",X"03",X"03",X"14",X"27",X"03",X"03",X"18",X"0B",X"22",X"1C",
		X"0A",X"08",X"0D",X"11",X"09",X"3E",X"00",X"00",X"15",X"2A",X"00",X"00",X"19",X"0B",X"23",X"1D",
		X"0A",X"08",X"0E",X"12",X"09",X"3F",X"00",X"00",X"16",X"2F",X"00",X"00",X"1A",X"0B",X"24",X"1E",
		X"0A",X"08",X"0F",X"13",X"09",X"5B",X"00",X"00",X"17",X"3B",X"00",X"00",X"1B",X"0B",X"26",X"1F",
		X"0A",X"08",X"00",X"00",X"09",X"00",X"60",X"C5",X"00",X"00",X"CB",X"C8",X"00",X"0B",X"00",X"00",
		X"0A",X"08",X"00",X"00",X"09",X"00",X"61",X"C6",X"00",X"00",X"CC",X"C9",X"00",X"0B",X"00",X"00",
		X"0A",X"08",X"00",X"00",X"09",X"00",X"C4",X"C7",X"00",X"00",X"CD",X"CA",X"00",X"0B",X"00",X"00",
		X"0A",X"BB",X"FF",X"77",X"E0",X"FF",X"7C",X"E0",X"FF",X"81",X"01",X"00",X"86",X"01",X"00",X"8B",
		X"01",X"00",X"8B",X"01",X"00",X"90",X"01",X"00",X"95",X"20",X"00",X"9A",X"20",X"00",X"9F",X"20",
		X"00",X"9F",X"20",X"00",X"A4",X"20",X"00",X"A9",X"FF",X"FF",X"AE",X"FF",X"FF",X"B3",X"FF",X"FF",
		X"B3",X"FF",X"FF",X"B8",X"FF",X"FF",X"BD",X"E0",X"FF",X"C2",X"E0",X"FF",X"77",X"62",X"6E",X"63",
		X"00",X"00",X"66",X"6A",X"00",X"00",X"66",X"6A",X"6D",X"00",X"66",X"6A",X"6D",X"00",X"62",X"6E",
		X"63",X"00",X"66",X"6A",X"6D",X"6A",X"00",X"00",X"00",X"6D",X"00",X"6B",X"00",X"00",X"6A",X"6B",
		X"6D",X"00",X"6A",X"6B",X"6D",X"00",X"6A",X"00",X"6D",X"00",X"6A",X"6B",X"6D",X"6A",X"00",X"00",
		X"00",X"6C",X"00",X"6C",X"00",X"00",X"6A",X"6B",X"6D",X"00",X"6A",X"6B",X"6D",X"00",X"6A",X"00",
		X"6D",X"00",X"6A",X"6B",X"6D",X"6A",X"00",X"00",X"00",X"6B",X"00",X"6D",X"00",X"00",X"6A",X"6C",
		X"6D",X"00",X"6A",X"6C",X"6D",X"00",X"6A",X"00",X"6D",X"00",X"6A",X"6C",X"6D",X"6A",X"00",X"00",
		X"00",X"66",X"6E",X"6E",X"6A",X"00",X"6A",X"6C",X"6D",X"00",X"6A",X"6C",X"6D",X"00",X"6A",X"00",
		X"6D",X"00",X"6A",X"6C",X"6D",X"64",X"71",X"65",X"6D",X"00",X"00",X"00",X"6B",X"00",X"6A",X"6D",
		X"69",X"00",X"6A",X"6D",X"69",X"00",X"64",X"71",X"65",X"00",X"6A",X"6D",X"69",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"56",X"00",X"47",X"41",X"4D",X"45",X"00",X"47",X"52",
		X"55",X"45",X"4E",X"42",X"45",X"52",X"47",X"00",X"31",X"39",X"38",X"35",X"00",X"00",X"00",X"00",
		X"00",X"66",X"6E",X"63",X"00",X"00",X"66",X"6A",X"00",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"00",X"6D",X"00",X"6D",X"00",X"6B",
		X"00",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"68",X"71",X"65",X"00",X"6C",X"00",X"6C",X"00",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"6E",X"63",X"00",X"6B",X"00",X"6D",
		X"00",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"6A",X"00",X"6D",X"00",X"66",X"6E",X"6E",X"6A",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"71",X"65",X"6D",X"00",X"00",X"00",
		X"6B",X"00",X"68",X"71",X"71",X"00",X"68",X"71",X"71",X"00",X"00",X"00",X"00",X"11",X"11",X"11",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"22",X"21",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"32",X"10",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"44",X"44",X"44",X"43",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"32",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",
		X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"32",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"32",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"32",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"32",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"32",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"32",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"32",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"40",X"00",X"03",X"21",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"03",
		X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"03",X"21",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"04",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"03",
		X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"03",X"21",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"44",X"40",X"00",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"10",X"00",
		X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"03",X"21",X"00",X"00",X"00",X"04",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"32",X"10",X"00",X"00",X"40",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"03",X"21",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"32",
		X"10",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"03",X"21",X"04",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"03",X"21",X"04",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"03",X"21",X"00",X"40",X"00",X"00",X"04",X"00",X"04",X"44",X"40",X"00",X"03",
		X"21",X"00",X"04",X"00",X"00",X"40",X"00",X"40",X"00",X"04",X"00",X"03",X"21",X"00",X"00",X"44",
		X"44",X"00",X"04",X"00",X"00",X"00",X"40",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"04",X"03",X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"03",
		X"21",X"52",X"41",X"4D",X"20",X"20",X"20",X"42",X"41",X"44",X"24",X"49",X"4E",X"54",X"20",X"20",
		X"20",X"42",X"41",X"44",X"24",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"58",X"20",X"52",X"45",
		X"41",X"44",X"59",X"24",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"58",X"24",X"54",X"49",X"44",
		X"45",X"52",X"43",X"24",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"48",X"49",X"2D",X"53",X"43",X"4F",X"52",X"45",X"20",X"20",
		X"24",X"50",X"55",X"53",X"48",X"24",X"52",X"41",X"4E",X"4B",X"20",X"20",X"53",X"43",X"4F",X"52",
		X"45",X"20",X"20",X"20",X"20",X"4E",X"41",X"4D",X"45",X"24",X"55",X"53",X"45",X"20",X"53",X"45",
		X"4C",X"45",X"43",X"54",X"2D",X"42",X"55",X"54",X"54",X"4F",X"4E",X"24",X"20",X"20",X"20",X"20",
		X"46",X"4F",X"52",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"4F",X"46",X"24",X"20",X"20",
		X"20",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"24",X"24",X"45",X"4E",X"44",X"20",X"53",
		X"45",X"4C",X"45",X"43",X"54",X"49",X"4F",X"4E",X"20",X"42",X"59",X"24",X"20",X"20",X"20",X"20",
		X"53",X"54",X"41",X"52",X"54",X"2D",X"42",X"55",X"54",X"54",X"4F",X"4E",X"24",X"46",X"4F",X"52",
		X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"4F",X"46",X"20",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"53",X"24",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"24",X"20",X"31",X"53",
		X"54",X"24",X"20",X"32",X"4E",X"44",X"24",X"20",X"33",X"52",X"44",X"24",X"20",X"34",X"54",X"48",
		X"24",X"20",X"35",X"54",X"48",X"24",X"20",X"36",X"54",X"48",X"24",X"20",X"37",X"54",X"48",X"24",
		X"20",X"38",X"54",X"48",X"24",X"20",X"39",X"54",X"48",X"24",X"31",X"30",X"54",X"48",X"24",X"31",
		X"31",X"54",X"48",X"24",X"31",X"32",X"54",X"48",X"24",X"31",X"33",X"54",X"48",X"24",X"31",X"34",
		X"54",X"48",X"24",X"31",X"35",X"54",X"48",X"24",X"31",X"36",X"54",X"48",X"24",X"31",X"37",X"54",
		X"48",X"24",X"31",X"38",X"54",X"48",X"24",X"31",X"39",X"54",X"48",X"24",X"32",X"30",X"54",X"48",
		X"24",X"55",X"53",X"45",X"20",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"20",X"54",X"4F",
		X"24",X"20",X"20",X"20",X"20",X"57",X"52",X"49",X"54",X"45",X"20",X"4E",X"41",X"4D",X"45",X"24",
		X"24",X"55",X"53",X"45",X"20",X"53",X"50",X"45",X"45",X"44",X"2D",X"42",X"55",X"54",X"54",X"4F",
		X"4E",X"24",X"20",X"20",X"20",X"20",X"54",X"4F",X"20",X"46",X"49",X"4E",X"49",X"53",X"48",X"24",
		X"20",X"20",X"20",X"20",X"45",X"4E",X"54",X"52",X"59",X"24",X"53",X"4C",X"4C",X"41",X"42",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"24",X"54",X"49",X"4D",X"45",
		X"24",X"54",X"56",X"20",X"47",X"41",X"4D",X"45",X"20",X"31",X"39",X"38",X"35",X"24",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"24",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"24",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",
		X"54",X"49",X"4F",X"4E",X"53",X"24",X"21",X"10",X"27",X"DD",X"21",X"0E",X"60",X"CD",X"C8",X"10",
		X"FD",X"21",X"0E",X"60",X"DD",X"21",X"5C",X"66",X"CD",X"96",X"10",X"FD",X"21",X"0E",X"60",X"DD",
		X"21",X"80",X"61",X"06",X"14",X"CD",X"96",X"10",X"11",X"0B",X"00",X"DD",X"19",X"10",X"F6",X"21",
		X"B1",X"93",X"11",X"2D",X"19",X"0E",X"01",X"CD",X"2B",X"0C",X"21",X"02",X"60",X"CB",X"46",X"11",
		X"34",X"19",X"21",X"A0",X"93",X"C4",X"17",X"0C",X"3E",X"02",X"ED",X"47",X"FB",X"AF",X"32",X"06",
		X"A0",X"32",X"03",X"A0",X"32",X"5F",X"66",X"3C",X"32",X"CD",X"60",X"CD",X"E9",X"0E",X"DD",X"21",
		X"FC",X"60",X"CD",X"C0",X"10",X"C2",X"91",X"1C",X"21",X"81",X"93",X"11",X"14",X"00",X"01",X"1C",
		X"1E",X"CD",X"FF",X"0B",X"06",X"0E",X"DD",X"21",X"64",X"93",X"FD",X"21",X"64",X"9F",X"21",X"DD",
		X"15",X"11",X"E0",X"FF",X"C5",X"DD",X"E5",X"FD",X"E5",X"06",X"18",X"7E",X"DD",X"77",X"00",X"78",
		X"E6",X"03",X"C6",X"04",X"00",X"00",X"00",X"23",X"DD",X"19",X"FD",X"19",X"10",X"ED",X"FD",X"E1",
		X"DD",X"E1",X"C1",X"DD",X"23",X"FD",X"23",X"10",X"DB",X"21",X"D9",X"92",X"11",X"AE",X"1A",X"0E",
		X"14",X"CD",X"17",X"0C",X"11",X"E0",X"FF",X"01",X"64",X"00",X"C5",X"21",X"07",X"00",X"CD",X"90",
		X"0F",X"06",X"0E",X"21",X"64",X"9F",X"C5",X"E5",X"06",X"18",X"CD",X"E0",X"32",X"00",X"00",X"00",
		X"00",X"19",X"10",X"F6",X"E1",X"C1",X"23",X"10",X"ED",X"DD",X"21",X"FC",X"60",X"CD",X"C0",X"10",
		X"C1",X"C2",X"91",X"1C",X"0B",X"78",X"B1",X"C2",X"9A",X"1B",X"AF",X"32",X"D4",X"60",X"32",X"71",
		X"61",X"3E",X"03",X"32",X"6F",X"61",X"3E",X"08",X"32",X"70",X"61",X"CD",X"DA",X"02",X"3E",X"01",
		X"32",X"CD",X"60",X"CD",X"01",X"0B",X"CD",X"00",X"26",X"CD",X"FA",X"20",X"CD",X"D6",X"2F",X"CD",
		X"22",X"0F",X"DD",X"21",X"FC",X"60",X"CD",X"C0",X"10",X"C2",X"91",X"1C",X"CD",X"44",X"28",X"38",
		X"16",X"06",X"0F",X"C5",X"21",X"14",X"00",X"CD",X"90",X"0F",X"DD",X"21",X"FC",X"60",X"CD",X"C0",
		X"10",X"C1",X"C2",X"91",X"1C",X"10",X"EC",X"21",X"81",X"93",X"11",X"00",X"00",X"01",X"1A",X"1E",
		X"CD",X"FF",X"0B",X"21",X"DE",X"92",X"0E",X"02",X"11",X"AE",X"1A",X"CD",X"17",X"0C",X"3E",X"64",
		X"32",X"C0",X"60",X"21",X"05",X"00",X"CD",X"90",X"0F",X"DD",X"21",X"FC",X"60",X"CD",X"C0",X"10",
		X"C2",X"91",X"1C",X"21",X"C0",X"60",X"35",X"CA",X"48",X"1B",X"7E",X"E6",X"03",X"4F",X"87",X"87",
		X"47",X"87",X"87",X"87",X"80",X"DD",X"21",X"02",X"29",X"5F",X"16",X"00",X"DD",X"19",X"06",X"09",
		X"FD",X"21",X"7F",X"1C",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"C5",X"DD",X"E5",X"FD",X"E5",X"CD",
		X"E5",X"28",X"FD",X"E1",X"FD",X"23",X"FD",X"23",X"DD",X"E1",X"C1",X"10",X"E7",X"18",X"B4",X"4E",
		X"92",X"46",X"92",X"88",X"91",X"4E",X"91",X"94",X"91",X"56",X"92",X"14",X"93",X"4E",X"93",X"08",
		X"93",X"3E",X"01",X"32",X"06",X"A0",X"CD",X"09",X"0F",X"AF",X"32",X"5F",X"66",X"32",X"01",X"A0",
		X"21",X"81",X"93",X"11",X"18",X"00",X"01",X"1A",X"1F",X"CD",X"FF",X"0B",X"21",X"F5",X"92",X"11",
		X"6A",X"19",X"01",X"19",X"06",X"CD",X"E0",X"0B",X"CD",X"95",X"0E",X"AF",X"32",X"D4",X"60",X"CD",
		X"92",X"29",X"21",X"01",X"60",X"CB",X"6E",X"CA",X"EF",X"1C",X"21",X"01",X"60",X"CB",X"76",X"20",
		X"F1",X"3A",X"D4",X"60",X"C6",X"11",X"32",X"D4",X"60",X"E6",X"0F",X"FE",X"06",X"28",X"DC",X"4F",
		X"3A",X"FD",X"60",X"B7",X"20",X"D9",X"3A",X"FC",X"60",X"3D",X"B9",X"38",X"CE",X"18",X"D0",X"3A",
		X"D4",X"60",X"E6",X"0F",X"3C",X"32",X"0E",X"60",X"21",X"00",X"00",X"22",X"0F",X"60",X"FD",X"21",
		X"0E",X"60",X"DD",X"21",X"FC",X"60",X"CD",X"66",X"10",X"21",X"05",X"93",X"11",X"19",X"00",X"01",
		X"12",X"17",X"CD",X"FF",X"0B",X"01",X"19",X"06",X"11",X"41",X"1A",X"21",X"F5",X"92",X"CD",X"E0",
		X"0B",X"21",X"2C",X"01",X"22",X"88",X"98",X"AF",X"32",X"ED",X"60",X"3A",X"ED",X"60",X"F5",X"21",
		X"06",X"93",X"87",X"5F",X"16",X"00",X"19",X"0E",X"04",X"11",X"24",X"19",X"CD",X"17",X"0C",X"11",
		X"20",X"00",X"19",X"F1",X"C6",X"31",X"77",X"11",X"C0",X"FF",X"19",X"22",X"E8",X"60",X"22",X"EA",
		X"60",X"CB",X"47",X"20",X"0B",X"21",X"02",X"60",X"CB",X"56",X"20",X"04",X"3E",X"01",X"18",X"01",
		X"AF",X"32",X"01",X"A0",X"32",X"5F",X"66",X"AF",X"32",X"FF",X"60",X"3A",X"ED",X"60",X"87",X"67",
		X"3A",X"FF",X"60",X"6F",X"29",X"29",X"29",X"EB",X"21",X"82",X"D4",X"AF",X"ED",X"52",X"22",X"C3",
		X"60",X"06",X"05",X"DD",X"21",X"A2",X"1D",X"C5",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E7",X"C1",
		X"28",X"09",X"11",X"04",X"00",X"DD",X"19",X"10",X"EE",X"18",X"E6",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"E9",X"00",X"07",X"06",X"1E",X"00",X"03",X"DE",X"1D",X"00",X"00",X"F3",X"1D",X"00",X"02",
		X"B6",X"1D",X"00",X"01",X"D5",X"1D",X"3A",X"FF",X"60",X"11",X"E0",X"FF",X"3C",X"E6",X"07",X"32",
		X"FF",X"60",X"2A",X"E8",X"60",X"19",X"CB",X"C4",X"CB",X"8C",X"22",X"E8",X"60",X"21",X"0F",X"00",
		X"CD",X"90",X"0F",X"18",X"96",X"3A",X"FF",X"60",X"3D",X"11",X"20",X"00",X"18",X"DF",X"2A",X"E8",
		X"60",X"35",X"7E",X"FE",X"FF",X"20",X"04",X"36",X"5A",X"18",X"E2",X"FE",X"41",X"30",X"DE",X"36",
		X"00",X"18",X"DA",X"2A",X"E8",X"60",X"34",X"7E",X"FE",X"01",X"20",X"04",X"36",X"41",X"18",X"CD",
		X"FE",X"5B",X"38",X"C9",X"18",X"E9",X"3A",X"ED",X"60",X"57",X"1E",X"00",X"CB",X"3A",X"CB",X"1B",
		X"DD",X"21",X"75",X"68",X"DD",X"19",X"2A",X"EA",X"60",X"11",X"E0",X"FF",X"06",X"08",X"7E",X"DD",
		X"77",X"00",X"19",X"DD",X"23",X"10",X"F7",X"21",X"14",X"00",X"CD",X"90",X"0F",X"3A",X"D4",X"60",
		X"21",X"ED",X"60",X"E6",X"0F",X"34",X"BE",X"D2",X"2B",X"1D",X"3A",X"D4",X"60",X"E6",X"F0",X"32",
		X"D4",X"60",X"CD",X"02",X"0F",X"DD",X"21",X"72",X"61",X"CD",X"38",X"10",X"AF",X"32",X"71",X"61",
		X"3E",X"08",X"32",X"70",X"61",X"3A",X"02",X"60",X"1F",X"1F",X"1F",X"E6",X"03",X"C6",X"03",X"32",
		X"6F",X"61",X"CD",X"DA",X"02",X"11",X"00",X"68",X"06",X"06",X"C5",X"21",X"00",X"61",X"01",X"75",
		X"00",X"ED",X"B0",X"21",X"0B",X"00",X"19",X"EB",X"C1",X"10",X"EF",X"AF",X"32",X"CD",X"60",X"3A",
		X"D4",X"60",X"E6",X"07",X"57",X"1E",X"00",X"CB",X"3A",X"CB",X"1B",X"21",X"00",X"68",X"19",X"11",
		X"00",X"61",X"01",X"80",X"00",X"ED",X"B0",X"CD",X"01",X"0B",X"11",X"8A",X"1A",X"21",X"50",X"90",
		X"0E",X"01",X"CD",X"2B",X"0C",X"3A",X"6F",X"61",X"47",X"21",X"4B",X"90",X"05",X"28",X"0E",X"36",
		X"72",X"CB",X"D4",X"00",X"00",X"CB",X"94",X"2D",X"7D",X"FE",X"B1",X"20",X"EF",X"21",X"A0",X"93",
		X"11",X"34",X"19",X"0E",X"01",X"CD",X"17",X"0C",X"3A",X"D4",X"60",X"E6",X"0F",X"CB",X"47",X"F5",
		X"C6",X"31",X"32",X"C0",X"92",X"06",X"08",X"21",X"F4",X"93",X"11",X"75",X"61",X"1A",X"77",X"2B",
		X"13",X"10",X"FA",X"F1",X"28",X"09",X"21",X"02",X"60",X"CB",X"56",X"3E",X"03",X"28",X"01",X"AF",
		X"32",X"5F",X"66",X"32",X"01",X"A0",X"11",X"15",X"19",X"21",X"DA",X"92",X"0E",X"04",X"CD",X"17",
		X"0C",X"3A",X"D4",X"60",X"E6",X"0F",X"C6",X"31",X"32",X"FA",X"91",X"CD",X"00",X"26",X"06",X"0E",
		X"21",X"DA",X"92",X"11",X"E0",X"FF",X"36",X"00",X"19",X"10",X"FB",X"CD",X"FA",X"20",X"21",X"32",
		X"00",X"CD",X"90",X"0F",X"CD",X"D6",X"2F",X"3A",X"EC",X"60",X"CB",X"47",X"20",X"14",X"21",X"71",
		X"61",X"34",X"7E",X"E6",X"03",X"FE",X"03",X"20",X"04",X"34",X"CD",X"53",X"2A",X"CD",X"DA",X"02",
		X"18",X"04",X"21",X"6F",X"61",X"35",X"CD",X"5F",X"20",X"3A",X"D4",X"60",X"E6",X"0F",X"57",X"1E",
		X"00",X"CB",X"3A",X"CB",X"1B",X"21",X"00",X"68",X"19",X"EB",X"01",X"80",X"00",X"21",X"00",X"61",
		X"ED",X"B0",X"3A",X"EC",X"60",X"CB",X"47",X"CA",X"7B",X"1E",X"06",X"06",X"3A",X"D4",X"60",X"3C",
		X"32",X"D4",X"60",X"5F",X"E6",X"0F",X"57",X"7B",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"BA",X"30",X"08",X"3A",X"D4",X"60",X"E6",X"F0",X"32",X"D4",X"60",X"3A",X"D4",X"60",X"E6",X"0F",
		X"57",X"1E",X"00",X"CB",X"3A",X"CB",X"1B",X"21",X"6F",X"68",X"19",X"7E",X"B7",X"C2",X"7B",X"1E",
		X"10",X"CA",X"21",X"81",X"93",X"11",X"18",X"00",X"01",X"1A",X"1F",X"CD",X"FF",X"0B",X"21",X"02",
		X"60",X"CB",X"46",X"CA",X"56",X"20",X"06",X"06",X"21",X"71",X"68",X"11",X"80",X"00",X"3E",X"31",
		X"77",X"3C",X"19",X"10",X"FB",X"06",X"06",X"C5",X"DD",X"21",X"72",X"68",X"FD",X"21",X"F2",X"68",
		X"06",X"05",X"CD",X"A9",X"10",X"30",X"1E",X"C5",X"DD",X"E5",X"FD",X"E5",X"06",X"0C",X"DD",X"5E",
		X"FF",X"FD",X"56",X"FF",X"DD",X"72",X"FF",X"FD",X"73",X"FF",X"DD",X"23",X"FD",X"23",X"10",X"EE",
		X"FD",X"E1",X"DD",X"E1",X"C1",X"11",X"80",X"00",X"DD",X"19",X"FD",X"19",X"10",X"D4",X"C1",X"10",
		X"C6",X"FD",X"21",X"72",X"68",X"06",X"06",X"21",X"65",X"93",X"FD",X"7E",X"00",X"FD",X"B6",X"01",
		X"FD",X"B6",X"02",X"28",X"38",X"C5",X"E5",X"FD",X"E5",X"11",X"24",X"19",X"0E",X"04",X"CD",X"17",
		X"0C",X"11",X"20",X"00",X"19",X"FD",X"7E",X"FF",X"77",X"E5",X"DD",X"E1",X"11",X"A0",X"FE",X"DD",
		X"19",X"11",X"18",X"00",X"CD",X"9D",X"02",X"11",X"C0",X"FF",X"19",X"11",X"E0",X"FF",X"06",X"08",
		X"FD",X"7E",X"03",X"77",X"FD",X"23",X"19",X"10",X"F7",X"FD",X"E1",X"E1",X"C1",X"11",X"80",X"00",
		X"FD",X"19",X"23",X"23",X"10",X"B4",X"21",X"18",X"01",X"CD",X"90",X"0F",X"C3",X"2D",X"1B",X"3A",
		X"6F",X"61",X"B7",X"C0",X"21",X"CD",X"60",X"CB",X"46",X"C0",X"11",X"24",X"19",X"21",X"7A",X"92",
		X"0E",X"04",X"CD",X"17",X"0C",X"3A",X"D4",X"60",X"E6",X"0F",X"C6",X"31",X"32",X"9A",X"91",X"11",
		X"D3",X"19",X"21",X"7B",X"92",X"CD",X"17",X"0C",X"21",X"82",X"00",X"CD",X"90",X"0F",X"21",X"02",
		X"60",X"CB",X"46",X"C8",X"FD",X"21",X"72",X"61",X"DD",X"21",X"80",X"61",X"06",X"14",X"11",X"0B",
		X"00",X"CD",X"A9",X"10",X"38",X"05",X"DD",X"19",X"10",X"F7",X"C9",X"11",X"5B",X"66",X"21",X"50",
		X"66",X"05",X"C5",X"28",X"0B",X"78",X"87",X"80",X"87",X"87",X"90",X"06",X"00",X"4F",X"ED",X"B8",
		X"CD",X"95",X"10",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"06",X"08",X"11",X"75",X"61",X"1A",X"DD",
		X"77",X"00",X"13",X"DD",X"23",X"10",X"F7",X"CD",X"44",X"28",X"C1",X"3E",X"13",X"90",X"FD",X"21",
		X"48",X"47",X"5F",X"16",X"00",X"FD",X"19",X"06",X"17",X"11",X"E0",X"FF",X"FD",X"36",X"00",X"19",
		X"FD",X"19",X"10",X"F8",X"21",X"C8",X"00",X"C3",X"90",X"0F",X"21",X"FF",X"60",X"35",X"20",X"13",
		X"2A",X"C0",X"60",X"E5",X"D1",X"06",X"06",X"CB",X"3A",X"CB",X"1B",X"10",X"FA",X"AF",X"ED",X"52",
		X"22",X"C0",X"60",X"2A",X"C0",X"60",X"3A",X"CD",X"60",X"CB",X"4F",X"C0",X"3A",X"EC",X"60",X"FE",
		X"04",X"28",X"08",X"2B",X"7C",X"B5",X"20",X"EE",X"C3",X"84",X"21",X"21",X"CD",X"60",X"CB",X"D6",
		X"21",X"00",X"00",X"CD",X"DF",X"2F",X"21",X"70",X"61",X"7E",X"CD",X"50",X"35",X"F5",X"CD",X"4C",
		X"14",X"F1",X"F5",X"87",X"4F",X"87",X"81",X"FD",X"21",X"D6",X"26",X"5F",X"16",X"00",X"FD",X"19",
		X"06",X"0C",X"00",X"00",X"00",X"FD",X"AE",X"00",X"32",X"80",X"98",X"FD",X"23",X"21",X"06",X"00",
		X"CD",X"90",X"0F",X"10",X"ED",X"F1",X"FE",X"02",X"28",X"12",X"CD",X"B2",X"26",X"AF",X"32",X"EC",
		X"60",X"CD",X"EB",X"07",X"21",X"CD",X"60",X"CB",X"96",X"C3",X"FA",X"20",X"3E",X"01",X"32",X"6F",
		X"61",X"C3",X"AC",X"23",X"2A",X"E2",X"60",X"AF",X"32",X"ED",X"60",X"CD",X"E3",X"25",X"38",X"1B",
		X"2A",X"E4",X"60",X"3E",X"0B",X"32",X"ED",X"60",X"CD",X"E3",X"25",X"38",X"0E",X"2A",X"E6",X"60",
		X"3E",X"16",X"32",X"ED",X"60",X"CD",X"E3",X"25",X"D2",X"A2",X"23",X"ED",X"43",X"E8",X"60",X"ED",
		X"53",X"EA",X"60",X"3E",X"14",X"BA",X"DA",X"F0",X"22",X"BB",X"DA",X"F0",X"22",X"21",X"CD",X"60",
		X"CB",X"D6",X"CD",X"28",X"0D",X"C6",X"18",X"21",X"5F",X"66",X"AE",X"32",X"FA",X"67",X"21",X"00",
		X"00",X"CD",X"DF",X"2F",X"3A",X"ED",X"60",X"5F",X"16",X"00",X"FD",X"21",X"4E",X"61",X"FD",X"19",
		X"06",X"0F",X"C5",X"FD",X"E5",X"21",X"64",X"00",X"DD",X"21",X"0E",X"60",X"CD",X"C8",X"10",X"CD",
		X"C2",X"26",X"FD",X"E1",X"06",X"04",X"C5",X"FD",X"E5",X"CD",X"70",X"35",X"78",X"87",X"87",X"4F",
		X"87",X"87",X"87",X"81",X"DD",X"21",X"DE",X"28",X"5F",X"16",X"00",X"DD",X"19",X"78",X"E6",X"01",
		X"C6",X"18",X"4F",X"CD",X"CC",X"28",X"FD",X"E1",X"C1",X"10",X"DB",X"C1",X"10",X"C4",X"FD",X"36",
		X"0A",X"00",X"21",X"58",X"61",X"06",X"03",X"11",X"0B",X"00",X"7E",X"B7",X"C2",X"C4",X"22",X"19",
		X"10",X"F8",X"21",X"98",X"3A",X"22",X"C0",X"60",X"21",X"81",X"93",X"06",X"1A",X"C5",X"E5",X"06",
		X"18",X"7E",X"B7",X"C4",X"6A",X"22",X"23",X"10",X"F8",X"E1",X"C1",X"11",X"E0",X"FF",X"19",X"10",
		X"EC",X"06",X"08",X"C5",X"78",X"CD",X"D7",X"01",X"21",X"0A",X"00",X"CD",X"90",X"0F",X"C1",X"10",
		X"F2",X"21",X"6F",X"61",X"34",X"3E",X"02",X"C3",X"AE",X"23",X"E5",X"C5",X"36",X"00",X"87",X"4F",
		X"87",X"87",X"81",X"6F",X"26",X"00",X"DD",X"21",X"0E",X"60",X"CD",X"C8",X"10",X"CD",X"C2",X"26",
		X"CD",X"80",X"35",X"2A",X"C0",X"60",X"7C",X"ED",X"44",X"28",X"04",X"5F",X"16",X"FF",X"19",X"22",
		X"C0",X"60",X"2B",X"7C",X"B5",X"20",X"FB",X"21",X"CC",X"60",X"3A",X"BF",X"60",X"CB",X"67",X"28",
		X"08",X"E6",X"0F",X"ED",X"44",X"C6",X"20",X"18",X"04",X"E6",X"0F",X"C6",X"10",X"77",X"E5",X"CD",
		X"28",X"0D",X"C6",X"14",X"4F",X"E1",X"7E",X"E6",X"04",X"81",X"21",X"5F",X"66",X"AE",X"32",X"FA",
		X"67",X"C1",X"E1",X"C9",X"3A",X"ED",X"60",X"FE",X"0B",X"20",X"06",X"DD",X"21",X"E4",X"60",X"18",
		X"0C",X"38",X"06",X"DD",X"21",X"E6",X"60",X"18",X"04",X"DD",X"21",X"E2",X"60",X"DD",X"36",X"00",
		X"00",X"DD",X"36",X"01",X"00",X"CD",X"EB",X"07",X"21",X"CD",X"60",X"CB",X"96",X"C3",X"BE",X"25",
		X"2A",X"EA",X"60",X"11",X"04",X"00",X"06",X"0B",X"DD",X"21",X"06",X"27",X"7C",X"DD",X"BE",X"00",
		X"30",X"10",X"DD",X"BE",X"01",X"38",X"0B",X"7D",X"DD",X"BE",X"02",X"30",X"05",X"DD",X"BE",X"03",
		X"30",X"07",X"DD",X"19",X"10",X"E6",X"C3",X"BE",X"25",X"05",X"78",X"87",X"2A",X"E8",X"60",X"CB",
		X"7C",X"28",X"02",X"C6",X"16",X"CB",X"7D",X"28",X"02",X"C6",X"2C",X"5F",X"16",X"00",X"DD",X"21",
		X"32",X"27",X"DD",X"19",X"DD",X"7E",X"00",X"CD",X"9E",X"27",X"DD",X"7E",X"01",X"DD",X"E5",X"CD",
		X"9E",X"27",X"DD",X"E1",X"DA",X"BE",X"25",X"DD",X"E5",X"DD",X"21",X"4E",X"61",X"3A",X"ED",X"60",
		X"5F",X"DD",X"19",X"DD",X"E1",X"DD",X"5E",X"01",X"DD",X"21",X"89",X"27",X"16",X"00",X"DD",X"19",
		X"0E",X"02",X"CD",X"0C",X"10",X"3A",X"AD",X"60",X"DD",X"86",X"00",X"E6",X"0F",X"CD",X"D6",X"27",
		X"21",X"64",X"00",X"DD",X"21",X"0E",X"60",X"CD",X"C8",X"10",X"CD",X"C2",X"26",X"CD",X"40",X"35",
		X"21",X"0C",X"02",X"22",X"F2",X"67",X"06",X"0A",X"21",X"05",X"00",X"CD",X"90",X"0F",X"3A",X"F3",
		X"67",X"3C",X"E6",X"03",X"32",X"F3",X"67",X"10",X"EF",X"21",X"04",X"02",X"22",X"F2",X"67",X"C3",
		X"BE",X"25",X"3A",X"C4",X"60",X"FE",X"0C",X"30",X"12",X"CD",X"6B",X"13",X"3E",X"01",X"32",X"EC",
		X"60",X"CD",X"22",X"0F",X"21",X"64",X"00",X"CD",X"90",X"0F",X"C9",X"2A",X"C3",X"60",X"7C",X"C6",
		X"FE",X"57",X"7D",X"C6",X"FA",X"5F",X"E6",X"07",X"28",X"12",X"FE",X"07",X"28",X"0E",X"7A",X"E6",
		X"07",X"28",X"05",X"FE",X"07",X"C2",X"A2",X"24",X"0E",X"02",X"18",X"17",X"7A",X"E6",X"07",X"28",
		X"08",X"FE",X"07",X"28",X"04",X"0E",X"03",X"18",X"0A",X"4F",X"7B",X"E6",X"07",X"B9",X"0E",X"00",
		X"28",X"01",X"0C",X"C5",X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"4F",X"00",X"00",X"00",X"3E",
		X"FF",X"00",X"E6",X"C0",X"6F",X"3E",X"FF",X"00",X"1F",X"1F",X"E6",X"30",X"B5",X"C6",X"30",X"91",
		X"4F",X"7B",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"00",X"90",X"11",X"20",X"00",X"3D",X"FA",
		X"25",X"24",X"19",X"18",X"F9",X"59",X"19",X"C1",X"7E",X"B7",X"28",X"76",X"C5",X"36",X"00",X"CD",
		X"00",X"32",X"E5",X"81",X"6F",X"26",X"00",X"DD",X"21",X"0E",X"60",X"CD",X"C8",X"10",X"CD",X"C2",
		X"26",X"CD",X"15",X"13",X"E1",X"CD",X"20",X"35",X"00",X"E6",X"07",X"3D",X"FA",X"53",X"24",X"CB",
		X"09",X"18",X"F8",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"7D",
		X"E6",X"03",X"47",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"EB",X"21",X"1C",X"02",X"AF",
		X"ED",X"52",X"E5",X"D1",X"29",X"19",X"58",X"19",X"11",X"00",X"61",X"19",X"79",X"A6",X"77",X"C1",
		X"79",X"FE",X"02",X"30",X"0D",X"B7",X"3E",X"14",X"28",X"02",X"3E",X"1C",X"21",X"CE",X"60",X"96",
		X"18",X"0B",X"3A",X"CE",X"60",X"20",X"02",X"EE",X"08",X"4F",X"3E",X"10",X"91",X"CD",X"D6",X"27",
		X"18",X"00",X"3A",X"C4",X"60",X"FE",X"1B",X"D2",X"5D",X"25",X"FE",X"17",X"DA",X"5D",X"25",X"3A",
		X"CE",X"60",X"FE",X"04",X"DA",X"7E",X"25",X"FE",X"0D",X"D2",X"7E",X"25",X"3A",X"70",X"61",X"FE",
		X"06",X"20",X"06",X"FD",X"21",X"2D",X"25",X"18",X"0C",X"38",X"06",X"FD",X"21",X"27",X"25",X"18",
		X"04",X"FD",X"21",X"33",X"25",X"3A",X"C3",X"60",X"21",X"CB",X"60",X"96",X"FD",X"BE",X"00",X"30",
		X"06",X"FD",X"21",X"39",X"25",X"18",X"2A",X"FD",X"BE",X"01",X"30",X"06",X"FD",X"21",X"42",X"25",
		X"18",X"1F",X"FD",X"BE",X"02",X"30",X"06",X"FD",X"21",X"4B",X"25",X"18",X"14",X"FD",X"BE",X"03",
		X"30",X"DF",X"FD",X"BE",X"04",X"30",X"E5",X"FD",X"BE",X"05",X"DA",X"7E",X"25",X"FD",X"21",X"54",
		X"25",X"3A",X"CE",X"60",X"D6",X"04",X"5F",X"16",X"00",X"FD",X"19",X"CD",X"30",X"35",X"CD",X"D6",
		X"27",X"CD",X"4D",X"13",X"C3",X"7E",X"25",X"05",X"08",X"0B",X"FB",X"F8",X"F5",X"03",X"06",X"09",
		X"FD",X"FA",X"F7",X"03",X"05",X"07",X"FD",X"FB",X"F9",X"03",X"03",X"02",X"01",X"00",X"0F",X"0E",
		X"0D",X"0D",X"00",X"01",X"03",X"02",X"01",X"0E",X"0D",X"0E",X"0F",X"0D",X"0D",X"0E",X"0F",X"00",
		X"0F",X"0E",X"0D",X"0D",X"03",X"03",X"02",X"01",X"00",X"01",X"02",X"03",X"03",X"3A",X"C4",X"60",
		X"FE",X"FE",X"38",X"1A",X"3A",X"CE",X"60",X"EE",X"08",X"4F",X"3E",X"10",X"91",X"FE",X"08",X"20",
		X"0A",X"0E",X"07",X"CD",X"0C",X"10",X"3A",X"AD",X"60",X"C6",X"05",X"CD",X"D6",X"27",X"3A",X"C3",
		X"60",X"FE",X"20",X"30",X"1B",X"3A",X"CE",X"60",X"FE",X"0A",X"30",X"32",X"B7",X"28",X"1E",X"FE",
		X"08",X"28",X"1A",X"4F",X"3E",X"10",X"91",X"4F",X"E6",X"03",X"20",X"01",X"0C",X"79",X"18",X"0E",
		X"3A",X"C3",X"60",X"FE",X"EC",X"38",X"17",X"3A",X"CE",X"60",X"B7",X"20",X"06",X"3C",X"CD",X"D6",
		X"27",X"18",X"0B",X"FE",X"08",X"20",X"03",X"3D",X"18",X"F4",X"38",X"02",X"18",X"D5",X"2A",X"C3",
		X"60",X"3A",X"CF",X"60",X"EE",X"01",X"32",X"CF",X"60",X"CB",X"47",X"20",X"06",X"ED",X"5B",X"D0",
		X"60",X"18",X"04",X"ED",X"5B",X"D2",X"60",X"7C",X"82",X"67",X"7D",X"83",X"6F",X"22",X"C3",X"60",
		X"C3",X"FA",X"20",X"7C",X"B5",X"C8",X"3A",X"C3",X"60",X"95",X"4F",X"30",X"02",X"ED",X"44",X"FE",
		X"1A",X"D0",X"5F",X"3A",X"C4",X"60",X"94",X"47",X"30",X"02",X"ED",X"44",X"57",X"FE",X"1A",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"06",X"32",X"81",X"98",
		X"CD",X"B2",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",
		X"88",X"10",X"00",X"22",X"CB",X"60",X"CD",X"85",X"26",X"3A",X"71",X"61",X"DD",X"21",X"55",X"26",
		X"87",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"22",X"C0",X"60",X"CD",
		X"EB",X"07",X"AF",X"32",X"EC",X"60",X"21",X"00",X"00",X"CD",X"DF",X"2F",X"CD",X"8C",X"0E",X"21",
		X"A0",X"00",X"C3",X"90",X"0F",X"40",X"01",X"40",X"01",X"54",X"01",X"00",X"00",X"18",X"01",X"18",
		X"01",X"40",X"01",X"00",X"00",X"FA",X"00",X"FA",X"00",X"2C",X"01",X"00",X"00",X"C8",X"00",X"C8",
		X"00",X"FA",X"00",X"00",X"00",X"96",X"00",X"96",X"00",X"C8",X"00",X"00",X"00",X"64",X"00",X"64",
		X"00",X"96",X"00",X"00",X"00",X"21",X"01",X"02",X"22",X"88",X"98",X"0E",X"08",X"CD",X"0C",X"10",
		X"3A",X"AD",X"60",X"DD",X"21",X"C3",X"60",X"C6",X"80",X"DD",X"77",X"00",X"DD",X"36",X"01",X"20",
		X"0E",X"06",X"CD",X"0C",X"10",X"3A",X"AD",X"60",X"3C",X"FE",X"04",X"38",X"02",X"C6",X"09",X"C3",
		X"D6",X"27",X"3A",X"70",X"61",X"87",X"4F",X"3E",X"14",X"91",X"21",X"5F",X"66",X"AE",X"32",X"80",
		X"98",X"C9",X"21",X"CD",X"60",X"CB",X"46",X"C0",X"DD",X"21",X"72",X"61",X"FD",X"21",X"0E",X"60",
		X"CD",X"46",X"10",X"DD",X"E5",X"FD",X"E1",X"DD",X"21",X"5C",X"66",X"CD",X"AA",X"10",X"D0",X"C3",
		X"96",X"10",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1E",X"00",X"1E",X"00",X"0D",X"10",
		X"0D",X"10",X"0D",X"10",X"0D",X"10",X"0D",X"10",X"0D",X"10",X"0D",X"10",X"0A",X"0A",X"07",X"0A",
		X"07",X"0A",X"07",X"0A",X"07",X"0A",X"18",X"14",X"03",X"00",X"18",X"14",X"07",X"02",X"18",X"14",
		X"0B",X"06",X"18",X"14",X"0F",X"0A",X"18",X"13",X"13",X"0E",X"16",X"10",X"16",X"10",X"13",X"0E",
		X"18",X"13",X"0F",X"0A",X"18",X"14",X"0B",X"06",X"18",X"14",X"07",X"02",X"18",X"14",X"03",X"00",
		X"18",X"14",X"0F",X"10",X"00",X"10",X"10",X"11",X"00",X"11",X"12",X"11",X"00",X"12",X"12",X"13",
		X"00",X"13",X"13",X"14",X"00",X"14",X"01",X"14",X"10",X"0F",X"00",X"0F",X"0E",X"0F",X"00",X"0E",
		X"0D",X"0E",X"00",X"0D",X"0D",X"0C",X"00",X"0C",X"0B",X"0C",X"00",X"0B",X"0A",X"0B",X"06",X"05",
		X"00",X"05",X"04",X"05",X"00",X"04",X"03",X"04",X"00",X"03",X"03",X"02",X"00",X"02",X"01",X"02",
		X"00",X"01",X"14",X"01",X"05",X"06",X"00",X"06",X"06",X"07",X"00",X"07",X"08",X"07",X"00",X"08",
		X"09",X"08",X"00",X"09",X"09",X"0A",X"00",X"0A",X"0B",X"0A",X"00",X"01",X"02",X"03",X"04",X"04",
		X"05",X"06",X"07",X"08",X"08",X"09",X"0A",X"0B",X"0C",X"0C",X"0D",X"0E",X"0F",X"00",X"DD",X"E5",
		X"B7",X"28",X"30",X"3D",X"CB",X"3F",X"0E",X"01",X"30",X"02",X"0E",X"10",X"21",X"ED",X"60",X"5E",
		X"83",X"5F",X"16",X"00",X"DD",X"21",X"4E",X"61",X"DD",X"19",X"79",X"FE",X"01",X"DD",X"7E",X"00",
		X"28",X"08",X"91",X"38",X"0E",X"DD",X"77",X"00",X"18",X"09",X"E6",X"0F",X"37",X"28",X"04",X"DD",
		X"35",X"00",X"AF",X"DD",X"E1",X"C9",X"E6",X"0F",X"32",X"CE",X"60",X"87",X"DD",X"21",X"04",X"28",
		X"87",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"7E",X"00",X"32",X"D0",X"60",X"DD",X"7E",X"01",X"32",
		X"D1",X"60",X"DD",X"7E",X"02",X"32",X"D2",X"60",X"DD",X"7E",X"03",X"32",X"D3",X"60",X"21",X"CF",
		X"60",X"CB",X"C6",X"C9",X"00",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",
		X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",
		X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"01",X"21",X"81",X"93",X"01",X"1A",X"1E",X"11",X"18",X"00",X"CD",X"FF",X"0B",
		X"0E",X"19",X"11",X"AE",X"1A",X"21",X"DD",X"92",X"CD",X"17",X"0C",X"21",X"02",X"60",X"CB",X"46",
		X"20",X"02",X"37",X"C9",X"11",X"DD",X"19",X"21",X"A4",X"28",X"06",X"14",X"CD",X"CD",X"0B",X"06",
		X"14",X"DD",X"21",X"68",X"91",X"21",X"83",X"61",X"11",X"04",X"00",X"C5",X"DD",X"E5",X"06",X"08",
		X"7E",X"DD",X"77",X"00",X"11",X"E0",X"FF",X"23",X"DD",X"19",X"10",X"F4",X"11",X"03",X"00",X"19",
		X"DD",X"E1",X"C1",X"DD",X"23",X"10",X"E4",X"11",X"56",X"19",X"21",X"46",X"93",X"0E",X"03",X"CD",
		X"17",X"0C",X"AF",X"C9",X"80",X"61",X"8B",X"61",X"96",X"61",X"A1",X"61",X"AC",X"61",X"B7",X"61",
		X"C2",X"61",X"CD",X"61",X"D8",X"61",X"E3",X"61",X"EE",X"61",X"F9",X"61",X"04",X"62",X"0F",X"62",
		X"1A",X"62",X"25",X"62",X"30",X"62",X"3B",X"62",X"46",X"62",X"51",X"62",X"FD",X"7E",X"0A",X"E6",
		X"07",X"FD",X"21",X"48",X"04",X"87",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",
		X"01",X"11",X"1F",X"00",X"19",X"11",X"E0",X"FF",X"06",X"06",X"C5",X"E5",X"06",X"06",X"DD",X"7E",
		X"00",X"77",X"CD",X"D0",X"32",X"00",X"00",X"19",X"DD",X"23",X"10",X"F2",X"E1",X"23",X"C1",X"10",
		X"E9",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EA",X"EB",X"00",X"00",X"00",X"00",X"EC",X"ED",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"EF",X"F0",X"F1",X"00",X"00",X"F2",X"01",X"01",X"F3",X"00",X"00",X"F4",X"01",X"01",
		X"F5",X"00",X"00",X"F6",X"F7",X"F8",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EF",
		X"EF",X"F0",X"F0",X"F1",X"F2",X"01",X"01",X"01",X"01",X"F3",X"F2",X"01",X"01",X"01",X"01",X"F3",
		X"F4",X"01",X"01",X"01",X"01",X"F5",X"F4",X"01",X"01",X"01",X"01",X"F5",X"F6",X"F7",X"F7",X"F8",
		X"F8",X"F9",X"06",X"06",X"3A",X"D4",X"60",X"E6",X"0F",X"F5",X"DD",X"21",X"07",X"2A",X"4F",X"C5",
		X"CB",X"79",X"0E",X"18",X"20",X"02",X"0E",X"07",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"21",
		X"13",X"2A",X"CD",X"EC",X"29",X"DD",X"23",X"DD",X"23",X"C1",X"0D",X"10",X"E2",X"F1",X"87",X"87",
		X"FD",X"21",X"23",X"2A",X"87",X"5F",X"16",X"00",X"FD",X"19",X"21",X"0B",X"92",X"0E",X"19",X"06",
		X"02",X"CD",X"EE",X"29",X"CD",X"10",X"35",X"E6",X"07",X"3C",X"47",X"3E",X"08",X"90",X"87",X"4F",
		X"CD",X"30",X"13",X"69",X"26",X"00",X"CD",X"90",X"0F",X"10",X"F5",X"C9",X"06",X"04",X"C5",X"06",
		X"04",X"FD",X"7E",X"00",X"77",X"CD",X"D0",X"32",X"00",X"00",X"23",X"FD",X"23",X"10",X"F2",X"11",
		X"DC",X"FF",X"19",X"C1",X"10",X"E8",X"C9",X"C6",X"91",X"6B",X"91",X"D0",X"91",X"90",X"92",X"EB",
		X"92",X"86",X"92",X"66",X"6A",X"6A",X"68",X"6E",X"00",X"00",X"71",X"6E",X"00",X"00",X"71",X"67",
		X"6D",X"6D",X"69",X"69",X"6D",X"6D",X"6D",X"00",X"00",X"00",X"00",X"6E",X"00",X"62",X"68",X"63",
		X"65",X"00",X"71",X"6E",X"71",X"00",X"71",X"63",X"65",X"63",X"65",X"6A",X"68",X"00",X"00",X"6D",
		X"69",X"6D",X"6D",X"66",X"6A",X"6E",X"71",X"6E",X"00",X"63",X"65",X"62",X"6A",X"66",X"64",X"63",
		X"00",X"63",X"65",X"21",X"00",X"00",X"22",X"F2",X"67",X"01",X"1A",X"1F",X"11",X"00",X"00",X"21",
		X"81",X"93",X"CD",X"FF",X"0B",X"CD",X"68",X"2C",X"3E",X"66",X"32",X"81",X"93",X"32",X"43",X"93",
		X"3C",X"32",X"61",X"90",X"32",X"A3",X"90",X"3C",X"32",X"5D",X"93",X"32",X"9F",X"93",X"3C",X"32",
		X"BD",X"90",X"32",X"7F",X"90",X"11",X"20",X"2F",X"01",X"02",X"02",X"21",X"23",X"92",X"CD",X"E0",
		X"0B",X"11",X"18",X"2E",X"01",X"1A",X"18",X"21",X"A5",X"92",X"CD",X"E0",X"0B",X"21",X"A5",X"92",
		X"06",X"0C",X"C5",X"06",X"18",X"7E",X"FE",X"02",X"20",X"03",X"AF",X"18",X"06",X"FE",X"72",X"20",
		X"07",X"3E",X"1B",X"CB",X"D4",X"77",X"CB",X"94",X"23",X"10",X"EA",X"11",X"C8",X"FF",X"19",X"C1",
		X"10",X"E0",X"11",X"2A",X"2F",X"21",X"24",X"93",X"01",X"03",X"04",X"C5",X"CD",X"E0",X"0B",X"C1",
		X"11",X"46",X"2F",X"21",X"84",X"91",X"CD",X"E0",X"0B",X"AF",X"32",X"EC",X"60",X"3E",X"01",X"32",
		X"CF",X"60",X"21",X"B8",X"0B",X"22",X"C0",X"60",X"21",X"63",X"2B",X"22",X"CB",X"60",X"22",X"D0",
		X"60",X"3E",X"04",X"32",X"D8",X"60",X"32",X"D9",X"60",X"32",X"DA",X"60",X"21",X"28",X"12",X"22",
		X"C5",X"60",X"22",X"DC",X"60",X"21",X"E5",X"12",X"22",X"C7",X"60",X"22",X"DE",X"60",X"21",X"86",
		X"F8",X"22",X"C9",X"60",X"22",X"E0",X"60",X"3E",X"02",X"32",X"FB",X"67",X"21",X"B8",X"0B",X"DD",
		X"21",X"0E",X"60",X"CD",X"C8",X"10",X"DD",X"21",X"11",X"60",X"CD",X"38",X"10",X"CD",X"83",X"0E",
		X"CD",X"8E",X"2C",X"2A",X"CB",X"60",X"11",X"83",X"D3",X"CD",X"03",X"10",X"28",X"33",X"CD",X"28",
		X"0D",X"C6",X"14",X"4F",X"3A",X"CF",X"60",X"CB",X"47",X"28",X"0F",X"CB",X"87",X"C6",X"0C",X"21",
		X"CB",X"60",X"CB",X"4E",X"28",X"02",X"C6",X"04",X"81",X"4F",X"79",X"21",X"5F",X"66",X"AE",X"32",
		X"FA",X"67",X"3A",X"0F",X"60",X"B7",X"28",X"09",X"3A",X"EC",X"60",X"CB",X"4F",X"28",X"C1",X"18",
		X"F1",X"21",X"14",X"00",X"CD",X"90",X"0F",X"21",X"00",X"00",X"E5",X"DD",X"E1",X"01",X"7B",X"1E",
		X"DD",X"5E",X"00",X"DD",X"56",X"01",X"19",X"DD",X"23",X"0B",X"78",X"B1",X"20",X"F2",X"3A",X"04",
		X"30",X"01",X"00",X"08",X"3A",X"01",X"30",X"E6",X"C0",X"A9",X"07",X"4F",X"10",X"F6",X"85",X"6F",
		X"11",X"15",X"0B",X"19",X"11",X"A9",X"2B",X"D5",X"E9",X"CD",X"D6",X"2F",X"06",X"18",X"21",X"A5",
		X"92",X"E5",X"21",X"05",X"00",X"CD",X"90",X"0F",X"E1",X"E5",X"0E",X"00",X"7E",X"FE",X"66",X"28",
		X"2A",X"FE",X"68",X"28",X"26",X"FE",X"6A",X"28",X"22",X"FE",X"67",X"28",X"22",X"FE",X"69",X"28",
		X"1E",X"FE",X"6D",X"28",X"1A",X"79",X"B7",X"28",X"08",X"36",X"00",X"CB",X"D4",X"36",X"00",X"CB",
		X"94",X"FE",X"02",X"28",X"12",X"11",X"E0",X"FF",X"19",X"18",X"D1",X"0E",X"01",X"18",X"E6",X"79",
		X"B7",X"28",X"F2",X"0E",X"02",X"18",X"DE",X"E1",X"23",X"10",X"B6",X"DD",X"21",X"06",X"92",X"FD",
		X"21",X"06",X"46",X"DD",X"36",X"00",X"5C",X"DD",X"36",X"01",X"5F",X"DD",X"36",X"E0",X"5D",X"DD",
		X"36",X"E1",X"5E",X"FD",X"36",X"00",X"02",X"FD",X"36",X"01",X"02",X"FD",X"36",X"E0",X"02",X"FD",
		X"36",X"E1",X"02",X"DD",X"21",X"0E",X"60",X"3A",X"0F",X"60",X"32",X"0E",X"60",X"AF",X"32",X"0F",
		X"60",X"CD",X"EC",X"10",X"45",X"78",X"B7",X"28",X"19",X"FD",X"21",X"11",X"60",X"DD",X"21",X"0E",
		X"60",X"CD",X"96",X"10",X"CD",X"C2",X"26",X"CD",X"6A",X"13",X"21",X"0D",X"00",X"CD",X"90",X"0F",
		X"10",X"E7",X"CD",X"F2",X"0E",X"21",X"2C",X"01",X"CD",X"90",X"0F",X"C3",X"1B",X"0F",X"77",X"CB",
		X"D4",X"71",X"CB",X"94",X"19",X"10",X"F7",X"C9",X"06",X"08",X"DD",X"21",X"E8",X"2D",X"16",X"00",
		X"C5",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"46",X"02",X"DD",X"4E",X"03",X"DD",X"7E",X"04",
		X"DD",X"5E",X"05",X"CD",X"5E",X"2C",X"C1",X"1E",X"06",X"DD",X"19",X"10",X"E3",X"C9",X"2A",X"C0",
		X"60",X"2B",X"7C",X"B5",X"20",X"FB",X"06",X"04",X"DD",X"21",X"C6",X"2F",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"C5",X"E7",X"C1",X"28",X"07",X"DD",X"23",X"DD",X"23",X"10",X"EF",X"C9",X"78",X"3D",
		X"F5",X"2A",X"D0",X"60",X"ED",X"5B",X"CB",X"60",X"CD",X"04",X"10",X"20",X"34",X"CD",X"B7",X"2D",
		X"79",X"87",X"DD",X"21",X"86",X"2F",X"87",X"5F",X"16",X"00",X"DD",X"19",X"F1",X"F5",X"5F",X"DD",
		X"19",X"DD",X"7E",X"00",X"FE",X"FF",X"28",X"75",X"DD",X"21",X"66",X"2F",X"87",X"5F",X"16",X"00",
		X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"22",X"D0",X"60",X"F1",X"32",X"CF",X"60",X"18",
		X"40",X"3A",X"CF",X"60",X"47",X"F1",X"B8",X"28",X"38",X"F5",X"4F",X"CD",X"D0",X"2D",X"C1",X"20",
		X"30",X"C5",X"2A",X"D0",X"60",X"CD",X"B7",X"2D",X"79",X"87",X"87",X"5F",X"16",X"00",X"DD",X"21",
		X"86",X"2F",X"F1",X"32",X"CF",X"60",X"83",X"5F",X"DD",X"19",X"DD",X"7E",X"00",X"DD",X"21",X"66",
		X"2F",X"87",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"22",X"D0",X"60",
		X"C9",X"3A",X"CF",X"60",X"DD",X"21",X"CE",X"2F",X"87",X"5F",X"16",X"00",X"DD",X"19",X"2A",X"CB",
		X"60",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"19",X"22",X"CB",X"60",X"18",X"02",X"F1",X"C9",X"06",
		X"08",X"3E",X"D3",X"BC",X"28",X"05",X"D6",X"18",X"10",X"F9",X"C9",X"48",X"7D",X"CB",X"41",X"28",
		X"02",X"C6",X"0C",X"06",X"0A",X"6F",X"3E",X"B8",X"BD",X"28",X"05",X"D6",X"08",X"10",X"F9",X"C9",
		X"05",X"68",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"11",X"86",X"91",X"19",X"3E",X"09",X"91",
		X"3D",X"28",X"05",X"2C",X"2C",X"2C",X"18",X"F8",X"7E",X"FE",X"72",X"C0",X"36",X"00",X"3A",X"0F",
		X"60",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",X"5F",X"AF",X"41",X"83",X"10",X"FD",
		X"F5",X"CD",X"7F",X"14",X"DD",X"21",X"11",X"60",X"CD",X"EC",X"10",X"F1",X"5F",X"16",X"00",X"19",
		X"DD",X"21",X"11",X"60",X"C3",X"C8",X"10",X"01",X"00",X"10",X"DD",X"21",X"66",X"2F",X"DD",X"5E",
		X"00",X"DD",X"56",X"01",X"CD",X"03",X"10",X"C8",X"0C",X"DD",X"23",X"DD",X"23",X"10",X"EF",X"C9",
		X"D5",X"DD",X"E5",X"59",X"16",X"00",X"DD",X"21",X"E4",X"2D",X"DD",X"19",X"DD",X"7E",X"00",X"B8",
		X"DD",X"E1",X"D1",X"C9",X"02",X"03",X"00",X"01",X"61",X"40",X"1A",X"02",X"6E",X"20",X"A3",X"40",
		X"16",X"02",X"6E",X"20",X"BD",X"40",X"16",X"02",X"71",X"20",X"7F",X"40",X"1A",X"02",X"71",X"20",
		X"62",X"40",X"1D",X"02",X"6D",X"01",X"A4",X"40",X"19",X"02",X"6D",X"01",X"44",X"43",X"19",X"02",
		X"6A",X"01",X"82",X"43",X"1D",X"02",X"6A",X"01",X"02",X"02",X"02",X"66",X"6E",X"6E",X"6E",X"67",
		X"24",X"02",X"02",X"02",X"6A",X"00",X"00",X"72",X"6D",X"24",X"02",X"02",X"02",X"6A",X"00",X"00",
		X"00",X"6D",X"24",X"02",X"02",X"02",X"6A",X"00",X"00",X"6E",X"6E",X"67",X"24",X"02",X"02",X"02",
		X"6A",X"72",X"72",X"00",X"00",X"6D",X"24",X"02",X"02",X"02",X"6A",X"00",X"00",X"00",X"00",X"6D",
		X"24",X"02",X"02",X"66",X"6E",X"6E",X"6E",X"00",X"00",X"6D",X"24",X"02",X"02",X"6A",X"00",X"00",
		X"72",X"72",X"72",X"6D",X"24",X"02",X"02",X"6A",X"00",X"00",X"00",X"00",X"00",X"6D",X"24",X"02",
		X"02",X"6A",X"00",X"00",X"6E",X"6E",X"6E",X"6E",X"67",X"24",X"02",X"02",X"6A",X"72",X"72",X"72",
		X"72",X"00",X"00",X"6D",X"24",X"02",X"02",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"24",
		X"02",X"66",X"6E",X"6E",X"6E",X"6E",X"6E",X"00",X"00",X"6D",X"24",X"02",X"6A",X"00",X"00",X"72",
		X"72",X"72",X"72",X"72",X"6D",X"24",X"02",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",
		X"24",X"02",X"6A",X"00",X"00",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"67",X"24",X"02",X"6A",X"72",
		X"72",X"72",X"72",X"72",X"72",X"00",X"00",X"6D",X"24",X"02",X"6A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6D",X"24",X"66",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"00",X"00",X"6D",
		X"24",X"6A",X"00",X"00",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"6D",X"24",X"6A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"24",X"6A",X"00",X"00",X"6E",X"6E",X"6E",X"6E",
		X"6E",X"6E",X"6E",X"6E",X"67",X"24",X"6A",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"00",
		X"00",X"6D",X"24",X"68",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"69",X"24",
		X"66",X"00",X"00",X"67",X"24",X"64",X"71",X"71",X"65",X"24",X"62",X"6E",X"6E",X"6E",X"6E",X"63",
		X"24",X"6A",X"54",X"49",X"4D",X"45",X"6D",X"24",X"6A",X"20",X"20",X"20",X"20",X"6D",X"24",X"64",
		X"71",X"71",X"71",X"71",X"65",X"24",X"62",X"6E",X"6E",X"6E",X"6E",X"6E",X"63",X"24",X"6A",X"42",
		X"4F",X"4E",X"55",X"53",X"6D",X"24",X"6A",X"20",X"20",X"20",X"20",X"20",X"6D",X"24",X"64",X"71",
		X"71",X"71",X"71",X"71",X"65",X"24",X"63",X"2B",X"AB",X"2B",X"AB",X"43",X"6B",X"43",X"6B",X"5B",
		X"A3",X"5B",X"A3",X"73",X"73",X"73",X"73",X"8B",X"9B",X"8B",X"9B",X"A3",X"7B",X"A3",X"7B",X"BB",
		X"93",X"BB",X"93",X"D3",X"83",X"D3",X"FF",X"FF",X"FF",X"01",X"02",X"00",X"FF",X"FF",X"FF",X"03",
		X"01",X"FF",X"04",X"FF",X"FF",X"02",X"FF",X"FF",X"03",X"05",X"06",X"04",X"FF",X"FF",X"FF",X"07",
		X"05",X"FF",X"08",X"FF",X"FF",X"06",X"FF",X"FF",X"07",X"09",X"0A",X"08",X"FF",X"FF",X"FF",X"0B",
		X"09",X"FF",X"0C",X"FF",X"FF",X"0A",X"FF",X"FF",X"0B",X"0D",X"0E",X"0C",X"FF",X"FF",X"FF",X"0F",
		X"0D",X"FF",X"FF",X"FF",X"FF",X"0E",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"00",X"00",X"01",
		X"FF",X"FF",X"00",X"FF",X"01",X"00",X"21",X"00",X"00",X"22",X"80",X"98",X"22",X"88",X"98",X"22",
		X"84",X"98",X"22",X"8C",X"98",X"22",X"90",X"98",X"C9",X"2B",X"AB",X"43",X"6B",X"43",X"6B",X"5B",
		X"A3",X"5B",X"A3",X"73",X"73",X"73",X"73",X"8B",X"9B",X"8B",X"9B",X"A3",X"7B",X"A3",X"7B",X"BB",
		X"06",X"08",X"21",X"00",X"60",X"AF",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",X"06",X"04",
		X"21",X"00",X"68",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",X"00",X"06",X"08",X"21",X"00",
		X"98",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",X"06",X"04",X"3E",X"20",X"21",X"00",X"90",
		X"0E",X"00",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F7",X"21",X"C0",X"60",X"06",X"40",X"3E",X"FF",
		X"77",X"23",X"10",X"FC",X"21",X"00",X"88",X"06",X"00",X"77",X"23",X"10",X"FC",X"31",X"C0",X"67",
		X"C3",X"1D",X"02",X"FF",X"FF",X"FF",X"5C",X"30",X"6D",X"00",X"D2",X"00",X"01",X"A0",X"03",X"21",
		X"00",X"60",X"36",X"00",X"23",X"0B",X"78",X"B1",X"20",X"F8",X"C3",X"9A",X"01",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D6",X"17",X"32",X"80",X"98",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"3A",X"5F",X"66",X"00",X"CB",X"47",X"28",X"03",X"C3",X"80",X"31",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"6B",X"2F",X"32",X"8A",X"98",X"3A",X"01",X"6B",X"2F",X"32",X"8B",X"98",X"3A",X"02",
		X"6B",X"2F",X"32",X"86",X"98",X"3A",X"03",X"6B",X"2F",X"32",X"87",X"98",X"3A",X"04",X"6B",X"2F",
		X"32",X"8E",X"98",X"3A",X"05",X"6B",X"2F",X"32",X"8F",X"98",X"3A",X"06",X"6B",X"2F",X"32",X"92",
		X"98",X"3A",X"07",X"6B",X"2F",X"32",X"93",X"98",X"3A",X"08",X"6B",X"2F",X"32",X"82",X"98",X"3A",
		X"09",X"6B",X"2F",X"32",X"83",X"98",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"00",X"6B",X"D6",X"10",X"32",X"8A",X"98",X"3A",X"01",X"6B",X"D6",X"10",X"32",X"8B",X"98",
		X"3A",X"02",X"6B",X"D6",X"10",X"32",X"86",X"98",X"3A",X"03",X"6B",X"D6",X"10",X"32",X"87",X"98",
		X"3A",X"04",X"6B",X"D6",X"10",X"32",X"8E",X"98",X"3A",X"05",X"6B",X"D6",X"10",X"32",X"8F",X"98",
		X"3A",X"06",X"6B",X"D6",X"10",X"32",X"92",X"98",X"3A",X"07",X"6B",X"D6",X"10",X"32",X"93",X"98",
		X"3A",X"08",X"6B",X"D6",X"10",X"32",X"82",X"98",X"3A",X"09",X"6B",X"D6",X"10",X"32",X"83",X"98",
		X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4F",X"87",X"87",X"F5",X"3E",X"B0",X"8C",X"67",X"F1",X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"AF",X"32",X"C5",X"60",X"32",X"C6",X"60",X"F1",X"21",X"06",X"00",X"C9",X"FF",X"FF",X"FF",
		X"F5",X"E5",X"DD",X"E5",X"E1",X"7D",X"FE",X"DC",X"20",X"03",X"01",X"A8",X"37",X"FE",X"DE",X"20",
		X"03",X"01",X"AE",X"37",X"FE",X"E0",X"20",X"03",X"01",X"B0",X"37",X"E1",X"F1",X"C9",X"FF",X"FF",
		X"F5",X"E5",X"FD",X"E5",X"E1",X"7D",X"FE",X"DC",X"20",X"03",X"11",X"A8",X"37",X"FE",X"DE",X"20",
		X"03",X"11",X"AE",X"37",X"FE",X"E0",X"20",X"03",X"11",X"B0",X"37",X"E1",X"F1",X"C9",X"FF",X"FF",
		X"F5",X"E5",X"00",X"00",X"00",X"7D",X"FE",X"DC",X"20",X"03",X"11",X"A8",X"37",X"FE",X"DE",X"20",
		X"03",X"11",X"AE",X"37",X"FE",X"E0",X"20",X"03",X"11",X"B0",X"37",X"E1",X"F1",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"3A",X"C5",X"60",X"2F",X"32",X"86",X"98",X"3A",X"C6",X"60",X"2F",X"32",X"87",X"98",X"3A",
		X"C7",X"60",X"2F",X"32",X"8E",X"98",X"3A",X"C8",X"60",X"2F",X"32",X"8F",X"98",X"3A",X"C9",X"60",
		X"2F",X"32",X"92",X"98",X"3A",X"CA",X"60",X"2F",X"32",X"93",X"98",X"F1",X"C9",X"FF",X"FF",X"FF",
		X"E5",X"F5",X"79",X"E6",X"0F",X"4F",X"00",X"3E",X"0C",X"84",X"67",X"71",X"F1",X"E1",X"C9",X"FF",
		X"C5",X"3A",X"BD",X"67",X"47",X"7E",X"3C",X"81",X"E6",X"0F",X"77",X"C1",X"C9",X"E5",X"F5",X"DD",
		X"E5",X"E1",X"3E",X"04",X"84",X"67",X"F1",X"E6",X"0F",X"77",X"E1",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"01",X"32",X"01",X"A0",X"AF",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"32",X"01",X"A0",X"3C",X"32",X"01",X"A0",X"3D",X"32",X"01",X"A0",X"3C",X"C9",X"FF",X"FF",
		X"6F",X"26",X"07",X"FD",X"7D",X"FE",X"F4",X"20",X"03",X"22",X"84",X"98",X"FE",X"F6",X"20",X"03",
		X"22",X"8C",X"98",X"FE",X"F8",X"20",X"03",X"22",X"90",X"98",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"3E",X"72",X"32",X"E6",X"69",X"32",X"09",X"6A",X"00",X"32",X"29",X"6A",X"32",X"CC",X"69",
		X"32",X"EC",X"69",X"32",X"0C",X"6A",X"32",X"EF",X"69",X"32",X"0F",X"6A",X"32",X"2F",X"6A",X"32",
		X"4F",X"6A",X"32",X"B2",X"69",X"32",X"D2",X"69",X"32",X"F2",X"69",X"32",X"12",X"6A",X"32",X"32",
		X"6A",X"32",X"D5",X"69",X"32",X"F5",X"69",X"32",X"15",X"6A",X"32",X"35",X"6A",X"32",X"55",X"6A",
		X"32",X"75",X"6A",X"32",X"98",X"69",X"32",X"B8",X"69",X"32",X"D8",X"69",X"32",X"F8",X"69",X"32",
		X"18",X"6A",X"32",X"38",X"6A",X"32",X"58",X"6A",X"32",X"BB",X"69",X"32",X"DB",X"69",X"32",X"FB",
		X"69",X"32",X"1B",X"6A",X"32",X"3B",X"6A",X"32",X"5B",X"6A",X"32",X"7B",X"6A",X"32",X"9B",X"6A",
		X"F1",X"00",X"21",X"A5",X"92",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E5",X"C5",X"3A",X"00",X"B8",X"32",X"00",X"60",X"21",X"00",X"60",X"CB",X"47",X"20",X"03",X"06",
		X"DF",X"70",X"CB",X"4F",X"20",X"03",X"06",X"BF",X"70",X"3A",X"00",X"B8",X"32",X"01",X"60",X"21",
		X"01",X"60",X"CB",X"57",X"20",X"03",X"06",X"DF",X"70",X"CB",X"5F",X"20",X"03",X"06",X"BF",X"70",
		X"3A",X"00",X"A8",X"2F",X"21",X"01",X"60",X"CB",X"7F",X"20",X"03",X"06",X"FB",X"70",X"CB",X"77",
		X"20",X"03",X"06",X"FD",X"70",X"CB",X"6F",X"20",X"03",X"06",X"F7",X"70",X"CB",X"67",X"20",X"03",
		X"06",X"FE",X"70",X"CB",X"5F",X"20",X"03",X"06",X"EF",X"70",X"FE",X"77",X"20",X"03",X"06",X"EB",
		X"70",X"FE",X"B7",X"20",X"03",X"06",X"ED",X"70",X"00",X"00",X"3A",X"00",X"A0",X"2F",X"21",X"00",
		X"60",X"CB",X"7F",X"20",X"03",X"06",X"FD",X"70",X"CB",X"77",X"20",X"03",X"06",X"FB",X"70",X"CB",
		X"6F",X"20",X"03",X"06",X"F7",X"70",X"CB",X"67",X"20",X"03",X"06",X"FE",X"70",X"CB",X"5F",X"20",
		X"03",X"06",X"7F",X"70",X"FE",X"77",X"20",X"03",X"06",X"7D",X"70",X"FE",X"B7",X"20",X"03",X"06",
		X"7B",X"70",X"C1",X"E1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E5",X"CB",X"BC",X"CB",X"A4",X"CB",X"EC",X"CB",X"F4",X"CB",X"DC",X"7E",X"FE",X"72",X"E1",X"C9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E5",X"CB",X"BC",X"CB",X"A4",X"CB",X"EC",X"CB",X"F4",X"CB",X"DC",X"36",X"00",X"E1",X"3A",X"0F",
		X"60",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DD",X"21",X"0B",X"60",X"F5",X"3E",X"00",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"D4",X"60",X"F5",X"3E",X"02",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2B",X"7D",X"0E",X"7F",X"F5",X"3E",X"04",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"7E",X"00",X"F5",X"3E",X"06",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"3E",X"0A",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D6",X"02",X"77",X"F5",X"3E",X"08",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"3E",X"0C",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"3E",X"0E",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"3E",X"10",X"CD",X"00",X"36",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"E5",X"D5",X"C5",X"00",X"00",X"00",X"21",X"00",X"37",X"6F",X"00",X"00",X"7E",X"32",X"00",
		X"A8",X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"C0",X"D3",X"09",X"3E",X"0E",X"D3",
		X"08",X"23",X"7E",X"D3",X"09",X"3E",X"0F",X"D3",X"08",X"3E",X"7F",X"D3",X"09",X"3E",X"07",X"32",
		X"00",X"B0",X"32",X"04",X"A0",X"AF",X"32",X"04",X"A0",X"C5",X"01",X"80",X"02",X"0D",X"20",X"FD",
		X"10",X"FB",X"C1",X"3E",X"FF",X"32",X"04",X"A0",X"C1",X"D1",X"E1",X"F1",X"C9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"79",X"28",X"70",X"C0",X"20",X"97",X"04",X"A4",X"70",X"C0",X"20",X"C0",X"40",X"40",X"20",X"85",
		X"35",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
