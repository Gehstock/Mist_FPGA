library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity k_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of k_rom is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"1C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"4C",X"DE",X"92",X"92",X"92",X"F6",X"64",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"E0",X"70",X"17",X"17",X"70",X"E0",X"00",X"00",
		X"82",X"44",X"28",X"10",X"28",X"44",X"82",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"0B",X"0A",X"0F",X"00",X"00",X"00",X"03",X"05",X"05",X"05",X"87",X"00",X"00",X"00",X"81",X"02",
		X"82",X"02",X"C3",X"00",X"00",X"00",X"C0",X"81",X"C0",X"80",X"E0",X"00",X"00",X"00",X"E0",X"40",
		X"09",X"05",X"03",X"00",X"00",X"00",X"05",X"0A",X"04",X"02",X"81",X"00",X"00",X"00",X"02",X"85",
		X"82",X"81",X"C0",X"00",X"00",X"00",X"81",X"42",X"40",X"40",X"E0",X"00",X"00",X"00",X"40",X"A0",
		X"0A",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"85",X"87",X"00",X"00",X"00",X"00",X"00",X"00",
		X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"50",X"7C",X"00",X"00",X"00",X"1C",X"28",
		X"2C",X"28",X"3E",X"00",X"00",X"00",X"0E",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"28",X"1C",X"00",X"00",X"00",X"28",X"54",
		X"24",X"14",X"0E",X"00",X"00",X"00",X"14",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"07",X"00",X"00",X"00",X"01",X"02",
		X"80",X"00",X"C0",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"02",X"05",
		X"80",X"80",X"C0",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"0F",X"FE",X"FF",X"FF",X"F7",X"F7",X"F3",X"FB",X"F9",
		X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"F9",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"7F",X"3F",X"0F",X"01",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"03",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"03",X"0F",
		X"00",X"00",X"00",X"01",X"8E",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"0F",X"03",X"03",X"03",X"03",X"02",X"00",
		X"E0",X"F0",X"F8",X"FC",X"8E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"F8",X"E0",
		X"00",X"00",X"E0",X"FC",X"FF",X"FF",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"0F",X"0F",X"1F",X"1E",X"1E",X"3C",X"3C",X"3C",X"80",X"00",X"03",X"0F",X"1F",X"1F",X"3F",X"3F",
		X"01",X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"F0",X"F0",X"F8",X"78",X"78",X"3C",X"3C",X"3C",
		X"3C",X"3C",X"3C",X"1E",X"1E",X"1F",X"0F",X"0F",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"00",X"80",
		X"FC",X"FC",X"F8",X"F8",X"F0",X"C0",X"00",X"01",X"3C",X"3C",X"3C",X"78",X"78",X"F8",X"F0",X"F0",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FF",X"FF",X"3F",X"07",X"00",X"00",
		X"07",X"1F",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",
		X"00",X"00",X"1B",X"1F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"07",X"1F",X"27",X"27",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"FC",
		X"27",X"27",X"1F",X"07",X"07",X"03",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"E7",X"7B",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FC",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"00",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"40",X"40",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"40",X"40",X"40",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"07",X"3F",X"FC",X"FB",X"FB",X"FC",
		X"00",X"00",X"E0",X"FC",X"3F",X"DF",X"DF",X"3E",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"B0",X"98",X"D8",X"D8",X"CC",X"CC",X"CC",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"CC",X"D8",X"D8",X"98",X"B0",X"70",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0B",X"1D",X"1F",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"D8",
		X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"00",X"D0",X"BC",X"FE",X"F6",X"FB",X"FB",X"FB",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"EC",X"EC",X"EC",X"EC",X"D8",X"F8",X"F0",X"C0",
		X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"FB",X"F6",X"FE",X"FC",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"04",X"08",X"08",X"08",X"08",X"04",X"03",X"C0",X"20",X"10",X"10",X"10",X"10",X"20",X"C0",
		X"01",X"01",X"01",X"01",X"FF",X"FF",X"01",X"01",X"80",X"80",X"80",X"80",X"FF",X"FF",X"80",X"80",
		X"01",X"01",X"FF",X"FF",X"01",X"01",X"01",X"01",X"80",X"80",X"FF",X"FF",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3C",X"1E",X"0F",X"07",X"0F",X"1E",X"3C",X"FF",
		X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F8",
		X"F8",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"00",X"00",X"FF",
		X"FF",X"03",X"07",X"0F",X"1E",X"3C",X"78",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"06",X"03",X"03",X"06",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F8",X"F8",X"E0",
		X"E3",X"E3",X"E1",X"E1",X"E1",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",
		X"01",X"FF",X"FF",X"00",X"00",X"F8",X"F8",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"00",X"00",X"3F",
		X"3F",X"27",X"27",X"07",X"07",X"07",X"07",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"3F",X"27",X"27",X"07",X"07",X"07",X"07",X"FF",X"FF",X"00",X"00",X"FF",
		X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",
		X"FF",X"1C",X"38",X"F0",X"C0",X"C0",X"F0",X"38",X"1C",X"FF",X"FF",X"00",X"00",X"1F",X"1F",X"07",
		X"E7",X"E7",X"C7",X"C7",X"C7",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"FF",X"FF",X"00",X"00",X"1F",X"1F",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
