library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"91",X"8D",X"92",X"8A",X"92",X"8D",X"92",X"8A",X"92",X"8D",X"91",X"88",X"91",X"8D",X"91",
		X"88",X"91",X"8F",X"94",X"FF",X"E7",X"AF",X"32",X"C8",X"42",X"3E",X"19",X"32",X"A3",X"42",X"F7",
		X"C3",X"61",X"09",X"E7",X"F7",X"C9",X"DD",X"21",X"80",X"42",X"C3",X"A1",X"07",X"DD",X"21",X"88",
		X"42",X"C3",X"A1",X"07",X"1F",X"0B",X"3F",X"0C",X"5F",X"05",X"B4",X"91",X"8D",X"B9",X"98",X"96",
		X"B4",X"99",X"91",X"8F",X"B4",X"80",X"80",X"94",X"94",X"94",X"94",X"91",X"8F",X"8D",X"80",X"99",
		X"99",X"99",X"9B",X"99",X"98",X"96",X"94",X"91",X"80",X"91",X"B9",X"B1",X"94",X"CF",X"80",X"A0",
		X"80",X"91",X"91",X"92",X"94",X"96",X"98",X"D6",X"C0",X"80",X"92",X"92",X"94",X"B6",X"98",X"99",
		X"D8",X"A0",X"B4",X"D9",X"99",X"98",X"96",X"94",X"D8",X"B6",X"B6",X"B4",X"BB",X"B9",X"B8",X"D9",
		X"C0",X"99",X"99",X"99",X"99",X"99",X"99",X"98",X"96",X"D9",X"B4",X"91",X"91",X"AF",X"8F",X"8F",
		X"99",X"99",X"98",X"96",X"D6",X"D4",X"94",X"91",X"91",X"91",X"B1",X"8F",X"8D",X"92",X"91",X"92",
		X"94",X"B6",X"A0",X"94",X"92",X"8F",X"8F",X"AF",X"8D",X"8C",X"8D",X"8C",X"8D",X"8F",X"D1",X"94",
		X"91",X"91",X"91",X"B1",X"8F",X"8D",X"92",X"91",X"92",X"94",X"B6",X"98",X"96",X"B4",X"94",X"96",
		X"94",X"92",X"91",X"8F",X"CA",X"AC",X"AF",X"CD",X"C0",X"FF",X"1F",X"05",X"5F",X"05",X"D9",X"D6",
		X"D9",X"D8",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",X"8D",X"92",X"8A",X"92",X"8D",X"92",
		X"8A",X"92",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",X"8F",X"94",X"88",X"94",X"8A",X"94",
		X"8C",X"94",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",X"8D",X"92",X"8A",X"92",X"8D",X"92",
		X"8A",X"92",X"8D",X"92",X"8A",X"92",X"8D",X"92",X"8A",X"92",X"8F",X"94",X"88",X"94",X"8F",X"94",
		X"88",X"94",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",X"8D",X"91",X"89",X"91",X"8A",X"92",
		X"8F",X"92",X"8F",X"94",X"88",X"94",X"8F",X"94",X"88",X"94",X"8D",X"91",X"88",X"91",X"AD",X"A0",
		X"D2",X"C0",X"D1",X"C0",X"DF",X"C0",X"D2",X"D2",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",
		X"8D",X"92",X"8A",X"92",X"8D",X"92",X"8A",X"92",X"8F",X"94",X"88",X"94",X"8F",X"94",X"88",X"94",
		X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",X"8D",X"91",X"88",X"91",
		X"8D",X"92",X"8A",X"92",X"8D",X"92",X"8A",X"92",X"8F",X"94",X"88",X"94",X"8F",X"94",X"88",X"94",
		X"D2",X"D4",X"8D",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"8F",X"60",X"6F",X"8F",X"60",X"6F",
		X"91",X"60",X"71",X"93",X"60",X"73",X"74",X"74",X"74",X"60",X"94",X"60",X"76",X"D8",X"B9",X"B9",
		X"98",X"60",X"B9",X"60",X"8F",X"60",X"6F",X"91",X"60",X"D2",X"60",X"94",X"60",X"76",X"94",X"60",
		X"72",X"91",X"60",X"71",X"92",X"60",X"D4",X"60",X"A0",X"74",X"76",X"78",X"60",X"B9",X"B9",X"98",
		X"60",X"B9",X"60",X"8F",X"60",X"6F",X"91",X"60",X"72",X"80",X"60",X"76",X"94",X"60",X"73",X"94",
		X"80",X"B2",X"B1",X"8F",X"60",X"CD",X"FF",X"1F",X"05",X"5F",X"06",X"B9",X"B9",X"B9",X"B9",X"B8",
		X"B2",X"B1",X"AF",X"AD",X"B4",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B8",X"B8",X"B8",X"B8",X"B4",
		X"B1",X"BD",X"B4",X"B4",X"B4",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"98",X"80",X"A0",X"B6",X"B4",
		X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"92",X"97",X"97",X"99",X"9B",X"97",X"9B",X"99",X"92",
		X"97",X"97",X"99",X"9B",X"B7",X"96",X"92",X"97",X"97",X"99",X"9B",X"9C",X"9B",X"99",X"97",X"96",
		X"92",X"94",X"96",X"B7",X"97",X"80",X"FF",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"94",X"60",
		X"76",X"94",X"92",X"94",X"96",X"B7",X"92",X"60",X"74",X"92",X"90",X"8F",X"90",X"92",X"80",X"94",
		X"60",X"76",X"94",X"92",X"94",X"96",X"97",X"94",X"94",X"97",X"96",X"99",X"B7",X"97",X"80",X"FF",
		X"1F",X"0B",X"5F",X"06",X"90",X"60",X"70",X"90",X"92",X"90",X"90",X"B0",X"8F",X"60",X"70",X"8F",
		X"8D",X"8B",X"8B",X"8B",X"80",X"90",X"60",X"70",X"90",X"92",X"90",X"90",X"90",X"90",X"8F",X"92",
		X"92",X"90",X"AF",X"8F",X"80",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"72",X"74",X"B6",X"96",
		X"B6",X"96",X"B7",X"96",X"B6",X"7B",X"7B",X"B9",X"96",X"96",X"94",X"92",X"B4",X"94",X"B4",X"80",
		X"B6",X"96",X"B6",X"96",X"B7",X"96",X"B6",X"9B",X"B9",X"96",X"94",X"96",X"94",X"B2",X"92",X"B2",
		X"80",X"FF",X"1F",X"0B",X"5F",X"06",X"72",X"74",X"B6",X"8D",X"8D",X"8F",X"8D",X"AF",X"92",X"B2",
		X"80",X"AD",X"8D",X"8F",X"91",X"92",X"B2",X"91",X"B1",X"72",X"74",X"B6",X"8D",X"8D",X"8F",X"8D",
		X"AF",X"92",X"B2",X"97",X"B6",X"92",X"91",X"92",X"9D",X"AA",X"8A",X"AA",X"80",X"FF",X"1F",X"0B",
		X"3F",X"0D",X"5F",X"06",X"8A",X"AF",X"8E",X"8C",X"AA",X"80",X"8A",X"AC",X"AE",X"AF",X"8A",X"8A",
		X"8C",X"8A",X"88",X"87",X"8C",X"8A",X"88",X"87",X"A5",X"AA",X"AA",X"80",X"FF",X"1F",X"0B",X"5F",
		X"06",X"8A",X"AF",X"8E",X"8C",X"AA",X"80",X"8A",X"A9",X"A8",X"A7",X"87",X"83",X"88",X"87",X"85",
		X"83",X"A3",X"A5",X"A1",X"80",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"8A",X"87",X"8A",X"8A",
		X"8A",X"8C",X"8A",X"8A",X"8A",X"87",X"8A",X"8A",X"8A",X"8C",X"8A",X"8A",X"8A",X"AF",X"B1",X"93",
		X"60",X"6F",X"8F",X"8F",X"B1",X"AE",X"AF",X"80",X"FF",X"1F",X"0B",X"5F",X"06",X"87",X"83",X"87",
		X"87",X"87",X"86",X"87",X"87",X"87",X"83",X"87",X"87",X"87",X"87",X"85",X"87",X"88",X"AA",X"AA",
		X"8A",X"60",X"67",X"87",X"8A",X"A8",X"A8",X"A7",X"80",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",
		X"8F",X"93",X"B6",X"B6",X"BB",X"9A",X"98",X"96",X"96",X"93",X"94",X"96",X"80",X"BA",X"98",X"98",
		X"94",X"98",X"96",X"96",X"9B",X"9B",X"9A",X"98",X"96",X"9A",X"9B",X"80",X"8F",X"93",X"B6",X"B6",
		X"BB",X"9A",X"98",X"96",X"96",X"93",X"94",X"96",X"80",X"BA",X"98",X"98",X"94",X"98",X"96",X"96",
		X"9B",X"9B",X"9A",X"98",X"96",X"9A",X"9B",X"80",X"A0",X"FF",X"1F",X"0B",X"5F",X"06",X"8F",X"8F",
		X"B3",X"B3",X"B8",X"96",X"94",X"93",X"93",X"8F",X"91",X"93",X"80",X"B6",X"94",X"94",X"8F",X"94",
		X"93",X"93",X"93",X"93",X"96",X"93",X"8F",X"91",X"93",X"80",X"8F",X"8F",X"B3",X"B3",X"B8",X"96",
		X"94",X"93",X"93",X"8F",X"91",X"93",X"80",X"B6",X"94",X"94",X"8F",X"94",X"93",X"93",X"93",X"93",
		X"96",X"93",X"8F",X"91",X"93",X"80",X"A0",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"8D",X"92",
		X"96",X"B9",X"99",X"96",X"B7",X"97",X"94",X"B6",X"B9",X"80",X"96",X"97",X"99",X"BB",X"9B",X"9B",
		X"9B",X"99",X"9B",X"9C",X"DD",X"A0",X"9D",X"9D",X"BD",X"9B",X"99",X"BB",X"99",X"97",X"9B",X"80",
		X"B9",X"A0",X"96",X"97",X"B9",X"98",X"99",X"BB",X"99",X"97",X"D6",X"FF",X"1F",X"0B",X"5F",X"06",
		X"8D",X"92",X"96",X"B6",X"96",X"92",X"B4",X"94",X"91",X"B2",X"B6",X"80",X"92",X"94",X"96",X"B7",
		X"97",X"97",X"97",X"96",X"97",X"98",X"D9",X"A0",X"99",X"99",X"B9",X"97",X"96",X"B7",X"96",X"94",
		X"97",X"80",X"B6",X"A0",X"92",X"94",X"B6",X"95",X"96",X"B7",X"96",X"94",X"D2",X"FF",X"1F",X"0B",
		X"3F",X"0D",X"5F",X"06",X"8C",X"B1",X"91",X"94",X"B8",X"80",X"8C",X"90",X"90",X"90",X"93",X"B6",
		X"A0",X"B6",X"98",X"96",X"94",X"94",X"93",X"91",X"93",X"93",X"94",X"96",X"B8",X"A0",X"96",X"76",
		X"74",X"96",X"76",X"74",X"AC",X"B0",X"D1",X"FF",X"1F",X"05",X"5F",X"06",X"80",X"B1",X"B1",X"B1",
		X"B1",X"AC",X"AC",X"AC",X"AC",X"AA",X"AA",X"AA",X"AA",X"AC",X"AC",X"AC",X"AC",X"8A",X"80",X"8A",
		X"80",X"AC",X"AC",X"B1",X"FF",X"E7",X"3E",X"01",X"32",X"C8",X"42",X"32",X"C3",X"42",X"F7",X"C3",
		X"70",X"16",X"DD",X"21",X"B0",X"42",X"DD",X"7E",X"00",X"FE",X"FF",X"28",X"25",X"CD",X"A9",X"14",
		X"AF",X"C9",X"E7",X"3E",X"00",X"32",X"C3",X"42",X"F7",X"C3",X"6B",X"16",X"3A",X"C8",X"42",X"A7",
		X"20",X"14",X"E7",X"DD",X"21",X"B0",X"42",X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"CD",X"A9",X"14",
		X"AF",X"C9",X"AF",X"32",X"C8",X"42",X"3E",X"FF",X"C9",X"DD",X"35",X"01",X"C0",X"3A",X"C2",X"42",
		X"DD",X"77",X"01",X"DD",X"7E",X"08",X"A7",X"28",X"16",X"21",X"C4",X"42",X"35",X"7E",X"A7",X"28",
		X"0B",X"CD",X"4D",X"02",X"ED",X"5B",X"C5",X"42",X"19",X"EF",X"18",X"03",X"DD",X"77",X"08",X"DD",
		X"CB",X"00",X"46",X"C2",X"E3",X"14",X"DD",X"7E",X"07",X"D6",X"01",X"FA",X"E3",X"14",X"DD",X"77",
		X"07",X"47",X"DF",X"DD",X"35",X"00",X"C0",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"47",X"E6",
		X"1F",X"CA",X"94",X"15",X"FE",X"1F",X"C2",X"AE",X"15",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",X"06",X"00",X"21",X"16",X"15",X"09",X"5E",X"23",
		X"56",X"2A",X"B2",X"42",X"D5",X"C9",X"26",X"15",X"39",X"15",X"49",X"15",X"52",X"15",X"8C",X"15",
		X"8C",X"15",X"8C",X"15",X"8C",X"15",X"4E",X"CB",X"21",X"CB",X"21",X"06",X"00",X"21",X"E3",X"15",
		X"09",X"DD",X"75",X"04",X"DD",X"74",X"05",X"18",X"43",X"4E",X"06",X"00",X"21",X"5B",X"16",X"09",
		X"7E",X"32",X"C2",X"42",X"DD",X"77",X"01",X"18",X"33",X"7E",X"DD",X"77",X"06",X"DD",X"77",X"07",
		X"18",X"2A",X"7E",X"DD",X"77",X"08",X"DD",X"77",X"09",X"A7",X"28",X"20",X"47",X"E6",X"E0",X"07",
		X"07",X"07",X"32",X"C4",X"42",X"78",X"16",X"00",X"21",X"00",X"00",X"E6",X"0F",X"87",X"5F",X"78",
		X"E6",X"10",X"20",X"04",X"ED",X"52",X"18",X"01",X"19",X"22",X"C5",X"42",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",X"E7",X"14",X"06",X"00",X"DF",X"DD",
		X"36",X"00",X"FF",X"C9",X"CD",X"9C",X"15",X"06",X"00",X"DF",X"18",X"39",X"78",X"E6",X"E0",X"07",
		X"07",X"07",X"47",X"3E",X"01",X"10",X"04",X"DD",X"77",X"00",X"C9",X"07",X"18",X"F7",X"C5",X"CD",
		X"9C",X"15",X"C1",X"78",X"E6",X"1F",X"3D",X"07",X"4F",X"06",X"00",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"09",X"5E",X"23",X"56",X"EB",X"EF",X"DD",X"7E",X"09",X"DD",X"77",X"08",X"DD",X"46",X"06",
		X"78",X"DD",X"77",X"07",X"DF",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",
		X"74",X"03",X"C9",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",X"06",X"F3",
		X"05",X"9E",X"05",X"4E",X"05",X"01",X"05",X"B9",X"04",X"76",X"04",X"36",X"04",X"F9",X"03",X"C0",
		X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",
		X"02",X"3B",X"02",X"1B",X"02",X"FD",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",X"01",X"7D",
		X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",
		X"00",X"E3",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",
		X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",
		X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"11",X"0F",X"0D",X"0B",X"0A",
		X"09",X"08",X"07",X"03",X"05",X"14",X"13",X"11",X"10",X"0F",X"0E",X"3A",X"C8",X"42",X"A7",X"C0",
		X"21",X"94",X"16",X"11",X"B0",X"42",X"01",X"0A",X"00",X"ED",X"B0",X"3A",X"C3",X"42",X"87",X"4F",
		X"87",X"81",X"4F",X"21",X"9E",X"16",X"09",X"11",X"B2",X"42",X"7E",X"12",X"CD",X"91",X"16",X"7E",
		X"12",X"23",X"13",X"C9",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"16",
		X"CD",X"16",X"CD",X"16",X"B8",X"16",X"CD",X"16",X"CD",X"16",X"1F",X"0F",X"3F",X"09",X"5F",X"09",
		X"7F",X"00",X"6D",X"71",X"74",X"79",X"D6",X"FF",X"1F",X"02",X"3F",X"07",X"5F",X"09",X"7F",X"00",
		X"94",X"8D",X"88",X"94",X"8D",X"88",X"94",X"8D",X"88",X"94",X"8D",X"C8",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
