library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity burnin_rubber_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of burnin_rubber_prog is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"2C",X"FF",X"C0",X"28",X"8A",X"28",X"98",X"28",X"B8",X"C5",X"02",X"F0",X"46",X"CD",X"01",X"10",
		X"29",X"FF",X"49",X"E0",X"85",X"03",X"2A",X"2A",X"2A",X"2A",X"2A",X"85",X"01",X"40",X"E4",X"C0",
		X"CD",X"04",X"10",X"29",X"FF",X"49",X"C0",X"F0",X"2A",X"85",X"04",X"40",X"E4",X"C0",X"CD",X"04",
		X"10",X"29",X"FF",X"45",X"04",X"F0",X"1C",X"40",X"E4",X"C0",X"CD",X"04",X"10",X"29",X"FF",X"45",
		X"04",X"F0",X"10",X"40",X"E4",X"C0",X"CD",X"04",X"10",X"29",X"FF",X"45",X"04",X"F0",X"04",X"C9",
		X"FF",X"85",X"00",X"8D",X"00",X"10",X"68",X"C8",X"68",X"CA",X"68",X"20",X"28",X"8A",X"28",X"98",
		X"28",X"C5",X"00",X"F0",X"40",X"CD",X"04",X"10",X"49",X"C0",X"45",X"04",X"F0",X"37",X"E6",X"06",
		X"C9",X"02",X"8D",X"02",X"10",X"C4",X"01",X"C5",X"03",X"A9",X"80",X"F0",X"2E",X"C2",X"00",X"CD",
		X"00",X"10",X"29",X"FF",X"49",X"0F",X"06",X"04",X"90",X"02",X"2A",X"2A",X"49",X"03",X"F0",X"3D",
		X"E8",X"A9",X"01",X"F0",X"38",X"E8",X"A9",X"02",X"F0",X"2B",X"E8",X"C5",X"06",X"A9",X"02",X"D0",
		X"1F",X"C9",X"00",X"85",X"00",X"68",X"C8",X"68",X"CA",X"68",X"60",X"C2",X"05",X"C5",X"04",X"A9",
		X"40",X"F0",X"1A",X"E8",X"A9",X"80",X"F0",X"15",X"E8",X"A9",X"C0",X"F0",X"DE",X"2C",X"A1",X"C0",
		X"A6",X"06",X"2C",X"CD",X"C0",X"C5",X"03",X"A9",X"60",X"B0",X"02",X"C2",X"04",X"C5",X"05",X"F8",
		X"18",X"7D",X"EF",X"C0",X"B9",X"F7",X"C0",X"90",X"03",X"D9",X"F7",X"C0",X"85",X"05",X"B8",X"A6",
		X"06",X"2C",X"A1",X"C0",X"C2",X"E7",X"C5",X"FF",X"C5",X"FF",X"EA",X"AA",X"B0",X"F8",X"60",X"01",
		X"02",X"03",X"01",X"06",X"08",X"03",X"01",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"78",
		X"B8",X"C2",X"FF",X"9A",X"C9",X"00",X"85",X"02",X"8D",X"01",X"10",X"8D",X"00",X"54",X"8D",X"00",
		X"58",X"8D",X"02",X"10",X"8D",X"00",X"10",X"38",X"40",X"AF",X"C2",X"40",X"BA",X"C2",X"40",X"CE",
		X"C2",X"40",X"11",X"C3",X"40",X"DE",X"C2",X"40",X"FE",X"E6",X"C9",X"FF",X"85",X"02",X"40",X"E5",
		X"E1",X"40",X"BA",X"C2",X"40",X"AB",X"D4",X"40",X"77",X"DC",X"40",X"DE",X"C2",X"C2",X"18",X"40",
		X"B2",X"C2",X"C2",X"00",X"40",X"C3",X"C2",X"40",X"5B",X"DB",X"AE",X"02",X"04",X"AE",X"22",X"04",
		X"C9",X"00",X"85",X"09",X"C5",X"08",X"85",X"12",X"40",X"07",X"D9",X"C5",X"12",X"A9",X"02",X"90",
		X"03",X"40",X"1D",X"D9",X"C2",X"31",X"C9",X"00",X"40",X"B2",X"C2",X"40",X"C3",X"C2",X"C9",X"00",
		X"8D",X"00",X"54",X"C5",X"09",X"8D",X"01",X"10",X"40",X"B7",X"DC",X"40",X"11",X"C3",X"40",X"B1",
		X"D3",X"40",X"16",X"DA",X"40",X"33",X"D5",X"40",X"F0",X"D5",X"C5",X"07",X"B0",X"42",X"40",X"8F",
		X"EB",X"2C",X"2E",X"C1",X"C5",X"05",X"F0",X"37",X"C9",X"00",X"85",X"08",X"85",X"12",X"CD",X"04",
		X"10",X"29",X"FF",X"49",X"18",X"F0",X"28",X"A9",X"08",X"F0",X"12",X"A9",X"10",X"B0",X"20",X"C5",
		X"05",X"A9",X"02",X"90",X"1A",X"E6",X"08",X"40",X"7F",X"EA",X"40",X"FB",X"DB",X"E6",X"08",X"40",
		X"75",X"EA",X"40",X"FB",X"DB",X"C9",X"01",X"85",X"07",X"C2",X"FF",X"9A",X"2C",X"31",X"C1",X"60",
		X"40",X"82",X"C2",X"40",X"F5",X"D8",X"40",X"33",X"C3",X"40",X"1B",X"C8",X"40",X"D2",X"D2",X"40",
		X"D0",X"C6",X"40",X"E1",X"C6",X"40",X"9E",X"CC",X"40",X"A6",X"CD",X"40",X"B2",X"CB",X"40",X"26",
		X"C4",X"40",X"0F",X"DC",X"40",X"29",X"DC",X"40",X"33",X"DB",X"40",X"5B",X"DB",X"40",X"F7",X"DA",
		X"40",X"BC",X"DA",X"40",X"50",X"DA",X"40",X"07",X"D9",X"C5",X"12",X"A9",X"02",X"90",X"03",X"40",
		X"1D",X"D9",X"40",X"9E",X"C2",X"C5",X"33",X"49",X"80",X"F0",X"B5",X"C5",X"18",X"49",X"5F",X"85",
		X"18",X"C2",X"60",X"C9",X"00",X"40",X"E1",X"C2",X"40",X"36",X"CC",X"40",X"05",X"DC",X"90",X"17",
		X"40",X"CB",X"DC",X"C5",X"08",X"A9",X"02",X"D0",X"03",X"2C",X"64",X"C1",X"E6",X"09",X"C5",X"09",
		X"49",X"01",X"85",X"09",X"2C",X"64",X"C1",X"40",X"CB",X"DC",X"40",X"E1",X"DC",X"C9",X"00",X"8D",
		X"00",X"54",X"40",X"3D",X"DA",X"A6",X"08",X"B0",X"E3",X"C9",X"00",X"85",X"12",X"CD",X"01",X"10",
		X"29",X"FF",X"49",X"08",X"F0",X"03",X"40",X"C3",X"E8",X"C9",X"00",X"8D",X"01",X"10",X"85",X"09",
		X"85",X"07",X"C9",X"00",X"8D",X"02",X"10",X"C2",X"02",X"40",X"A6",X"DC",X"2C",X"2E",X"C1",X"2C",
		X"31",X"C1",X"CD",X"00",X"10",X"10",X"FB",X"40",X"D7",X"D4",X"40",X"19",X"D6",X"40",X"36",X"CC",
		X"40",X"5D",X"D4",X"E6",X"30",X"CD",X"00",X"10",X"50",X"FB",X"40",X"18",X"EB",X"60",X"C5",X"33",
		X"49",X"40",X"F0",X"0A",X"C5",X"30",X"A9",X"80",X"90",X"04",X"C9",X"80",X"85",X"33",X"60",X"C9",
		X"00",X"CA",X"95",X"00",X"E8",X"E0",X"F1",X"B0",X"F9",X"60",X"C9",X"00",X"CA",X"9D",X"00",X"04",
		X"E8",X"B0",X"FA",X"CA",X"9D",X"00",X"03",X"9D",X"00",X"02",X"E8",X"B0",X"F7",X"60",X"C9",X"00",
		X"CA",X"9D",X"00",X"05",X"9D",X"00",X"06",X"9D",X"00",X"07",X"E8",X"B0",X"F4",X"60",X"C9",X"00",
		X"CA",X"9D",X"00",X"40",X"9D",X"00",X"44",X"E8",X"B0",X"F7",X"C9",X"00",X"9D",X"00",X"41",X"9D",
		X"00",X"45",X"E8",X"B0",X"F7",X"9D",X"00",X"42",X"9D",X"00",X"46",X"9D",X"00",X"43",X"9D",X"00",
		X"47",X"E8",X"B0",X"F1",X"C0",X"00",X"C9",X"00",X"99",X"80",X"04",X"A8",X"A0",X"20",X"90",X"F8",
		X"60",X"C2",X"07",X"DD",X"23",X"C3",X"9D",X"00",X"5C",X"DD",X"2B",X"C3",X"9D",X"08",X"5C",X"AA",
		X"10",X"F1",X"60",X"FF",X"F8",X"FF",X"C0",X"3F",X"C7",X"E3",X"00",X"FF",X"C7",X"E1",X"93",X"49",
		X"3F",X"7F",X"00",X"C5",X"33",X"49",X"C0",X"B0",X"26",X"C5",X"18",X"49",X"20",X"B0",X"06",X"40",
		X"60",X"C3",X"40",X"92",X"C3",X"40",X"5B",X"C4",X"C2",X"40",X"40",X"1B",X"D4",X"40",X"D8",X"C4",
		X"40",X"8C",X"CE",X"40",X"CC",X"C8",X"40",X"30",X"D4",X"40",X"A2",X"CA",X"40",X"99",X"C6",X"60",
		X"C5",X"7A",X"B0",X"2D",X"C9",X"80",X"85",X"7A",X"C9",X"03",X"85",X"8E",X"C9",X"14",X"85",X"8F",
		X"85",X"91",X"C9",X"80",X"85",X"7B",X"C9",X"00",X"85",X"39",X"40",X"7F",X"D4",X"A9",X"06",X"B0",
		X"04",X"C9",X"38",X"85",X"7B",X"C9",X"E0",X"85",X"7C",X"C5",X"07",X"B0",X"04",X"C9",X"90",X"85",
		X"7B",X"60",X"C5",X"7A",X"49",X"68",X"B0",X"51",X"C5",X"37",X"49",X"03",X"CA",X"C5",X"7B",X"18",
		X"7D",X"EA",X"C3",X"85",X"7B",X"C5",X"7A",X"49",X"10",X"B0",X"1E",X"C5",X"37",X"49",X"04",X"F0",
		X"03",X"40",X"FB",X"C3",X"C5",X"37",X"49",X"08",X"F0",X"0F",X"CA",X"C5",X"7C",X"18",X"7D",X"EA",
		X"C3",X"A9",X"E0",X"90",X"02",X"C9",X"E0",X"85",X"7C",X"C5",X"7C",X"A9",X"70",X"D0",X"02",X"C9",
		X"70",X"2A",X"2A",X"2A",X"2A",X"58",X"E9",X"07",X"CA",X"DD",X"F3",X"C3",X"85",X"CD",X"25",X"F0",
		X"F0",X"07",X"C5",X"CD",X"85",X"F0",X"40",X"44",X"DA",X"60",X"00",X"02",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"02",X"12",X"11",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"A6",X"8E",X"B0",X"26",X"C9",
		X"03",X"85",X"8E",X"C5",X"7C",X"A9",X"7D",X"90",X"1C",X"A6",X"7C",X"C5",X"7C",X"A9",X"9A",X"50",
		X"14",X"A6",X"7C",X"C5",X"7C",X"A9",X"B8",X"50",X"0C",X"A6",X"7C",X"C5",X"7C",X"A9",X"7C",X"D0",
		X"04",X"C9",X"7C",X"85",X"7C",X"60",X"C5",X"33",X"49",X"C0",X"B0",X"2E",X"C5",X"18",X"49",X"A0",
		X"B0",X"28",X"C5",X"2C",X"F0",X"04",X"49",X"10",X"F0",X"20",X"C5",X"7A",X"49",X"10",X"F0",X"06",
		X"C5",X"80",X"A9",X"10",X"D0",X"14",X"C9",X"03",X"85",X"96",X"C9",X"E0",X"58",X"E5",X"7C",X"A9",
		X"0A",X"90",X"07",X"E6",X"96",X"58",X"E9",X"14",X"D0",X"F9",X"60",X"C5",X"7A",X"49",X"FB",X"85",
		X"7A",X"49",X"48",X"B0",X"32",X"C9",X"2C",X"85",X"7F",X"C5",X"7A",X"49",X"10",X"B0",X"1D",X"25",
		X"37",X"49",X"10",X"F0",X"22",X"C5",X"18",X"49",X"20",X"B0",X"1C",X"C5",X"90",X"F0",X"18",X"C9",
		X"90",X"85",X"7A",X"C9",X"3F",X"85",X"80",X"C9",X"03",X"40",X"44",X"DA",X"A6",X"80",X"40",X"B6",
		X"C4",X"40",X"98",X"C4",X"40",X"A1",X"C4",X"60",X"C5",X"80",X"A9",X"2F",X"90",X"02",X"A6",X"7C",
		X"60",X"C5",X"80",X"A9",X"20",X"D0",X"0E",X"A9",X"10",X"D0",X"08",X"C5",X"80",X"B0",X"04",X"C9",
		X"84",X"85",X"7A",X"E6",X"7C",X"60",X"C2",X"06",X"C5",X"80",X"A9",X"08",X"B0",X"05",X"C9",X"04",
		X"40",X"44",X"DA",X"58",X"E9",X"08",X"90",X"05",X"AA",X"A9",X"08",X"D0",X"F7",X"C9",X"29",X"18",
		X"69",X"04",X"AA",X"10",X"FA",X"85",X"7F",X"60",X"C5",X"97",X"49",X"58",X"B0",X"34",X"C2",X"06",
		X"8A",X"28",X"C5",X"98",X"18",X"7D",X"77",X"C5",X"10",X"02",X"29",X"0F",X"85",X"38",X"C5",X"99",
		X"18",X"7D",X"78",X"C5",X"85",X"39",X"40",X"87",X"C5",X"40",X"3A",X"C6",X"68",X"CA",X"C5",X"18",
		X"50",X"10",X"AA",X"AA",X"10",X"DA",X"40",X"0A",X"CD",X"C5",X"97",X"49",X"02",X"F0",X"03",X"40",
		X"73",X"C6",X"60",X"C5",X"97",X"49",X"40",X"B0",X"5D",X"C9",X"00",X"85",X"D4",X"C0",X"06",X"C5",
		X"98",X"18",X"79",X"7F",X"C5",X"10",X"02",X"29",X"0F",X"85",X"38",X"C5",X"99",X"18",X"79",X"80",
		X"C5",X"85",X"39",X"40",X"87",X"C5",X"C5",X"8C",X"A9",X"05",X"B0",X"06",X"C5",X"8D",X"A9",X"07",
		X"F0",X"09",X"C5",X"8D",X"A9",X"01",X"F0",X"03",X"58",X"D0",X"01",X"18",X"46",X"D4",X"88",X"88",
		X"10",X"CD",X"C5",X"D4",X"F0",X"20",X"85",X"9E",X"C5",X"97",X"49",X"20",X"F0",X"12",X"C9",X"41",
		X"85",X"97",X"E6",X"21",X"C9",X"20",X"85",X"9D",X"C9",X"06",X"40",X"44",X"DA",X"2C",X"76",X"C5",
		X"C5",X"97",X"09",X"08",X"85",X"97",X"60",X"FC",X"04",X"04",X"04",X"04",X"FC",X"FC",X"FC",X"F6",
		X"0A",X"0A",X"0A",X"0A",X"F6",X"F6",X"F6",X"8A",X"28",X"98",X"28",X"C5",X"23",X"18",X"65",X"39",
		X"49",X"F0",X"85",X"CD",X"40",X"7F",X"D4",X"85",X"CE",X"C5",X"38",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"26",X"CD",X"18",X"65",X"CD",X"C8",X"26",X"CE",X"C9",X"9D",X"90",X"03",X"18",X"69",X"80",X"85",
		X"D5",X"C9",X"EE",X"65",X"CE",X"85",X"D6",X"C5",X"38",X"49",X"10",X"08",X"D1",X"D5",X"48",X"B0",
		X"04",X"2A",X"2A",X"2A",X"2A",X"49",X"0F",X"85",X"8C",X"C9",X"40",X"85",X"C9",X"C5",X"8C",X"85",
		X"C7",X"40",X"3B",X"D4",X"C9",X"00",X"18",X"65",X"CB",X"85",X"D5",X"C9",X"F7",X"65",X"CC",X"85",
		X"D6",X"C5",X"39",X"49",X"0C",X"0A",X"0A",X"18",X"65",X"D5",X"85",X"D5",X"C5",X"38",X"49",X"0F",
		X"C8",X"C5",X"39",X"49",X"03",X"CA",X"C9",X"00",X"85",X"8D",X"D1",X"D5",X"5D",X"32",X"C6",X"F0",
		X"04",X"C9",X"01",X"85",X"8D",X"C5",X"D6",X"18",X"69",X"04",X"85",X"D6",X"D1",X"D5",X"5D",X"32",
		X"C6",X"F0",X"07",X"C5",X"8D",X"18",X"69",X"04",X"85",X"8D",X"8A",X"18",X"69",X"04",X"CA",X"D1",
		X"D5",X"5D",X"32",X"C6",X"F0",X"07",X"C5",X"8D",X"18",X"69",X"02",X"85",X"8D",X"68",X"C8",X"68",
		X"CA",X"60",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"C5",X"8C",X"C6",X"8D",X"E0",X"01",
		X"F0",X"56",X"E0",X"07",X"B0",X"08",X"A9",X"05",X"F0",X"4E",X"A9",X"09",X"F0",X"4A",X"A9",X"06",
		X"90",X"21",X"A9",X"0E",X"D0",X"1D",X"A9",X"08",X"F0",X"19",X"A9",X"09",X"F0",X"15",X"E0",X"06",
		X"F0",X"04",X"E0",X"05",X"B0",X"32",X"C9",X"08",X"85",X"97",X"C2",X"01",X"40",X"A6",X"DC",X"C9",
		X"05",X"B0",X"0B",X"C9",X"40",X"85",X"97",X"C2",X"01",X"40",X"A6",X"DC",X"C9",X"01",X"40",X"44",
		X"DA",X"C2",X"01",X"40",X"A6",X"DC",X"C9",X"20",X"85",X"9D",X"C5",X"18",X"09",X"80",X"85",X"18",
		X"C5",X"38",X"85",X"29",X"C5",X"39",X"85",X"2A",X"60",X"C5",X"7A",X"49",X"48",X"F0",X"28",X"28",
		X"A6",X"80",X"B0",X"0C",X"C5",X"33",X"09",X"40",X"85",X"33",X"C9",X"00",X"85",X"7A",X"85",X"30",
		X"C5",X"80",X"2A",X"2A",X"2A",X"49",X"03",X"CA",X"68",X"A9",X"08",X"B0",X"05",X"8A",X"18",X"69",
		X"04",X"CA",X"DD",X"C8",X"C6",X"85",X"7F",X"60",X"66",X"62",X"5E",X"5A",X"76",X"72",X"6E",X"6A",
		X"C5",X"36",X"49",X"20",X"B0",X"06",X"C5",X"7A",X"49",X"48",X"F0",X"04",X"C9",X"00",X"85",X"96",
		X"60",X"40",X"EE",X"C6",X"40",X"2B",X"C7",X"40",X"68",X"C7",X"40",X"8F",X"C7",X"60",X"C5",X"18",
		X"49",X"A0",X"B0",X"36",X"C5",X"96",X"F0",X"32",X"C5",X"7A",X"F0",X"2E",X"49",X"10",X"F0",X"06",
		X"C5",X"80",X"A9",X"10",X"D0",X"23",X"C9",X"20",X"85",X"8F",X"C9",X"00",X"85",X"90",X"C9",X"E0",
		X"58",X"E5",X"7C",X"85",X"CD",X"F0",X"12",X"F8",X"C5",X"8F",X"18",X"69",X"02",X"85",X"8F",X"C5",
		X"90",X"69",X"00",X"85",X"90",X"A6",X"CD",X"B0",X"EF",X"B8",X"60",X"C2",X"04",X"40",X"17",X"DB",
		X"C9",X"5D",X"85",X"CF",X"C0",X"02",X"C5",X"18",X"49",X"A0",X"B0",X"24",X"C5",X"2C",X"F0",X"04",
		X"49",X"10",X"F0",X"1C",X"C0",X"00",X"C5",X"90",X"B0",X"02",X"C9",X"0A",X"18",X"65",X"CF",X"91",
		X"DD",X"E6",X"DD",X"C2",X"8F",X"40",X"7D",X"DB",X"A6",X"DD",X"A6",X"DD",X"D1",X"DD",X"B0",X"07",
		X"C9",X"5D",X"91",X"DD",X"88",X"10",X"F9",X"60",X"C0",X"00",X"C9",X"67",X"85",X"CD",X"C5",X"90",
		X"F0",X"0A",X"C5",X"30",X"49",X"04",X"F0",X"04",X"C9",X"01",X"85",X"CD",X"C5",X"CD",X"99",X"82",
		X"40",X"C5",X"CD",X"A9",X"67",X"F0",X"02",X"E6",X"CD",X"A8",X"A0",X"08",X"90",X"EE",X"60",X"E6",
		X"E3",X"C4",X"24",X"C2",X"01",X"C5",X"7C",X"85",X"39",X"40",X"81",X"D4",X"85",X"8C",X"A9",X"0F",
		X"F0",X"07",X"40",X"D7",X"D5",X"C5",X"D4",X"F0",X"0A",X"C9",X"00",X"85",X"39",X"88",X"AA",X"10",
		X"E4",X"50",X"32",X"C5",X"E3",X"49",X"08",X"F0",X"2C",X"C5",X"E8",X"F0",X"0B",X"C5",X"7A",X"49",
		X"10",X"B0",X"05",X"C9",X"09",X"40",X"44",X"DA",X"C0",X"00",X"84",X"E8",X"C2",X"00",X"DD",X"03",
		X"C8",X"85",X"CE",X"E8",X"DD",X"03",X"C8",X"85",X"CD",X"E8",X"DD",X"03",X"C8",X"91",X"CD",X"E8",
		X"E0",X"18",X"B0",X"EA",X"60",X"C9",X"55",X"85",X"E8",X"C0",X"00",X"C2",X"00",X"DD",X"03",X"C8",
		X"85",X"CE",X"E8",X"DD",X"03",X"C8",X"85",X"CD",X"E8",X"C9",X"00",X"91",X"CD",X"E8",X"E0",X"18",
		X"B0",X"EB",X"60",X"44",X"AF",X"01",X"44",X"B0",X"01",X"44",X"CF",X"01",X"44",X"D0",X"01",X"40",
		X"AF",X"F0",X"40",X"B0",X"F1",X"40",X"CF",X"F2",X"40",X"D0",X"F3",X"C5",X"18",X"49",X"20",X"B0",
		X"51",X"C5",X"35",X"50",X"39",X"C2",X"00",X"86",X"E9",X"D5",X"3A",X"B0",X"03",X"40",X"56",X"C9",
		X"D5",X"3A",X"F0",X"20",X"D5",X"44",X"0A",X"C8",X"D9",X"73",X"C8",X"85",X"D9",X"D9",X"74",X"C8",
		X"85",X"DA",X"C9",X"C8",X"28",X"C9",X"50",X"28",X"40",X"1B",X"D4",X"40",X"13",X"C5",X"6C",X"D9",
		X"00",X"40",X"30",X"D4",X"C5",X"E9",X"18",X"69",X"10",X"CA",X"A9",X"40",X"90",X"C9",X"C5",X"35",
		X"49",X"40",X"F0",X"0E",X"C5",X"3A",X"05",X"4A",X"05",X"5A",X"05",X"6A",X"B0",X"04",X"C9",X"80",
		X"85",X"35",X"60",X"87",X"C8",X"97",X"C8",X"97",X"C8",X"97",X"C8",X"87",X"C8",X"A0",X"C8",X"A9",
		X"C8",X"B2",X"C8",X"87",X"C8",X"87",X"C8",X"40",X"BB",X"C8",X"40",X"7E",X"D0",X"40",X"DA",X"C8",
		X"40",X"83",X"CD",X"40",X"3A",X"C9",X"60",X"40",X"BB",X"C8",X"40",X"1B",X"CF",X"2C",X"8D",X"C8",
		X"40",X"BB",X"C8",X"40",X"86",X"CF",X"2C",X"8D",X"C8",X"40",X"45",X"CD",X"40",X"AC",X"CF",X"2C",
		X"8D",X"C8",X"40",X"E7",X"CF",X"40",X"42",X"CC",X"2C",X"90",X"C8",X"40",X"04",X"CD",X"C5",X"97",
		X"49",X"02",X"F0",X"07",X"C9",X"40",X"85",X"97",X"40",X"64",X"C5",X"60",X"C5",X"97",X"49",X"20",
		X"F0",X"63",X"C0",X"00",X"C5",X"99",X"A9",X"7E",X"90",X"45",X"C5",X"97",X"49",X"20",X"F0",X"55",
		X"C0",X"00",X"C5",X"99",X"A9",X"DE",X"D0",X"37",X"A9",X"40",X"90",X"33",X"C0",X"01",X"C5",X"9E",
		X"2A",X"2A",X"49",X"03",X"CA",X"DD",X"36",X"C9",X"85",X"CD",X"C5",X"A1",X"A9",X"05",X"F0",X"04",
		X"A9",X"06",X"B0",X"0F",X"C5",X"9D",X"2A",X"C5",X"CD",X"90",X"08",X"29",X"FF",X"10",X"02",X"09",
		X"02",X"85",X"CD",X"C5",X"CD",X"18",X"79",X"98",X"00",X"99",X"98",X"00",X"88",X"50",X"08",X"C5",
		X"9E",X"49",X"03",X"CA",X"2C",X"F5",X"C8",X"A6",X"9D",X"B0",X"0A",X"C5",X"97",X"49",X"DF",X"85",
		X"97",X"C9",X"00",X"85",X"9E",X"60",X"FE",X"FE",X"02",X"02",X"C5",X"97",X"49",X"40",X"F0",X"15",
		X"A6",X"9D",X"B0",X"03",X"40",X"F9",X"D1",X"C5",X"9D",X"2A",X"2A",X"2A",X"85",X"CD",X"C9",X"59",
		X"58",X"E5",X"CD",X"85",X"9C",X"60",X"C5",X"18",X"50",X"1C",X"C5",X"35",X"49",X"C0",X"B0",X"16",
		X"8A",X"18",X"69",X"3A",X"85",X"D9",X"C9",X"00",X"85",X"DA",X"C0",X"0F",X"C9",X"00",X"91",X"D9",
		X"88",X"10",X"FB",X"40",X"04",X"CA",X"60",X"01",X"02",X"06",X"02",X"02",X"09",X"06",X"02",X"09",
		X"06",X"02",X"02",X"03",X"02",X"05",X"06",X"07",X"09",X"05",X"02",X"09",X"07",X"02",X"06",X"09",
		X"06",X"01",X"01",X"02",X"08",X"03",X"09",X"02",X"01",X"02",X"08",X"02",X"09",X"03",X"09",X"02",
		X"01",X"08",X"09",X"09",X"09",X"02",X"06",X"07",X"02",X"09",X"03",X"04",X"06",X"07",X"07",X"07",
		X"02",X"09",X"06",X"04",X"04",X"07",X"02",X"09",X"09",X"03",X"04",X"05",X"08",X"07",X"07",X"01",
		X"02",X"04",X"04",X"08",X"03",X"09",X"06",X"01",X"01",X"02",X"02",X"04",X"04",X"06",X"09",X"08",
		X"03",X"04",X"02",X"04",X"08",X"09",X"01",X"02",X"04",X"04",X"01",X"04",X"04",X"07",X"01",X"08",
		X"04",X"04",X"05",X"09",X"02",X"07",X"01",X"08",X"04",X"05",X"04",X"09",X"02",X"07",X"04",X"04",
		X"04",X"05",X"01",X"07",X"04",X"04",X"05",X"07",X"02",X"04",X"01",X"07",X"08",X"09",X"05",X"01",
		X"07",X"06",X"05",X"07",X"C9",X"00",X"85",X"92",X"C5",X"18",X"49",X"40",X"B0",X"06",X"C5",X"22",
		X"A9",X"06",X"90",X"1E",X"8A",X"B0",X"1B",X"85",X"39",X"40",X"7F",X"D4",X"A9",X"04",X"90",X"12",
		X"A9",X"07",X"90",X"08",X"A9",X"0B",X"F0",X"04",X"A9",X"0E",X"90",X"06",X"E6",X"92",X"C9",X"30",
		X"B0",X"0E",X"C5",X"17",X"A9",X"C0",X"90",X"02",X"C9",X"C0",X"A9",X"40",X"D0",X"02",X"C9",X"80",
		X"85",X"98",X"C9",X"08",X"85",X"99",X"C9",X"00",X"85",X"97",X"85",X"9E",X"40",X"13",X"C5",X"C5",
		X"9E",X"B0",X"44",X"C9",X"80",X"95",X"3A",X"C5",X"98",X"95",X"3B",X"C5",X"99",X"95",X"3C",X"C5",
		X"92",X"F0",X"0A",X"C5",X"17",X"49",X"03",X"C8",X"D9",X"00",X"CA",X"10",X"22",X"C5",X"90",X"F0",
		X"0E",X"C5",X"35",X"49",X"20",X"B0",X"08",X"09",X"20",X"85",X"35",X"C9",X"00",X"F0",X"10",X"C4",
		X"1F",X"E6",X"1F",X"A0",X"88",X"90",X"05",X"C9",X"2E",X"85",X"1F",X"C8",X"D9",X"77",X"C9",X"95",
		X"44",X"C8",X"D9",X"98",X"CA",X"95",X"3F",X"60",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",
		X"54",X"55",X"C5",X"18",X"49",X"20",X"B0",X"0A",X"C9",X"40",X"85",X"E9",X"C5",X"7A",X"49",X"58",
		X"F0",X"01",X"60",X"C9",X"00",X"85",X"CD",X"CA",X"8A",X"28",X"E4",X"E9",X"F0",X"3B",X"C9",X"00",
		X"85",X"CF",X"D5",X"3A",X"F0",X"33",X"49",X"40",X"B0",X"2F",X"D5",X"3B",X"85",X"92",X"D5",X"3C",
		X"85",X"93",X"D5",X"44",X"A9",X"06",X"90",X"0A",X"C9",X"0E",X"85",X"94",X"C9",X"10",X"85",X"95",
		X"B0",X"14",X"A9",X"09",X"90",X"0A",X"C9",X"0E",X"85",X"94",X"C9",X"0C",X"85",X"95",X"B0",X"06",
		X"C9",X"10",X"85",X"94",X"85",X"95",X"40",X"3F",X"CB",X"68",X"CA",X"C5",X"CF",X"F0",X"2C",X"95",
		X"41",X"C9",X"A0",X"85",X"CE",X"D4",X"44",X"D9",X"35",X"CB",X"95",X"40",X"F0",X"06",X"C5",X"7A",
		X"49",X"04",X"F0",X"0E",X"C9",X"41",X"85",X"CE",X"C9",X"20",X"95",X"40",X"E6",X"21",X"C9",X"06",
		X"B0",X"02",X"C9",X"07",X"40",X"44",X"DA",X"C5",X"CE",X"95",X"3A",X"8A",X"18",X"69",X"10",X"CA",
		X"A9",X"40",X"90",X"84",X"60",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"00",X"10",X"10",X"C5",
		X"7B",X"58",X"E5",X"92",X"CA",X"10",X"11",X"29",X"FF",X"CA",X"C5",X"CD",X"09",X"01",X"85",X"CD",
		X"C5",X"CF",X"09",X"02",X"85",X"CF",X"B0",X"0C",X"C5",X"CD",X"09",X"02",X"85",X"CD",X"C5",X"CF",
		X"09",X"01",X"85",X"CF",X"E0",X"10",X"50",X"02",X"10",X"41",X"C5",X"7C",X"58",X"E5",X"93",X"C8",
		X"10",X"11",X"29",X"FF",X"C8",X"C5",X"CD",X"09",X"04",X"85",X"CD",X"C5",X"CF",X"09",X"08",X"85",
		X"CF",X"B0",X"0C",X"C5",X"CD",X"09",X"08",X"85",X"CD",X"C5",X"CF",X"09",X"04",X"85",X"CF",X"A0",
		X"10",X"10",X"18",X"E4",X"94",X"10",X"14",X"A4",X"95",X"10",X"10",X"C5",X"7A",X"09",X"20",X"85",
		X"7A",X"C5",X"CD",X"85",X"81",X"C9",X"10",X"85",X"80",X"B0",X"89",X"C9",X"00",X"85",X"CF",X"85",
		X"CD",X"60",X"C2",X"00",X"C0",X"00",X"D5",X"3A",X"F0",X"2D",X"49",X"60",X"F0",X"04",X"C9",X"00",
		X"F0",X"03",X"C5",X"30",X"2A",X"58",X"4A",X"49",X"03",X"99",X"80",X"04",X"D5",X"3F",X"99",X"81",
		X"04",X"D5",X"3B",X"18",X"69",X"08",X"29",X"FF",X"99",X"82",X"04",X"D5",X"3C",X"58",X"E9",X"08",
		X"99",X"83",X"04",X"A8",X"A8",X"A8",X"A8",X"8A",X"18",X"69",X"10",X"CA",X"A9",X"40",X"90",X"C6",
		X"A9",X"50",X"D0",X"36",X"C5",X"7A",X"49",X"58",X"F0",X"BC",X"C2",X"00",X"C5",X"7F",X"85",X"CD",
		X"C9",X"01",X"99",X"80",X"04",X"C5",X"CD",X"99",X"81",X"04",X"C5",X"7B",X"18",X"7D",X"2E",X"CC",
		X"29",X"FF",X"99",X"82",X"04",X"E8",X"C5",X"7C",X"18",X"7D",X"2E",X"CC",X"99",X"83",X"04",X"E6",
		X"CD",X"A8",X"A8",X"A8",X"A8",X"E8",X"E0",X"08",X"B0",X"D6",X"40",X"06",X"C3",X"60",X"00",X"F0",
		X"10",X"F0",X"00",X"00",X"10",X"00",X"C0",X"20",X"D9",X"80",X"04",X"99",X"00",X"48",X"88",X"10",
		X"F7",X"60",X"C5",X"97",X"49",X"10",X"F0",X"32",X"C9",X"80",X"85",X"97",X"C9",X"0A",X"40",X"44",
		X"DA",X"C6",X"8B",X"F0",X"10",X"DD",X"FE",X"01",X"9D",X"00",X"02",X"DD",X"FF",X"01",X"9D",X"01",
		X"02",X"AA",X"AA",X"B0",X"F0",X"C5",X"98",X"49",X"07",X"29",X"07",X"18",X"65",X"98",X"8D",X"00",
		X"02",X"C5",X"99",X"8D",X"01",X"02",X"E6",X"8B",X"E6",X"8B",X"60",X"C0",X"00",X"C9",X"00",X"91",
		X"DD",X"A8",X"91",X"DD",X"98",X"18",X"69",X"1F",X"C8",X"A0",X"A0",X"90",X"F0",X"8A",X"C8",X"A4",
		X"8B",X"B0",X"01",X"60",X"D9",X"00",X"02",X"99",X"FE",X"01",X"A8",X"2C",X"8F",X"CC",X"C6",X"8B",
		X"F0",X"59",X"DD",X"FE",X"01",X"F0",X"50",X"85",X"38",X"DD",X"FF",X"01",X"18",X"65",X"96",X"9D",
		X"FF",X"01",X"58",X"E9",X"08",X"85",X"39",X"40",X"63",X"CD",X"C5",X"39",X"A9",X"E0",X"90",X"0A",
		X"40",X"7B",X"CC",X"A6",X"8B",X"A6",X"8B",X"2C",X"F7",X"CC",X"49",X"07",X"C8",X"D9",X"FC",X"CC",
		X"85",X"CD",X"C9",X"00",X"C8",X"91",X"DD",X"A8",X"91",X"DD",X"C0",X"20",X"91",X"DD",X"A8",X"91",
		X"DD",X"98",X"18",X"69",X"1F",X"C8",X"C5",X"CD",X"91",X"DD",X"A8",X"E6",X"CD",X"C5",X"CD",X"91",
		X"DD",X"E6",X"CD",X"A0",X"80",X"90",X"EA",X"AA",X"AA",X"B0",X"A7",X"60",X"80",X"86",X"8C",X"92",
		X"98",X"9E",X"A4",X"AA",X"C5",X"97",X"49",X"40",X"B0",X"0B",X"C6",X"8B",X"F0",X"07",X"40",X"16",
		X"CD",X"AA",X"AA",X"B0",X"F9",X"60",X"DD",X"FE",X"01",X"85",X"38",X"49",X"F8",X"18",X"69",X"08",
		X"58",X"E5",X"98",X"D0",X"02",X"29",X"FF",X"A9",X"0C",X"D0",X"19",X"DD",X"FF",X"01",X"85",X"39",
		X"18",X"69",X"08",X"58",X"E5",X"99",X"D0",X"02",X"29",X"FF",X"A9",X"0C",X"D0",X"06",X"C5",X"97",
		X"09",X"02",X"85",X"97",X"60",X"C6",X"8B",X"F0",X"19",X"40",X"16",X"CD",X"C5",X"97",X"49",X"02",
		X"F0",X"0C",X"40",X"63",X"CD",X"40",X"7B",X"CC",X"C5",X"97",X"49",X"FD",X"85",X"97",X"AA",X"AA",
		X"B0",X"E7",X"60",X"C5",X"38",X"2A",X"2A",X"2A",X"85",X"CD",X"C9",X"00",X"85",X"CE",X"C5",X"39",
		X"49",X"F8",X"0A",X"46",X"CE",X"0A",X"46",X"CE",X"05",X"CD",X"85",X"DD",X"C5",X"CE",X"09",X"40",
		X"85",X"DE",X"60",X"C5",X"97",X"49",X"40",X"F0",X"1C",X"C5",X"99",X"A9",X"40",X"90",X"09",X"18",
		X"65",X"96",X"85",X"99",X"A9",X"E8",X"90",X"0D",X"C5",X"A1",X"B0",X"06",X"C5",X"35",X"49",X"DF",
		X"85",X"35",X"40",X"F9",X"D1",X"60",X"C2",X"00",X"D5",X"3A",X"2A",X"90",X"07",X"C9",X"40",X"95",
		X"3A",X"40",X"CB",X"CD",X"8A",X"18",X"69",X"10",X"CA",X"A9",X"40",X"90",X"EB",X"C5",X"8A",X"F0",
		X"09",X"40",X"4A",X"CE",X"40",X"1F",X"CE",X"40",X"78",X"CE",X"60",X"C4",X"8A",X"F0",X"1E",X"D9",
		X"FC",X"02",X"99",X"00",X"03",X"D9",X"FD",X"02",X"99",X"01",X"03",X"D9",X"FE",X"02",X"99",X"02",
		X"03",X"D9",X"FF",X"02",X"99",X"03",X"03",X"88",X"88",X"88",X"88",X"B0",X"E2",X"D5",X"3B",X"8D",
		X"00",X"03",X"D5",X"3C",X"18",X"69",X"10",X"8D",X"01",X"03",X"D4",X"44",X"D9",X"15",X"CE",X"8D",
		X"02",X"03",X"58",X"E9",X"01",X"40",X"C5",X"DB",X"C9",X"20",X"8D",X"03",X"03",X"C5",X"8A",X"18",
		X"69",X"04",X"85",X"8A",X"60",X"0D",X"0A",X"0A",X"0A",X"0D",X"0A",X"07",X"0A",X"07",X"07",X"C4",
		X"8A",X"D9",X"FF",X"02",X"B0",X"23",X"D9",X"FC",X"02",X"85",X"38",X"D9",X"FD",X"02",X"85",X"39",
		X"C9",X"00",X"28",X"99",X"FE",X"02",X"40",X"63",X"CD",X"68",X"C8",X"91",X"DD",X"A8",X"91",X"DD",
		X"C5",X"8A",X"58",X"E9",X"04",X"85",X"8A",X"B0",X"D6",X"60",X"C4",X"8A",X"98",X"F0",X"28",X"28",
		X"D9",X"FC",X"02",X"85",X"38",X"D9",X"FD",X"02",X"85",X"39",X"40",X"63",X"CD",X"D9",X"FE",X"02",
		X"C8",X"D9",X"DF",X"DB",X"18",X"69",X"75",X"C0",X"00",X"91",X"DD",X"A8",X"C9",X"74",X"91",X"DD",
		X"68",X"58",X"E9",X"04",X"C8",X"B0",X"D5",X"60",X"C4",X"8A",X"F0",X"0F",X"D9",X"FF",X"02",X"58",
		X"E9",X"01",X"99",X"FF",X"02",X"88",X"88",X"88",X"88",X"B0",X"F1",X"60",X"C5",X"97",X"49",X"4C",
		X"F0",X"58",X"49",X"48",X"B0",X"54",X"C5",X"99",X"85",X"39",X"18",X"65",X"23",X"85",X"CE",X"40",
		X"7F",X"D4",X"85",X"CD",X"A9",X"0B",X"F0",X"04",X"A9",X"0E",X"B0",X"0C",X"C5",X"98",X"A9",X"60",
		X"90",X"38",X"C5",X"CE",X"A9",X"60",X"D0",X"16",X"C5",X"CD",X"A9",X"0C",X"B0",X"2C",X"C4",X"24",
		X"A8",X"C5",X"CE",X"50",X"02",X"88",X"88",X"40",X"81",X"D4",X"A9",X"0C",X"B0",X"1C",X"C9",X"20",
		X"85",X"EF",X"C5",X"98",X"85",X"38",X"C5",X"99",X"85",X"39",X"40",X"63",X"CD",X"C5",X"DD",X"85",
		X"ED",X"C5",X"DE",X"85",X"EE",X"C9",X"0F",X"40",X"C5",X"DB",X"C5",X"EF",X"F0",X"24",X"C2",X"02",
		X"DD",X"EE",X"DB",X"95",X"F1",X"AA",X"10",X"F8",X"C5",X"ED",X"85",X"DD",X"C5",X"EE",X"85",X"DE",
		X"C0",X"05",X"C9",X"00",X"91",X"DD",X"88",X"10",X"FB",X"A6",X"EF",X"F0",X"05",X"C2",X"F3",X"40",
		X"71",X"DB",X"60",X"04",X"04",X"04",X"05",X"07",X"04",X"05",X"04",X"40",X"46",X"D2",X"50",X"54",
		X"C5",X"A3",X"B0",X"20",X"C5",X"9D",X"B0",X"1C",X"C5",X"96",X"2A",X"85",X"CE",X"C5",X"17",X"49",
		X"01",X"18",X"65",X"CE",X"CA",X"DD",X"13",X"CF",X"85",X"9F",X"C2",X"01",X"C5",X"98",X"10",X"02",
		X"C2",X"FF",X"86",X"A3",X"E6",X"9D",X"58",X"C5",X"96",X"E5",X"9F",X"85",X"CE",X"D0",X"19",X"C5",
		X"CE",X"29",X"FF",X"18",X"69",X"01",X"85",X"CE",X"58",X"C5",X"99",X"CA",X"E5",X"CE",X"85",X"99",
		X"8A",X"F0",X"1B",X"D0",X"19",X"2C",X"F6",X"D1",X"18",X"C5",X"99",X"65",X"CE",X"85",X"99",X"90",
		X"0D",X"2C",X"F6",X"D1",X"C5",X"A3",X"29",X"FF",X"18",X"69",X"01",X"85",X"A3",X"60",X"18",X"C5",
		X"98",X"65",X"A3",X"85",X"98",X"60",X"40",X"46",X"D2",X"50",X"14",X"E6",X"9D",X"40",X"E0",X"D1",
		X"C6",X"96",X"AA",X"AA",X"AA",X"8A",X"50",X"08",X"18",X"65",X"99",X"85",X"99",X"D0",X"0A",X"60",
		X"C5",X"99",X"58",X"E9",X"03",X"85",X"99",X"D0",X"F6",X"2C",X"F6",X"D1",X"40",X"46",X"D2",X"50",
		X"29",X"C5",X"9D",X"B0",X"0A",X"C2",X"01",X"C5",X"98",X"10",X"02",X"C2",X"FF",X"86",X"A4",X"E6",
		X"9D",X"40",X"E0",X"D1",X"C6",X"96",X"AA",X"AA",X"AA",X"8A",X"50",X"0F",X"18",X"65",X"99",X"85",
		X"99",X"D0",X"11",X"18",X"C5",X"98",X"65",X"A4",X"85",X"98",X"60",X"C5",X"99",X"58",X"E9",X"03",
		X"85",X"99",X"D0",X"F6",X"2C",X"F6",X"D1",X"40",X"46",X"D2",X"50",X"38",X"C5",X"96",X"B0",X"0A",
		X"C5",X"99",X"58",X"E9",X"03",X"85",X"99",X"90",X"EB",X"60",X"C5",X"A2",X"B0",X"09",X"C5",X"96",
		X"85",X"9F",X"C5",X"17",X"2A",X"85",X"A2",X"E6",X"9D",X"40",X"A2",X"D1",X"C5",X"9C",X"A9",X"53",
		X"F0",X"13",X"C5",X"99",X"A5",X"A2",X"90",X"08",X"E6",X"9C",X"C5",X"99",X"69",X"04",X"85",X"A2",
		X"E6",X"99",X"F0",X"C0",X"60",X"A6",X"99",X"F0",X"BB",X"C5",X"07",X"F0",X"1B",X"CD",X"01",X"10",
		X"49",X"10",X"F0",X"14",X"C5",X"22",X"49",X"07",X"A9",X"03",X"F0",X"E8",X"C5",X"18",X"49",X"40",
		X"B0",X"06",X"C5",X"22",X"A9",X"01",X"90",X"28",X"C5",X"99",X"A5",X"A2",X"D0",X"D6",X"C5",X"97",
		X"09",X"10",X"85",X"97",X"C2",X"FF",X"C5",X"18",X"49",X"40",X"F0",X"09",X"C5",X"22",X"49",X"07",
		X"CA",X"DD",X"76",X"D0",X"CA",X"86",X"CD",X"C5",X"99",X"58",X"E5",X"CD",X"90",X"03",X"85",X"A2",
		X"60",X"C9",X"01",X"85",X"A2",X"60",X"3E",X"32",X"30",X"2A",X"21",X"1B",X"14",X"0D",X"40",X"46",
		X"D2",X"50",X"20",X"C5",X"96",X"A9",X"05",X"D0",X"03",X"2C",X"20",X"CF",X"C5",X"A6",X"F0",X"1E",
		X"C5",X"9D",X"F0",X"1A",X"A6",X"9D",X"18",X"C9",X"7E",X"65",X"A6",X"CA",X"C9",X"D0",X"69",X"00",
		X"28",X"8A",X"28",X"60",X"73",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"9E",X"AF",X"C5",X"96",
		X"85",X"9F",X"C5",X"19",X"2A",X"2A",X"2A",X"85",X"CE",X"C6",X"A1",X"DD",X"A4",X"D0",X"58",X"E5",
		X"CE",X"85",X"9D",X"C5",X"18",X"49",X"40",X"F0",X"0D",X"C5",X"22",X"49",X"0F",X"0A",X"85",X"CE",
		X"C5",X"9D",X"E5",X"CE",X"85",X"9D",X"C5",X"7C",X"A5",X"99",X"90",X"35",X"E9",X"08",X"A5",X"99",
		X"90",X"26",X"E9",X"15",X"A5",X"99",X"90",X"0E",X"40",X"A2",X"D1",X"C9",X"69",X"85",X"A6",X"E6",
		X"99",X"B0",X"48",X"2C",X"F6",X"D1",X"40",X"A2",X"D1",X"C5",X"9D",X"2A",X"D0",X"04",X"E6",X"99",
		X"F0",X"F1",X"C9",X"77",X"85",X"A6",X"B0",X"33",X"40",X"A2",X"D1",X"C9",X"89",X"85",X"A6",X"B0",
		X"2A",X"69",X"08",X"A5",X"99",X"D0",X"F1",X"69",X"15",X"A5",X"99",X"D0",X"0E",X"40",X"A2",X"D1",
		X"C9",X"9E",X"85",X"A6",X"A6",X"99",X"B0",X"13",X"2C",X"F6",X"D1",X"40",X"A2",X"D1",X"C5",X"9D",
		X"2A",X"D0",X"04",X"A6",X"99",X"F0",X"BC",X"C9",X"AC",X"85",X"A6",X"C5",X"A4",X"F0",X"14",X"C5",
		X"A2",X"F0",X"10",X"A6",X"A2",X"18",X"C9",X"3B",X"65",X"A4",X"CA",X"C9",X"D1",X"69",X"00",X"28",
		X"8A",X"28",X"60",X"C9",X"50",X"85",X"A2",X"C5",X"7B",X"A5",X"98",X"90",X"26",X"E9",X"08",X"A5",
		X"98",X"90",X"1B",X"E9",X"15",X"A5",X"98",X"90",X"07",X"C9",X"2D",X"85",X"A4",X"E6",X"98",X"60",
		X"C5",X"9D",X"2A",X"D0",X"02",X"E6",X"98",X"C9",X"34",X"85",X"A4",X"E6",X"98",X"60",X"C9",X"42",
		X"85",X"A4",X"60",X"69",X"08",X"A5",X"98",X"D0",X"F5",X"69",X"15",X"A5",X"98",X"D0",X"07",X"C9",
		X"53",X"85",X"A4",X"A6",X"98",X"60",X"C5",X"9D",X"2A",X"D0",X"02",X"A6",X"98",X"C9",X"5A",X"85",
		X"A4",X"60",X"C2",X"04",X"CD",X"01",X"10",X"49",X"10",X"F0",X"02",X"C2",X"20",X"86",X"CE",X"C5",
		X"9D",X"45",X"CE",X"A5",X"A0",X"85",X"A0",X"F0",X"04",X"C5",X"96",X"85",X"9F",X"C5",X"96",X"58",
		X"E5",X"9F",X"85",X"CE",X"90",X"0A",X"18",X"C5",X"99",X"65",X"CE",X"85",X"99",X"D0",X"0D",X"60",
		X"C5",X"CE",X"29",X"FF",X"18",X"69",X"01",X"85",X"CE",X"2C",X"C6",X"D1",X"2C",X"F6",X"D1",X"60",
		X"58",X"C5",X"96",X"E9",X"03",X"B0",X"0E",X"C5",X"9D",X"2A",X"90",X"09",X"18",X"C5",X"99",X"69",
		X"01",X"85",X"99",X"D0",X"01",X"60",X"C6",X"9A",X"9A",X"C9",X"00",X"C8",X"99",X"97",X"00",X"A8",
		X"A0",X"10",X"B0",X"F8",X"60",X"C2",X"00",X"E0",X"40",X"B0",X"01",X"60",X"C0",X"00",X"C5",X"98",
		X"58",X"F5",X"3B",X"D0",X"06",X"C0",X"80",X"29",X"FF",X"69",X"01",X"85",X"CD",X"C5",X"99",X"58",
		X"F5",X"3C",X"D0",X"04",X"29",X"FF",X"69",X"01",X"28",X"8A",X"18",X"69",X"10",X"CA",X"68",X"18",
		X"65",X"CD",X"F0",X"D3",X"D0",X"D1",X"A9",X"20",X"D0",X"CD",X"98",X"F0",X"04",X"A6",X"98",X"A6",
		X"98",X"E6",X"98",X"2C",X"07",X"D2",X"DA",X"E8",X"E8",X"86",X"9A",X"C5",X"97",X"CA",X"49",X"40",
		X"B0",X"23",X"8A",X"49",X"20",X"F0",X"22",X"C2",X"0F",X"D5",X"7A",X"28",X"D5",X"97",X"95",X"7A",
		X"AA",X"10",X"F6",X"40",X"B3",X"CA",X"C2",X"00",X"C0",X"0F",X"D5",X"7A",X"95",X"97",X"68",X"95",
		X"7A",X"E8",X"88",X"10",X"F5",X"C6",X"9A",X"9A",X"60",X"C5",X"97",X"49",X"08",X"B0",X"04",X"C9",
		X"00",X"85",X"9E",X"C5",X"97",X"49",X"F7",X"85",X"97",X"C5",X"9E",X"49",X"0F",X"F0",X"3D",X"A9",
		X"0F",X"F0",X"0D",X"A9",X"0C",X"90",X"0C",X"C5",X"99",X"18",X"65",X"96",X"85",X"99",X"90",X"11",
		X"2C",X"F6",X"D1",X"C5",X"96",X"2A",X"85",X"CD",X"C5",X"99",X"18",X"65",X"CD",X"85",X"99",X"D0",
		X"EF",X"C5",X"9E",X"49",X"06",X"F0",X"04",X"A6",X"98",X"A6",X"98",X"C5",X"9E",X"49",X"09",X"F0",
		X"04",X"E6",X"98",X"E6",X"98",X"C9",X"00",X"85",X"9D",X"C9",X"80",X"60",X"40",X"05",X"D2",X"C9",
		X"00",X"60",X"40",X"E7",X"D2",X"C5",X"18",X"50",X"0D",X"49",X"20",X"F0",X"09",X"40",X"20",X"D3",
		X"40",X"52",X"D3",X"40",X"F2",X"D3",X"60",X"C5",X"19",X"49",X"3F",X"A9",X"3F",X"90",X"30",X"C5",
		X"18",X"49",X"A0",X"B0",X"2A",X"C5",X"7A",X"49",X"68",X"B0",X"24",X"C9",X"80",X"85",X"7A",X"C9",
		X"03",X"85",X"96",X"C5",X"18",X"09",X"20",X"85",X"18",X"C9",X"00",X"85",X"8F",X"85",X"90",X"C9",
		X"13",X"85",X"F0",X"40",X"44",X"DA",X"C2",X"3F",X"C9",X"00",X"95",X"3A",X"AA",X"10",X"FB",X"60",
		X"C5",X"7A",X"49",X"10",X"B0",X"2B",X"C2",X"00",X"C5",X"7C",X"F0",X"0D",X"A9",X"7C",X"F0",X"09",
		X"E8",X"A6",X"7C",X"D0",X"04",X"E6",X"7C",X"E6",X"7C",X"C5",X"7B",X"A9",X"5C",X"F0",X"09",X"E8",
		X"A6",X"7B",X"D0",X"04",X"E6",X"7B",X"E6",X"7B",X"8A",X"B0",X"06",X"C5",X"36",X"09",X"80",X"85",
		X"36",X"60",X"C5",X"36",X"49",X"40",X"B0",X"33",X"C5",X"24",X"49",X"3F",X"B0",X"52",X"58",X"C9",
		X"7C",X"E5",X"23",X"90",X"4B",X"85",X"4C",X"85",X"5C",X"C9",X"39",X"85",X"4B",X"C9",X"4C",X"85",
		X"5B",X"C5",X"22",X"49",X"03",X"0A",X"18",X"69",X"7D",X"85",X"4F",X"85",X"5F",X"E6",X"5F",X"C9",
		X"C0",X"85",X"4A",X"85",X"5A",X"C5",X"36",X"09",X"40",X"85",X"36",X"C5",X"36",X"49",X"20",X"B0",
		X"1F",X"C5",X"4C",X"18",X"65",X"96",X"85",X"4C",X"85",X"5C",X"A9",X"7C",X"90",X"12",X"C9",X"7C",
		X"85",X"4C",X"85",X"5C",X"E6",X"22",X"C5",X"36",X"09",X"20",X"85",X"36",X"C9",X"00",X"85",X"96",
		X"60",X"C5",X"18",X"49",X"04",X"F0",X"1A",X"C5",X"22",X"49",X"03",X"0A",X"0A",X"0A",X"CA",X"C0",
		X"07",X"DD",X"D2",X"D3",X"99",X"08",X"5C",X"E8",X"88",X"10",X"F6",X"C5",X"36",X"49",X"DF",X"85",
		X"36",X"60",X"00",X"9B",X"7F",X"49",X"00",X"00",X"E2",X"FF",X"00",X"56",X"1C",X"49",X"DD",X"C7",
		X"50",X"FF",X"00",X"DD",X"3F",X"49",X"41",X"83",X"E1",X"FF",X"00",X"2F",X"7F",X"49",X"FF",X"C0",
		X"F0",X"FF",X"C5",X"36",X"A9",X"E0",X"B0",X"22",X"40",X"45",X"E7",X"C5",X"18",X"49",X"DF",X"85",
		X"18",X"C5",X"36",X"49",X"20",X"85",X"36",X"C9",X"00",X"85",X"35",X"85",X"7A",X"85",X"4A",X"85",
		X"5A",X"C5",X"18",X"09",X"04",X"85",X"18",X"40",X"B1",X"D3",X"60",X"8A",X"18",X"69",X"3A",X"85",
		X"E1",X"C9",X"00",X"85",X"E2",X"C0",X"0F",X"D1",X"E1",X"99",X"97",X"00",X"88",X"10",X"F8",X"60",
		X"C0",X"0F",X"D9",X"97",X"00",X"91",X"E1",X"88",X"10",X"F8",X"60",X"C9",X"00",X"85",X"CB",X"85",
		X"CC",X"85",X"CA",X"26",X"C7",X"90",X"0D",X"18",X"C5",X"CB",X"65",X"C9",X"85",X"CB",X"C5",X"CC",
		X"65",X"CA",X"85",X"CC",X"06",X"C9",X"46",X"CA",X"C5",X"C7",X"B0",X"E7",X"60",X"C0",X"04",X"E6",
		X"13",X"E6",X"15",X"66",X"14",X"66",X"15",X"66",X"16",X"D0",X"06",X"C5",X"15",X"65",X"13",X"85",
		X"15",X"88",X"B0",X"EF",X"C5",X"14",X"65",X"16",X"85",X"16",X"65",X"15",X"85",X"17",X"60",X"C4",
		X"24",X"C5",X"25",X"85",X"28",X"C5",X"23",X"18",X"65",X"39",X"90",X"11",X"A8",X"C5",X"18",X"49",
		X"40",X"F0",X"0A",X"C5",X"28",X"F0",X"06",X"A0",X"40",X"90",X"02",X"C0",X"3F",X"C9",X"F5",X"85",
		X"A7",X"C9",X"D6",X"18",X"65",X"28",X"85",X"A8",X"D1",X"A7",X"60",X"C9",X"0C",X"8D",X"12",X"04",
		X"8D",X"32",X"04",X"C9",X"00",X"8D",X"0B",X"04",X"8D",X"2B",X"04",X"C9",X"FF",X"8D",X"0C",X"04",
		X"8D",X"2C",X"04",X"C9",X"01",X"8D",X"0D",X"04",X"8D",X"2D",X"04",X"C5",X"07",X"B0",X"07",X"85",
		X"96",X"C9",X"7F",X"8D",X"0C",X"04",X"60",X"C5",X"2C",X"F0",X"04",X"49",X"10",X"F0",X"3E",X"C5",
		X"23",X"58",X"E5",X"96",X"85",X"23",X"D0",X"35",X"A6",X"24",X"C5",X"24",X"A9",X"FF",X"B0",X"12",
		X"C5",X"25",X"29",X"01",X"85",X"25",X"F0",X"0A",X"C9",X"3F",X"85",X"24",X"C5",X"18",X"09",X"40",
		X"85",X"18",X"C5",X"24",X"28",X"29",X"FF",X"85",X"19",X"68",X"F0",X"11",X"49",X"3F",X"A9",X"04",
		X"D0",X"06",X"C5",X"35",X"09",X"40",X"85",X"35",X"C9",X"00",X"40",X"C5",X"DB",X"60",X"E6",X"D5",
		X"B0",X"02",X"E6",X"D6",X"E6",X"DF",X"B0",X"02",X"E6",X"E0",X"C5",X"31",X"B0",X"02",X"A6",X"32",
		X"A6",X"31",X"60",X"C5",X"2B",X"49",X"F7",X"85",X"2B",X"C9",X"00",X"85",X"39",X"C9",X"02",X"85",
		X"CD",X"C4",X"24",X"C5",X"23",X"18",X"65",X"2A",X"90",X"01",X"A8",X"84",X"24",X"84",X"D2",X"98",
		X"49",X"3F",X"F0",X"69",X"A9",X"3F",X"F0",X"65",X"40",X"7F",X"D4",X"85",X"8C",X"40",X"D7",X"D5",
		X"C4",X"D2",X"C5",X"D4",X"B0",X"20",X"C2",X"03",X"A6",X"CD",X"E6",X"D2",X"C4",X"D2",X"98",X"49",
		X"3F",X"A9",X"3F",X"F0",X"48",X"40",X"81",X"D4",X"85",X"8C",X"40",X"D7",X"D5",X"C5",X"D4",X"F0",
		X"E5",X"AA",X"B0",X"E4",X"F0",X"37",X"C9",X"FD",X"85",X"D3",X"C2",X"00",X"A6",X"D2",X"C4",X"D2",
		X"98",X"49",X"3F",X"A9",X"3F",X"F0",X"26",X"40",X"81",X"D4",X"85",X"8C",X"40",X"D7",X"D5",X"E6",
		X"D3",X"C5",X"D4",X"B0",X"08",X"C2",X"04",X"C9",X"05",X"85",X"CD",X"B0",X"BB",X"E8",X"E0",X"03",
		X"90",X"DA",X"C5",X"D3",X"50",X"07",X"C5",X"CD",X"58",X"E5",X"D3",X"85",X"CD",X"C9",X"00",X"85",
		X"23",X"85",X"26",X"C5",X"24",X"58",X"E5",X"CD",X"85",X"24",X"85",X"27",X"C9",X"03",X"85",X"96",
		X"C5",X"07",X"B0",X"02",X"85",X"96",X"60",X"C9",X"00",X"85",X"D4",X"C5",X"8C",X"A9",X"04",X"F0",
		X"0E",X"A9",X"0B",X"F0",X"0A",X"A9",X"0C",X"F0",X"06",X"A9",X"0E",X"D0",X"02",X"E6",X"D4",X"60",
		X"C9",X"00",X"85",X"31",X"C9",X"02",X"85",X"32",X"E6",X"23",X"B0",X"02",X"E6",X"24",X"40",X"19",
		X"D6",X"C5",X"31",X"B0",X"02",X"A6",X"32",X"A6",X"31",X"C5",X"32",X"05",X"31",X"B0",X"E9",X"C5",
		X"2B",X"09",X"08",X"85",X"2B",X"8D",X"00",X"54",X"60",X"C5",X"25",X"85",X"28",X"58",X"C5",X"23",
		X"E5",X"26",X"CA",X"F0",X"48",X"50",X"23",X"18",X"C5",X"26",X"69",X"80",X"85",X"D9",X"C5",X"27",
		X"69",X"01",X"85",X"DA",X"90",X"06",X"C5",X"25",X"29",X"01",X"85",X"28",X"40",X"8B",X"D6",X"E6",
		X"D9",X"B0",X"02",X"E6",X"DA",X"AA",X"B0",X"F4",X"F0",X"23",X"58",X"C5",X"26",X"E9",X"80",X"85",
		X"D9",X"C5",X"27",X"E9",X"00",X"85",X"DA",X"D0",X"06",X"C5",X"25",X"29",X"01",X"85",X"28",X"40",
		X"8B",X"D6",X"C5",X"D9",X"B0",X"02",X"A6",X"DA",X"A6",X"D9",X"E8",X"B0",X"F2",X"C5",X"24",X"85",
		X"27",X"0A",X"49",X"02",X"09",X"01",X"85",X"CD",X"C5",X"2B",X"49",X"F8",X"05",X"CD",X"85",X"2B",
		X"8D",X"00",X"54",X"C5",X"23",X"8D",X"00",X"58",X"85",X"26",X"60",X"C4",X"DA",X"40",X"9D",X"D4",
		X"85",X"D6",X"C5",X"D9",X"26",X"D6",X"6A",X"18",X"69",X"9D",X"85",X"D5",X"C5",X"D6",X"69",X"EE",
		X"85",X"D6",X"C5",X"D9",X"49",X"0F",X"C8",X"C5",X"D9",X"2A",X"49",X"78",X"18",X"19",X"E5",X"D6",
		X"69",X"00",X"85",X"DF",X"C5",X"DA",X"49",X"01",X"69",X"F7",X"85",X"E0",X"C5",X"D9",X"2A",X"C0",
		X"00",X"D1",X"D5",X"90",X"04",X"0A",X"0A",X"0A",X"0A",X"49",X"F0",X"85",X"CD",X"D1",X"DF",X"49",
		X"0F",X"05",X"CD",X"28",X"58",X"C5",X"DF",X"E9",X"00",X"85",X"DF",X"C5",X"E0",X"E9",X"A7",X"85",
		X"E0",X"68",X"91",X"DF",X"60",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"80",X"81",X"82",
		X"83",X"84",X"85",X"86",X"87",X"00",X"00",X"0B",X"04",X"03",X"06",X"0F",X"05",X"06",X"05",X"06",
		X"05",X"06",X"0F",X"05",X"0A",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"08",X"0B",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"04",X"03",X"01",X"0A",X"0C",X"0C",X"09",X"09",X"09",X"0C",X"0C",X"0C",X"08",
		X"0D",X"07",X"07",X"06",X"05",X"06",X"0F",X"0F",X"0F",X"05",X"0D",X"0B",X"0E",X"0E",X"0E",X"0E",
		X"04",X"03",X"01",X"06",X"05",X"00",X"00",X"0B",X"04",X"03",X"06",X"05",X"01",X"01",X"02",X"06",
		X"05",X"06",X"0F",X"0F",X"05",X"0A",X"09",X"09",X"0C",X"09",X"0C",X"09",X"0C",X"08",X"0D",X"0D",
		X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"01",X"0A",X"09",X"08",X"00",X"06",X"0F",X"05",X"06",X"0F",
		X"0F",X"05",X"07",X"07",X"0A",X"08",X"0B",X"0E",X"0E",X"04",X"03",X"02",X"02",X"02",X"0A",X"0C",
		X"09",X"09",X"0C",X"08",X"00",X"00",X"00",X"0E",X"02",X"02",X"0D",X"0D",X"01",X"01",X"0A",X"09",
		X"09",X"03",X"06",X"04",X"03",X"06",X"0F",X"0F",X"0F",X"0F",X"05",X"0A",X"0C",X"08",X"0B",X"0E",
		X"0E",X"07",X"07",X"06",X"05",X"07",X"00",X"00",X"0D",X"02",X"0D",X"02",X"0A",X"0C",X"09",X"09",
		X"08",X"0D",X"0D",X"06",X"0F",X"04",X"03",X"01",X"06",X"0E",X"0E",X"00",X"0E",X"00",X"0B",X"00",
		X"02",X"02",X"02",X"02",X"07",X"00",X"00",X"0C",X"09",X"0C",X"0C",X"08",X"00",X"00",X"0B",X"04",
		X"03",X"06",X"0F",X"05",X"0A",X"09",X"09",X"09",X"09",X"09",X"09",X"0C",X"09",X"0C",X"09",X"08",
		X"0D",X"0D",X"06",X"0F",X"0F",X"05",X"06",X"05",X"06",X"04",X"03",X"00",X"0B",X"0E",X"04",X"03",
		X"06",X"0F",X"05",X"0D",X"0D",X"02",X"02",X"0D",X"0D",X"0B",X"0E",X"04",X"03",X"06",X"0F",X"05",
		X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"0C",X"09",X"0C",X"0C",X"08",X"00",X"00",X"0B",X"04",
		X"03",X"06",X"0F",X"05",X"0A",X"09",X"09",X"09",X"09",X"09",X"09",X"0C",X"09",X"0C",X"09",X"08",
		X"0D",X"0D",X"00",X"00",X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"0B",X"0E",X"04",X"03",
		X"06",X"0F",X"05",X"0D",X"0D",X"00",X"00",X"00",X"00",X"0B",X"0E",X"04",X"03",X"06",X"0F",X"05",
		X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"0B",X"04",X"03",X"0D",X"02",X"02",X"02",X"01",X"01",
		X"0A",X"09",X"09",X"09",X"0C",X"08",X"0D",X"07",X"07",X"0A",X"09",X"08",X"07",X"06",X"05",X"02",
		X"02",X"02",X"02",X"01",X"00",X"00",X"0D",X"0D",X"0D",X"01",X"07",X"07",X"0A",X"0C",X"09",X"08",
		X"00",X"00",X"00",X"00",X"0B",X"0E",X"0E",X"04",X"03",X"01",X"07",X"07",X"0A",X"08",X"0D",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"04",X"03",X"01",X"0A",X"0C",X"09",X"08",
		X"00",X"00",X"00",X"02",X"0B",X"0E",X"0E",X"04",X"03",X"01",X"07",X"07",X"0A",X"08",X"0D",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",X"01",X"07",X"07",X"0A",X"0C",X"09",X"08",
		X"00",X"00",X"00",X"00",X"01",X"02",X"0B",X"04",X"03",X"01",X"07",X"07",X"0A",X"08",X"0D",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0C",X"08",X"07",X"00",X"07",X"00",X"07",X"00",X"0D",
		X"0D",X"0D",X"0B",X"04",X"03",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",
		X"0B",X"04",X"03",X"01",X"01",X"01",X"01",X"01",X"07",X"07",X"07",X"0A",X"0C",X"09",X"09",X"09",
		X"09",X"09",X"09",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"C6",X"09",X"CD",X"00",X"10",X"49",X"40",X"B0",X"01",X"CA",X"DD",
		X"02",X"10",X"29",X"FF",X"85",X"37",X"60",X"C2",X"00",X"2C",X"C3",X"D9",X"26",X"40",X"2C",X"6F",
		X"6A",X"FE",X"2C",X"40",X"62",X"63",X"20",X"6D",X"5D",X"69",X"6C",X"5F",X"FF",X"C2",X"02",X"2C",
		X"C3",X"D9",X"38",X"40",X"2D",X"6F",X"6A",X"FF",X"C2",X"04",X"2C",X"C3",X"D9",X"83",X"43",X"6A",
		X"5B",X"6E",X"6E",X"5F",X"6C",X"68",X"FF",X"C2",X"06",X"2C",X"C3",X"D9",X"C7",X"41",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"20",X"20",X"47",X"45",X"54",X"20",X"52",X"45",X"41",X"44",X"59",
		X"FF",X"C2",X"08",X"2C",X"C3",X"D9",X"C7",X"41",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"20",
		X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"FF",X"C2",X"0A",X"2C",X"C3",X"D9",
		X"09",X"42",X"54",X"49",X"4D",X"45",X"FF",X"C2",X"0C",X"2C",X"C3",X"D9",X"0B",X"42",X"47",X"41",
		X"4D",X"45",X"20",X"20",X"4F",X"56",X"45",X"52",X"FF",X"C2",X"0E",X"2C",X"C3",X"D9",X"C5",X"42",
		X"73",X"69",X"6F",X"6C",X"20",X"5D",X"5B",X"6C",X"20",X"5D",X"5B",X"68",X"20",X"69",X"68",X"66",
		X"73",X"20",X"64",X"6F",X"67",X"6A",X"FE",X"03",X"43",X"71",X"62",X"5F",X"68",X"20",X"6D",X"6A",
		X"5F",X"5F",X"5E",X"20",X"63",X"6D",X"20",X"69",X"70",X"5F",X"6C",X"20",X"36",X"35",X"35",X"67",
		X"6A",X"62",X"FF",X"DD",X"06",X"DA",X"85",X"D5",X"DD",X"07",X"DA",X"85",X"D6",X"C0",X"FF",X"A8",
		X"D1",X"D5",X"85",X"D9",X"85",X"DB",X"A8",X"D1",X"D5",X"85",X"DA",X"09",X"04",X"85",X"DC",X"A8",
		X"98",X"18",X"65",X"D5",X"85",X"D5",X"C9",X"00",X"65",X"D6",X"85",X"D6",X"C0",X"00",X"D1",X"D5",
		X"A9",X"FF",X"F0",X"11",X"A9",X"FE",X"F0",X"D7",X"58",X"E9",X"20",X"91",X"D9",X"C9",X"00",X"91",
		X"DB",X"A8",X"2C",X"EE",X"D9",X"60",X"0C",X"D9",X"22",X"D9",X"2D",X"D9",X"3C",X"D9",X"56",X"D9",
		X"70",X"D9",X"7C",X"D9",X"8E",X"D9",X"C5",X"18",X"49",X"08",X"B0",X"20",X"C9",X"80",X"40",X"44",
		X"DA",X"40",X"37",X"D9",X"C5",X"09",X"18",X"69",X"16",X"8D",X"CE",X"41",X"C2",X"40",X"40",X"A6",
		X"DC",X"C2",X"20",X"40",X"EA",X"C2",X"C5",X"18",X"09",X"08",X"85",X"18",X"60",X"40",X"51",X"D9",
		X"40",X"24",X"DA",X"60",X"28",X"C5",X"07",X"F0",X"05",X"68",X"28",X"8D",X"02",X"10",X"68",X"60",
		X"C9",X"61",X"85",X"D9",X"C9",X"40",X"85",X"DA",X"C2",X"00",X"C0",X"00",X"DD",X"B3",X"DA",X"91",
		X"D9",X"E8",X"A8",X"DD",X"B3",X"DA",X"F0",X"02",X"91",X"D9",X"A0",X"08",X"90",X"F4",X"E8",X"A8",
		X"DD",X"B3",X"DA",X"91",X"D9",X"E8",X"C5",X"D9",X"18",X"69",X"20",X"85",X"D9",X"A9",X"C1",X"90",
		X"D9",X"E6",X"D9",X"C2",X"00",X"C0",X"00",X"DD",X"B3",X"DA",X"91",X"D9",X"E8",X"A8",X"DD",X"B3",
		X"DA",X"F0",X"02",X"91",X"D9",X"A0",X"03",X"90",X"F4",X"E8",X"A8",X"DD",X"B3",X"DA",X"91",X"D9",
		X"E8",X"C5",X"D9",X"18",X"69",X"20",X"85",X"D9",X"90",X"02",X"E6",X"DA",X"C5",X"D9",X"A9",X"22",
		X"B0",X"D3",X"60",X"6A",X"6D",X"6B",X"6E",X"00",X"6C",X"68",X"6F",X"69",X"40",X"28",X"D9",X"C5",
		X"22",X"18",X"69",X"01",X"85",X"CD",X"C9",X"00",X"85",X"CE",X"C5",X"CD",X"58",X"E9",X"0A",X"90",
		X"0D",X"85",X"CD",X"F8",X"C5",X"CE",X"69",X"00",X"85",X"CE",X"B8",X"2C",X"CA",X"DA",X"06",X"CE",
		X"06",X"CE",X"06",X"CE",X"06",X"CE",X"C5",X"CE",X"05",X"CD",X"85",X"F1",X"C2",X"08",X"40",X"17",
		X"DB",X"C2",X"F1",X"40",X"79",X"DB",X"60",X"C4",X"1A",X"A0",X"05",X"90",X"02",X"C0",X"05",X"A0",
		X"00",X"F0",X"0F",X"C9",X"63",X"85",X"CD",X"C9",X"43",X"85",X"CE",X"C9",X"73",X"91",X"CD",X"88",
		X"B0",X"F9",X"60",X"21",X"40",X"3A",X"40",X"DD",X"29",X"DB",X"85",X"DD",X"DD",X"2A",X"DB",X"85",
		X"DE",X"C9",X"01",X"85",X"CD",X"0A",X"85",X"CE",X"60",X"53",X"42",X"23",X"40",X"E3",X"40",X"BB",
		X"43",X"A6",X"43",X"C5",X"12",X"A9",X"02",X"90",X"1E",X"C5",X"09",X"29",X"01",X"49",X"01",X"28",
		X"CA",X"DC",X"DF",X"DC",X"C2",X"00",X"D9",X"03",X"04",X"95",X"F1",X"A8",X"E8",X"E0",X"03",X"B0",
		X"F5",X"C2",X"F3",X"68",X"40",X"67",X"DB",X"40",X"61",X"DB",X"60",X"C2",X"0C",X"C0",X"02",X"B0",
		X"07",X"C2",X"1D",X"C5",X"09",X"49",X"01",X"C8",X"D9",X"91",X"DB",X"85",X"DD",X"C9",X"40",X"85",
		X"DE",X"C9",X"03",X"85",X"CD",X"C9",X"05",X"85",X"CE",X"C9",X"0B",X"85",X"CF",X"D5",X"00",X"28",
		X"2A",X"2A",X"2A",X"2A",X"40",X"94",X"DB",X"68",X"40",X"94",X"DB",X"AA",X"A6",X"CD",X"B0",X"ED",
		X"60",X"44",X"56",X"4D",X"49",X"0F",X"B0",X"0E",X"C4",X"CE",X"F0",X"0E",X"A6",X"CE",X"B0",X"0D",
		X"C0",X"00",X"84",X"CE",X"F0",X"04",X"C4",X"CE",X"B0",X"F6",X"18",X"65",X"CF",X"C0",X"00",X"91",
		X"DD",X"E6",X"DD",X"B0",X"02",X"E6",X"DE",X"60",X"C4",X"96",X"F0",X"08",X"C9",X"00",X"40",X"C5",
		X"DB",X"88",X"B0",X"F8",X"60",X"C8",X"F8",X"C5",X"1B",X"18",X"79",X"DF",X"DB",X"85",X"1B",X"C5",
		X"1C",X"79",X"E0",X"DB",X"85",X"1C",X"C5",X"1D",X"79",X"E1",X"DB",X"85",X"1D",X"B8",X"60",X"08",
		X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"05",X"00",X"00",X"10",
		X"00",X"F8",X"C5",X"05",X"18",X"69",X"01",X"85",X"05",X"B8",X"60",X"F8",X"C5",X"05",X"58",X"E9",
		X"01",X"85",X"05",X"B8",X"60",X"F8",X"C5",X"1A",X"58",X"E9",X"01",X"85",X"1A",X"B8",X"60",X"F8",
		X"58",X"C5",X"1B",X"E5",X"0A",X"C5",X"1C",X"E5",X"0B",X"C5",X"1D",X"E5",X"0C",X"90",X"09",X"C2",
		X"02",X"D5",X"1B",X"95",X"0A",X"AA",X"10",X"F9",X"60",X"F8",X"C5",X"18",X"2A",X"D0",X"46",X"CD",
		X"01",X"10",X"49",X"06",X"A9",X"04",X"D0",X"17",X"58",X"C5",X"0D",X"E5",X"1B",X"C5",X"0E",X"E5",
		X"1C",X"C5",X"0F",X"E5",X"1D",X"D0",X"2E",X"C5",X"18",X"09",X"01",X"85",X"18",X"B0",X"1A",X"C0",
		X"00",X"C5",X"1D",X"58",X"E5",X"0F",X"90",X"1D",X"A8",X"A4",X"1E",X"90",X"F6",X"F0",X"F4",X"28",
		X"40",X"69",X"DC",X"84",X"1E",X"68",X"2C",X"53",X"DC",X"C5",X"1A",X"18",X"69",X"01",X"85",X"1A",
		X"C9",X"08",X"40",X"44",X"DA",X"B8",X"60",X"CD",X"01",X"10",X"29",X"FF",X"28",X"49",X"01",X"CA",
		X"DD",X"9C",X"DC",X"8D",X"02",X"04",X"8D",X"22",X"04",X"68",X"49",X"06",X"CA",X"C9",X"00",X"85",
		X"0D",X"DD",X"9E",X"DC",X"85",X"0E",X"DD",X"9F",X"DC",X"85",X"0F",X"60",X"03",X"05",X"00",X"03",
		X"00",X"07",X"00",X"02",X"00",X"03",X"CD",X"00",X"10",X"10",X"FB",X"CD",X"00",X"10",X"50",X"FB",
		X"40",X"18",X"EB",X"AA",X"B0",X"F0",X"60",X"C4",X"09",X"DE",X"DF",X"DC",X"C0",X"00",X"DD",X"00",
		X"04",X"99",X"18",X"00",X"E8",X"A8",X"A0",X"18",X"90",X"F4",X"60",X"C4",X"09",X"DE",X"DF",X"DC",
		X"C0",X"00",X"D9",X"18",X"00",X"9D",X"00",X"04",X"E8",X"A8",X"A0",X"18",X"90",X"F4",X"60",X"00",
		X"20",X"C9",X"00",X"CA",X"85",X"9E",X"85",X"A0",X"85",X"A1",X"C9",X"45",X"85",X"9F",X"C0",X"02",
		X"D9",X"1B",X"00",X"95",X"A2",X"E8",X"88",X"10",X"F7",X"C9",X"00",X"85",X"99",X"8D",X"00",X"54",
		X"C9",X"00",X"85",X"9A",X"C9",X"05",X"85",X"9B",X"C2",X"01",X"C0",X"02",X"58",X"C5",X"A4",X"F1",
		X"9A",X"88",X"C5",X"A3",X"F1",X"9A",X"88",X"C5",X"A2",X"F1",X"9A",X"D0",X"19",X"C5",X"9A",X"18",
		X"69",X"03",X"85",X"9A",X"C5",X"9B",X"69",X"00",X"85",X"9B",X"8A",X"F8",X"18",X"69",X"01",X"CA",
		X"B8",X"E0",X"01",X"B0",X"D5",X"60",X"86",X"A7",X"86",X"D1",X"40",X"58",X"DD",X"40",X"CF",X"DD",
		X"40",X"A2",X"DE",X"40",X"51",X"DE",X"40",X"FC",X"DE",X"40",X"69",X"DF",X"40",X"6B",X"D9",X"40",
		X"95",X"DF",X"40",X"A9",X"DF",X"2C",X"40",X"DD",X"C9",X"29",X"85",X"CD",X"C9",X"06",X"85",X"CE",
		X"C9",X"2C",X"85",X"9A",X"C9",X"06",X"85",X"9B",X"40",X"9B",X"DD",X"C0",X"02",X"D9",X"A2",X"00",
		X"91",X"CD",X"88",X"10",X"F8",X"C2",X"01",X"D5",X"CD",X"95",X"CF",X"AA",X"10",X"F9",X"C9",X"69",
		X"85",X"CD",X"C9",X"07",X"85",X"CE",X"C9",X"6C",X"85",X"9A",X"C9",X"07",X"85",X"9B",X"40",X"9B",
		X"DD",X"C0",X"02",X"C9",X"00",X"91",X"CD",X"88",X"10",X"F9",X"60",X"C2",X"00",X"C0",X"02",X"D1",
		X"CD",X"91",X"9A",X"88",X"10",X"F9",X"E4",X"A7",X"F0",X"24",X"8A",X"F8",X"58",X"E9",X"01",X"CA",
		X"B8",X"C5",X"CD",X"58",X"E9",X"03",X"85",X"CD",X"C5",X"CE",X"E9",X"00",X"85",X"CE",X"C5",X"9A",
		X"58",X"E9",X"03",X"85",X"9A",X"C5",X"9B",X"E9",X"00",X"85",X"9B",X"2C",X"9D",X"DD",X"60",X"C5",
		X"A7",X"B0",X"09",X"C0",X"05",X"C9",X"0C",X"85",X"97",X"40",X"01",X"DE",X"A9",X"06",X"D0",X"0B",
		X"C8",X"CA",X"D9",X"DE",X"DE",X"85",X"97",X"E8",X"40",X"01",X"DE",X"A9",X"99",X"B0",X"09",X"C0",
		X"04",X"C9",X"09",X"85",X"97",X"40",X"01",X"DE",X"C0",X"03",X"C9",X"06",X"85",X"97",X"40",X"01",
		X"DE",X"88",X"F0",X"26",X"C5",X"A7",X"F8",X"58",X"E9",X"01",X"85",X"A7",X"B8",X"C5",X"CD",X"58",
		X"E9",X"03",X"85",X"CD",X"C5",X"CE",X"E9",X"00",X"85",X"CE",X"C5",X"CF",X"58",X"E9",X"03",X"85",
		X"CF",X"C5",X"D0",X"E9",X"00",X"85",X"D0",X"2C",X"01",X"DE",X"C0",X"00",X"C5",X"A7",X"99",X"A0",
		X"07",X"F8",X"C5",X"A7",X"18",X"69",X"01",X"85",X"A7",X"B8",X"A8",X"A0",X"05",X"B0",X"ED",X"C0",
		X"0E",X"D1",X"CD",X"99",X"90",X"07",X"D1",X"CF",X"99",X"80",X"07",X"88",X"10",X"F3",X"68",X"68",
		X"60",X"98",X"28",X"C2",X"00",X"C0",X"00",X"DD",X"A0",X"07",X"A5",X"D1",X"B0",X"05",X"CD",X"0F",
		X"42",X"F0",X"34",X"DD",X"A0",X"07",X"B0",X"0F",X"C9",X"16",X"99",X"D3",X"48",X"C9",X"15",X"99",
		X"F3",X"48",X"99",X"13",X"49",X"B0",X"16",X"28",X"2A",X"2A",X"2A",X"2A",X"F0",X"06",X"18",X"69",
		X"15",X"99",X"F3",X"48",X"68",X"49",X"0F",X"18",X"69",X"15",X"99",X"13",X"49",X"A8",X"A8",X"E8",
		X"E0",X"05",X"B0",X"C3",X"68",X"C8",X"60",X"99",X"F3",X"48",X"99",X"13",X"49",X"99",X"D3",X"48",
		X"F0",X"EB",X"C9",X"80",X"85",X"9A",X"C9",X"40",X"85",X"9B",X"C2",X"3B",X"C0",X"06",X"8A",X"91",
		X"9A",X"E8",X"E0",X"59",X"F0",X"16",X"A8",X"A8",X"A0",X"1A",X"B0",X"F2",X"C5",X"9A",X"18",X"69",
		X"60",X"85",X"9A",X"C5",X"9B",X"69",X"00",X"85",X"9B",X"2C",X"AC",X"DE",X"C2",X"0B",X"DD",X"E4",
		X"DE",X"9D",X"A6",X"41",X"DD",X"F0",X"DE",X"9D",X"4A",X"42",X"AA",X"10",X"F1",X"60",X"00",X"00",
		X"03",X"06",X"09",X"0C",X"4D",X"4A",X"3B",X"00",X"4C",X"4F",X"3C",X"00",X"3F",X"48",X"3E",X"00",
		X"2E",X"21",X"2D",X"25",X"00",X"00",X"00",X"33",X"23",X"2F",X"32",X"25",X"C9",X"42",X"85",X"9B",
		X"C9",X"70",X"85",X"9A",X"C2",X"00",X"C0",X"00",X"84",X"A5",X"DD",X"80",X"07",X"28",X"2A",X"2A",
		X"2A",X"2A",X"28",X"B0",X"08",X"C5",X"A5",X"50",X"04",X"68",X"2C",X"27",X"DF",X"C9",X"80",X"85",
		X"A5",X"68",X"18",X"69",X"15",X"91",X"9A",X"A8",X"68",X"49",X"0F",X"28",X"B0",X"08",X"C5",X"A5",
		X"50",X"04",X"68",X"2C",X"40",X"DF",X"C9",X"80",X"85",X"A5",X"68",X"18",X"69",X"15",X"91",X"9A",
		X"E8",X"A8",X"A0",X"06",X"B0",X"C4",X"C5",X"A5",X"50",X"06",X"C0",X"05",X"C9",X"15",X"91",X"9A",
		X"E0",X"0F",X"F0",X"14",X"C5",X"9A",X"18",X"69",X"40",X"85",X"9A",X"C5",X"9B",X"69",X"00",X"85",
		X"9B",X"C9",X"00",X"85",X"A5",X"2C",X"06",X"DF",X"60",X"C9",X"42",X"85",X"9B",X"C9",X"6A",X"85",
		X"9A",X"C2",X"00",X"C0",X"00",X"DD",X"90",X"07",X"91",X"9A",X"A8",X"E8",X"E0",X"0F",X"F0",X"14",
		X"A0",X"03",X"B0",X"F1",X"C5",X"9A",X"18",X"69",X"40",X"85",X"9A",X"C5",X"9B",X"69",X"00",X"85",
		X"9B",X"2C",X"73",X"DF",X"60",X"C9",X"00",X"85",X"98",X"C2",X"03",X"DD",X"A5",X"DF",X"9D",X"00",
		X"48",X"AA",X"10",X"F7",X"60",X"01",X"7A",X"C4",X"28",X"40",X"8D",X"E1",X"C6",X"09",X"CD",X"00",
		X"10",X"49",X"40",X"B0",X"02",X"C2",X"00",X"DD",X"02",X"10",X"29",X"FF",X"28",X"49",X"10",X"A5",
		X"A0",X"85",X"A0",X"F0",X"62",X"90",X"60",X"68",X"C5",X"98",X"A9",X"1E",X"90",X"1E",X"58",X"E9",
		X"1E",X"0A",X"CA",X"DD",X"E0",X"DF",X"85",X"9A",X"DD",X"E1",X"DF",X"85",X"9B",X"6C",X"9A",X"00",
		X"27",X"E1",X"27",X"E1",X"0D",X"E1",X"0D",X"E1",X"41",X"E1",X"41",X"E1",X"C6",X"97",X"C4",X"99",
		X"A0",X"03",X"B0",X"03",X"2C",X"41",X"E1",X"C9",X"03",X"8D",X"02",X"10",X"C0",X"00",X"CD",X"02",
		X"48",X"29",X"FF",X"85",X"9A",X"CD",X"03",X"48",X"58",X"E9",X"04",X"85",X"9B",X"2A",X"2A",X"2A",
		X"2A",X"66",X"9A",X"2A",X"66",X"9A",X"2A",X"66",X"9A",X"18",X"69",X"40",X"85",X"9B",X"A6",X"9A",
		X"C9",X"00",X"91",X"9A",X"2C",X"83",X"E0",X"68",X"49",X"0F",X"CA",X"DD",X"46",X"E0",X"A5",X"A1",
		X"85",X"A1",X"F0",X"0F",X"18",X"65",X"98",X"10",X"02",X"C9",X"00",X"A9",X"24",X"90",X"02",X"C9",
		X"23",X"85",X"98",X"2C",X"58",X"E0",X"00",X"01",X"FF",X"00",X"F6",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C5",X"98",X"58",X"E9",X"0A",X"A8",
		X"D0",X"FB",X"69",X"0A",X"88",X"CA",X"DD",X"75",X"E0",X"8D",X"02",X"48",X"D9",X"7F",X"E0",X"8D",
		X"03",X"48",X"2C",X"A9",X"DF",X"C4",X"B4",X"A4",X"94",X"84",X"74",X"64",X"54",X"44",X"34",X"28",
		X"40",X"58",X"70",X"40",X"E3",X"E0",X"C0",X"08",X"40",X"8D",X"E1",X"AE",X"03",X"48",X"88",X"B0",
		X"F7",X"C9",X"00",X"EE",X"01",X"48",X"40",X"8D",X"E1",X"C2",X"04",X"CD",X"02",X"48",X"A5",X"9A",
		X"F0",X"0C",X"90",X"02",X"C2",X"FC",X"8A",X"18",X"6D",X"02",X"48",X"8D",X"02",X"48",X"CD",X"03",
		X"48",X"A5",X"9B",X"D0",X"0C",X"CD",X"03",X"48",X"18",X"69",X"02",X"8D",X"03",X"48",X"2C",X"96",
		X"E0",X"C9",X"04",X"8D",X"02",X"10",X"AE",X"01",X"48",X"C0",X"08",X"40",X"8D",X"E1",X"EE",X"03",
		X"48",X"88",X"B0",X"F7",X"C6",X"97",X"C5",X"98",X"18",X"69",X"3B",X"9D",X"90",X"07",X"E6",X"97",
		X"E6",X"99",X"60",X"C0",X"00",X"C5",X"97",X"A9",X"03",X"90",X"06",X"A8",X"E9",X"03",X"2C",X"E7",
		X"E0",X"CA",X"DD",X"FD",X"E0",X"85",X"9A",X"D9",X"00",X"E1",X"85",X"9B",X"60",X"A4",X"9C",X"94",
		X"98",X"A8",X"B8",X"C8",X"D8",X"D0",X"D0",X"D0",X"98",X"A8",X"B8",X"C8",X"D8",X"C6",X"97",X"C4",
		X"99",X"88",X"50",X"10",X"C9",X"09",X"8D",X"02",X"10",X"AA",X"C9",X"00",X"9D",X"90",X"07",X"A6",
		X"99",X"A6",X"97",X"60",X"2C",X"A9",X"DF",X"C6",X"97",X"C4",X"99",X"A0",X"03",X"F0",X"12",X"C9",
		X"09",X"8D",X"02",X"10",X"C9",X"00",X"9D",X"90",X"07",X"E6",X"97",X"E6",X"99",X"60",X"2C",X"A9",
		X"DF",X"C9",X"02",X"8D",X"02",X"10",X"68",X"68",X"40",X"A2",X"DE",X"40",X"FC",X"DE",X"40",X"69",
		X"DF",X"C9",X"56",X"8D",X"0F",X"42",X"40",X"51",X"DE",X"C5",X"99",X"F0",X"02",X"A6",X"97",X"40",
		X"E3",X"E0",X"C9",X"7A",X"8D",X"01",X"48",X"DD",X"05",X"E1",X"8D",X"02",X"48",X"D9",X"08",X"E1",
		X"8D",X"03",X"48",X"C2",X"40",X"40",X"A6",X"DC",X"C2",X"60",X"C9",X"00",X"8D",X"00",X"48",X"40",
		X"E1",X"C2",X"C0",X"0E",X"D9",X"90",X"07",X"91",X"CD",X"88",X"10",X"F8",X"60",X"CD",X"00",X"10",
		X"50",X"FB",X"CD",X"00",X"10",X"10",X"FB",X"40",X"18",X"EB",X"E6",X"9E",X"C5",X"9E",X"A9",X"20",
		X"B0",X"14",X"C9",X"00",X"85",X"9E",X"C5",X"9F",X"F8",X"58",X"E9",X"01",X"85",X"9F",X"B8",X"10",
		X"05",X"68",X"68",X"2C",X"41",X"E1",X"C5",X"9E",X"C2",X"00",X"49",X"08",X"F0",X"02",X"C2",X"56",
		X"8E",X"0F",X"42",X"40",X"51",X"DE",X"C5",X"9F",X"28",X"2A",X"2A",X"2A",X"2A",X"18",X"69",X"15",
		X"8D",X"10",X"42",X"68",X"49",X"0F",X"69",X"15",X"8D",X"11",X"42",X"CD",X"04",X"10",X"29",X"FF",
		X"49",X"18",X"B0",X"CD",X"60",X"CD",X"00",X"10",X"10",X"FB",X"40",X"18",X"EB",X"C9",X"00",X"8D",
		X"00",X"54",X"85",X"E6",X"85",X"C1",X"40",X"FD",X"E1",X"40",X"2B",X"E2",X"60",X"C9",X"20",X"85",
		X"CD",X"40",X"BA",X"E8",X"40",X"3C",X"EE",X"40",X"89",X"EA",X"40",X"6D",X"EA",X"40",X"BA",X"E8",
		X"40",X"C8",X"E6",X"C6",X"E5",X"DC",X"62",X"E2",X"40",X"6E",X"E2",X"40",X"C8",X"E6",X"E6",X"E5",
		X"C5",X"E5",X"A9",X"02",X"B0",X"ED",X"C9",X"00",X"85",X"E5",X"60",X"C9",X"20",X"85",X"CD",X"C6",
		X"E5",X"DC",X"64",X"E2",X"40",X"6E",X"E2",X"C6",X"E5",X"DC",X"69",X"E2",X"40",X"E9",X"E5",X"40",
		X"C8",X"E6",X"E6",X"E5",X"C5",X"E5",X"A9",X"05",X"B0",X"E1",X"40",X"60",X"E6",X"40",X"BA",X"E8",
		X"C9",X"20",X"85",X"CD",X"40",X"C8",X"E6",X"40",X"C8",X"E6",X"40",X"C8",X"E6",X"C9",X"00",X"85",
		X"E5",X"60",X"0C",X"1D",X"32",X"37",X"3C",X"41",X"46",X"00",X"03",X"06",X"09",X"0C",X"D1",X"97",
		X"85",X"DD",X"A8",X"D1",X"97",X"A8",X"28",X"49",X"07",X"CA",X"F0",X"0A",X"18",X"C5",X"DD",X"69",
		X"20",X"85",X"DD",X"AA",X"B0",X"F6",X"68",X"2A",X"2A",X"2A",X"CA",X"DD",X"DF",X"E2",X"85",X"DE",
		X"C2",X"00",X"D1",X"97",X"F0",X"12",X"A9",X"FF",X"F0",X"14",X"58",X"E5",X"CD",X"81",X"DD",X"E6",
		X"DD",X"B0",X"02",X"E6",X"DE",X"A8",X"B0",X"EA",X"60",X"68",X"48",X"2C",X"C0",X"E2",X"C5",X"B7",
		X"28",X"2A",X"2A",X"2A",X"2A",X"CA",X"08",X"28",X"C5",X"C1",X"B0",X"ED",X"68",X"48",X"F0",X"0C",
		X"58",X"DD",X"E3",X"E2",X"E9",X"1B",X"C2",X"00",X"81",X"DD",X"E6",X"DD",X"68",X"49",X"0F",X"CA",
		X"58",X"DD",X"E3",X"E2",X"E9",X"1B",X"C2",X"00",X"81",X"DD",X"A8",X"E6",X"DD",X"B0",X"B3",X"40",
		X"41",X"42",X"43",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"41",X"42",X"43",
		X"44",X"45",X"46",X"02",X"1C",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"90",X"FF",X"00",X"09",
		X"04",X"42",X"55",X"52",X"4E",X"49",X"4E",X"3F",X"20",X"52",X"55",X"42",X"42",X"45",X"52",X"00",
		X"07",X"06",X"40",X"20",X"42",X"45",X"53",X"54",X"20",X"3A",X"20",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"53",X"20",X"40",X"00",X"09",X"09",X"36",X"20",X"00",X"09",X"0B",X"37",X"20",X"00",X"09",
		X"0D",X"38",X"20",X"00",X"09",X"0F",X"39",X"20",X"00",X"09",X"11",X"3A",X"20",X"00",X"05",X"15",
		X"42",X"4F",X"4E",X"55",X"53",X"20",X"43",X"41",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"02",X"15",X"42",X"4F",X"4E",X"55",X"53",X"20",X"43",
		X"41",X"52",X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"50",
		X"4F",X"49",X"4E",X"54",X"53",X"00",X"0F",X"15",X"32",X"30",X"30",X"30",X"30",X"00",X"0F",X"15",
		X"33",X"30",X"30",X"30",X"30",X"00",X"12",X"15",X"37",X"30",X"30",X"30",X"30",X"00",X"12",X"15",
		X"33",X"30",X"30",X"30",X"30",X"00",X"08",X"09",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",
		X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"5B",X"00",X"07",X"14",X"4E",X"45",X"58",X"54",X"06",
		X"57",X"41",X"59",X"06",X"49",X"53",X"06",X"53",X"50",X"52",X"49",X"4E",X"47",X"00",X"07",X"14",
		X"4E",X"45",X"58",X"54",X"06",X"57",X"41",X"59",X"06",X"49",X"53",X"06",X"53",X"55",X"4D",X"4D",
		X"45",X"52",X"00",X"08",X"14",X"4E",X"45",X"58",X"54",X"06",X"57",X"41",X"59",X"06",X"49",X"53",
		X"06",X"46",X"41",X"4C",X"4C",X"00",X"07",X"14",X"4E",X"45",X"58",X"54",X"06",X"57",X"41",X"59",
		X"06",X"49",X"53",X"06",X"57",X"49",X"4E",X"54",X"45",X"52",X"00",X"0B",X"16",X"47",X"4F",X"4F",
		X"44",X"06",X"4C",X"55",X"43",X"4B",X"5B",X"00",X"06",X"0B",X"59",X"4F",X"55",X"06",X"53",X"4D",
		X"41",X"53",X"48",X"45",X"44",X"06",X"FF",X"06",X"43",X"41",X"52",X"53",X"5E",X"00",X"08",X"0D",
		X"42",X"4F",X"4E",X"55",X"53",X"06",X"50",X"4F",X"49",X"4E",X"54",X"53",X"06",X"41",X"52",X"45",
		X"5C",X"00",X"08",X"12",X"14",X"11",X"11",X"06",X"10",X"06",X"FF",X"06",X"0F",X"06",X"00",X"0A",
		X"12",X"45",X"58",X"54",X"52",X"41",X"06",X"06",X"00",X"08",X"12",X"15",X"11",X"11",X"06",X"10",
		X"06",X"FF",X"06",X"0F",X"06",X"00",X"08",X"12",X"16",X"11",X"11",X"06",X"10",X"06",X"FF",X"06",
		X"0F",X"06",X"00",X"08",X"09",X"54",X"4F",X"06",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",X"45",
		X"06",X"50",X"4C",X"41",X"59",X"00",X"0B",X"0B",X"49",X"4E",X"53",X"45",X"52",X"54",X"06",X"43",
		X"4F",X"49",X"4E",X"00",X"07",X"0D",X"57",X"49",X"54",X"48",X"49",X"4E",X"06",X"06",X"FF",X"06",
		X"53",X"45",X"43",X"4F",X"4E",X"44",X"53",X"00",X"0B",X"0B",X"50",X"55",X"53",X"48",X"06",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"00",X"03",X"17",X"1C",X"55",X"50",X"06",X"FF",X"06",X"43",X"52",
		X"45",X"44",X"49",X"54",X"53",X"06",X"00",X"03",X"19",X"1D",X"55",X"50",X"06",X"FF",X"06",X"43",
		X"52",X"45",X"44",X"49",X"54",X"53",X"06",X"00",X"05",X"14",X"50",X"52",X"45",X"53",X"45",X"4E",
		X"54",X"45",X"44",X"20",X"42",X"59",X"20",X"44",X"41",X"54",X"41",X"20",X"45",X"41",X"53",X"54",
		X"00",X"03",X"16",X"79",X"20",X"43",X"4F",X"50",X"52",X"92",X"36",X"3E",X"3D",X"37",X"20",X"44",
		X"41",X"54",X"41",X"20",X"45",X"41",X"53",X"54",X"20",X"49",X"4E",X"43",X"92",X"00",X"04",X"06",
		X"53",X"43",X"4F",X"52",X"45",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"20",X"42",X"59",X"90",
		X"00",X"02",X"09",X"36",X"92",X"43",X"52",X"41",X"53",X"48",X"49",X"4E",X"47",X"20",X"43",X"41",
		X"52",X"53",X"20",X"49",X"4E",X"54",X"4F",X"20",X"42",X"41",X"52",X"52",X"49",X"45",X"52",X"53",
		X"00",X"02",X"0B",X"37",X"92",X"4A",X"55",X"4D",X"50",X"49",X"4E",X"47",X"20",X"41",X"4E",X"44",
		X"20",X"4C",X"41",X"4E",X"44",X"49",X"4E",X"47",X"20",X"4F",X"4E",X"20",X"43",X"41",X"52",X"53",
		X"00",X"02",X"0D",X"38",X"92",X"42",X"4F",X"4E",X"55",X"53",X"20",X"50",X"4F",X"49",X"4E",X"54",
		X"53",X"20",X"46",X"4F",X"52",X"20",X"46",X"49",X"4E",X"49",X"53",X"48",X"49",X"4E",X"47",X"00",
		X"0F",X"0D",X"7A",X"7B",X"7C",X"00",X"04",X"0E",X"43",X"4F",X"55",X"52",X"53",X"45",X"00",X"12",
		X"17",X"FF",X"06",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"53",X"00",X"12",X"19",X"FF",X"06",
		X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"53",X"00",X"02",X"10",X"39",X"92",X"38",X"37",X"20",
		X"43",X"4F",X"55",X"52",X"53",X"45",X"53",X"20",X"41",X"52",X"45",X"20",X"41",X"56",X"41",X"49",
		X"4C",X"41",X"42",X"4C",X"45",X"00",X"04",X"11",X"54",X"52",X"59",X"20",X"43",X"4F",X"4E",X"54",
		X"49",X"4E",X"55",X"4F",X"55",X"53",X"20",X"50",X"4C",X"41",X"59",X"20",X"54",X"4F",X"20",X"53",
		X"45",X"45",X"00",X"04",X"12",X"4D",X"4F",X"52",X"45",X"20",X"43",X"4F",X"55",X"52",X"53",X"45",
		X"53",X"00",X"0E",X"0F",X"54",X"49",X"4C",X"54",X"00",X"98",X"28",X"C9",X"03",X"85",X"E4",X"C2",
		X"00",X"D9",X"40",X"06",X"81",X"DD",X"A8",X"E6",X"DD",X"A6",X"E4",X"B0",X"F4",X"C9",X"03",X"85",
		X"E4",X"C9",X"00",X"81",X"DD",X"E6",X"DD",X"A6",X"E4",X"B0",X"F8",X"C9",X"03",X"85",X"E4",X"68",
		X"C8",X"D9",X"00",X"05",X"28",X"2A",X"2A",X"2A",X"2A",X"CA",X"F0",X"08",X"C5",X"E6",X"09",X"01",
		X"85",X"E6",X"B0",X"06",X"C5",X"E6",X"49",X"01",X"F0",X"06",X"58",X"DD",X"E3",X"E2",X"E9",X"1B",
		X"C2",X"00",X"81",X"DD",X"E6",X"DD",X"68",X"49",X"0F",X"CA",X"F0",X"08",X"C5",X"E6",X"09",X"01",
		X"85",X"E6",X"B0",X"06",X"C5",X"E6",X"49",X"01",X"F0",X"06",X"58",X"DD",X"E3",X"E2",X"E9",X"1B",
		X"C2",X"00",X"81",X"DD",X"A8",X"E6",X"DD",X"A6",X"E4",X"B0",X"B6",X"C9",X"00",X"85",X"E6",X"60",
		X"C9",X"20",X"85",X"CD",X"C0",X"00",X"CD",X"01",X"10",X"29",X"FF",X"28",X"49",X"04",X"B0",X"2C",
		X"C9",X"57",X"85",X"97",X"C9",X"E3",X"85",X"98",X"40",X"6E",X"E2",X"C9",X"25",X"85",X"CD",X"C0",
		X"00",X"68",X"49",X"02",X"B0",X"0A",X"C9",X"8E",X"85",X"97",X"C9",X"E3",X"85",X"98",X"B0",X"08",
		X"C9",X"86",X"85",X"97",X"C9",X"E3",X"85",X"98",X"40",X"6E",X"E2",X"60",X"C9",X"3E",X"85",X"97",
		X"C9",X"E3",X"85",X"98",X"40",X"6E",X"E2",X"C9",X"25",X"85",X"CD",X"C0",X"00",X"68",X"49",X"02",
		X"B0",X"0A",X"C9",X"76",X"85",X"97",X"C9",X"E3",X"85",X"98",X"B0",X"08",X"C9",X"7E",X"85",X"97",
		X"C9",X"E3",X"85",X"98",X"40",X"6E",X"E2",X"60",X"C2",X"40",X"CD",X"00",X"10",X"10",X"FB",X"8A",
		X"28",X"C5",X"05",X"85",X"B7",X"C0",X"00",X"40",X"6E",X"E2",X"40",X"94",X"C1",X"68",X"CA",X"CD",
		X"00",X"10",X"50",X"FB",X"40",X"18",X"EB",X"AA",X"10",X"E0",X"60",X"C2",X"01",X"CD",X"00",X"10",
		X"10",X"FB",X"CD",X"00",X"10",X"50",X"FB",X"40",X"18",X"EB",X"AA",X"B0",X"F0",X"60",X"CD",X"27",
		X"E7",X"85",X"0C",X"CD",X"28",X"E7",X"85",X"0B",X"CD",X"29",X"E7",X"85",X"0A",X"C2",X"0E",X"DD",
		X"27",X"E7",X"9D",X"00",X"05",X"AA",X"10",X"F7",X"C2",X"0E",X"58",X"DD",X"36",X"E7",X"E9",X"06",
		X"9D",X"40",X"06",X"AA",X"10",X"F4",X"60",X"01",X"00",X"12",X"00",X"76",X"84",X"00",X"53",X"28",
		X"00",X"32",X"36",X"00",X"19",X"82",X"53",X"41",X"57",X"4B",X"49",X"53",X"53",X"55",X"5A",X"4B",
		X"49",X"54",X"59",X"4F",X"53",X"C9",X"82",X"40",X"44",X"DA",X"C9",X"06",X"85",X"CD",X"C9",X"96",
		X"85",X"97",X"C9",X"E3",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"C2",X"30",X"40",X"ED",X"E6",
		X"40",X"A4",X"E7",X"40",X"D2",X"E7",X"C9",X"06",X"85",X"CD",X"C5",X"22",X"49",X"03",X"0A",X"CA",
		X"DD",X"9C",X"E7",X"85",X"97",X"DD",X"9D",X"E7",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"C2",
		X"30",X"40",X"ED",X"E6",X"C9",X"FB",X"85",X"97",X"C9",X"E3",X"85",X"98",X"C0",X"00",X"40",X"6E",
		X"E2",X"C2",X"60",X"40",X"ED",X"E6",X"C2",X"20",X"40",X"EA",X"C2",X"60",X"E6",X"E3",X"A9",X"E3",
		X"BE",X"E3",X"D3",X"E3",X"C9",X"00",X"85",X"B7",X"C5",X"21",X"85",X"CF",X"F0",X"11",X"C9",X"06",
		X"85",X"CD",X"F8",X"18",X"C5",X"B7",X"69",X"01",X"85",X"B7",X"A6",X"CF",X"B0",X"F5",X"B8",X"C9",
		X"08",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"C2",X"30",X"40",X"ED",
		X"E6",X"60",X"C9",X"1E",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"C2",
		X"30",X"40",X"ED",X"E6",X"C5",X"21",X"F0",X"32",X"C5",X"22",X"A9",X"01",X"B0",X"0E",X"C9",X"32",
		X"85",X"97",X"C9",X"E4",X"85",X"98",X"C9",X"03",X"85",X"D2",X"B0",X"2A",X"C5",X"22",X"A9",X"02",
		X"B0",X"0E",X"C9",X"49",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C9",X"04",X"85",X"D2",X"B0",X"16",
		X"C9",X"56",X"85",X"97",X"C9",X"E4",X"85",X"98",X"B0",X"08",X"C9",X"3F",X"85",X"97",X"C9",X"E4",
		X"85",X"98",X"C9",X"05",X"85",X"D2",X"C0",X"00",X"40",X"6E",X"E2",X"C9",X"00",X"85",X"CE",X"85",
		X"CF",X"85",X"E6",X"C5",X"21",X"B0",X"04",X"C9",X"64",X"85",X"21",X"F8",X"18",X"C5",X"CE",X"65",
		X"D2",X"85",X"CE",X"C5",X"CF",X"69",X"00",X"85",X"CF",X"A6",X"21",X"B0",X"EF",X"B8",X"C5",X"CF",
		X"40",X"83",X"E8",X"C5",X"CE",X"40",X"83",X"E8",X"C0",X"02",X"C2",X"00",X"58",X"C9",X"30",X"E9",
		X"1B",X"81",X"DD",X"E6",X"DD",X"88",X"B0",X"F2",X"C2",X"30",X"40",X"ED",X"E6",X"F8",X"18",X"C5",
		X"1C",X"65",X"CE",X"85",X"1C",X"C5",X"1D",X"65",X"CF",X"85",X"1D",X"B8",X"40",X"61",X"DB",X"40",
		X"29",X"DC",X"60",X"28",X"2A",X"2A",X"2A",X"2A",X"CA",X"F0",X"04",X"C9",X"FF",X"85",X"E6",X"C5",
		X"E6",X"F0",X"0C",X"58",X"DD",X"E3",X"E2",X"E9",X"1B",X"C2",X"00",X"81",X"DD",X"E6",X"DD",X"68",
		X"49",X"0F",X"CA",X"F0",X"04",X"C9",X"FF",X"85",X"E6",X"C5",X"E6",X"F0",X"0C",X"58",X"DD",X"E3",
		X"E2",X"E9",X"1B",X"C2",X"00",X"81",X"DD",X"E6",X"DD",X"60",X"C9",X"F3",X"85",X"97",X"C9",X"E2",
		X"85",X"98",X"60",X"40",X"6D",X"EA",X"8D",X"01",X"10",X"C9",X"06",X"85",X"B6",X"C9",X"06",X"85",
		X"CD",X"C9",X"63",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"C5",X"10",
		X"85",X"B7",X"C9",X"A6",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"CD",
		X"0A",X"04",X"40",X"42",X"E9",X"C9",X"7F",X"85",X"97",X"C9",X"E5",X"85",X"98",X"C0",X"00",X"40",
		X"6E",X"E2",X"C5",X"11",X"F0",X"22",X"85",X"B7",X"C9",X"B7",X"85",X"97",X"C9",X"E4",X"85",X"98",
		X"C0",X"00",X"40",X"6E",X"E2",X"CD",X"2A",X"04",X"40",X"42",X"E9",X"C9",X"8C",X"85",X"97",X"C9",
		X"E5",X"85",X"98",X"C0",X"00",X"40",X"6E",X"E2",X"C9",X"09",X"8D",X"02",X"10",X"40",X"5F",X"E9",
		X"F8",X"C5",X"B6",X"E9",X"01",X"85",X"B6",X"B8",X"10",X"EE",X"C2",X"60",X"C9",X"00",X"40",X"E1",
		X"C2",X"60",X"28",X"C9",X"00",X"85",X"B7",X"68",X"CA",X"F0",X"06",X"40",X"55",X"E9",X"AA",X"B0",
		X"FA",X"40",X"55",X"E9",X"60",X"F8",X"18",X"C5",X"B7",X"69",X"01",X"85",X"B7",X"B8",X"60",X"C2",
		X"40",X"CD",X"00",X"10",X"10",X"FB",X"8A",X"28",X"C5",X"05",X"B0",X"0A",X"C9",X"76",X"85",X"97",
		X"C9",X"E4",X"85",X"98",X"B0",X"08",X"C9",X"98",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C0",X"00",
		X"40",X"6E",X"E2",X"C9",X"01",X"85",X"C1",X"C9",X"84",X"85",X"97",X"C9",X"E4",X"85",X"98",X"C5",
		X"B6",X"85",X"B7",X"C0",X"00",X"40",X"6E",X"E2",X"C9",X"00",X"85",X"C1",X"40",X"BA",X"E8",X"C9",
		X"20",X"85",X"CD",X"C5",X"05",X"85",X"B7",X"C0",X"00",X"40",X"6E",X"E2",X"40",X"C1",X"E9",X"C9",
		X"06",X"85",X"CD",X"68",X"CA",X"CD",X"00",X"10",X"10",X"FB",X"40",X"18",X"EB",X"AA",X"10",X"A1",
		X"60",X"C5",X"05",X"F0",X"56",X"CD",X"04",X"10",X"29",X"FF",X"49",X"18",X"F0",X"4D",X"A9",X"08",
		X"F0",X"19",X"A9",X"10",X"B0",X"45",X"C5",X"05",X"A9",X"02",X"90",X"3F",X"C9",X"00",X"85",X"08",
		X"E6",X"08",X"40",X"7F",X"EA",X"40",X"FB",X"DB",X"2C",X"EF",X"E9",X"C9",X"00",X"85",X"08",X"E6",
		X"08",X"40",X"75",X"EA",X"40",X"FB",X"DB",X"C9",X"01",X"85",X"07",X"C2",X"FF",X"9A",X"40",X"CB",
		X"DC",X"40",X"1C",X"EA",X"C2",X"01",X"40",X"A6",X"DC",X"C9",X"00",X"8D",X"02",X"10",X"C2",X"01",
		X"40",X"A6",X"DC",X"C9",X"00",X"40",X"C3",X"C2",X"2C",X"37",X"C1",X"60",X"C2",X"2C",X"C9",X"00",
		X"95",X"00",X"E8",X"E0",X"F1",X"B0",X"F9",X"85",X"1A",X"85",X"1B",X"85",X"1C",X"85",X"1D",X"85",
		X"1E",X"85",X"1F",X"85",X"21",X"C2",X"07",X"9D",X"02",X"04",X"9D",X"22",X"04",X"AA",X"10",X"F7",
		X"8D",X"11",X"04",X"8D",X"12",X"04",X"8D",X"31",X"04",X"8D",X"32",X"04",X"CD",X"0C",X"04",X"09",
		X"3F",X"8D",X"0C",X"04",X"CD",X"2C",X"04",X"09",X"3F",X"8D",X"2C",X"04",X"CD",X"00",X"04",X"49",
		X"44",X"8D",X"00",X"04",X"CD",X"20",X"04",X"49",X"44",X"8D",X"20",X"04",X"60",X"C2",X"60",X"C9",
		X"00",X"40",X"E1",X"C2",X"60",X"F8",X"18",X"C5",X"10",X"69",X"01",X"85",X"10",X"B8",X"60",X"F8",
		X"18",X"C5",X"11",X"69",X"01",X"85",X"11",X"B8",X"60",X"C9",X"00",X"85",X"C6",X"40",X"E2",X"EA",
		X"E6",X"C6",X"C5",X"C6",X"0A",X"CA",X"E0",X"06",X"90",X"F3",X"8A",X"28",X"40",X"BA",X"E8",X"40",
		X"F2",X"EA",X"40",X"6D",X"EA",X"68",X"CA",X"40",X"E2",X"EA",X"40",X"BA",X"E8",X"40",X"C8",X"E6",
		X"E6",X"C6",X"C5",X"C6",X"0A",X"CA",X"E0",X"0C",X"90",X"ED",X"40",X"E2",X"EA",X"E6",X"C6",X"C5",
		X"C6",X"0A",X"CA",X"E0",X"10",X"90",X"F3",X"8A",X"28",X"40",X"BA",X"E8",X"40",X"C8",X"E6",X"68",
		X"CA",X"40",X"E2",X"EA",X"E6",X"C6",X"C5",X"C6",X"0A",X"CA",X"E0",X"16",X"90",X"F3",X"40",X"F2",
		X"EA",X"60",X"DD",X"02",X"EB",X"85",X"97",X"DD",X"03",X"EB",X"85",X"98",X"C0",X"00",X"40",X"6E",
		X"E2",X"60",X"40",X"BA",X"E8",X"40",X"C8",X"E6",X"40",X"C8",X"E6",X"40",X"C8",X"E6",X"40",X"C8",
		X"E6",X"60",X"C8",X"E4",X"E1",X"E4",X"70",X"E5",X"FE",X"E4",X"11",X"E5",X"31",X"E5",X"51",X"E5",
		X"76",X"E5",X"99",X"E5",X"B6",X"E5",X"D3",X"E5",X"40",X"5C",X"C0",X"CD",X"04",X"10",X"2A",X"90",
		X"01",X"60",X"40",X"DE",X"C2",X"85",X"09",X"85",X"08",X"85",X"07",X"C2",X"18",X"40",X"B2",X"C2",
		X"40",X"BA",X"C2",X"C9",X"20",X"85",X"CD",X"C9",X"E2",X"85",X"97",X"C9",X"E5",X"85",X"98",X"C0",
		X"00",X"40",X"6E",X"E2",X"C9",X"00",X"8D",X"00",X"54",X"8D",X"02",X"10",X"C5",X"05",X"F0",X"09",
		X"F8",X"C5",X"05",X"58",X"E9",X"01",X"85",X"05",X"B8",X"C2",X"00",X"CD",X"00",X"10",X"10",X"FB",
		X"8A",X"28",X"40",X"BA",X"E8",X"C5",X"05",X"85",X"B7",X"C0",X"00",X"40",X"6E",X"E2",X"68",X"CA",
		X"CD",X"00",X"10",X"50",X"FB",X"40",X"5C",X"C0",X"AA",X"B0",X"E0",X"40",X"6D",X"EA",X"C9",X"00",
		X"8D",X"01",X"10",X"C2",X"FF",X"9A",X"2C",X"2E",X"C1",X"40",X"33",X"D5",X"40",X"F0",X"D5",X"40",
		X"82",X"C2",X"40",X"94",X"C1",X"40",X"2B",X"EE",X"40",X"DD",X"EB",X"40",X"33",X"C3",X"40",X"47",
		X"EC",X"40",X"B2",X"CB",X"40",X"32",X"ED",X"40",X"D0",X"C6",X"40",X"9E",X"CC",X"40",X"E1",X"C6",
		X"40",X"A6",X"CD",X"40",X"26",X"C4",X"40",X"50",X"DA",X"40",X"9E",X"C2",X"C5",X"33",X"10",X"CF",
		X"C9",X"00",X"85",X"18",X"85",X"33",X"E6",X"2C",X"C5",X"2C",X"49",X"03",X"A9",X"03",X"B0",X"B9",
		X"C9",X"00",X"85",X"2C",X"85",X"2D",X"85",X"2E",X"85",X"2F",X"85",X"1F",X"60",X"C5",X"2C",X"49",
		X"10",X"F0",X"3B",X"C5",X"7A",X"49",X"68",X"B0",X"35",X"C5",X"2D",X"B0",X"2F",X"C5",X"2E",X"0A",
		X"CA",X"DD",X"1F",X"EC",X"85",X"37",X"DD",X"20",X"EC",X"85",X"2D",X"E6",X"2E",X"C5",X"2E",X"A9",
		X"06",X"B0",X"19",X"40",X"89",X"D9",X"C2",X"7F",X"40",X"CA",X"E6",X"C2",X"40",X"40",X"CA",X"E6",
		X"C9",X"00",X"CA",X"9D",X"00",X"42",X"9D",X"00",X"43",X"E8",X"B0",X"F7",X"A6",X"2D",X"60",X"04",
		X"40",X"00",X"40",X"06",X"15",X"10",X"01",X"00",X"20",X"05",X"10",X"00",X"18",X"05",X"10",X"06",
		X"50",X"04",X"90",X"10",X"10",X"06",X"24",X"10",X"10",X"05",X"30",X"00",X"3C",X"05",X"20",X"02",
		X"28",X"04",X"00",X"04",X"00",X"00",X"00",X"C5",X"2C",X"49",X"20",X"B0",X"2A",X"C2",X"00",X"86",
		X"E9",X"40",X"1B",X"D4",X"40",X"78",X"EC",X"C5",X"97",X"F0",X"09",X"40",X"13",X"C5",X"40",X"0B",
		X"ED",X"40",X"8D",X"C8",X"40",X"30",X"D4",X"C5",X"2C",X"49",X"10",X"F0",X"0A",X"C5",X"E9",X"18",
		X"69",X"10",X"CA",X"A9",X"40",X"90",X"D8",X"60",X"C5",X"2C",X"49",X"10",X"F0",X"34",X"C5",X"97",
		X"B0",X"30",X"40",X"F9",X"D1",X"C5",X"2F",X"0A",X"0A",X"CA",X"DD",X"B5",X"EC",X"A5",X"24",X"B0",
		X"21",X"DD",X"B6",X"EC",X"A5",X"23",X"90",X"1A",X"C9",X"80",X"85",X"97",X"DD",X"B4",X"EC",X"85",
		X"98",X"C9",X"08",X"85",X"99",X"DD",X"B3",X"EC",X"85",X"A1",X"CA",X"DD",X"98",X"CA",X"85",X"9C",
		X"E6",X"2F",X"60",X"00",X"88",X"7E",X"F0",X"02",X"B0",X"7E",X"F0",X"01",X"48",X"7D",X"80",X"07",
		X"80",X"7D",X"10",X"07",X"78",X"7C",X"78",X"02",X"98",X"7C",X"10",X"05",X"80",X"7A",X"E0",X"04",
		X"70",X"79",X"10",X"00",X"50",X"77",X"F0",X"09",X"90",X"75",X"E0",X"08",X"34",X"71",X"10",X"04",
		X"90",X"6E",X"E0",X"01",X"58",X"6E",X"80",X"08",X"80",X"6D",X"A0",X"04",X"88",X"6A",X"40",X"00",
		X"88",X"6B",X"10",X"05",X"B8",X"6A",X"E0",X"04",X"88",X"6A",X"40",X"06",X"A0",X"6A",X"80",X"07",
		X"88",X"6A",X"E0",X"07",X"70",X"6A",X"C0",X"FF",X"FF",X"FF",X"FF",X"C5",X"97",X"49",X"60",X"B0",
		X"20",X"C5",X"A1",X"A9",X"07",X"B0",X"0B",X"C5",X"98",X"85",X"17",X"40",X"E7",X"CF",X"40",X"42",
		X"CC",X"60",X"C5",X"99",X"18",X"69",X"02",X"85",X"99",X"A9",X"F8",X"90",X"04",X"C9",X"00",X"85",
		X"97",X"60",X"C5",X"2C",X"49",X"10",X"B0",X"06",X"40",X"3F",X"ED",X"40",X"7A",X"ED",X"60",X"C5",
		X"2C",X"49",X"08",X"B0",X"31",X"C9",X"80",X"85",X"3A",X"C9",X"50",X"85",X"3B",X"C9",X"08",X"85",
		X"3C",X"C6",X"1F",X"DD",X"77",X"ED",X"85",X"44",X"CA",X"DD",X"98",X"CA",X"85",X"3F",X"C9",X"80",
		X"85",X"2F",X"C9",X"04",X"85",X"37",X"C9",X"58",X"85",X"7B",X"C9",X"00",X"85",X"96",X"E6",X"1F",
		X"C5",X"2C",X"09",X"08",X"85",X"2C",X"60",X"00",X"02",X"08",X"C5",X"3A",X"F0",X"01",X"60",X"C6",
		X"1F",X"DD",X"18",X"EE",X"85",X"D5",X"DD",X"27",X"EE",X"85",X"3C",X"E8",X"DD",X"18",X"EE",X"85",
		X"D4",X"C9",X"00",X"85",X"D3",X"C9",X"A0",X"85",X"3B",X"C6",X"D5",X"C5",X"3C",X"18",X"69",X"18",
		X"85",X"3C",X"DD",X"1D",X"EE",X"85",X"44",X"C5",X"2C",X"49",X"04",X"B0",X"0A",X"C2",X"00",X"40",
		X"CB",X"CD",X"C9",X"FF",X"8D",X"03",X"03",X"C4",X"D3",X"C9",X"01",X"99",X"84",X"04",X"C6",X"44",
		X"DD",X"98",X"CA",X"99",X"85",X"04",X"C5",X"3B",X"29",X"FF",X"99",X"86",X"04",X"C5",X"3C",X"99",
		X"87",X"04",X"C5",X"D3",X"18",X"69",X"04",X"85",X"D3",X"E6",X"D5",X"C5",X"D5",X"A5",X"D4",X"90",
		X"B8",X"C5",X"2C",X"09",X"04",X"85",X"2C",X"40",X"C1",X"CD",X"A6",X"2F",X"B0",X"29",X"C2",X"60",
		X"C9",X"20",X"85",X"CD",X"40",X"BA",X"E8",X"40",X"CA",X"E6",X"40",X"04",X"C3",X"C5",X"2C",X"49",
		X"F3",X"85",X"2C",X"C9",X"E0",X"85",X"7C",X"C5",X"1F",X"A9",X"03",X"90",X"0A",X"C5",X"2C",X"09",
		X"10",X"85",X"2C",X"C9",X"90",X"85",X"7B",X"60",X"00",X"00",X"02",X"07",X"0A",X"00",X"04",X"01",
		X"02",X"03",X"05",X"07",X"06",X"08",X"09",X"00",X"68",X"38",X"58",X"40",X"BA",X"E8",X"C9",X"20",
		X"85",X"CD",X"C5",X"05",X"85",X"B7",X"C0",X"00",X"40",X"6E",X"E2",X"60",X"C2",X"60",X"C9",X"00",
		X"85",X"10",X"85",X"11",X"40",X"E1",X"C2",X"C0",X"1A",X"D9",X"67",X"EE",X"99",X"03",X"41",X"F0",
		X"05",X"C9",X"02",X"99",X"03",X"45",X"D9",X"82",X"EE",X"99",X"23",X"41",X"F0",X"05",X"C9",X"02",
		X"99",X"23",X"45",X"88",X"10",X"E3",X"60",X"20",X"21",X"24",X"25",X"28",X"29",X"2C",X"2D",X"30",
		X"2C",X"2D",X"38",X"00",X"28",X"29",X"24",X"25",X"20",X"21",X"20",X"21",X"34",X"35",X"28",X"29",
		X"48",X"49",X"22",X"23",X"26",X"27",X"2A",X"2B",X"2E",X"2F",X"32",X"2E",X"2F",X"3A",X"00",X"2A",
		X"2B",X"26",X"27",X"22",X"23",X"22",X"23",X"36",X"37",X"2A",X"2B",X"00",X"00",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"33",X"3F",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"3F",X"00",X"00",X"00",X"00",X"83",X"33",X"33",X"3F",X"00",
		X"00",X"00",X"08",X"33",X"33",X"33",X"3F",X"00",X"00",X"00",X"04",X"33",X"33",X"33",X"40",X"00",
		X"00",X"00",X"00",X"43",X"33",X"33",X"80",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"38",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"33",X"80",X"00",X"00",X"00",X"04",X"33",X"33",X"33",X"3F",
		X"00",X"00",X"00",X"08",X"33",X"33",X"33",X"3F",X"00",X"00",X"00",X"04",X"33",X"33",X"33",X"3F",
		X"00",X"00",X"00",X"08",X"33",X"33",X"33",X"3F",X"00",X"00",X"00",X"04",X"33",X"33",X"33",X"40",
		X"00",X"00",X"00",X"08",X"33",X"33",X"34",X"00",X"00",X"00",X"00",X"F3",X"33",X"33",X"3F",X"00",
		X"00",X"00",X"00",X"83",X"33",X"33",X"3F",X"00",X"00",X"00",X"00",X"43",X"33",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"18",X"00",X"00",X"00",X"00",X"81",X"22",X"22",X"13",X"F0",
		X"00",X"00",X"08",X"31",X"22",X"22",X"13",X"F0",X"00",X"00",X"F3",X"31",X"22",X"22",X"13",X"F0",
		X"00",X"00",X"F3",X"31",X"22",X"22",X"13",X"F0",X"00",X"00",X"F3",X"31",X"22",X"22",X"13",X"F0",
		X"00",X"00",X"F3",X"31",X"22",X"22",X"14",X"00",X"00",X"00",X"F3",X"31",X"22",X"22",X"18",X"00",
		X"00",X"00",X"F3",X"31",X"22",X"22",X"13",X"80",X"00",X"00",X"04",X"31",X"22",X"22",X"13",X"38",
		X"00",X"00",X"00",X"41",X"22",X"22",X"13",X"33",X"F0",X"00",X"00",X"F1",X"22",X"22",X"13",X"33",
		X"F0",X"00",X"00",X"F1",X"22",X"22",X"13",X"34",X"00",X"00",X"00",X"01",X"22",X"22",X"13",X"40",
		X"00",X"00",X"00",X"01",X"22",X"22",X"14",X"00",X"00",X"00",X"00",X"01",X"22",X"33",X"33",X"38",
		X"00",X"00",X"83",X"33",X"33",X"33",X"33",X"34",X"00",X"00",X"43",X"33",X"33",X"33",X"33",X"40",
		X"00",X"00",X"83",X"33",X"33",X"33",X"33",X"F0",X"00",X"00",X"43",X"33",X"33",X"66",X"63",X"F0",
		X"00",X"00",X"83",X"33",X"33",X"DD",X"C3",X"F0",X"00",X"00",X"43",X"33",X"33",X"DD",X"C3",X"F0",
		X"00",X"00",X"83",X"33",X"33",X"DD",X"C3",X"F0",X"00",X"00",X"43",X"33",X"33",X"AA",X"A3",X"F0",
		X"00",X"00",X"83",X"33",X"33",X"33",X"33",X"F0",X"00",X"0F",X"33",X"33",X"33",X"33",X"33",X"F0",
		X"00",X"08",X"33",X"33",X"33",X"33",X"33",X"F0",X"00",X"04",X"33",X"33",X"33",X"33",X"33",X"F0",
		X"00",X"00",X"43",X"33",X"33",X"33",X"33",X"F0",X"00",X"00",X"04",X"33",X"33",X"33",X"34",X"00",
		X"00",X"00",X"00",X"43",X"33",X"33",X"3F",X"00",X"00",X"00",X"00",X"F3",X"33",X"DD",X"59",X"AD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"AA",X"50",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",X"33",X"F0",X"00",
		X"00",X"E0",X"00",X"0F",X"33",X"33",X"F0",X"00",X"00",X"00",X"00",X"0F",X"33",X"33",X"F0",X"00",
		X"00",X"00",X"00",X"0F",X"33",X"33",X"F0",X"00",X"00",X"00",X"00",X"0F",X"33",X"33",X"F0",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"F0",X"00",X"00",X"00",X"00",X"83",X"33",X"33",X"F0",X"00",
		X"00",X"00",X"08",X"33",X"33",X"33",X"33",X"3F",X"00",X"00",X"F3",X"33",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"83",X"33",X"33",X"F0",X"33",X"3F",X"00",X"00",X"43",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"F3",X"33",X"33",X"F0",X"33",X"3F",X"00",X"00",X"04",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"08",X"33",X"33",X"F0",X"33",X"3F",X"00",X"00",X"04",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"08",X"33",X"33",X"F0",X"33",X"3F",X"00",X"00",X"E4",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"08",X"33",X"33",X"F0",X"33",X"40",X"00",X"00",X"83",X"33",X"33",X"F0",X"34",
		X"00",X"00",X"08",X"33",X"33",X"33",X"F0",X"4E",X"00",X"00",X"83",X"33",X"33",X"33",X"F0",X"00",
		X"00",X"00",X"43",X"33",X"33",X"33",X"F0",X"00",X"00",X"00",X"04",X"33",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"43",X"33",X"33",X"3F",X"00",X"00",X"00",X"00",X"F3",X"33",X"33",X"3F",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"3F",X"00",X"00",X"00",X"E0",X"F3",X"33",X"33",X"40",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"80",X"00",X"00",X"00",X"00",X"F3",X"33",X"33",X"40",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"8E",X"00",X"00",X"00",X"00",X"F3",X"33",X"33",X"30",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"F0",X"00",X"00",X"00",X"00",X"F3",X"33",X"33",X"F0",X"08",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"F0",X"03",X"80",X"00",X"00",X"F3",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"F3",X"33",X"33",X"F0",X"33",X"3F",X"00",X"00",X"04",X"33",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"00",X"43",X"33",X"F0",X"33",X"3F",X"00",X"00",X"00",X"83",X"33",X"F0",X"33",
		X"3F",X"00",X"00",X"08",X"33",X"33",X"F0",X"33",X"3F",X"00",X"00",X"04",X"33",X"33",X"3F",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"40",X"00",X"00",X"00",X"00",X"04",X"33",X"33",X"80",X"00",
		X"00",X"00",X"00",X"08",X"33",X"33",X"3F",X"00",X"00",X"00",X"00",X"F3",X"33",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"AA",X"AA",X"B1",X"00",X"00",X"00",X"01",X"BA",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"10",X"00",X"00",X"00",X"00",X"01",X"22",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C0",X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C0",
		X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"C0",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C0",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"33",X"3F",X"00",
		X"00",X"00",X"00",X"83",X"33",X"33",X"38",X"00",X"00",X"00",X"00",X"43",X"33",X"33",X"34",X"00",
		X"00",X"00",X"00",X"83",X"33",X"33",X"38",X"00",X"00",X"00",X"00",X"43",X"33",X"33",X"34",X"E0",
		X"00",X"00",X"00",X"83",X"33",X"33",X"38",X"00",X"00",X"00",X"00",X"43",X"33",X"33",X"34",X"00",
		X"00",X"00",X"00",X"83",X"33",X"33",X"38",X"00",X"00",X"00",X"00",X"43",X"33",X"33",X"34",X"00",
		X"00",X"00",X"00",X"83",X"33",X"33",X"38",X"00",X"00",X"00",X"00",X"43",X"33",X"33",X"34",X"00",
		X"00",X"00",X"00",X"83",X"33",X"33",X"3F",X"00",X"00",X"00",X"00",X"43",X"33",X"33",X"38",X"00",
		X"00",X"00",X"00",X"F3",X"33",X"66",X"66",X"71",X"00",X"00",X"00",X"01",X"76",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"22",X"10",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"E0",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"01",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"01",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"01",X"22",X"66",X"59",X"66",X"66",X"66",X"66",X"66",X"66",X"DD",X"50",X"9D",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",
		X"DA",X"AA",X"DD",X"DD",X"DD",X"DD",X"50",X"9D",X"C0",X"00",X"CD",X"DD",X"DD",X"DD",X"59",X"6D",
		X"C0",X"00",X"CD",X"DD",X"DD",X"DD",X"59",X"DD",X"C0",X"00",X"CD",X"DD",X"DD",X"DD",X"59",X"DD",
		X"C0",X"00",X"CD",X"DD",X"DD",X"DD",X"59",X"DD",X"C0",X"00",X"CD",X"DD",X"DD",X"DD",X"59",X"DD",
		X"C0",X"00",X"CD",X"DD",X"DD",X"DD",X"59",X"DD",X"D6",X"66",X"DD",X"DD",X"DD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"D6",X"66",X"66",X"66",X"66",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DA",X"AA",X"AA",X"AA",X"AA",X"DD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",
		X"00",X"00",X"00",X"01",X"CD",X"DD",X"DD",X"C1",X"00",X"00",X"00",X"01",X"CD",X"22",X"10",X"00",
		X"00",X"00",X"00",X"81",X"22",X"22",X"10",X"00",X"00",X"00",X"08",X"31",X"22",X"22",X"10",X"00",
		X"00",X"00",X"F3",X"31",X"22",X"22",X"10",X"00",X"00",X"00",X"F3",X"31",X"22",X"22",X"1F",X"00",
		X"00",X"00",X"F3",X"31",X"22",X"22",X"1F",X"00",X"00",X"00",X"F3",X"31",X"22",X"22",X"1F",X"00",
		X"00",X"00",X"F3",X"31",X"22",X"22",X"1F",X"00",X"00",X"00",X"04",X"31",X"22",X"22",X"18",X"00",
		X"00",X"00",X"00",X"41",X"22",X"22",X"13",X"80",X"00",X"00",X"00",X"F1",X"22",X"22",X"13",X"38",
		X"00",X"00",X"00",X"01",X"22",X"22",X"13",X"33",X"F0",X"00",X"00",X"E1",X"22",X"22",X"13",X"33",
		X"F0",X"00",X"00",X"01",X"22",X"22",X"13",X"34",X"00",X"00",X"00",X"01",X"22",X"22",X"13",X"40",
		X"00",X"00",X"00",X"01",X"22",X"22",X"14",X"00",X"00",X"00",X"00",X"01",X"22",X"DA",X"59",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"09",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"09",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"09",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"09",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"09",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"09",X"DD",
		X"AA",X"AA",X"AA",X"AA",X"DD",X"D5",X"09",X"DD",X"50",X"00",X"00",X"00",X"5D",X"D5",X"09",X"DD",
		X"50",X"00",X"00",X"00",X"5D",X"D5",X"09",X"DD",X"50",X"00",X"00",X"00",X"5D",X"D5",X"09",X"DD",
		X"50",X"00",X"00",X"00",X"5D",X"D5",X"09",X"DD",X"50",X"00",X"00",X"00",X"5D",X"D5",X"09",X"DD",
		X"D6",X"90",X"00",X"00",X"5D",X"D5",X"09",X"DD",X"DD",X"90",X"00",X"00",X"5D",X"D5",X"09",X"DD",
		X"DD",X"D6",X"66",X"66",X"DD",X"D6",X"59",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"34",X"00",X"33",
		X"3F",X"E0",X"00",X"08",X"33",X"40",X"00",X"33",X"3F",X"00",X"00",X"04",X"33",X"80",X"00",X"33",
		X"38",X"00",X"00",X"00",X"43",X"40",X"00",X"33",X"34",X"00",X"00",X"00",X"04",X"80",X"00",X"33",
		X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"66",X"66",X"66",X"33",X"00",X"00",X"33",
		X"33",X"AA",X"AA",X"AA",X"33",X"00",X"00",X"33",X"34",X"00",X"00",X"0F",X"33",X"80",X"00",X"33",
		X"38",X"00",X"00",X"0F",X"33",X"3F",X"00",X"33",X"34",X"00",X"00",X"08",X"33",X"3F",X"00",X"33",
		X"38",X"00",X"00",X"83",X"33",X"3F",X"00",X"33",X"34",X"00",X"00",X"43",X"33",X"3F",X"00",X"33",
		X"3F",X"00",X"00",X"83",X"33",X"38",X"00",X"33",X"3F",X"E0",X"00",X"43",X"33",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"CF",X"FF",X"EF",X"FF",X"AF",X"AF",X"AF",X"AF",
		X"6F",X"DF",X"6F",X"DF",X"EF",X"FF",X"CF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"7F",X"0F",X"6F",X"FF",X"6F",X"CF",X"7F",
		X"CF",X"7F",X"CF",X"6F",X"FF",X"6F",X"FF",X"7F",X"8F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"02",X"02",X"06",X"06",X"0E",X"0E",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"86",X"0E",X"CF",X"04",X"C8",X"00",X"4F",X"0F",X"C0",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"09",X"0A",X"02",X"06",X"00",X"00",X"0F",X"0F",X"00",X"03",X"00",
		X"00",X"08",X"E0",X"02",X"F0",X"30",X"F4",X"74",X"04",X"C6",X"A6",X"87",X"A7",X"A6",X"A6",X"A6",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"C2",X"00",X"C0",X"02",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"D0",X"50",X"D0",X"40",X"90",X"01",X"C0",X"F0",X"70",X"F0",X"30",X"E0",X"08",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"30",X"F0",X"FA",X"D0",X"B0",X"10",X"D0",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",
		X"18",X"D0",X"D0",X"B0",X"F8",X"F0",X"F0",X"32",X"04",X"04",X"02",X"02",X"00",X"00",X"00",X"08",
		X"00",X"01",X"00",X"01",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"21",X"20",X"80",X"30",X"00",X"10",X"00",X"40",X"00",X"00",X"0C",X"1E",X"0E",X"0F",X"0F",X"0F",
		X"50",X"00",X"00",X"08",X"00",X"08",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0B",X"0A",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",
		X"C7",X"F5",X"E5",X"FF",X"6F",X"0F",X"EF",X"7F",X"6F",X"FF",X"6F",X"CF",X"6F",X"CF",X"6F",X"1F",
		X"0F",X"0A",X"0A",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",
		X"FF",X"35",X"F5",X"FF",X"FF",X"FF",X"0F",X"FF",X"AF",X"8F",X"AF",X"AF",X"FF",X"BF",X"6F",X"8F",
		X"60",X"10",X"62",X"C2",X"68",X"C1",X"6A",X"F0",X"E8",X"71",X"61",X"04",X"E0",X"F1",X"C0",X"F4",
		X"0C",X"C9",X"0A",X"0D",X"04",X"0D",X"04",X"0E",X"0D",X"0A",X"05",X"09",X"04",X"0A",X"05",X"0E",
		X"6F",X"8D",X"FD",X"BF",X"AF",X"A7",X"AF",X"8F",X"0F",X"FF",X"FF",X"FE",X"FF",X"FB",X"FF",X"3F",
		X"1F",X"0E",X"0D",X"0E",X"0F",X"0F",X"0F",X"0E",X"0E",X"0B",X"0F",X"0F",X"0D",X"0F",X"0F",X"0D",
		X"08",X"02",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"00",X"00",X"00",X"00",
		X"02",X"05",X"0B",X"02",X"F4",X"30",X"F9",X"F0",X"90",X"10",X"10",X"12",X"51",X"3E",X"70",X"B0",
		X"07",X"0E",X"0D",X"0D",X"0F",X"0B",X"0F",X"05",X"04",X"00",X"09",X"00",X"0D",X"42",X"08",X"00",
		X"0F",X"0B",X"87",X"06",X"0B",X"03",X"1D",X"03",X"11",X"0C",X"1B",X"82",X"9A",X"10",X"15",X"68",
		X"70",X"B0",X"50",X"31",X"13",X"13",X"93",X"17",X"FF",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"10",X"60",X"90",X"10",X"10",X"80",X"10",X"00",X"10",X"01",X"03",X"03",X"87",X"0F",X"0F",X"0F",
		X"00",X"01",X"02",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"0F",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"EA",X"CB",X"FE",
		X"EF",X"FF",X"7F",X"8F",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"6F",X"CF",X"4F",X"C5",X"05",X"07",
		X"3F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"0A",X"FA",X"0F",
		X"FF",X"FF",X"1F",X"EF",X"4F",X"8F",X"2F",X"9F",X"AF",X"8F",X"AF",X"AF",X"FF",X"B5",X"05",X"9F",
		X"0B",X"0D",X"4F",X"CF",X"6D",X"CD",X"76",X"FE",X"FD",X"FF",X"7F",X"FF",X"7B",X"8D",X"EF",X"F7",
		X"CF",X"FE",X"07",X"EF",X"06",X"0F",X"0F",X"07",X"0F",X"05",X"0F",X"0E",X"07",X"0B",X"0F",X"EE",
		X"0F",X"96",X"FB",X"B7",X"AD",X"AF",X"A5",X"8F",X"2B",X"9B",X"47",X"8D",X"1B",X"EB",X"F7",X"FF",
		X"F7",X"03",X"31",X"00",X"00",X"00",X"0B",X"08",X"00",X"05",X"09",X"09",X"00",X"02",X"38",X"03",
		X"0B",X"87",X"0F",X"CD",X"07",X"0A",X"0E",X"07",X"0B",X"05",X"0A",X"07",X"03",X"00",X"70",X"00",
		X"FF",X"83",X"FE",X"FD",X"03",X"0F",X"00",X"02",X"0E",X"80",X"22",X"C1",X"F0",X"F0",X"B0",X"F0",
		X"3F",X"0F",X"76",X"07",X"0B",X"04",X"0D",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"30",
		X"B1",X"30",X"F2",X"10",X"E1",X"10",X"F0",X"10",X"B0",X"10",X"B0",X"10",X"D0",X"10",X"D0",X"10",
		X"BF",X"FF",X"FE",X"F7",X"2F",X"CF",X"0F",X"8B",X"0B",X"0E",X"05",X"09",X"F0",X"F0",X"F0",X"80",
		X"73",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"07",X"0D",X"0B",X"00",X"08",X"00",X"C0",X"00",X"80",
		X"DF",X"1F",X"DB",X"17",X"BF",X"1B",X"BF",X"1B",X"F7",X"1C",X"EA",X"14",X"F0",X"10",X"B0",X"30",
		X"0F",X"3F",X"0B",X"0F",X"0F",X"0D",X"0E",X"07",X"0F",X"0D",X"0E",X"09",X"74",X"08",X"30",X"00",
		X"0F",X"0F",X"0F",X"0D",X"0F",X"07",X"0F",X"0F",X"0E",X"0F",X"0B",X"07",X"0E",X"0B",X"0B",X"0F",
		X"0D",X"07",X"0E",X"0D",X"0F",X"FF",X"0F",X"1E",X"0B",X"D5",X"0D",X"F7",X"0B",X"DD",X"0B",X"1E",
		X"0F",X"0B",X"0B",X"0F",X"0E",X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"07",X"0E",X"0F",
		X"0F",X"0D",X"EB",X"0D",X"FF",X"1E",X"8F",X"FD",X"5D",X"C7",X"5F",X"1F",X"FB",X"5F",X"0F",X"7B",
		X"0F",X"1F",X"07",X"D3",X"01",X"F0",X"00",X"D0",X"01",X"13",X"01",X"F1",X"00",X"05",X"0F",X"0F",
		X"0B",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0F",
		X"0F",X"7F",X"F6",X"50",X"50",X"10",X"50",X"C0",X"80",X"F0",X"F0",X"10",X"E0",X"00",X"05",X"0F",
		X"0F",X"0E",X"0C",X"08",X"0C",X"08",X"00",X"00",X"08",X"08",X"00",X"00",X"08",X"08",X"0C",X"0E",
		X"00",X"00",X"01",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"C0",X"90",X"C0",X"F3",X"7F",X"7F",X"1F",X"EF",X"1F",X"CF",X"5F",X"8F",X"FF",X"FF",X"7F",X"FF",
		X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"06",X"FF",X"0F",X"EF",X"1F",X"CF",X"1F",X"9F",X"1F",X"9F",X"1F",X"BF",X"1F",X"AF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"68",X"78",X"5A",X"87",X"0D",X"A2",X"2A",X"22",X"66",X"66",X"EE",X"EE",X"66",X"66",X"66",
		X"F0",X"E0",X"3C",X"28",X"0F",X"69",X"E1",X"F0",X"C3",X"87",X"00",X"FF",X"FF",X"00",X"96",X"00",
		X"C1",X"2D",X"C3",X"0B",X"1E",X"D2",X"A1",X"2D",X"69",X"0F",X"00",X"FF",X"FF",X"00",X"78",X"00",
		X"F0",X"F0",X"C1",X"B0",X"2D",X"0B",X"45",X"45",X"44",X"66",X"66",X"77",X"77",X"66",X"66",X"66",
		X"F0",X"F0",X"34",X"F0",X"F0",X"E0",X"F0",X"34",X"F0",X"78",X"B0",X"F0",X"92",X"34",X"F0",X"F0",
		X"F0",X"F0",X"16",X"F0",X"F0",X"D0",X"F0",X"92",X"F0",X"E0",X"F0",X"92",X"F0",X"F0",X"34",X"F0",
		X"78",X"F0",X"78",X"F0",X"92",X"34",X"D0",X"F0",X"F0",X"F0",X"92",X"C1",X"F0",X"F0",X"F0",X"F0",
		X"D0",X"F0",X"E0",X"34",X"92",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"92",X"F0",X"E0",X"F0",X"F0",
		X"03",X"90",X"08",X"87",X"41",X"0F",X"0B",X"2D",X"07",X"02",X"08",X"41",X"09",X"0D",X"0F",X"0A",
		X"0E",X"0A",X"01",X"00",X"0C",X"0C",X"0F",X"43",X"94",X"0B",X"03",X"A1",X"07",X"03",X"28",X"05",
		X"07",X"0F",X"C2",X"07",X"03",X"04",X"02",X"41",X"02",X"01",X"09",X"08",X"0E",X"43",X"0E",X"09",
		X"0B",X"03",X"00",X"10",X"08",X"48",X"02",X"0F",X"09",X"03",X"25",X"4B",X"09",X"09",X"08",X"0E",
		X"83",X"07",X"0F",X"07",X"83",X"0F",X"0F",X"2C",X"41",X"41",X"29",X"29",X"0F",X"07",X"03",X"01",
		X"07",X"70",X"0F",X"1C",X"49",X"83",X"41",X"20",X"0F",X"07",X"0D",X"07",X"02",X"03",X"02",X"00",
		X"1C",X"0F",X"83",X"0F",X"0B",X"0A",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"02",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"EF",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"BF",X"FF",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"CF",X"FF",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"3F",X"FF",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0F",X"8F",X"AD",X"AD",X"0F",X"5E",X"2D",X"8F",X"4F",X"DE",X"9E",X"AF",X"8F",X"5E",X"8F",X"4B",
		X"3F",X"6F",X"5F",X"2F",X"BF",X"2F",X"BF",X"1F",X"2F",X"5F",X"AF",X"6F",X"BF",X"5F",X"AF",X"1F",
		X"0F",X"2F",X"2F",X"0F",X"0F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",X"4F",X"0F",X"0F",
		X"0F",X"1F",X"2F",X"1F",X"0F",X"0F",X"0F",X"1F",X"1F",X"4F",X"0F",X"0F",X"2F",X"0F",X"0F",X"2F",
		X"1E",X"3C",X"96",X"5A",X"38",X"34",X"1E",X"3C",X"34",X"1E",X"50",X"F0",X"3C",X"D2",X"34",X"F0",
		X"DF",X"AF",X"4F",X"CF",X"8F",X"8F",X"5E",X"8E",X"0F",X"0D",X"4B",X"2D",X"50",X"F0",X"F0",X"D0",
		X"8F",X"1F",X"2F",X"2F",X"0F",X"4F",X"0F",X"AF",X"BF",X"EF",X"1E",X"0F",X"D2",X"A0",X"F0",X"F0",
		X"0F",X"4F",X"8F",X"9F",X"4F",X"CF",X"2F",X"CF",X"EF",X"3F",X"4F",X"CF",X"0F",X"0F",X"58",X"F0",
		X"0F",X"4A",X"0C",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A5",X"4B",X"0D",X"87",X"07",X"0B",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"5A",X"4B",X"0F",X"09",X"86",X"0F",X"0B",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1C",X"29",X"1C",X"4B",X"A5",X"1A",X"06",X"04",X"0F",X"0F",X"07",X"0E",X"0C",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"EF",X"DF",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"BF",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"FF",X"CF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"3F",
		X"4F",X"2F",X"0F",X"0F",X"2F",X"2F",X"9F",X"1F",X"2F",X"0F",X"0F",X"0F",X"4F",X"2F",X"0F",X"8F",
		X"0F",X"1F",X"8F",X"0F",X"9F",X"0F",X"0F",X"8F",X"0F",X"AF",X"0F",X"1F",X"8F",X"4F",X"0F",X"1F",
		X"0F",X"9F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"0F",X"0F",X"0F",X"4F",X"8F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"87",X"97",X"0F",X"4B",X"A7",X"87",X"0F",X"0F",X"A7",X"0F",
		X"4F",X"8F",X"0F",X"2F",X"8F",X"5F",X"1F",X"8F",X"4F",X"2F",X"1F",X"0F",X"0F",X"1F",X"0F",X"C1",
		X"0F",X"CF",X"1F",X"2F",X"CF",X"0F",X"BF",X"1F",X"1F",X"2F",X"0F",X"0F",X"0F",X"60",X"06",X"F0",
		X"0F",X"0F",X"1F",X"0F",X"4F",X"1F",X"0F",X"3F",X"2F",X"0B",X"07",X"07",X"0B",X"C1",X"F0",X"F0",
		X"87",X"85",X"87",X"B7",X"07",X"D3",X"43",X"C3",X"A1",X"C2",X"C1",X"F0",X"E0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"1F",X"8F",X"0F",X"0F",X"0F",X"4F",X"4F",X"1F",X"AF",X"6F",X"FF",X"1F",X"2D",X"B0",
		X"CF",X"0F",X"8F",X"0F",X"0F",X"0F",X"8F",X"8F",X"2F",X"4F",X"FF",X"4F",X"87",X"0A",X"61",X"F0",
		X"0F",X"0F",X"4F",X"8F",X"0F",X"4F",X"0F",X"4F",X"8F",X"3F",X"5F",X"BF",X"9F",X"1C",X"0D",X"E0",
		X"0F",X"0F",X"4F",X"0F",X"0F",X"2F",X"1F",X"8F",X"0F",X"2F",X"1F",X"6F",X"BF",X"4F",X"8F",X"94",
		X"0F",X"0F",X"0F",X"2F",X"0F",X"8F",X"0F",X"0F",X"1F",X"0F",X"4F",X"8F",X"1F",X"4F",X"4F",X"0F",
		X"2F",X"8F",X"1F",X"2F",X"0F",X"0F",X"0F",X"1F",X"4F",X"AF",X"2F",X"8F",X"4F",X"2F",X"4F",X"1F",
		X"0F",X"4F",X"4F",X"0F",X"1F",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"8F",X"1F",X"0F",
		X"0F",X"2F",X"4F",X"2F",X"0F",X"1F",X"0F",X"2F",X"2F",X"8F",X"0F",X"0F",X"4F",X"0F",X"0F",X"4F",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0C",X"08",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0D",X"0F",X"0F",X"0D",X"05",X"03",X"0E",X"0E",X"09",X"0B",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"07",X"0F",X"0F",X"0E",X"0D",X"09",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"01",X"07",X"02",X"03",X"07",X"03",X"01",X"00",X"00",X"00",
		X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"28",X"CD",X"00",X"10",X"49",X"10",X"B0",X"0B",X"CD",X"00",X"A0",X"A9",X"2C",X"B0",X"04",X"68",
		X"2C",X"00",X"A0",X"68",X"2C",X"03",X"C0",X"78",X"B8",X"C2",X"FF",X"9A",X"CD",X"00",X"10",X"49",
		X"10",X"B0",X"0A",X"CD",X"00",X"A0",X"A9",X"2C",X"B0",X"03",X"2C",X"03",X"A0",X"2C",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"17",X"FF",X"17",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
