library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_0 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"C6",X"C6",X"82",X"C6",X"C6",X"7C",X"00",X"00",X"06",X"FE",X"FE",X"86",X"00",X"00",
		X"00",X"66",X"F2",X"BA",X"9E",X"8E",X"C6",X"62",X"00",X"7C",X"FE",X"92",X"92",X"92",X"C6",X"44",
		X"00",X"18",X"FE",X"1E",X"1A",X"D8",X"F8",X"F8",X"00",X"9C",X"BE",X"B2",X"B2",X"B2",X"F6",X"F6",
		X"00",X"4C",X"DE",X"92",X"92",X"92",X"FE",X"7C",X"00",X"E0",X"F0",X"98",X"8E",X"86",X"C2",X"E0",
		X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"7C",X"FE",X"92",X"92",X"92",X"F6",X"64",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"28",X"02",X"A4",X"25",X"A4",X"19",X"40",X"14",
		X"00",X"00",X"00",X"18",X"18",X"04",X"03",X"02",X"00",X"00",X"00",X"18",X"18",X"20",X"C0",X"40",
		X"02",X"03",X"04",X"18",X"18",X"00",X"00",X"00",X"40",X"C0",X"20",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"D6",X"D0",X"D0",X"D0",X"D6",X"7E",
		X"00",X"44",X"EE",X"BA",X"92",X"82",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"7C",X"FE",X"82",X"82",X"BA",X"FE",X"FE",X"00",X"C6",X"C6",X"92",X"92",X"92",X"FE",X"FE",
		X"00",X"C0",X"C0",X"90",X"92",X"96",X"FE",X"FE",X"00",X"6C",X"EE",X"8A",X"8A",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"D0",X"10",X"16",X"FE",X"FE",X"00",X"00",X"C6",X"FE",X"FE",X"FE",X"C6",X"00",
		X"00",X"FC",X"FE",X"C2",X"06",X"0E",X"0C",X"08",X"00",X"82",X"C6",X"EE",X"38",X"92",X"FE",X"FE",
		X"00",X"1E",X"0E",X"06",X"02",X"E2",X"FE",X"FE",X"00",X"FE",X"C6",X"60",X"30",X"60",X"C6",X"FE",
		X"00",X"FE",X"CE",X"9C",X"38",X"72",X"E6",X"FE",X"00",X"7C",X"EE",X"C6",X"C6",X"C6",X"EE",X"7C",
		X"00",X"60",X"F0",X"90",X"90",X"92",X"FE",X"FE",X"00",X"06",X"7E",X"F6",X"CE",X"C6",X"DE",X"7C",
		X"00",X"62",X"F6",X"9E",X"90",X"96",X"FE",X"FE",X"00",X"C4",X"8E",X"9A",X"9A",X"B2",X"F2",X"66",
		X"00",X"F0",X"C2",X"FE",X"FE",X"FE",X"C2",X"F0",X"00",X"FC",X"FE",X"FA",X"02",X"02",X"FE",X"FC",
		X"00",X"C0",X"F8",X"FC",X"0E",X"FC",X"F8",X"C0",X"00",X"FE",X"C6",X"0C",X"18",X"0C",X"C6",X"FE",
		X"00",X"C6",X"C6",X"28",X"10",X"28",X"C6",X"C6",X"00",X"FE",X"FE",X"D2",X"12",X"16",X"F6",X"F6",
		X"00",X"CE",X"E2",X"F2",X"BA",X"9E",X"8E",X"E6",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"C0",X"C0",X"80",X"C0",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"00",X"00",X"08",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"08",X"1C",X"34",X"08",X"00",X"00",X"00",X"00",X"0C",X"28",X"04",X"2E",X"14",X"00",
		X"00",X"08",X"A0",X"88",X"7C",X"20",X"48",X"00",X"38",X"60",X"8A",X"8A",X"22",X"58",X"38",X"00",
		X"10",X"24",X"00",X"40",X"44",X"42",X"28",X"10",X"02",X"10",X"04",X"02",X"00",X"20",X"02",X"0C",
		X"01",X"08",X"00",X"01",X"00",X"10",X"01",X"06",X"04",X"01",X"00",X"01",X"00",X"09",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"EE",X"E0",X"EE",X"0E",X"EE",X"E0",X"EE",X"0E",X"EE",X"E0",X"EE",X"0E",X"EE",X"00",X"00",
		X"0E",X"EE",X"E0",X"EE",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3B",X"44",X"92",X"BA",X"92",X"44",X"B8",X"81",X"F0",X"08",X"04",X"02",X"C1",X"21",X"11",X"91",
		X"89",X"88",X"84",X"83",X"40",X"20",X"10",X"0F",X"91",X"11",X"21",X"C1",X"02",X"04",X"08",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"08",X"04",X"04",X"04",X"08",X"F0",X"E0",
		X"03",X"07",X"3F",X"7F",X"FC",X"FC",X"78",X"30",X"C0",X"80",X"00",X"00",X"80",X"40",X"40",X"80",
		X"00",X"00",X"00",X"00",X"0F",X"1B",X"38",X"3F",X"00",X"00",X"3C",X"1C",X"08",X"88",X"F8",X"40",
		X"2F",X"09",X"0D",X"00",X"00",X"00",X"00",X"00",X"24",X"2C",X"1C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"3C",X"1C",X"08",X"88",X"F8",X"C0",
		X"2E",X"0B",X"0B",X"03",X"02",X"00",X"00",X"00",X"64",X"6C",X"3C",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3D",X"00",X"00",X"3C",X"1C",X"08",X"88",X"F8",X"40",
		X"2E",X"0B",X"0D",X"01",X"00",X"00",X"00",X"00",X"64",X"6C",X"BC",X"84",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"FF",X"11",X"11",X"11",X"11",X"FF",X"00",
		X"7E",X"81",X"81",X"81",X"81",X"81",X"81",X"00",X"00",X"81",X"81",X"81",X"81",X"81",X"81",X"7E",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"7E",X"7E",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"81",X"81",X"81",X"81",X"81",X"81",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",
		X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",
		X"12",X"0C",X"02",X"12",X"0A",X"00",X"34",X"0A",X"20",X"12",X"04",X"00",X"48",X"15",X"42",X"94",
		X"00",X"92",X"00",X"14",X"52",X"20",X"0A",X"01",X"80",X"50",X"45",X"32",X"0C",X"20",X"94",X"08",
		X"07",X"41",X"33",X"07",X"1B",X"01",X"07",X"1B",X"01",X"63",X"17",X"03",X"01",X"1B",X"23",X"05",
		X"87",X"8B",X"71",X"01",X"2B",X"17",X"03",X"C1",X"0B",X"07",X"03",X"37",X"0B",X"11",X"47",X"09",
		X"FF",X"6D",X"44",X"28",X"20",X"10",X"10",X"08",X"FF",X"EE",X"94",X"44",X"22",X"40",X"20",X"10",
		X"FF",X"DD",X"48",X"48",X"89",X"15",X"11",X"08",X"FF",X"E6",X"42",X"84",X"0A",X"09",X"10",X"08",
		X"00",X"00",X"85",X"4A",X"52",X"42",X"67",X"FF",X"00",X"00",X"05",X"92",X"62",X"11",X"3B",X"FF",
		X"10",X"90",X"60",X"24",X"28",X"44",X"EE",X"FF",X"20",X"10",X"14",X"08",X"6A",X"11",X"3B",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0E",X"1C",X"04",X"02",X"02",X"02",X"00",X"00",X"80",X"00",
		X"1A",X"10",X"20",X"1C",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4D",X"13",X"20",X"40",X"00",X"00",X"00",X"00",
		X"0D",X"2D",X"1D",X"0D",X"0D",X"0D",X"1D",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",
		X"04",X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"07",X"04",X"04",X"04",X"04",X"01",X"03",X"07",X"3F",X"3F",X"3E",X"3C",X"BF",X"03",X"03",X"80",
		X"04",X"04",X"04",X"27",X"24",X"24",X"04",X"04",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"04",X"34",X"07",X"04",X"04",X"04",X"04",X"04",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"06",X"05",X"04",X"04",X"08",X"04",X"08",X"30",X"30",X"38",X"3C",X"3E",
		X"04",X"04",X"04",X"04",X"07",X"04",X"04",X"34",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FC",X"B8",X"1F",X"15",X"7F",X"DC",X"7E",
		X"70",X"FE",X"1F",X"0A",X"1F",X"F4",X"7B",X"FF",X"FF",X"ED",X"FF",X"FB",X"FF",X"BD",X"FF",X"F7",
		X"18",X"3C",X"06",X"7C",X"81",X"F7",X"FD",X"BF",X"FF",X"39",X"1F",X"3C",X"FF",X"5E",X"74",X"3C",
		X"EC",X"E0",X"F0",X"FF",X"DF",X"E0",X"7C",X"F8",X"08",X"04",X"08",X"10",X"10",X"08",X"04",X"08",
		X"1F",X"0B",X"87",X"CD",X"FF",X"FF",X"DE",X"07",X"5F",X"3C",X"99",X"C3",X"E1",X"FD",X"EF",X"FF",
		X"FD",X"FF",X"B7",X"FF",X"FB",X"BF",X"FB",X"7F",X"1F",X"81",X"FD",X"F3",X"B7",X"BB",X"FF",X"FF",
		X"F7",X"A5",X"C7",X"87",X"83",X"41",X"00",X"00",X"FF",X"EB",X"7F",X"EF",X"FD",X"FC",X"70",X"38",
		X"FF",X"FB",X"CF",X"83",X"03",X"87",X"85",X"03",X"FF",X"FF",X"77",X"E5",X"CF",X"5F",X"5C",X"00",
		X"60",X"6E",X"E7",X"C3",X"73",X"FF",X"F6",X"FF",X"06",X"4E",X"82",X"C3",X"E5",X"F7",X"FF",X"FF",
		X"00",X"83",X"83",X"C7",X"E7",X"BF",X"FF",X"EF",X"3C",X"3E",X"77",X"7F",X"FD",X"FF",X"7B",X"EF",
		X"00",X"1F",X"20",X"40",X"90",X"99",X"9D",X"81",X"00",X"F0",X"08",X"44",X"A4",X"14",X"94",X"34",
		X"81",X"91",X"99",X"9C",X"40",X"20",X"1F",X"00",X"14",X"94",X"34",X"A4",X"44",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"40",X"84",X"8C",X"9C",X"80",X"00",X"F0",X"08",X"44",X"A4",X"A4",X"A4",X"A4",
		X"80",X"84",X"8C",X"9C",X"40",X"20",X"1F",X"00",X"A4",X"A4",X"A4",X"A4",X"44",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"40",X"9C",X"8C",X"84",X"80",X"00",X"F0",X"08",X"44",X"44",X"44",X"44",X"44",
		X"80",X"9C",X"8C",X"84",X"40",X"20",X"1F",X"00",X"44",X"44",X"44",X"44",X"44",X"08",X"F0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"08",X"04",X"04",X"04",X"04",X"03",X"00",X"00",X"60",X"90",X"90",X"90",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"60",X"90",X"90",X"90",X"92",X"0C",X"00",
		X"00",X"61",X"92",X"12",X"12",X"12",X"0C",X"00",X"00",X"06",X"09",X"09",X"09",X"01",X"00",X"00",
		X"00",X"10",X"20",X"20",X"20",X"20",X"C0",X"00",X"00",X"06",X"09",X"09",X"09",X"49",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"86",X"49",X"48",X"48",X"48",X"30",X"00",
		X"02",X"02",X"3C",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"40",X"40",X"3C",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"02",X"3C",X"40",X"40",X"3C",
		X"40",X"3C",X"02",X"02",X"3C",X"40",X"40",X"20",X"3C",X"40",X"40",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"3C",X"02",X"02",X"3C",X"40",X"40",X"3C",X"02",X"02",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"20",X"40",X"40",X"3C",X"02",X"02",X"3C",X"40",
		X"3C",X"06",X"03",X"01",X"01",X"03",X"07",X"3E",X"00",X"00",X"40",X"C0",X"C0",X"40",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"07",X"00",X"03",X"00",X"00",X"98",X"70",X"70",X"98",X"00",X"00",
		X"00",X"00",X"01",X"E3",X"FF",X"03",X"61",X"00",X"00",X"00",X"02",X"03",X"03",X"02",X"00",X"00",
		X"3C",X"60",X"C0",X"80",X"80",X"C0",X"E0",X"7C",X"00",X"00",X"19",X"0E",X"0E",X"19",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"E0",X"00",X"C0",X"00",X"00",X"80",X"CE",X"FF",X"C0",X"86",X"00",
		X"7C",X"E6",X"C3",X"81",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"18",
		X"A4",X"A4",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"3C",X"18",X"18",X"24",
		X"7C",X"38",X"10",X"10",X"18",X"58",X"58",X"10",X"18",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"81",X"81",X"81",X"C3",X"E6",X"7C",X"24",X"18",X"18",X"3C",X"24",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"A4",X"A4",X"10",X"58",X"58",X"18",X"10",X"10",X"38",X"7C",
		X"00",X"00",X"06",X"3E",X"3E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"07",X"01",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"C0",X"40",X"00",
		X"20",X"60",X"E0",X"E0",X"E0",X"E0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"7C",X"7C",X"60",X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"03",X"02",X"00",
		X"00",X"00",X"80",X"E0",X"E0",X"80",X"00",X"00",X"04",X"06",X"07",X"07",X"07",X"07",X"06",X"04",
		X"00",X"3C",X"3C",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"18",X"18",X"3C",X"3C",X"00",X"3C",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"3C",X"3C",X"7E",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"26",X"02",X"03",X"07",X"3E",X"04",X"00",X"00",X"00",X"40",X"E0",X"20",X"00",X"00",X"00",
		X"00",X"07",X"08",X"00",X"0F",X"01",X"00",X"00",X"00",X"88",X"48",X"F8",X"90",X"10",X"00",X"00",
		X"00",X"01",X"73",X"FE",X"FE",X"13",X"01",X"00",X"00",X"00",X"00",X"04",X"07",X"02",X"00",X"00",
		X"00",X"20",X"7C",X"E0",X"C0",X"40",X"64",X"38",X"00",X"00",X"08",X"09",X"1F",X"13",X"11",X"00",
		X"00",X"00",X"80",X"F0",X"80",X"10",X"E0",X"00",X"00",X"80",X"C8",X"7F",X"7F",X"CE",X"80",X"00",
		X"30",X"7C",X"E6",X"42",X"42",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"10",
		X"64",X"24",X"24",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"70",X"10",X"18",X"3C",
		X"E7",X"3C",X"18",X"18",X"3C",X"1C",X"1C",X"18",X"10",X"18",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"42",X"42",X"E6",X"7C",X"30",X"3C",X"18",X"10",X"70",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"28",X"24",X"24",X"74",X"18",X"1C",X"1C",X"3C",X"18",X"18",X"3C",X"66",
		X"01",X"03",X"07",X"05",X"0C",X"0E",X"0C",X"0E",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"01",X"03",X"07",X"05",X"0C",X"0E",X"0C",X"0E",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"10",X"00",
		X"01",X"03",X"07",X"05",X"0C",X"0E",X"0C",X"0E",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0C",X"0E",X"0C",X"05",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"04",X"00",X"00",X"00",X"0C",X"00",X"10",X"10",X"20",X"00",X"00",X"00",X"00",
		X"0E",X"0C",X"0E",X"0C",X"05",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"0C",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"00",
		X"0E",X"0C",X"0E",X"0C",X"05",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"56",X"0F",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"56",X"0F",
		X"00",X"00",X"08",X"30",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"56",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"3F",X"6A",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"3F",X"6A",X"F0",X"00",X"00",X"00",X"00",X"0C",X"10",X"00",X"00",
		X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"3F",X"6A",X"F0",X"00",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"00",
		X"00",X"00",X"18",X"3C",X"3C",X"58",X"20",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"1D",X"0E",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",
		X"00",X"00",X"18",X"3C",X"3C",X"58",X"20",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"1D",X"0E",X"07",X"02",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"20",X"10",X"10",
		X"00",X"00",X"18",X"3C",X"3C",X"58",X"20",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"1D",X"0E",X"07",X"02",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"02",X"07",X"0E",X"1D",X"18",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"14",X"20",X"58",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"07",X"0E",X"1D",X"18",X"10",X"10",X"20",X"00",X"00",X"02",X"0C",X"00",
		X"14",X"20",X"58",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"07",X"0E",X"1D",X"18",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"07",
		X"14",X"20",X"58",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"1C",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"30",X"F8",X"78",X"30",X"00",
		X"08",X"04",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"1C",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"30",X"F8",X"78",X"30",X"00",
		X"02",X"01",X"01",X"00",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"1C",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"30",X"F8",X"78",X"30",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0E",X"1C",X"0A",X"00",X"30",X"78",X"F8",X"30",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0E",X"1C",X"0A",X"00",X"30",X"78",X"F8",X"30",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"80",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0E",X"1C",X"0A",X"00",X"30",X"78",X"F8",X"30",X"80",X"00",X"00",
		X"00",X"00",X"20",X"C0",X"00",X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"40",X"10",X"20",X"40",X"00",X"00",X"00",X"00",X"08",
		X"20",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"02",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"40",X"00",X"00",X"00",X"00",X"10",
		X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"80",X"40",X"80",X"00",X"00",
		X"02",X"03",X"01",X"00",X"00",X"00",X"10",X"10",X"40",X"C0",X"80",X"00",X"00",X"00",X"10",X"10",
		X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"80",X"20",X"80",X"20",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",
		X"40",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"40",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"10",X"00",X"00",X"80",X"40",X"80",X"00",X"20",X"10",
		X"20",X"00",X"00",X"00",X"00",X"02",X"04",X"04",X"10",X"00",X"00",X"00",X"00",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"10",X"00",X"80",X"20",X"80",X"20",X"80",X"20",X"20",
		X"10",X"10",X"00",X"00",X"00",X"01",X"03",X"02",X"10",X"10",X"00",X"00",X"00",X"80",X"C0",X"40",
		X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"00",X"40",X"40",X"40",X"40",X"00",X"1E",X"00",
		X"20",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"20",X"00",X"00",X"20",X"40",X"40",X"04",X"18",X"00",
		X"20",X"00",X"00",X"01",X"04",X"08",X"10",X"00",X"00",X"00",X"20",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"10",X"10",X"20",X"00",X"00",X"10",X"20",X"24",X"58",X"20",X"00",
		X"20",X"00",X"00",X"09",X"10",X"24",X"08",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"1E",X"00",X"40",X"40",X"40",X"40",X"00",
		X"00",X"10",X"08",X"04",X"01",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"C0",X"20",X"00",X"00",
		X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"18",X"04",X"40",X"40",X"20",X"00",X"00",
		X"00",X"08",X"24",X"10",X"09",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",
		X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"58",X"24",X"20",X"10",X"00",X"00",
		X"00",X"02",X"02",X"02",X"02",X"00",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"04",X"02",X"02",X"20",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"10",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"00",X"00",X"10",X"00",X"08",X"04",X"02",X"80",X"00",X"00",
		X"00",X"00",X"08",X"04",X"24",X"1A",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",
		X"00",X"00",X"00",X"08",X"06",X"01",X"00",X"00",X"10",X"00",X"04",X"12",X"08",X"84",X"00",X"00",
		X"00",X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"10",
		X"00",X"78",X"00",X"02",X"02",X"02",X"02",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"02",X"04",X"08",X"00",X"10",
		X"00",X"18",X"20",X"02",X"02",X"04",X"00",X"00",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"06",X"08",X"00",X"00",X"00",X"00",X"00",X"84",X"08",X"12",X"04",X"00",X"10",
		X"00",X"04",X"1A",X"24",X"04",X"08",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"06",X"06",X"06",X"07",X"04",X"00",X"00",X"80",X"40",X"20",X"20",X"30",X"F8",X"68",
		X"00",X"04",X"07",X"06",X"06",X"02",X"02",X"01",X"68",X"F8",X"30",X"20",X"20",X"40",X"80",X"00",
		X"06",X"09",X"70",X"D0",X"88",X"18",X"13",X"00",X"00",X"00",X"80",X"40",X"20",X"30",X"F8",X"48",
		X"00",X"13",X"18",X"88",X"D0",X"70",X"09",X"06",X"48",X"F8",X"30",X"20",X"40",X"80",X"00",X"00",
		X"00",X"01",X"01",X"06",X"09",X"1F",X"09",X"00",X"80",X"40",X"40",X"00",X"20",X"B0",X"78",X"78",
		X"00",X"09",X"1F",X"09",X"06",X"01",X"01",X"00",X"78",X"78",X"B0",X"20",X"00",X"40",X"40",X"80",
		X"0F",X"06",X"03",X"00",X"03",X"02",X"03",X"1E",X"E0",X"C0",X"80",X"00",X"80",X"80",X"80",X"F0",
		X"0F",X"06",X"03",X"03",X"03",X"03",X"03",X"01",X"E0",X"C0",X"80",X"80",X"80",X"80",X"80",X"00",
		X"06",X"06",X"02",X"01",X"02",X"0B",X"0E",X"0F",X"C0",X"C0",X"80",X"00",X"80",X"A0",X"E0",X"E0",
		X"06",X"03",X"07",X"06",X"06",X"06",X"06",X"02",X"C0",X"80",X"40",X"20",X"20",X"20",X"20",X"40",
		X"06",X"03",X"02",X"01",X"02",X"0B",X"0A",X"0B",X"C0",X"80",X"80",X"00",X"80",X"A0",X"A0",X"A0",
		X"06",X"03",X"06",X"0C",X"0C",X"0C",X"0C",X"04",X"C0",X"80",X"70",X"08",X"04",X"04",X"04",X"04",
		X"01",X"03",X"03",X"03",X"03",X"03",X"06",X"0F",X"00",X"80",X"80",X"80",X"80",X"80",X"C0",X"E0",
		X"1E",X"03",X"02",X"03",X"00",X"03",X"06",X"0F",X"F0",X"80",X"80",X"80",X"00",X"80",X"C0",X"E0",
		X"02",X"06",X"06",X"06",X"06",X"07",X"03",X"06",X"40",X"20",X"20",X"20",X"20",X"40",X"80",X"C0",
		X"0F",X"0E",X"0B",X"02",X"01",X"02",X"06",X"06",X"E0",X"E0",X"A0",X"80",X"00",X"80",X"C0",X"C0",
		X"04",X"0C",X"0C",X"0C",X"0C",X"06",X"03",X"06",X"04",X"04",X"04",X"04",X"08",X"70",X"80",X"C0",
		X"0B",X"0A",X"0B",X"02",X"01",X"02",X"03",X"06",X"A0",X"A0",X"A0",X"80",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"10",X"18",X"1C",X"16",X"6F",X"D0",X"B0",X"60",
		X"06",X"0F",X"1F",X"3E",X"3C",X"38",X"00",X"00",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"0F",X"00",X"18",X"98",X"96",X"EE",X"D0",X"B0",X"7C",
		X"1A",X"31",X"21",X"01",X"02",X"0C",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"0D",X"1F",X"00",X"08",X"88",X"16",X"68",X"D0",X"B0",X"64",
		X"32",X"61",X"41",X"01",X"01",X"01",X"02",X"04",X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"3C",X"3E",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",
		X"03",X"03",X"03",X"02",X"00",X"00",X"00",X"00",X"60",X"B0",X"D0",X"7F",X"16",X"1C",X"18",X"10",
		X"00",X"00",X"0C",X"02",X"01",X"21",X"31",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"0F",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"7C",X"B0",X"D0",X"EE",X"96",X"98",X"18",X"00",
		X"04",X"02",X"01",X"01",X"01",X"41",X"61",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",
		X"1F",X"0D",X"01",X"01",X"01",X"00",X"00",X"00",X"64",X"B0",X"D0",X"68",X"16",X"88",X"08",X"00",
		X"08",X"18",X"38",X"68",X"F6",X"0B",X"0D",X"06",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",
		X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F8",X"7C",X"3C",X"1C",X"00",X"00",
		X"00",X"18",X"19",X"69",X"77",X"0B",X"0D",X"3E",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"1F",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"70",X"88",X"04",X"84",X"C0",X"60",X"00",X"00",
		X"00",X"10",X"11",X"68",X"16",X"1B",X"0D",X"26",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",
		X"1F",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"FC",X"82",X"01",X"00",X"80",X"C0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"00",X"00",X"1C",X"3C",X"7C",X"F8",X"F0",X"60",
		X"06",X"0D",X"0B",X"F6",X"68",X"38",X"18",X"08",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"1F",X"00",X"00",X"60",X"C0",X"84",X"04",X"88",X"70",
		X"3E",X"0D",X"0B",X"77",X"69",X"19",X"18",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"01",X"1F",X"26",X"60",X"C0",X"80",X"00",X"00",X"81",X"C2",X"FC",
		X"0D",X"0B",X"16",X"68",X"10",X"11",X"00",X"00",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"C0",
		X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"40",X"00",X"00",X"80",X"C0",
		X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"40",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"03",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"03",X"01",X"00",X"00",X"02",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"02",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",
		X"03",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",
		X"03",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",
		X"03",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"C0",
		X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"C0",
		X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"C0",
		X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"82",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"38",X"3C",X"3E",X"7F",X"FF",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"70",X"F8",X"7C",X"3C",X"1E",X"07",X"03",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"BE",X"BF",X"AF",X"BF",X"AB",X"BB",X"FF",X"9F",
		X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"9F",X"FB",X"BB",X"AF",X"BF",X"AB",X"AB",X"BE",
		X"00",X"00",X"00",X"3C",X"3E",X"14",X"15",X"3E",X"00",X"00",X"00",X"00",X"60",X"00",X"03",X"00",
		X"15",X"14",X"3E",X"3C",X"00",X"00",X"00",X"00",X"03",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"02",X"04",X"04",X"24",X"3C",X"07",X"C0",X"E0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",
		X"07",X"03",X"03",X"01",X"01",X"00",X"07",X"00",X"B0",X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"40",X"20",X"18",X"04",X"23",X"00",X"20",X"C0",X"40",X"82",X"84",X"38",X"C4",
		X"21",X"00",X"01",X"02",X"01",X"03",X"04",X"00",X"84",X"A0",X"20",X"10",X"08",X"88",X"04",X"00",
		X"02",X"02",X"01",X"01",X"01",X"00",X"40",X"2B",X"00",X"04",X"08",X"08",X"08",X"90",X"E0",X"20",
		X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"CE",X"41",X"80",X"40",X"20",X"10",X"20",
		X"00",X"00",X"00",X"20",X"20",X"11",X"0E",X"06",X"00",X"00",X"04",X"08",X"30",X"C0",X"C0",X"20",
		X"04",X"06",X"19",X"E0",X"01",X"02",X"04",X"04",X"38",X"44",X"83",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"09",X"00",X"20",X"20",X"34",X"82",X"84",X"E4",X"08",X"38",X"04",X"04",X"00",
		X"68",X"A0",X"20",X"11",X"00",X"07",X"00",X"00",X"04",X"04",X"0C",X"04",X"94",X"E2",X"81",X"40",
		X"09",X"10",X"20",X"10",X"80",X"00",X"80",X"00",X"B0",X"00",X"45",X"46",X"01",X"11",X"21",X"00",
		X"20",X"40",X"80",X"80",X"48",X"04",X"10",X"0D",X"00",X"00",X"01",X"09",X"0A",X"04",X"08",X"30",
		X"00",X"00",X"07",X"0B",X"1F",X"2D",X"3B",X"3F",X"00",X"00",X"E0",X"D0",X"F8",X"B4",X"DC",X"FC",
		X"3F",X"3B",X"2D",X"1F",X"0B",X"07",X"00",X"00",X"FC",X"DC",X"B4",X"F8",X"D0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
