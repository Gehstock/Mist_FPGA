library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity exerion_06 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;


architecture prom of exerion_06 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"E0",X"30",X"FF",X"FF",X"FF",X"FF",X"00",X"EE",X"33",X"00",X"88",X"FF",X"0F",X"07",
		X"00",X"EE",X"33",X"00",X"FF",X"FF",X"33",X"00",X"0F",X"0F",X"03",X"00",X"00",X"00",X"88",X"33",
		X"00",X"00",X"10",X"40",X"FF",X"FF",X"FF",X"FF",X"88",X"5B",X"CF",X"00",X"CC",X"FF",X"0F",X"07",
		X"80",X"FF",X"FF",X"00",X"3D",X"0F",X"CF",X"00",X"87",X"1E",X"0F",X"00",X"00",X"00",X"CC",X"31",
		X"00",X"00",X"10",X"40",X"FF",X"FF",X"FF",X"FF",X"4C",X"4B",X"0F",X"11",X"EE",X"FF",X"E1",X"34",
		X"C4",X"11",X"CC",X"11",X"D3",X"0F",X"0F",X"11",X"4B",X"0F",X"0F",X"01",X"00",X"00",X"EE",X"31",
		X"00",X"00",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"0F",X"32",X"EE",X"FF",X"2D",X"25",
		X"E6",X"30",X"00",X"33",X"D3",X"3C",X"07",X"23",X"87",X"F0",X"1E",X"03",X"00",X"00",X"FF",X"33",
		X"00",X"00",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"D2",X"32",X"E2",X"F8",X"E1",X"34",
		X"E6",X"F0",X"10",X"33",X"97",X"0E",X"0B",X"23",X"0F",X"0F",X"3C",X"03",X"00",X"08",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"E1",X"F0",X"47",X"EA",X"FB",X"0F",X"07",
		X"B3",X"F0",X"70",X"66",X"97",X"0D",X"0D",X"47",X"C3",X"3C",X"E1",X"34",X"00",X"EE",X"FF",X"71",
		X"00",X"00",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"97",X"F0",X"78",X"CF",X"F3",X"F8",X"E1",X"BC",
		X"B3",X"C0",X"F0",X"76",X"1F",X"0B",X"0E",X"47",X"E1",X"F0",X"78",X"25",X"CC",X"F3",X"FE",X"71",
		X"00",X"00",X"00",X"70",X"FF",X"FF",X"FF",X"FF",X"F1",X"F0",X"3C",X"CF",X"FF",X"FF",X"2D",X"AD",
		X"33",X"00",X"E0",X"70",X"1F",X"07",X"0F",X"47",X"E5",X"D2",X"F0",X"07",X"0F",X"F1",X"FC",X"33",
		X"FF",X"FF",X"C0",X"10",X"FF",X"FF",X"FF",X"FF",X"97",X"F0",X"78",X"CF",X"FB",X"F8",X"E1",X"BC",
		X"B3",X"C0",X"F0",X"76",X"1F",X"0B",X"0E",X"47",X"69",X"D2",X"B4",X"07",X"CC",X"F3",X"FE",X"71",
		X"FF",X"FF",X"70",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"E1",X"F0",X"47",X"EA",X"FA",X"0F",X"07",
		X"B3",X"F0",X"70",X"66",X"1F",X"49",X"0D",X"47",X"4B",X"C3",X"96",X"16",X"00",X"EE",X"FF",X"71",
		X"FF",X"FF",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"D2",X"32",X"E2",X"FA",X"A5",X"34",
		X"E6",X"F0",X"10",X"33",X"1F",X"68",X"0B",X"23",X"0F",X"69",X"1E",X"12",X"00",X"08",X"0F",X"03",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"0F",X"32",X"EE",X"FF",X"A5",X"25",
		X"E6",X"30",X"00",X"33",X"17",X"78",X"07",X"23",X"87",X"3C",X"1E",X"03",X"00",X"00",X"FF",X"31",
		X"FF",X"FF",X"90",X"40",X"FF",X"FF",X"FF",X"FF",X"4C",X"4B",X"0F",X"11",X"EE",X"FF",X"E1",X"25",
		X"C4",X"11",X"CC",X"11",X"93",X"3C",X"0F",X"11",X"87",X"96",X"1E",X"01",X"00",X"00",X"EE",X"31",
		X"FF",X"FF",X"90",X"40",X"FF",X"FF",X"FF",X"FF",X"88",X"5B",X"CF",X"00",X"CC",X"FF",X"0F",X"07",
		X"80",X"FF",X"FF",X"00",X"F1",X"1E",X"CF",X"00",X"0F",X"87",X"0F",X"00",X"00",X"00",X"CC",X"33",
		X"FF",X"FF",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"00",X"EE",X"33",X"00",X"88",X"FF",X"0F",X"07",
		X"00",X"EE",X"33",X"00",X"FF",X"FF",X"33",X"00",X"0F",X"0F",X"03",X"00",X"00",X"00",X"88",X"33",
		X"FF",X"FF",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B0",X"78",X"44",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"30",X"00",X"F0",X"F0",X"30",X"00",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"90",X"B2",X"EA",X"00",X"08",X"0F",X"00",X"70",X"F4",X"F0",X"78",X"00",X"FE",X"FF",X"F0",X"00",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"75",X"F4",X"11",X"0E",X"0F",X"03",X"72",X"FE",X"F0",X"3C",X"01",X"FE",X"FF",X"F3",X"10",
		X"00",X"00",X"80",X"10",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E8",X"32",X"E8",X"32",X"8F",X"FF",X"07",X"72",X"F4",X"F2",X"1E",X"21",X"FC",X"FF",X"F7",X"30",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"11",X"C0",X"75",X"9E",X"88",X"07",X"72",X"F0",X"F7",X"0F",X"30",X"F0",X"FF",X"FF",X"30",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"00",X"80",X"B2",X"8F",X"FF",X"0F",X"72",X"F4",X"7A",X"87",X"71",X"FC",X"FC",X"F3",X"52",
		X"00",X"00",X"80",X"10",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"00",X"B0",X"78",X"0F",X"0F",X"0F",X"72",X"FE",X"3C",X"CB",X"73",X"FE",X"FF",X"7F",X"43",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"E1",X"38",X"8F",X"FF",X"0F",X"72",X"F4",X"1E",X"E1",X"71",X"BE",X"FF",X"F7",X"70",
		X"C0",X"10",X"00",X"40",X"60",X"60",X"60",X"30",X"00",X"10",X"00",X"30",X"20",X"30",X"70",X"00",
		X"60",X"30",X"E0",X"30",X"8F",X"88",X"0F",X"72",X"F0",X"0F",X"F2",X"70",X"FE",X"FC",X"7F",X"43",
		X"E0",X"30",X"00",X"40",X"F0",X"40",X"F0",X"70",X"F0",X"70",X"90",X"70",X"B0",X"70",X"F0",X"00",
		X"F0",X"70",X"F0",X"70",X"8F",X"FF",X"0F",X"72",X"78",X"87",X"F7",X"70",X"F6",X"FE",X"F3",X"52",
		X"F0",X"70",X"F0",X"70",X"F0",X"50",X"F0",X"70",X"F0",X"70",X"90",X"70",X"90",X"70",X"F0",X"10",
		X"F0",X"70",X"F0",X"70",X"1E",X"0F",X"07",X"72",X"3C",X"C3",X"F2",X"30",X"F0",X"FF",X"FF",X"30",
		X"10",X"40",X"F0",X"70",X"90",X"70",X"90",X"40",X"F0",X"70",X"90",X"40",X"90",X"40",X"90",X"70",
		X"90",X"40",X"90",X"40",X"8F",X"FF",X"07",X"72",X"1E",X"E5",X"F0",X"30",X"FC",X"FF",X"F7",X"30",
		X"F0",X"70",X"F0",X"70",X"10",X"70",X"90",X"40",X"10",X"10",X"F0",X"40",X"F0",X"70",X"30",X"70",
		X"F0",X"70",X"F0",X"40",X"0E",X"0F",X"03",X"72",X"0F",X"FE",X"F0",X"10",X"FE",X"FF",X"F3",X"10",
		X"E0",X"30",X"20",X"40",X"30",X"60",X"30",X"60",X"20",X"10",X"F0",X"40",X"F0",X"70",X"30",X"60",
		X"F0",X"70",X"F0",X"60",X"08",X"0F",X"00",X"70",X"87",X"F4",X"F0",X"00",X"FE",X"FF",X"F0",X"00",
		X"C0",X"10",X"40",X"40",X"20",X"40",X"20",X"20",X"C0",X"10",X"F0",X"40",X"E0",X"30",X"30",X"00",
		X"60",X"30",X"60",X"20",X"00",X"00",X"00",X"70",X"C3",X"F0",X"30",X"00",X"F0",X"F0",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"70",X"60",X"30",X"20",X"20",X"E0",X"30",X"D0",X"50",X"D0",X"10",X"20",X"70",
		X"F0",X"70",X"10",X"40",X"10",X"00",X"10",X"60",X"00",X"60",X"E0",X"70",X"F0",X"70",X"E0",X"30",
		X"00",X"00",X"90",X"00",X"90",X"40",X"30",X"60",X"10",X"40",X"90",X"40",X"90",X"00",X"30",X"70",
		X"80",X"00",X"10",X"40",X"F0",X"30",X"20",X"30",X"00",X"40",X"10",X"00",X"00",X"60",X"10",X"40",
		X"00",X"00",X"90",X"00",X"90",X"40",X"10",X"40",X"10",X"40",X"90",X"40",X"90",X"00",X"10",X"50",
		X"80",X"00",X"F0",X"70",X"F0",X"70",X"C0",X"10",X"00",X"40",X"E0",X"70",X"80",X"10",X"10",X"40",
		X"00",X"00",X"90",X"00",X"F0",X"70",X"10",X"40",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"10",X"40",
		X"80",X"00",X"F0",X"70",X"F0",X"70",X"80",X"00",X"00",X"40",X"10",X"00",X"60",X"00",X"10",X"40",
		X"00",X"00",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"F0",X"70",X"F0",X"70",X"10",X"40",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"00",X"00",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"F0",X"70",X"10",X"40",X"10",X"60",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"00",X"00",X"E0",X"70",X"10",X"40",X"E0",X"30",X"10",X"40",X"10",X"40",X"10",X"00",X"E0",X"30",
		X"F0",X"70",X"10",X"40",X"10",X"20",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"E0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"E0",X"70",X"60",X"40",X"20",X"30",X"30",X"00",X"F0",X"30",X"F0",X"00",X"F0",X"30",
		X"30",X"60",X"30",X"00",X"30",X"40",X"00",X"00",X"00",X"40",X"60",X"60",X"CC",X"33",X"00",X"00",
		X"10",X"10",X"10",X"60",X"90",X"20",X"B0",X"70",X"10",X"00",X"00",X"40",X"00",X"30",X"00",X"40",
		X"40",X"70",X"C0",X"00",X"70",X"40",X"00",X"00",X"00",X"40",X"F0",X"40",X"62",X"64",X"00",X"00",
		X"10",X"10",X"10",X"50",X"90",X"10",X"90",X"70",X"F0",X"70",X"00",X"40",X"00",X"40",X"C0",X"70",
		X"80",X"70",X"00",X"70",X"F0",X"40",X"00",X"00",X"F0",X"70",X"F0",X"50",X"31",X"C8",X"00",X"00",
		X"F0",X"70",X"10",X"40",X"F0",X"70",X"90",X"40",X"F0",X"70",X"00",X"40",X"00",X"70",X"00",X"40",
		X"C0",X"10",X"C0",X"70",X"D0",X"50",X"00",X"00",X"F0",X"70",X"90",X"70",X"31",X"C8",X"66",X"33",
		X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"40",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"F0",X"00",X"F0",X"70",X"90",X"70",X"00",X"00",X"F0",X"70",X"10",X"70",X"F1",X"F8",X"66",X"33",
		X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"60",X"10",X"00",X"F0",X"70",X"F0",X"30",X"F0",X"70",
		X"70",X"10",X"F0",X"00",X"10",X"70",X"00",X"60",X"20",X"40",X"30",X"60",X"F1",X"F8",X"00",X"00",
		X"10",X"00",X"E0",X"30",X"10",X"00",X"60",X"20",X"30",X"00",X"F0",X"30",X"F0",X"00",X"F0",X"30",
		X"30",X"60",X"30",X"00",X"10",X"60",X"00",X"60",X"40",X"40",X"20",X"40",X"E2",X"74",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"33",X"00",X"00",
		X"BD",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"00",X"BD",X"FF",X"FF",X"F9",
		X"F9",X"F3",X"D5",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"F0",X"F0",X"F8",X"00",X"00",X"00",X"F9",X"CC",X"FF",X"FF",X"FF",X"1F",X"F0",X"F0",X"F8",
		X"F9",X"E2",X"D5",X"33",X"FF",X"00",X"EE",X"33",X"00",X"00",X"07",X"00",X"FF",X"FF",X"FF",X"FF",
		X"B5",X"F0",X"F0",X"F8",X"00",X"00",X"00",X"F9",X"E2",X"F0",X"F0",X"F8",X"A6",X"F0",X"F0",X"74",
		X"F9",X"EE",X"DD",X"00",X"F9",X"00",X"F1",X"74",X"00",X"00",X"02",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F9",X"F1",X"F0",X"F0",X"F8",X"CC",X"FF",X"FF",X"33",
		X"F9",X"00",X"00",X"00",X"F9",X"88",X"F0",X"F8",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F9",X"F9",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"04",
		X"BD",X"FF",X"FF",X"FF",X"F9",X"C4",X"FC",X"F9",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"F1",X"F0",X"F0",X"F8",X"FF",X"00",X"88",X"74",X"77",X"00",X"00",X"0E",
		X"1F",X"F0",X"F0",X"F8",X"F9",X"C4",X"32",X"F9",X"CC",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"F1",X"F0",X"F0",X"74",X"00",X"00",X"88",X"74",X"F9",X"33",X"00",X"04",
		X"B5",X"F0",X"F0",X"F8",X"F9",X"C4",X"32",X"F9",X"E2",X"F8",X"00",X"F9",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"33",X"FF",X"00",X"88",X"74",X"F1",X"FC",X"11",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F9",X"C4",X"32",X"F9",X"F1",X"F0",X"11",X"F9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"BD",X"FF",X"FF",X"FC",X"F7",X"F0",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"BD",X"F3",X"32",X"F9",X"F1",X"F3",X"32",X"F9",X"00",X"00",X"00",X"00",
		X"F1",X"F0",X"F0",X"F8",X"CC",X"FF",X"00",X"00",X"1F",X"F0",X"F0",X"F8",X"88",X"F3",X"F0",X"F8",
		X"FF",X"CC",X"33",X"FF",X"1F",X"F0",X"11",X"F9",X"F9",X"C4",X"32",X"F9",X"00",X"00",X"02",X"00",
		X"B5",X"F0",X"F0",X"F8",X"E2",X"F0",X"11",X"02",X"A6",X"F0",X"F0",X"F8",X"00",X"CC",X"F1",X"F8",
		X"F9",X"C4",X"32",X"F9",X"A6",X"F8",X"00",X"F9",X"F9",X"C4",X"32",X"F9",X"00",X"00",X"07",X"00",
		X"1F",X"FF",X"FF",X"FF",X"F1",X"F0",X"32",X"07",X"CC",X"FF",X"FF",X"FF",X"CC",X"77",X"EE",X"FF",
		X"F9",X"C4",X"32",X"F9",X"CC",X"77",X"04",X"FF",X"F9",X"C4",X"32",X"F9",X"00",X"00",X"02",X"00",
		X"B5",X"11",X"00",X"00",X"F9",X"F7",X"32",X"02",X"00",X"00",X"00",X"00",X"B7",X"74",X"00",X"00",
		X"F9",X"C4",X"32",X"F9",X"00",X"00",X"0E",X"00",X"BD",X"D5",X"FE",X"F9",X"00",X"00",X"00",X"00",
		X"E2",X"11",X"00",X"00",X"F9",X"C4",X"32",X"00",X"00",X"00",X"01",X"FF",X"1F",X"74",X"00",X"00",
		X"F9",X"C4",X"32",X"F9",X"CC",X"77",X"04",X"CC",X"1F",X"99",X"F0",X"F8",X"CC",X"77",X"00",X"CC",
		X"CC",X"11",X"00",X"00",X"F9",X"CC",X"33",X"00",X"00",X"08",X"03",X"F9",X"BD",X"33",X"00",X"00",
		X"F9",X"CC",X"33",X"F9",X"E2",X"F8",X"00",X"FB",X"B5",X"11",X"F1",X"F8",X"E2",X"F8",X"00",X"FB",
		X"00",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"00",X"00",X"01",X"F9",X"77",X"00",X"00",X"00",
		X"F9",X"00",X"00",X"F9",X"F1",X"F0",X"DD",X"F8",X"EE",X"11",X"EE",X"FF",X"F1",X"F0",X"DD",X"F8",
		X"87",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"E1",X"F0",X"F0",X"F0",X"78",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"C3",X"F0",X"F0",X"F0",X"3C",X"CF",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"87",X"F0",X"F0",X"F0",X"1E",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"1F",X"E1",X"F0",X"78",X"8F",X"3F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"3F",X"C3",X"F0",X"3C",X"CF",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"EF",X"87",X"F0",X"1E",X"7F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"8F",X"FF",X"77",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"CF",X"1F",X"69",X"8F",X"3F",X"2D",X"FF",X"FF",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"F0",
		X"F0",X"78",X"CF",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"0F",X"3F",X"0F",X"CF",X"0F",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"08",X"C3",X"F0",X"F0",
		X"F0",X"3C",X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"C3",X"1E",X"EF",X"0F",X"7F",X"87",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"87",X"F0",X"F0",
		X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"C3",X"78",X"CF",X"9F",X"3F",X"E1",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",
		X"F0",X"8F",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"87",X"F0",X"0F",X"FF",X"0F",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",
		X"0F",X"CF",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"0E",X"F0",X"3C",X"6F",X"C3",X"F0",X"8F",X"FF",X"77",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",
		X"0F",X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",
		X"0C",X"C3",X"78",X"0F",X"E1",X"3C",X"CF",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",
		X"00",X"87",X"F0",X"96",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",
		X"00",X"0E",X"E1",X"F0",X"78",X"8F",X"FF",X"77",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",
		X"00",X"08",X"C3",X"F0",X"3C",X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"87",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"C3",X"F0",X"3C",X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"E1",X"F0",X"78",X"8F",X"FF",X"77",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"87",X"F0",X"96",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"FF",
		X"0C",X"C3",X"78",X"0F",X"E1",X"3C",X"CF",X"FF",X"33",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"FF",
		X"0E",X"F0",X"3C",X"6F",X"C3",X"F0",X"8F",X"FF",X"77",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"3C",X"FF",
		X"87",X"F0",X"0F",X"FF",X"0F",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"3C",X"FF",
		X"C3",X"78",X"CF",X"FF",X"3F",X"E1",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"FF",
		X"FF",X"00",X"08",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"3C",X"EF",X"FF",X"19",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"08",X"0F",X"0F",X"EF",
		X"FF",X"11",X"0C",X"FF",X"FF",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"3C",X"FF",X"FF",X"00",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0C",X"E1",X"78",X"CF",
		X"FF",X"33",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"3C",X"FF",X"FF",X"00",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"8F",
		X"FF",X"7F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"FF",X"FF",X"00",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"87",X"F0",X"F0",X"1E",
		X"FF",X"1F",X"2D",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"FF",X"FF",X"00",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"3C",
		X"FF",X"0F",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"0F",X"3C",
		X"3F",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"3F",X"0F",X"CF",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"0F",X"3C",
		X"1F",X"E1",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"3F",X"0F",X"CF",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"3C",
		X"87",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"3C",
		X"C3",X"78",X"8F",X"FF",X"77",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"3C",
		X"E1",X"3C",X"CF",X"FF",X"33",X"00",X"00",X"00",X"0F",X"0F",X"87",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"F0",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"87",X"F0",X"F0",X"F0",X"1E",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"78",X"8F",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"8F",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"1E",X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"08",X"C3",X"F0",X"F0",X"78",X"CF",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"F0",X"3C",X"EF",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"0F",
		X"CF",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"F0",X"1E",X"FF",X"FF",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"0F",
		X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"8F",X"FF",X"77",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"C3",X"F0",X"F0",X"78",X"CF",X"FF",X"33",
		X"C3",X"3C",X"3F",X"F0",X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"F0",X"3C",X"EF",X"FF",X"11",
		X"C3",X"3C",X"0F",X"F0",X"0F",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"F0",X"1E",X"FF",X"FF",X"00",
		X"C3",X"3C",X"0F",X"F0",X"0F",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"1E",X"0F",X"0F",X"FF",
		X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"1E",X"0F",X"0F",X"FF",
		X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"3F",X"0F",
		X"CF",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"87",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"3F",X"0F",
		X"CF",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"8F",X"FF",X"77",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",
		X"0C",X"E1",X"F0",X"F0",X"F0",X"78",X"CF",X"FF",X"33",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",
		X"08",X"C3",X"F0",X"F0",X"F0",X"3C",X"EF",X"FF",X"11",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"87",X"F0",X"F0",X"F0",X"1E",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"0F",X"EF",X"FF",X"11",
		X"00",X"0E",X"F0",X"F0",X"F0",X"8F",X"FF",X"77",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"CF",X"FF",X"33",
		X"00",X"0C",X"E1",X"F0",X"78",X"CF",X"FF",X"33",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"F0",X"8F",X"FF",X"77",
		X"00",X"08",X"0F",X"0F",X"0F",X"EF",X"FF",X"11",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"1E",X"FF",X"FF",
		X"00",X"00",X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"08",X"C3",X"F0",X"F0",X"F0",X"3C",X"EF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"F0",X"F0",X"78",X"CF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"3F",X"F0",
		X"CF",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"8F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"0F",X"F0",
		X"0F",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"0F",X"F0",
		X"0F",X"C3",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"FF",X"FF",X"00",X"00",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"FF",
		X"00",X"00",X"E0",X"30",X"FF",X"FF",X"FF",X"FF",X"00",X"EE",X"33",X"00",X"88",X"FF",X"0F",X"07",
		X"00",X"EE",X"33",X"00",X"FF",X"FF",X"33",X"00",X"0F",X"0F",X"03",X"00",X"00",X"00",X"88",X"33",
		X"00",X"00",X"10",X"40",X"FF",X"FF",X"FF",X"FF",X"88",X"5B",X"CF",X"00",X"CC",X"FF",X"0F",X"07",
		X"80",X"FF",X"FF",X"00",X"3D",X"0F",X"CF",X"00",X"87",X"1E",X"0F",X"00",X"00",X"00",X"CC",X"31",
		X"00",X"00",X"10",X"40",X"FF",X"FF",X"FF",X"FF",X"4C",X"4B",X"0F",X"11",X"EE",X"FF",X"E1",X"34",
		X"C4",X"11",X"CC",X"11",X"D3",X"0F",X"0F",X"11",X"4B",X"0F",X"0F",X"01",X"00",X"00",X"EE",X"31",
		X"00",X"00",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"0F",X"32",X"EE",X"FF",X"2D",X"25",
		X"E6",X"30",X"00",X"33",X"D3",X"3C",X"07",X"23",X"87",X"F0",X"1E",X"03",X"00",X"00",X"FF",X"33",
		X"00",X"00",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"D2",X"32",X"E2",X"F8",X"E1",X"34",
		X"E6",X"F0",X"10",X"33",X"97",X"0E",X"0B",X"23",X"0F",X"0F",X"3C",X"03",X"00",X"08",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"E1",X"F0",X"47",X"EA",X"FB",X"0F",X"07",
		X"B3",X"F0",X"70",X"66",X"97",X"0D",X"0D",X"47",X"C3",X"3C",X"E1",X"34",X"00",X"EE",X"FF",X"71",
		X"00",X"00",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"97",X"F0",X"78",X"CF",X"F3",X"F8",X"E1",X"BC",
		X"B3",X"C0",X"F0",X"76",X"1F",X"0B",X"0E",X"47",X"E1",X"F0",X"78",X"25",X"CC",X"F3",X"FE",X"71",
		X"00",X"00",X"00",X"70",X"FF",X"FF",X"FF",X"FF",X"F1",X"F0",X"3C",X"CF",X"FF",X"FF",X"2D",X"AD",
		X"33",X"00",X"E0",X"70",X"1F",X"07",X"0F",X"47",X"E5",X"D2",X"F0",X"07",X"0F",X"F1",X"FC",X"33",
		X"FF",X"FF",X"C0",X"10",X"FF",X"FF",X"FF",X"FF",X"97",X"F0",X"78",X"CF",X"FB",X"F8",X"E1",X"BC",
		X"B3",X"C0",X"F0",X"76",X"1F",X"0B",X"0E",X"47",X"69",X"D2",X"B4",X"07",X"CC",X"F3",X"FE",X"71",
		X"FF",X"FF",X"70",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"E1",X"F0",X"47",X"EA",X"FA",X"0F",X"07",
		X"B3",X"F0",X"70",X"66",X"1F",X"49",X"0D",X"47",X"4B",X"C3",X"96",X"16",X"00",X"EE",X"FF",X"71",
		X"FF",X"FF",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"D2",X"32",X"E2",X"FA",X"A5",X"34",
		X"E6",X"F0",X"10",X"33",X"1F",X"68",X"0B",X"23",X"0F",X"69",X"1E",X"12",X"00",X"08",X"0F",X"03",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"2E",X"C3",X"0F",X"32",X"EE",X"FF",X"A5",X"25",
		X"E6",X"30",X"00",X"33",X"17",X"78",X"07",X"23",X"87",X"3C",X"1E",X"03",X"00",X"00",X"FF",X"31",
		X"FF",X"FF",X"90",X"40",X"FF",X"FF",X"FF",X"FF",X"4C",X"4B",X"0F",X"11",X"EE",X"FF",X"E1",X"25",
		X"C4",X"11",X"CC",X"11",X"93",X"3C",X"0F",X"11",X"87",X"96",X"1E",X"01",X"00",X"00",X"EE",X"31",
		X"FF",X"FF",X"90",X"40",X"FF",X"FF",X"FF",X"FF",X"88",X"5B",X"CF",X"00",X"CC",X"FF",X"0F",X"07",
		X"80",X"FF",X"FF",X"00",X"F1",X"1E",X"CF",X"00",X"0F",X"87",X"0F",X"00",X"00",X"00",X"CC",X"33",
		X"FF",X"FF",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"00",X"EE",X"33",X"00",X"88",X"FF",X"0F",X"07",
		X"00",X"EE",X"33",X"00",X"FF",X"FF",X"33",X"00",X"0F",X"0F",X"03",X"00",X"00",X"00",X"88",X"33",
		X"FF",X"FF",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B0",X"78",X"44",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"30",X"00",X"F0",X"F0",X"30",X"00",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"90",X"B2",X"EA",X"00",X"08",X"0F",X"00",X"70",X"F4",X"F0",X"78",X"00",X"FE",X"FF",X"F0",X"00",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"75",X"F4",X"11",X"0E",X"0F",X"03",X"72",X"FE",X"F0",X"3C",X"01",X"FE",X"FF",X"F3",X"10",
		X"00",X"00",X"80",X"10",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E8",X"32",X"E8",X"32",X"8F",X"FF",X"07",X"72",X"F4",X"F2",X"1E",X"21",X"FC",X"FF",X"F7",X"30",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"11",X"C0",X"75",X"9E",X"88",X"07",X"72",X"F0",X"F7",X"0F",X"30",X"F0",X"FF",X"FF",X"30",
		X"00",X"00",X"80",X"10",X"F0",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"00",X"80",X"B2",X"8F",X"FF",X"0F",X"72",X"F4",X"7A",X"87",X"71",X"FC",X"FC",X"F3",X"52",
		X"00",X"00",X"80",X"10",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"00",X"B0",X"78",X"0F",X"0F",X"0F",X"72",X"FE",X"3C",X"CB",X"73",X"FE",X"FF",X"7F",X"43",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"E1",X"38",X"8F",X"FF",X"0F",X"72",X"F4",X"1E",X"E1",X"71",X"BE",X"FF",X"F7",X"70",
		X"C0",X"10",X"00",X"40",X"60",X"60",X"60",X"30",X"00",X"10",X"00",X"30",X"20",X"30",X"70",X"00",
		X"60",X"30",X"E0",X"30",X"8F",X"88",X"0F",X"72",X"F0",X"0F",X"F2",X"70",X"FE",X"FC",X"7F",X"43",
		X"E0",X"30",X"00",X"40",X"F0",X"40",X"F0",X"70",X"F0",X"70",X"90",X"70",X"B0",X"70",X"F0",X"00",
		X"F0",X"70",X"F0",X"70",X"8F",X"FF",X"0F",X"72",X"78",X"87",X"F7",X"70",X"F6",X"FE",X"F3",X"52",
		X"F0",X"70",X"F0",X"70",X"F0",X"50",X"F0",X"70",X"F0",X"70",X"90",X"70",X"90",X"70",X"F0",X"10",
		X"F0",X"70",X"F0",X"70",X"1E",X"0F",X"07",X"72",X"3C",X"C3",X"F2",X"30",X"F0",X"FF",X"FF",X"30",
		X"10",X"40",X"F0",X"70",X"90",X"70",X"90",X"40",X"F0",X"70",X"90",X"40",X"90",X"40",X"90",X"70",
		X"90",X"40",X"90",X"40",X"8F",X"FF",X"07",X"72",X"1E",X"E5",X"F0",X"30",X"FC",X"FF",X"F7",X"30",
		X"F0",X"70",X"F0",X"70",X"10",X"70",X"90",X"40",X"10",X"10",X"F0",X"40",X"F0",X"70",X"30",X"70",
		X"F0",X"70",X"F0",X"40",X"0E",X"0F",X"03",X"72",X"0F",X"FE",X"F0",X"10",X"FE",X"FF",X"F3",X"10",
		X"E0",X"30",X"20",X"40",X"30",X"60",X"30",X"60",X"20",X"10",X"F0",X"40",X"F0",X"70",X"30",X"60",
		X"F0",X"70",X"F0",X"60",X"08",X"0F",X"00",X"70",X"87",X"F4",X"F0",X"00",X"FE",X"FF",X"F0",X"00",
		X"C0",X"10",X"40",X"40",X"20",X"40",X"20",X"20",X"C0",X"10",X"F0",X"40",X"E0",X"30",X"30",X"00",
		X"60",X"30",X"60",X"20",X"00",X"00",X"00",X"70",X"C3",X"F0",X"30",X"00",X"F0",X"F0",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"70",X"60",X"30",X"20",X"20",X"E0",X"30",X"D0",X"50",X"D0",X"10",X"20",X"70",
		X"F0",X"70",X"10",X"40",X"10",X"00",X"10",X"60",X"00",X"60",X"E0",X"70",X"F0",X"70",X"E0",X"30",
		X"00",X"00",X"90",X"00",X"90",X"40",X"30",X"60",X"10",X"40",X"90",X"40",X"90",X"00",X"30",X"70",
		X"80",X"00",X"10",X"40",X"F0",X"30",X"20",X"30",X"00",X"40",X"10",X"00",X"00",X"60",X"10",X"40",
		X"00",X"00",X"90",X"00",X"90",X"40",X"10",X"40",X"10",X"40",X"90",X"40",X"90",X"00",X"10",X"50",
		X"80",X"00",X"F0",X"70",X"F0",X"70",X"C0",X"10",X"00",X"40",X"E0",X"70",X"80",X"10",X"10",X"40",
		X"00",X"00",X"90",X"00",X"F0",X"70",X"10",X"40",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"10",X"40",
		X"80",X"00",X"F0",X"70",X"F0",X"70",X"80",X"00",X"00",X"40",X"10",X"00",X"60",X"00",X"10",X"40",
		X"00",X"00",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"F0",X"70",X"F0",X"70",X"10",X"40",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"00",X"00",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"F0",X"70",X"10",X"40",X"10",X"60",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"00",X"00",X"E0",X"70",X"10",X"40",X"E0",X"30",X"10",X"40",X"10",X"40",X"10",X"00",X"E0",X"30",
		X"F0",X"70",X"10",X"40",X"10",X"20",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"E0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"E0",X"70",X"60",X"40",X"20",X"30",X"30",X"00",X"F0",X"30",X"F0",X"00",X"F0",X"30",
		X"30",X"60",X"30",X"00",X"30",X"40",X"00",X"00",X"00",X"40",X"60",X"60",X"CC",X"33",X"00",X"00",
		X"10",X"10",X"10",X"60",X"90",X"20",X"B0",X"70",X"10",X"00",X"00",X"40",X"00",X"30",X"00",X"40",
		X"40",X"70",X"C0",X"00",X"70",X"40",X"00",X"00",X"00",X"40",X"F0",X"40",X"62",X"64",X"00",X"00",
		X"10",X"10",X"10",X"50",X"90",X"10",X"90",X"70",X"F0",X"70",X"00",X"40",X"00",X"40",X"C0",X"70",
		X"80",X"70",X"00",X"70",X"F0",X"40",X"00",X"00",X"F0",X"70",X"F0",X"50",X"31",X"C8",X"00",X"00",
		X"F0",X"70",X"10",X"40",X"F0",X"70",X"90",X"40",X"F0",X"70",X"00",X"40",X"00",X"70",X"00",X"40",
		X"C0",X"10",X"C0",X"70",X"D0",X"50",X"00",X"00",X"F0",X"70",X"90",X"70",X"31",X"C8",X"66",X"33",
		X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"40",X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"70",
		X"F0",X"00",X"F0",X"70",X"90",X"70",X"00",X"00",X"F0",X"70",X"10",X"70",X"F1",X"F8",X"66",X"33",
		X"F0",X"70",X"F0",X"70",X"F0",X"70",X"F0",X"60",X"10",X"00",X"F0",X"70",X"F0",X"30",X"F0",X"70",
		X"70",X"10",X"F0",X"00",X"10",X"70",X"00",X"60",X"20",X"40",X"30",X"60",X"F1",X"F8",X"00",X"00",
		X"10",X"00",X"E0",X"30",X"10",X"00",X"60",X"20",X"30",X"00",X"F0",X"30",X"F0",X"00",X"F0",X"30",
		X"30",X"60",X"30",X"00",X"10",X"60",X"00",X"60",X"40",X"40",X"20",X"40",X"E2",X"74",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"33",X"00",X"00",
		X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"70",X"00",X"00",X"F0",X"50",X"80",X"70",X"00",X"10",X"90",X"70",X"B0",X"70",X"F0",X"70",
		X"80",X"70",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"FF",X"FF",X"FF",X"FF",
		X"90",X"70",X"00",X"00",X"10",X"50",X"F0",X"70",X"F0",X"70",X"90",X"70",X"90",X"70",X"90",X"70",
		X"F0",X"70",X"10",X"70",X"00",X"00",X"88",X"00",X"88",X"00",X"80",X"00",X"FF",X"FF",X"FF",X"FF",
		X"10",X"40",X"F0",X"70",X"10",X"50",X"90",X"40",X"10",X"70",X"90",X"40",X"90",X"40",X"10",X"00",
		X"90",X"40",X"10",X"10",X"C4",X"11",X"C4",X"11",X"E2",X"32",X"E2",X"32",X"FF",X"FF",X"FF",X"FF",
		X"10",X"40",X"80",X"70",X"10",X"50",X"90",X"40",X"10",X"10",X"90",X"40",X"90",X"40",X"10",X"00",
		X"90",X"40",X"10",X"10",X"00",X"00",X"88",X"00",X"88",X"00",X"80",X"00",X"FF",X"FF",X"FF",X"FF",
		X"10",X"40",X"00",X"00",X"10",X"70",X"90",X"40",X"10",X"10",X"90",X"40",X"90",X"40",X"10",X"00",
		X"F0",X"40",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"70",X"00",X"00",X"70",X"70",X"30",X"60",X"F0",X"10",X"F0",X"60",X"F0",X"70",X"10",X"00",
		X"80",X"70",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"70",X"00",X"00",X"E0",X"50",X"00",X"70",X"00",X"10",X"A0",X"70",X"A0",X"70",X"E0",X"70",
		X"80",X"70",X"E0",X"70",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A0",X"70",X"00",X"00",X"20",X"50",X"E0",X"70",X"E0",X"70",X"A0",X"70",X"A0",X"70",X"A0",X"70",
		X"E0",X"70",X"A0",X"70",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"40",X"E0",X"70",X"20",X"50",X"A0",X"40",X"20",X"70",X"A0",X"40",X"A0",X"40",X"20",X"00",
		X"A0",X"40",X"A0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"40",X"00",X"70",X"20",X"70",X"A0",X"40",X"20",X"10",X"A0",X"40",X"A0",X"40",X"20",X"00",
		X"E0",X"40",X"A0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"70",X"00",X"00",X"60",X"70",X"A0",X"40",X"E0",X"10",X"E0",X"60",X"E0",X"70",X"20",X"00",
		X"80",X"70",X"E0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"30",X"00",X"00",X"E0",X"20",X"E0",X"30",X"00",X"10",X"A0",X"30",X"A0",X"30",X"E0",X"30",
		X"E0",X"30",X"E0",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"20",X"E0",X"30",X"A0",X"20",X"A0",X"20",X"E0",X"30",X"A0",X"20",X"A0",X"20",X"20",X"30",
		X"A0",X"20",X"A0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"30",X"80",X"30",X"A0",X"30",X"A0",X"20",X"20",X"10",X"E0",X"20",X"E0",X"30",X"20",X"00",
		X"E0",X"30",X"E0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"30",X"00",X"20",X"90",X"00",X"00",X"40",X"30",X"00",
		X"10",X"C0",X"70",X"80",X"40",X"00",X"00",X"00",X"00",X"C0",X"40",X"00",X"00",X"C0",X"70",X"00",
		X"00",X"00",X"C0",X"70",X"00",X"00",X"F0",X"30",X"00",X"20",X"90",X"00",X"00",X"C0",X"30",X"00",
		X"10",X"80",X"30",X"80",X"C0",X"70",X"00",X"00",X"00",X"20",X"30",X"00",X"00",X"C0",X"70",X"00",
		X"00",X"80",X"F0",X"F0",X"00",X"F0",X"F0",X"20",X"00",X"E0",X"F0",X"00",X"00",X"C0",X"30",X"00",
		X"10",X"00",X"10",X"80",X"40",X"C0",X"F0",X"00",X"00",X"20",X"10",X"00",X"00",X"40",X"50",X"00",
		X"00",X"F0",X"F0",X"10",X"C0",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"30",X"00",
		X"10",X"00",X"10",X"80",X"00",X"00",X"80",X"30",X"00",X"E0",X"70",X"00",X"00",X"C0",X"70",X"00",
		X"C0",X"F0",X"30",X"00",X"C0",X"10",X"10",X"00",X"00",X"E0",X"F0",X"00",X"00",X"C0",X"30",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"E0",X"30",X"00",X"20",X"40",X"00",X"00",X"C0",X"70",X"00",
		X"F0",X"70",X"00",X"00",X"C0",X"F0",X"10",X"20",X"00",X"80",X"30",X"00",X"00",X"C0",X"30",X"00",
		X"F0",X"F0",X"F0",X"F0",X"40",X"E0",X"F0",X"00",X"00",X"20",X"50",X"00",X"00",X"80",X"30",X"00",
		X"F0",X"00",X"00",X"80",X"00",X"80",X"F0",X"30",X"00",X"80",X"30",X"00",X"00",X"40",X"20",X"00",
		X"F0",X"F0",X"F0",X"F0",X"C0",X"F0",X"10",X"00",X"00",X"E0",X"70",X"00",X"00",X"C0",X"60",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"20",X"00",X"E0",X"F0",X"00",X"00",X"C0",X"30",X"00",
		X"10",X"00",X"00",X"80",X"C0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"80",X"10",
		X"10",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"10",X"F0",X"30",X"00",X"C0",X"F0",X"00",X"00",X"90",X"30",X"10",
		X"70",X"00",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"F0",X"C0",X"10",
		X"00",X"00",X"C0",X"F0",X"C0",X"00",X"10",X"30",X"00",X"60",X"10",X"00",X"00",X"10",X"10",X"10",
		X"D0",X"30",X"00",X"00",X"80",X"F0",X"F0",X"10",X"00",X"00",X"70",X"00",X"00",X"90",X"30",X"00",
		X"00",X"C0",X"F0",X"F0",X"40",X"00",X"00",X"20",X"00",X"C0",X"F0",X"00",X"00",X"F0",X"F0",X"10",
		X"10",X"E0",X"10",X"00",X"C0",X"10",X"80",X"30",X"00",X"E0",X"00",X"00",X"00",X"10",X"10",X"00",
		X"80",X"F0",X"F0",X"90",X"40",X"00",X"00",X"30",X"00",X"40",X"10",X"00",X"00",X"F0",X"F0",X"10",
		X"00",X"00",X"F0",X"00",X"40",X"00",X"00",X"20",X"00",X"C0",X"30",X"00",X"00",X"F0",X"F0",X"10",
		X"E0",X"F0",X"30",X"00",X"C0",X"00",X"80",X"10",X"00",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"30",X"C0",X"10",X"80",X"30",X"00",X"20",X"40",X"00",X"00",X"F0",X"F0",X"10",
		X"F0",X"30",X"10",X"00",X"80",X"F0",X"F0",X"00",X"00",X"20",X"80",X"00",X"00",X"F0",X"F0",X"10",
		X"00",X"00",X"80",X"F0",X"80",X"F0",X"F0",X"10",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"10",X"00",X"00",X"F0",X"70",X"00",X"00",X"C0",X"70",X"00",X"00",X"C0",X"30",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"E0",X"70",X"00",X"00",X"C0",X"30",X"00",X"00",X"30",X"80",X"10",
		X"F0",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"C0",X"10",X"80",X"30",X"00",X"00",X"E0",X"00",
		X"00",X"80",X"F0",X"F0",X"C0",X"30",X"00",X"C0",X"00",X"70",X"00",X"20",X"00",X"90",X"30",X"10",
		X"80",X"F0",X"10",X"80",X"F0",X"00",X"80",X"F0",X"C0",X"00",X"00",X"30",X"00",X"80",X"F0",X"10",
		X"10",X"F0",X"F0",X"10",X"E0",X"70",X"C0",X"F0",X"80",X"F0",X"C0",X"30",X"00",X"10",X"10",X"10",
		X"00",X"80",X"F0",X"B0",X"70",X"00",X"00",X"E0",X"40",X"80",X"30",X"20",X"00",X"F0",X"10",X"00",
		X"F0",X"F0",X"30",X"00",X"F0",X"F0",X"E0",X"70",X"C0",X"C0",X"F0",X"10",X"00",X"F0",X"F0",X"10",
		X"00",X"00",X"00",X"E0",X"30",X"00",X"00",X"C0",X"40",X"00",X"10",X"20",X"00",X"F0",X"F0",X"10",
		X"F0",X"70",X"00",X"00",X"30",X"C0",X"F0",X"30",X"40",X"80",X"30",X"00",X"00",X"F0",X"F0",X"10",
		X"00",X"00",X"00",X"80",X"10",X"C0",X"70",X"80",X"40",X"00",X"10",X"20",X"00",X"00",X"80",X"10",
		X"F0",X"00",X"00",X"00",X"10",X"80",X"30",X"00",X"40",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"10",X"10",X"00",X"10",X"80",X"30",X"80",X"C0",X"F0",X"F0",X"30",X"00",X"C0",X"F0",X"10",
		X"10",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"40",X"00",X"10",X"20",X"00",X"F0",X"70",X"00",
		X"60",X"00",X"F0",X"F0",X"10",X"00",X"10",X"80",X"C0",X"F0",X"F0",X"30",X"00",X"F0",X"70",X"00",
		X"10",X"F0",X"F0",X"00",X"10",X"00",X"10",X"00",X"C0",X"F0",X"F0",X"30",X"00",X"00",X"C0",X"10",
		X"30",X"00",X"F0",X"70",X"10",X"00",X"10",X"80",X"40",X"00",X"00",X"20",X"00",X"70",X"20",X"10",
		X"C0",X"F0",X"F0",X"30",X"10",X"00",X"10",X"80",X"C0",X"F0",X"F0",X"30",X"00",X"80",X"F0",X"10",
		X"10",X"00",X"10",X"60",X"F0",X"F0",X"F0",X"F0",X"C0",X"F0",X"F0",X"30",X"00",X"C0",X"F0",X"10",
		X"E0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"40",X"00",X"00",X"20",X"00",X"F0",X"30",X"00",
		X"10",X"00",X"10",X"C0",X"F0",X"F0",X"F0",X"F0",X"80",X"F0",X"F0",X"30",X"00",X"00",X"00",X"10",
		X"30",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"C0",X"10",X"80",X"30",X"00",X"70",X"00",X"00",
		X"10",X"00",X"00",X"80",X"F0",X"F0",X"F0",X"F0",X"00",X"E0",X"10",X"20",X"00",X"60",X"F0",X"00",
		X"10",X"00",X"00",X"80",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"30",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"C0",X"10",X"00",X"00",X"80",X"00",X"80",X"70",X"00",X"00",X"10",X"90",X"10",
		X"10",X"00",X"00",X"80",X"10",X"00",X"00",X"80",X"40",X"C0",X"70",X"20",X"00",X"E0",X"F0",X"00",
		X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"80",X"00",X"00",X"F0",X"10",X"00",X"10",X"00",X"10",
		X"30",X"00",X"00",X"C0",X"00",X"00",X"00",X"F0",X"40",X"80",X"30",X"20",X"00",X"F0",X"F0",X"10",
		X"E0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"00",X"E0",X"70",X"00",X"00",X"30",X"80",X"10",
		X"E0",X"F0",X"F0",X"70",X"70",X"00",X"00",X"C0",X"40",X"00",X"10",X"20",X"00",X"10",X"00",X"10",
		X"C0",X"F0",X"F0",X"30",X"C0",X"F0",X"F0",X"F0",X"C0",X"F0",X"00",X"00",X"00",X"E0",X"F0",X"00",
		X"C0",X"F0",X"F0",X"30",X"30",X"00",X"00",X"80",X"C0",X"F0",X"F0",X"30",X"00",X"F0",X"F0",X"10",
		X"00",X"F0",X"F0",X"00",X"00",X"E0",X"10",X"80",X"C0",X"F0",X"F0",X"30",X"00",X"C0",X"70",X"00",
		X"00",X"F0",X"F0",X"00",X"10",X"00",X"00",X"80",X"C0",X"F0",X"F0",X"30",X"00",X"E0",X"F0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
