library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity domino_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of domino_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"92",X"99",X"90",
		X"90",X"92",X"11",X"99",X"99",X"92",X"94",X"19",X"41",X"72",X"95",X"19",X"41",X"72",X"96",X"99",
		X"99",X"92",X"11",X"19",X"00",X"92",X"11",X"99",X"00",X"92",X"91",X"19",X"00",X"92",X"91",X"99",
		X"00",X"09",X"99",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"9A",X"00",X"00",X"09",X"9A",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"CC",X"00",X"00",
		X"09",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"90",X"00",X"99",X"CC",X"99",X"00",X"94",X"99",X"49",X"00",X"44",X"44",X"44",X"00",
		X"44",X"94",X"94",X"00",X"99",X"99",X"94",X"00",X"99",X"44",X"44",X"00",X"90",X"94",X"44",X"00",
		X"90",X"94",X"99",X"00",X"90",X"99",X"44",X"00",X"90",X"22",X"99",X"00",X"90",X"92",X"C9",X"00",
		X"99",X"99",X"C9",X"00",X"09",X"92",X"90",X"00",X"09",X"99",X"00",X"00",X"09",X"09",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"A9",X"90",X"00",X"00",X"A9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"9C",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"44",X"CC",X"90",X"00",X"44",X"99",X"99",X"00",X"49",X"44",X"49",X"00",
		X"49",X"94",X"44",X"00",X"49",X"99",X"94",X"00",X"99",X"44",X"94",X"00",X"C9",X"94",X"44",X"00",
		X"C9",X"94",X"44",X"00",X"99",X"99",X"99",X"00",X"00",X"22",X"44",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"49",X"00",X"99",X"99",X"49",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"94",X"99",X"00",X"99",X"94",X"99",X"00",
		X"99",X"94",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"91",X"00",X"29",X"00",
		X"91",X"00",X"91",X"00",X"99",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",
		X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"44",X"00",X"00",X"99",X"44",X"00",X"99",X"99",X"49",X"00",
		X"99",X"9D",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"C9",X"99",X"00",X"99",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"99",X"00",
		X"99",X"9D",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"09",X"44",X"99",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",
		X"09",X"49",X"49",X"00",X"09",X"99",X"99",X"00",X"09",X"22",X"99",X"00",X"09",X"99",X"29",X"00",
		X"00",X"19",X"29",X"00",X"00",X"11",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"11",X"19",X"00",X"00",X"11",X"19",X"00",X"00",X"19",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"44",X"44",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"49",X"49",X"00",
		X"09",X"99",X"99",X"00",X"09",X"22",X"29",X"00",X"09",X"92",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"22",X"19",X"00",X"00",X"99",X"11",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"19",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9A",X"00",X"00",X"99",X"9A",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"99",X"9A",X"00",X"00",X"C9",X"99",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"49",X"C9",X"00",X"00",X"99",X"99",X"00",X"90",X"44",X"44",X"00",
		X"90",X"44",X"44",X"00",X"90",X"99",X"99",X"00",X"99",X"99",X"49",X"00",X"29",X"44",X"99",X"00",
		X"29",X"44",X"92",X"90",X"99",X"99",X"29",X"99",X"29",X"99",X"99",X"19",X"22",X"00",X"99",X"19",
		X"92",X"00",X"99",X"99",X"99",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9A",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"C9",X"CC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"90",
		X"00",X"9C",X"99",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"CC",X"90",X"00",X"49",X"99",X"90",
		X"00",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"00",X"00",
		X"09",X"44",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"92",X"00",X"00",X"92",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"19",X"99",X"00",X"00",X"11",X"19",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"CC",X"90",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",
		X"09",X"C9",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"CC",X"00",X"00",
		X"99",X"C9",X"90",X"00",X"09",X"99",X"00",X"00",X"00",X"49",X"90",X"00",X"09",X"9F",X"90",X"00",
		X"09",X"99",X"90",X"00",X"99",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"49",X"44",X"99",X"00",
		X"49",X"49",X"99",X"00",X"49",X"99",X"99",X"00",X"44",X"49",X"99",X"00",X"99",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"09",X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"C9",X"99",X"00",X"00",X"C9",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"C9",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"94",X"CC",X"00",
		X"00",X"94",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"19",X"00",
		X"00",X"22",X"11",X"00",X"00",X"29",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"19",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"09",X"CC",X"99",X"00",X"09",X"CC",X"99",X"00",X"09",X"99",X"9C",X"00",X"09",X"44",X"CC",X"00",
		X"09",X"44",X"9C",X"00",X"09",X"44",X"99",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"99",X"49",X"00",
		X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"19",X"29",X"00",
		X"00",X"11",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"19",X"00",
		X"00",X"11",X"99",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"CC",X"99",X"00",X"09",X"CC",X"CC",X"00",X"09",X"99",X"CC",X"00",X"09",X"44",X"9C",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"49",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"9A",X"99",X"00",
		X"DD",X"92",X"99",X"00",X"99",X"99",X"CC",X"00",X"99",X"CC",X"9C",X"00",X"99",X"CC",X"CC",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"C9",X"00",X"99",X"99",X"99",X"00",X"99",X"CC",X"90",X"00",
		X"99",X"9C",X"99",X"00",X"99",X"99",X"49",X"00",X"99",X"49",X"49",X"00",X"99",X"99",X"44",X"00",
		X"99",X"94",X"49",X"00",X"DD",X"94",X"49",X"00",X"99",X"99",X"99",X"00",X"99",X"44",X"99",X"00",
		X"99",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"29",X"00",X"99",X"22",X"29",X"00",
		X"99",X"22",X"29",X"00",X"99",X"22",X"29",X"00",X"99",X"92",X"99",X"00",X"99",X"22",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"DD",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"9F",X"9C",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"94",X"00",X"00",X"99",X"94",X"00",X"00",X"9F",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"DD",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"91",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"99",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",
		X"00",X"99",X"49",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"09",X"99",X"90",X"00",X"09",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"49",X"49",X"90",X"00",X"99",X"44",X"90",X"00",
		X"90",X"44",X"90",X"00",X"90",X"44",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",
		X"00",X"22",X"19",X"00",X"00",X"22",X"19",X"00",X"00",X"22",X"19",X"00",X"00",X"92",X"19",X"00",
		X"00",X"99",X"19",X"00",X"00",X"09",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",
		X"09",X"99",X"00",X"00",X"09",X"CC",X"99",X"99",X"09",X"99",X"49",X"C9",X"09",X"99",X"49",X"99",
		X"09",X"44",X"99",X"00",X"09",X"44",X"00",X"00",X"09",X"49",X"90",X"00",X"09",X"94",X"90",X"00",
		X"09",X"99",X"90",X"00",X"09",X"11",X"90",X"00",X"99",X"11",X"99",X"00",X"99",X"11",X"22",X"00",
		X"C9",X"11",X"22",X"00",X"CC",X"11",X"99",X"00",X"C9",X"99",X"00",X"00",X"99",X"11",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"0A",X"00",X"00",X"CC",X"0A",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"99",X"00",
		X"09",X"CC",X"C9",X"00",X"09",X"C9",X"C9",X"00",X"09",X"C9",X"99",X"00",X"09",X"CC",X"49",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"49",X"00",X"00",X"94",X"49",X"00",X"00",X"44",X"49",X"00",
		X"09",X"49",X"49",X"00",X"09",X"99",X"99",X"00",X"09",X"CC",X"90",X"00",X"09",X"99",X"00",X"00",
		X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"49",X"90",X"00",X"09",X"94",X"90",X"00",
		X"09",X"99",X"90",X"00",X"09",X"11",X"90",X"00",X"99",X"11",X"99",X"00",X"99",X"11",X"22",X"00",
		X"C9",X"11",X"22",X"00",X"CC",X"11",X"99",X"00",X"C9",X"99",X"00",X"00",X"99",X"11",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",
		X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"D9",X"00",X"00",
		X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"00",
		X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"9F",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"9F",X"99",X"9F",X"00",X"DD",X"DD",X"DD",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"D9",X"00",
		X"00",X"99",X"9D",X"00",X"00",X"99",X"DD",X"00",X"00",X"D9",X"D9",X"00",X"00",X"DD",X"99",X"00",
		X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"DD",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"F9",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"D9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"C9",X"00",X"99",X"4E",X"C9",X"00",
		X"9C",X"4C",X"CC",X"00",X"9C",X"CC",X"C9",X"00",X"9C",X"9C",X"CC",X"00",X"99",X"99",X"C9",X"00",
		X"99",X"CC",X"C9",X"00",X"99",X"99",X"C9",X"00",X"99",X"F9",X"C9",X"90",X"99",X"99",X"C9",X"90",
		X"99",X"9F",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"44",X"99",X"90",X"99",X"CC",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"99",X"90",
		X"CC",X"49",X"9C",X"90",X"CC",X"49",X"9C",X"90",X"CC",X"44",X"9C",X"90",X"CC",X"44",X"99",X"90",
		X"CC",X"94",X"99",X"90",X"C9",X"99",X"9C",X"90",X"99",X"99",X"CC",X"00",X"C9",X"CC",X"CC",X"00",
		X"C9",X"CC",X"CC",X"00",X"C9",X"CC",X"EC",X"00",X"C9",X"CC",X"CE",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"BB",X"00",X"C9",X"BB",X"BB",X"00",X"C9",X"BB",X"BB",X"00",
		X"C9",X"BB",X"BB",X"00",X"C9",X"B9",X"BB",X"00",X"C9",X"99",X"BB",X"00",X"9B",X"B9",X"BB",X"00",
		X"BB",X"99",X"BB",X"00",X"BB",X"90",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"B9",X"00",X"BB",X"00",X"99",X"00",X"BB",X"00",X"EE",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",
		X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"99",X"00",X"BB",X"00",X"77",X"09",X"BB",X"00",
		X"97",X"09",X"99",X"00",X"99",X"09",X"BB",X"00",X"00",X"09",X"BB",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"09",X"00",X"00",X"79",X"99",X"00",X"00",X"79",X"95",X"00",X"00",X"79",X"55",X"00",X"00",
		X"99",X"55",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"99",X"99",X"00",X"55",X"99",X"55",X"00",
		X"55",X"95",X"55",X"00",X"55",X"55",X"95",X"90",X"59",X"55",X"95",X"90",X"59",X"55",X"95",X"90",
		X"99",X"55",X"55",X"90",X"00",X"59",X"55",X"90",X"00",X"59",X"55",X"90",X"00",X"55",X"55",X"90",
		X"00",X"55",X"95",X"90",X"00",X"55",X"95",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"55",X"00",
		X"00",X"95",X"55",X"00",X"00",X"99",X"59",X"00",X"00",X"79",X"99",X"00",X"00",X"97",X"99",X"00",
		X"00",X"99",X"59",X"00",X"00",X"59",X"55",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"79",X"90",X"00",X"00",X"79",X"99",X"00",X"90",X"99",X"59",X"00",X"90",
		X"55",X"59",X"00",X"90",X"55",X"59",X"00",X"90",X"55",X"59",X"99",X"90",X"55",X"59",X"55",X"90",
		X"55",X"55",X"55",X"90",X"59",X"55",X"55",X"90",X"59",X"95",X"95",X"00",X"99",X"95",X"95",X"00",
		X"09",X"99",X"95",X"00",X"09",X"55",X"55",X"00",X"99",X"59",X"55",X"00",X"77",X"59",X"55",X"90",
		X"79",X"55",X"95",X"99",X"99",X"55",X"95",X"79",X"95",X"99",X"99",X"99",X"59",X"00",X"09",X"99",
		X"59",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"44",X"99",X"00",X"00",X"49",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",
		X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"94",X"99",X"00",X"99",X"99",X"9F",X"00",X"99",X"49",X"99",X"00",X"99",X"94",X"99",X"00",
		X"99",X"44",X"99",X"00",X"99",X"9C",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"44",X"90",X"00",X"00",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"C9",X"00",X"00",X"94",X"CC",X"00",X"00",X"94",X"99",X"99",X"00",X"44",X"99",X"99",X"00",
		X"44",X"44",X"F9",X"00",X"49",X"44",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"99",X"00",
		X"99",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"92",X"99",X"00",
		X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"11",X"90",X"99",X"00",
		X"11",X"00",X"91",X"00",X"91",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"90",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"44",X"9C",X"90",X"00",X"94",X"CC",X"90",X"00",
		X"99",X"44",X"90",X"00",X"49",X"49",X"00",X"00",X"44",X"99",X"00",X"00",X"49",X"99",X"00",X"00",
		X"44",X"C9",X"00",X"00",X"94",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"90",X"29",X"00",X"99",X"90",X"29",X"00",X"11",X"90",X"99",X"00",
		X"11",X"00",X"91",X"00",X"91",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"30",X"00",X"F9",X"99",X"00",X"99",X"F9",X"99",X"00",
		X"9C",X"F9",X"9C",X"00",X"9C",X"F9",X"99",X"00",X"9C",X"9C",X"CC",X"00",X"99",X"9C",X"C9",X"00",
		X"99",X"C9",X"C9",X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",X"C9",X"00",X"99",X"99",X"C9",X"00",
		X"99",X"94",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"C9",X"99",X"90",X"99",X"CC",X"9D",X"90",
		X"99",X"99",X"9D",X"90",X"99",X"99",X"9D",X"90",X"C9",X"99",X"9D",X"90",X"CC",X"99",X"99",X"90",
		X"CC",X"49",X"99",X"90",X"CC",X"49",X"99",X"90",X"CC",X"44",X"99",X"90",X"99",X"99",X"99",X"90",
		X"00",X"99",X"90",X"99",X"09",X"90",X"99",X"09",X"99",X"90",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"A4",X"99",X"00",X"00",X"AA",X"49",X"00",X"99",X"9A",X"99",X"00",
		X"94",X"AA",X"94",X"00",X"94",X"44",X"49",X"00",X"94",X"94",X"44",X"00",X"99",X"99",X"49",X"00",
		X"99",X"44",X"49",X"00",X"99",X"99",X"49",X"00",X"99",X"9F",X"49",X"90",X"99",X"99",X"49",X"90",
		X"99",X"9F",X"99",X"90",X"99",X"9F",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"44",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"99",X"90",
		X"CC",X"49",X"9C",X"90",X"CC",X"49",X"9C",X"90",X"CC",X"44",X"9C",X"90",X"CC",X"44",X"99",X"90",
		X"CC",X"94",X"99",X"90",X"C9",X"99",X"9C",X"90",X"99",X"99",X"CC",X"00",X"C9",X"CC",X"CC",X"00",
		X"C9",X"CC",X"CC",X"00",X"C9",X"CC",X"EC",X"00",X"C9",X"CC",X"CE",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"FF",X"00",X"C9",X"44",X"F4",X"00",X"C9",X"FF",X"F4",X"00",
		X"C9",X"FF",X"FF",X"00",X"C9",X"9F",X"FF",X"00",X"C9",X"99",X"F4",X"00",X"99",X"99",X"F4",X"00",
		X"99",X"90",X"99",X"00",X"EE",X"90",X"EE",X"00",X"CC",X"99",X"EC",X"00",X"CC",X"C9",X"CE",X"00",
		X"9C",X"C9",X"C9",X"00",X"99",X"E9",X"E9",X"00",X"09",X"C9",X"CC",X"00",X"99",X"90",X"CE",X"00",
		X"9C",X"90",X"EC",X"00",X"99",X"00",X"CE",X"00",X"B9",X"00",X"EC",X"00",X"3B",X"00",X"9C",X"90",
		X"BB",X"90",X"99",X"90",X"BB",X"99",X"99",X"B0",X"99",X"BB",X"31",X"90",X"9B",X"BB",X"BB",X"90",
		X"99",X"B9",X"B9",X"90",X"99",X"99",X"99",X"00",X"BB",X"9B",X"9B",X"00",X"99",X"B9",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"09",X"00",X"91",X"00",X"99",X"00",X"99",X"90",X"2C",X"00",X"E9",X"90",X"2A",X"00",X"EE",X"90",
		X"2C",X"99",X"EE",X"99",X"CC",X"55",X"99",X"99",X"CC",X"99",X"45",X"49",X"CC",X"00",X"45",X"49",
		X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"69",X"00",X"45",X"49",
		X"66",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"66",X"00",X"45",X"09",
		X"99",X"00",X"47",X"99",X"AA",X"00",X"47",X"90",X"AA",X"00",X"47",X"00",X"AA",X"00",X"99",X"00",
		X"AA",X"00",X"59",X"00",X"AA",X"00",X"59",X"00",X"AA",X"00",X"99",X"00",X"AA",X"00",X"99",X"90",
		X"AA",X"00",X"95",X"99",X"99",X"00",X"95",X"B9",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"09",X"00",X"91",X"00",X"99",X"00",X"99",X"90",X"2C",X"00",X"E9",X"90",X"2A",X"00",X"EE",X"90",
		X"2C",X"99",X"99",X"99",X"CC",X"55",X"45",X"49",X"CC",X"99",X"45",X"49",X"CC",X"00",X"45",X"49",
		X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"69",X"00",X"45",X"49",
		X"66",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"66",X"00",X"47",X"99",
		X"66",X"00",X"47",X"90",X"99",X"00",X"47",X"00",X"AA",X"00",X"99",X"00",X"AA",X"00",X"59",X"00",
		X"AA",X"99",X"59",X"00",X"9A",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"99",X"00",
		X"90",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"90",X"00",X"99",X"00",X"90",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"4C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"09",X"00",X"09",X"CC",X"9A",X"00",X"99",X"CC",X"AA",X"00",X"9A",X"9C",X"AA",X"00",
		X"C9",X"99",X"AA",X"00",X"CC",X"AA",X"99",X"00",X"CC",X"A9",X"99",X"90",X"CC",X"99",X"99",X"90",
		X"C9",X"92",X"92",X"90",X"C9",X"AA",X"A2",X"90",X"99",X"AA",X"AA",X"99",X"00",X"AA",X"A9",X"09",
		X"99",X"AA",X"99",X"49",X"55",X"22",X"29",X"99",X"55",X"AA",X"AA",X"59",X"55",X"99",X"99",X"59",
		X"45",X"C9",X"90",X"59",X"45",X"90",X"90",X"59",X"45",X"00",X"90",X"59",X"59",X"00",X"90",X"59",
		X"59",X"00",X"90",X"59",X"99",X"00",X"90",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"A2",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"99",X"00",
		X"09",X"4C",X"9A",X"00",X"99",X"99",X"9A",X"00",X"9A",X"4C",X"9A",X"00",X"C9",X"CC",X"9A",X"00",
		X"CC",X"99",X"99",X"00",X"CC",X"AA",X"A9",X"90",X"CC",X"A9",X"99",X"90",X"C9",X"99",X"99",X"90",
		X"C9",X"92",X"92",X"90",X"99",X"AA",X"22",X"90",X"00",X"AA",X"A2",X"99",X"99",X"AA",X"AA",X"49",
		X"55",X"AA",X"AA",X"99",X"55",X"22",X"29",X"59",X"55",X"AA",X"AA",X"59",X"45",X"99",X"99",X"59",
		X"45",X"00",X"C9",X"59",X"45",X"00",X"C9",X"59",X"55",X"00",X"C9",X"59",X"55",X"00",X"99",X"59",
		X"99",X"00",X"22",X"99",X"00",X"00",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"09",X"44",X"99",X"00",
		X"99",X"44",X"AA",X"00",X"9A",X"44",X"AA",X"00",X"9A",X"94",X"AA",X"00",X"C9",X"99",X"AA",X"00",
		X"CC",X"99",X"99",X"00",X"CC",X"A9",X"A9",X"90",X"99",X"AA",X"A9",X"90",X"90",X"AA",X"AA",X"90",
		X"90",X"99",X"AA",X"90",X"90",X"AA",X"9A",X"90",X"00",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"09",
		X"55",X"AA",X"AA",X"99",X"55",X"AA",X"A9",X"59",X"55",X"AA",X"AA",X"59",X"45",X"99",X"99",X"59",
		X"45",X"00",X"C9",X"59",X"45",X"00",X"C9",X"59",X"55",X"00",X"C9",X"59",X"55",X"00",X"99",X"59",
		X"99",X"00",X"22",X"59",X"00",X"00",X"99",X"99",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"95",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"90",X"00",X"09",X"99",X"90",X"00",
		X"09",X"FF",X"99",X"00",X"99",X"FF",X"59",X"00",X"95",X"FF",X"55",X"00",X"95",X"FF",X"95",X"00",
		X"95",X"99",X"95",X"00",X"95",X"44",X"95",X"00",X"95",X"44",X"95",X"00",X"95",X"44",X"95",X"00",
		X"95",X"99",X"95",X"00",X"95",X"FF",X"95",X"00",X"95",X"FF",X"55",X"00",X"99",X"FF",X"59",X"00",
		X"09",X"FF",X"99",X"00",X"00",X"FF",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"29",X"09",X"00",X"09",X"92",X"99",X"00",X"09",X"99",X"94",X"00",
		X"09",X"A9",X"94",X"00",X"09",X"9C",X"99",X"00",X"09",X"C9",X"CC",X"00",X"09",X"C9",X"C9",X"00",
		X"D0",X"99",X"9C",X"00",X"D0",X"4C",X"99",X"00",X"00",X"CC",X"39",X"00",X"00",X"C9",X"99",X"00",
		X"90",X"99",X"90",X"00",X"99",X"39",X"00",X"00",X"55",X"39",X"00",X"00",X"55",X"39",X"90",X"00",
		X"99",X"33",X"99",X"00",X"96",X"39",X"66",X"00",X"96",X"99",X"66",X"00",X"96",X"39",X"66",X"00",
		X"66",X"99",X"66",X"90",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"99",X"22",X"99",X"99",
		X"97",X"22",X"77",X"29",X"77",X"66",X"75",X"D9",X"77",X"66",X"79",X"D9",X"79",X"66",X"9D",X"99",
		X"47",X"99",X"79",X"90",X"77",X"00",X"77",X"00",X"97",X"00",X"77",X"00",X"99",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"92",X"99",X"00",X"09",X"99",X"44",X"00",
		X"09",X"A9",X"54",X"00",X"09",X"CC",X"99",X"00",X"09",X"C9",X"C9",X"00",X"09",X"99",X"99",X"00",
		X"D0",X"45",X"90",X"00",X"D0",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"C9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"90",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"55",X"39",X"00",X"00",
		X"55",X"33",X"90",X"00",X"99",X"39",X"99",X"00",X"96",X"99",X"66",X"00",X"96",X"33",X"66",X"00",
		X"96",X"39",X"66",X"00",X"66",X"99",X"66",X"90",X"99",X"22",X"99",X"99",X"97",X"22",X"77",X"99",
		X"77",X"22",X"77",X"99",X"77",X"22",X"79",X"D9",X"79",X"66",X"9D",X"D9",X"79",X"66",X"99",X"69",
		X"57",X"66",X"79",X"99",X"55",X"99",X"77",X"90",X"95",X"00",X"77",X"00",X"99",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"99",X"00",
		X"09",X"99",X"EE",X"00",X"09",X"EE",X"AE",X"00",X"09",X"99",X"EE",X"00",X"09",X"EE",X"99",X"00",
		X"09",X"EE",X"EE",X"00",X"00",X"EE",X"E9",X"00",X"09",X"EE",X"99",X"00",X"99",X"EE",X"F9",X"00",
		X"9E",X"9E",X"F9",X"00",X"EE",X"9E",X"99",X"00",X"EE",X"99",X"90",X"00",X"EE",X"09",X"99",X"00",
		X"EE",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"EE",X"99",X"EE",X"00",
		X"9E",X"EE",X"AE",X"00",X"99",X"99",X"AE",X"00",X"09",X"EE",X"99",X"00",X"09",X"EE",X"E9",X"00",
		X"09",X"EE",X"E9",X"00",X"09",X"EE",X"99",X"00",X"00",X"9E",X"F9",X"00",X"00",X"9E",X"F9",X"00",
		X"00",X"9E",X"99",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9F",X"00",X"00",X"09",X"9F",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"9E",X"99",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"99",X"00",X"00",
		X"9E",X"99",X"00",X"00",X"9E",X"E9",X"00",X"00",X"9E",X"E9",X"00",X"00",X"EE",X"99",X"00",X"00",
		X"9E",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"40",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"D9",X"9A",X"00",X"A9",X"FD",X"99",X"90",X"AA",X"99",X"AA",X"90",
		X"99",X"99",X"2A",X"90",X"9A",X"99",X"99",X"90",X"AA",X"55",X"00",X"00",X"99",X"99",X"00",X"00",
		X"90",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",
		X"0F",X"A9",X"00",X"00",X"00",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"44",X"00",X"00",X"09",X"9C",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"55",X"90",X"00",
		X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"29",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"90",X"00",
		X"09",X"92",X"E9",X"00",X"09",X"99",X"E9",X"00",X"09",X"09",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",
		X"00",X"9C",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"77",X"90",X"00",X"00",X"77",X"90",X"00",
		X"00",X"97",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"2F",X"90",X"00",X"00",X"2F",X"90",X"00",
		X"00",X"9F",X"90",X"00",X"00",X"0F",X"90",X"00",X"00",X"0F",X"90",X"00",X"00",X"0F",X"90",X"00",
		X"99",X"99",X"00",X"00",X"C9",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"C9",X"00",X"00",X"90",X"C9",X"00",X"00",X"90",X"CC",X"00",X"00",X"90",X"99",X"00",X"00",
		X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",
		X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",
		X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"91",X"96",X"00",X"00",X"91",X"96",X"00",X"00",
		X"91",X"99",X"00",X"00",X"91",X"91",X"00",X"00",X"99",X"91",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"99",X"9C",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"92",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"99",X"92",X"99",X"99",X"99",X"92",X"99",X"99",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"69",X"00",
		X"00",X"99",X"66",X"99",X"00",X"66",X"66",X"99",X"00",X"99",X"99",X"19",X"00",X"99",X"99",X"19",
		X"00",X"66",X"09",X"99",X"00",X"66",X"00",X"90",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"99",X"00",X"00",X"77",X"99",X"00",X"00",X"74",X"99",X"90",
		X"00",X"44",X"49",X"90",X"00",X"99",X"49",X"90",X"00",X"49",X"99",X"90",X"00",X"44",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"9C",X"99",X"90",X"00",X"99",X"29",X"90",
		X"00",X"22",X"92",X"90",X"00",X"22",X"92",X"90",X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"29",X"99",X"00",
		X"00",X"99",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"69",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"96",X"99",X"00",X"00",X"96",X"11",X"00",X"00",X"96",X"11",X"00",X"00",X"96",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"99",X"99",X"00",X"00",X"9C",X"44",X"00",X"00",X"9C",X"44",X"99",X"99",X"99",X"94",X"99",X"99",
		X"09",X"A9",X"09",X"00",X"09",X"99",X"09",X"00",X"09",X"CC",X"09",X"00",X"09",X"C4",X"09",X"00",
		X"09",X"94",X"09",X"00",X"99",X"CC",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"92",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"19",X"00",X"00",X"09",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"66",X"00",X"44",X"00",X"66",X"00",X"44",X"00",X"66",X"00",X"44",X"00",X"99",X"00",
		X"99",X"00",X"77",X"00",X"EE",X"90",X"77",X"00",X"EE",X"90",X"77",X"00",X"4C",X"90",X"99",X"00",
		X"49",X"00",X"09",X"00",X"CC",X"00",X"90",X"00",X"9C",X"00",X"99",X"00",X"99",X"00",X"11",X"00",
		X"99",X"00",X"99",X"00",X"59",X"00",X"90",X"00",X"55",X"00",X"00",X"00",X"95",X"90",X"00",X"00",
		X"99",X"99",X"09",X"00",X"59",X"9C",X"99",X"00",X"55",X"CC",X"99",X"99",X"55",X"CC",X"77",X"49",
		X"99",X"99",X"44",X"49",X"11",X"00",X"44",X"49",X"11",X"09",X"44",X"99",X"11",X"99",X"44",X"90",
		X"11",X"99",X"94",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"09",X"00",X"00",X"90",X"09",X"00",X"90",X"00",X"09",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"09",X"99",X"44",X"00",X"97",X"79",X"44",X"00",X"77",X"79",X"44",X"90",X"77",X"79",
		X"99",X"90",X"77",X"79",X"EE",X"99",X"77",X"99",X"EE",X"C9",X"99",X"00",X"44",X"99",X"00",X"00",
		X"44",X"00",X"00",X"00",X"CC",X"00",X"90",X"99",X"99",X"00",X"99",X"39",X"59",X"00",X"33",X"19",
		X"59",X"00",X"11",X"39",X"55",X"00",X"99",X"99",X"95",X"90",X"00",X"00",X"95",X"99",X"99",X"00",
		X"99",X"9C",X"99",X"90",X"55",X"CC",X"99",X"99",X"55",X"CC",X"77",X"49",X"99",X"99",X"44",X"49",
		X"11",X"00",X"44",X"49",X"11",X"00",X"44",X"99",X"11",X"00",X"44",X"90",X"11",X"00",X"94",X"00",
		X"11",X"00",X"99",X"00",X"91",X"00",X"09",X"00",X"91",X"00",X"99",X"00",X"11",X"00",X"95",X"00",
		X"11",X"00",X"95",X"00",X"99",X"00",X"95",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",
		X"00",X"92",X"99",X"00",X"99",X"99",X"CC",X"00",X"9C",X"CC",X"9C",X"00",X"9C",X"CC",X"CC",X"00",
		X"CC",X"99",X"99",X"00",X"C9",X"99",X"C9",X"00",X"99",X"99",X"99",X"00",X"99",X"CC",X"90",X"00",
		X"09",X"9C",X"99",X"00",X"00",X"99",X"49",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"94",X"00",
		X"00",X"44",X"94",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"29",X"00",X"09",X"22",X"29",X"00",
		X"09",X"92",X"29",X"00",X"09",X"99",X"29",X"00",X"09",X"99",X"99",X"00",X"00",X"29",X"29",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"90",X"11",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",
		X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"97",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"94",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"D9",X"00",
		X"00",X"99",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
