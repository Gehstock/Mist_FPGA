library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"8C",X"4C",X"22",X"EE",X"4C",X"88",X"00",X"00",X"11",X"46",X"26",X"33",X"4C",X"9D",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"01",X"01",X"01",X"01",X"01",X"01",X"E1",X"E1",X"08",X"08",X"08",X"08",X"08",X"08",X"78",X"78",
		X"01",X"01",X"01",X"01",X"E1",X"E1",X"E1",X"E1",X"08",X"08",X"08",X"08",X"78",X"78",X"78",X"78",
		X"01",X"01",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"08",X"08",X"78",X"78",X"78",X"78",X"78",X"78",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",
		X"E1",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",X"78",X"78",X"08",X"08",X"08",X"08",X"08",X"08",
		X"E1",X"E1",X"E1",X"E1",X"01",X"01",X"01",X"01",X"78",X"78",X"78",X"78",X"08",X"08",X"08",X"08",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",X"01",X"78",X"78",X"78",X"78",X"78",X"78",X"08",X"08",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"FF",X"FF",X"44",X"44",X"44",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"66",X"33",X"11",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"77",X"00",
		X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"33",X"11",X"11",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"44",X"77",X"77",X"00",
		X"11",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"44",X"44",X"44",X"44",X"77",X"77",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"FF",X"FF",X"00",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"00",
		X"8F",X"8F",X"8F",X"CF",X"CF",X"8F",X"8F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"8F",X"CF",X"CF",X"8F",X"8F",X"0F",X"FF",X"FF",X"FF",X"77",X"BB",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"8F",X"CF",X"CF",X"8F",X"8F",X"0F",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"C7",X"EB",X"EB",X"C7",X"CF",X"CF",X"77",X"7E",X"3F",X"1F",X"1F",X"3F",X"76",X"77",
		X"CF",X"CF",X"8F",X"8F",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",
		X"00",X"00",X"00",X"01",X"8F",X"8F",X"CF",X"CF",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"30",X"70",X"78",X"3C",X"3C",X"78",X"70",X"30",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"1E",X"1E",X"1A",X"1E",X"1A",X"1E",X"F0",X"30",X"43",X"42",X"87",X"85",X"43",X"43",X"30",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"33",X"77",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"EE",X"CC",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"77",X"33",X"CC",X"EE",X"77",X"33",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"77",X"33",X"CC",X"EE",X"77",X"33",X"11",X"00",X"00",X"00",
		X"33",X"77",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"EE",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"88",X"22",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"33",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"EE",X"22",X"22",X"00",X"11",X"22",X"22",X"22",X"33",
		X"AA",X"AA",X"AA",X"22",X"00",X"00",X"00",X"EE",X"22",X"22",X"22",X"11",X"00",X"22",X"22",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"08",X"08",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",X"08",X"00",X"00",X"00",X"00",X"0F",X"0F",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"00",X"77",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"EE",X"EE",X"CC",X"88",X"00",
		X"00",X"00",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"BB",X"FF",X"11",X"11",X"33",X"11",X"22",X"33",X"33",X"33",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"55",X"BB",X"FF",X"11",X"11",X"33",X"11",X"22",X"33",X"33",X"33",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"0F",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"FF",X"FF",
		X"FF",X"EE",X"DD",X"BB",X"77",X"77",X"33",X"11",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"11",X"33",X"77",X"77",X"BB",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"FF",X"FF",X"FF",X"33",X"00",X"77",X"FF",X"FF",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"11",
		X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"EE",X"CC",X"CC",X"88",X"00",
		X"00",X"00",X"11",X"11",X"33",X"32",X"77",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"CF",X"8F",X"8F",X"01",X"00",X"00",X"00",X"FD",X"FA",X"FB",X"FD",X"F7",X"EE",X"88",X"00",
		X"00",X"00",X"00",X"01",X"8F",X"8F",X"CF",X"C7",X"00",X"88",X"EE",X"F7",X"FB",X"FD",X"FA",X"FD",
		X"61",X"34",X"1E",X"0F",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"02",X"00",X"00",X"00",
		X"C3",X"87",X"87",X"DF",X"DF",X"87",X"87",X"C3",X"00",X"00",X"30",X"F1",X"F1",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"1E",X"34",X"61",X"00",X"00",X"00",X"02",X"03",X"03",X"02",X"00",
		X"8F",X"0F",X"0F",X"8F",X"8F",X"0F",X"0F",X"8F",X"3F",X"0F",X"0F",X"BF",X"BF",X"0F",X"0F",X"3F",
		X"08",X"08",X"0F",X"0F",X"0F",X"88",X"88",X"CC",X"0A",X"0F",X"0F",X"0F",X"19",X"19",X"77",X"11",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"00",X"00",X"88",X"CC",X"EE",X"EE",X"77",X"BB",
		X"FF",X"77",X"32",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"88",X"88",X"0F",X"0F",X"0F",X"08",X"08",X"11",X"77",X"19",X"19",X"0F",X"0F",X"0F",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"22",X"33",X"00",X"33",X"77",X"FF",X"66",X"60",X"30",X"10",X"00",X"44",X"66",X"CC",X"44",
		X"00",X"00",X"88",X"F3",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"00",X"00",X"10",X"13",X"43",X"70",
		X"E1",X"E1",X"C0",X"C8",X"EC",X"C8",X"80",X"00",X"70",X"30",X"10",X"31",X"73",X"73",X"30",X"00",
		X"00",X"00",X"00",X"62",X"62",X"62",X"48",X"08",X"00",X"00",X"66",X"60",X"60",X"60",X"69",X"69",
		X"00",X"08",X"0C",X"60",X"62",X"44",X"00",X"00",X"69",X"69",X"69",X"60",X"60",X"66",X"00",X"00",
		X"00",X"00",X"08",X"C0",X"80",X"88",X"C0",X"E1",X"00",X"70",X"F4",X"E3",X"53",X"34",X"70",X"F0",
		X"E1",X"A0",X"A0",X"80",X"C4",X"00",X"00",X"00",X"F0",X"F6",X"F6",X"30",X"10",X"11",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"08",X"79",X"79",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"69",
		X"79",X"19",X"08",X"08",X"08",X"00",X"00",X"00",X"69",X"3C",X"34",X"30",X"33",X"00",X"00",X"00",
		X"33",X"22",X"77",X"C0",X"C0",X"C0",X"C0",X"C0",X"33",X"66",X"CC",X"CC",X"F0",X"F0",X"F0",X"40",
		X"99",X"88",X"00",X"00",X"00",X"00",X"CC",X"88",X"00",X"11",X"00",X"00",X"00",X"66",X"CC",X"99",
		X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"00",X"88",X"CC",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"8F",X"03",X"03",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"CC",X"EE",X"44",X"01",X"07",X"0F",X"0F",X"0F",
		X"77",X"7B",X"7B",X"7B",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"01",X"03",X"03",X"30",X"30",X"70",
		X"00",X"00",X"00",X"44",X"66",X"66",X"66",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"33",X"00",X"00",X"33",X"77",X"FF",X"66",X"60",X"30",X"10",X"00",X"44",X"66",X"CC",X"44",
		X"88",X"00",X"33",X"E6",X"C3",X"C0",X"C0",X"F3",X"77",X"77",X"CC",X"CC",X"F0",X"F0",X"F0",X"40",
		X"88",X"88",X"00",X"33",X"77",X"EE",X"CC",X"CC",X"00",X"11",X"00",X"00",X"00",X"00",X"11",X"33",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"8F",X"03",X"8B",X"07",X"07",X"0F",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"7B",X"7B",X"7B",X"33",X"70",X"30",X"30",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",
		X"88",X"CC",X"44",X"00",X"00",X"00",X"88",X"99",X"99",X"CC",X"66",X"00",X"00",X"00",X"11",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"77",X"22",X"33",X"40",X"F0",X"F0",X"F0",X"CC",X"CC",X"66",X"33",
		X"66",X"FF",X"77",X"33",X"00",X"33",X"22",X"77",X"44",X"CC",X"66",X"44",X"00",X"10",X"30",X"60",
		X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"01",X"44",X"EE",X"CC",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"8F",X"07",X"0F",
		X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"00",X"CC",X"88",X"01",X"07",X"0F",X"0F",X"0F",
		X"77",X"66",X"66",X"66",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"7B",X"7B",X"7B",X"77",X"70",X"30",X"30",X"03",X"03",X"01",X"00",X"00",
		X"CC",X"CC",X"EE",X"77",X"33",X"00",X"88",X"99",X"33",X"11",X"00",X"00",X"00",X"00",X"11",X"00",
		X"F3",X"C0",X"C0",X"F3",X"E6",X"33",X"00",X"88",X"40",X"F0",X"F0",X"F0",X"CC",X"EE",X"77",X"77",
		X"66",X"FF",X"77",X"33",X"00",X"00",X"33",X"66",X"44",X"CC",X"66",X"44",X"00",X"10",X"30",X"60",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"8B",X"03",X"8F",X"07",X"0F",
		X"00",X"40",X"F0",X"F0",X"3C",X"1E",X"1E",X"3C",X"50",X"50",X"50",X"70",X"E1",X"C3",X"C3",X"E1",
		X"70",X"70",X"70",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"00",X"80",X"D0",X"F0",X"F0",X"F0",
		X"F0",X"F7",X"F7",X"FF",X"FF",X"FF",X"11",X"00",X"F0",X"F0",X"F0",X"70",X"31",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"EE",X"FF",X"00",X"E0",X"80",X"88",X"EE",X"FF",X"FF",X"FF",X"00",
		X"33",X"33",X"11",X"11",X"11",X"11",X"11",X"33",X"88",X"CC",X"CC",X"CC",X"EE",X"EE",X"EE",X"7F",
		X"FF",X"FF",X"CC",X"FF",X"FF",X"CC",X"FF",X"FF",X"00",X"88",X"88",X"88",X"88",X"88",X"99",X"BB",
		X"FF",X"FE",X"F0",X"F0",X"F0",X"10",X"00",X"00",X"3F",X"3D",X"3C",X"F0",X"F0",X"B0",X"90",X"90",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F3",X"F3",X"F0",X"F0",X"F0",X"F0",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"77",X"77",X"33",
		X"11",X"33",X"77",X"EE",X"EE",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"DD",X"FF",X"FF",X"F3",X"F0",X"F0",X"30",X"90",X"33",X"11",X"16",X"1E",X"3C",X"F0",X"B0",X"90",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"EC",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"88",X"88",X"CC",X"CC",X"EE",X"FF",X"FF",X"77",
		X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"FE",X"FC",X"66",X"33",X"11",X"00",X"00",X"00",X"11",X"33",
		X"FF",X"FF",X"F0",X"87",X"87",X"F0",X"70",X"10",X"73",X"71",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F8",X"F0",X"F0",X"80",X"F0",X"C0",X"00",X"F0",X"FF",X"FF",X"F0",X"F0",X"78",X"F0",X"F0",X"F0",
		X"33",X"33",X"11",X"11",X"11",X"11",X"11",X"33",X"88",X"CC",X"CC",X"CC",X"EE",X"EE",X"EE",X"7F",
		X"FF",X"FF",X"CC",X"FF",X"FF",X"CC",X"FF",X"FF",X"00",X"88",X"88",X"88",X"88",X"88",X"99",X"BB",
		X"FF",X"FE",X"F0",X"F0",X"F0",X"10",X"00",X"00",X"3F",X"3D",X"3C",X"F0",X"F0",X"B0",X"90",X"90",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F3",X"F3",X"F0",X"F0",X"F0",X"F0",X"30",X"00",
		X"66",X"33",X"11",X"11",X"11",X"33",X"77",X"FF",X"33",X"66",X"66",X"EE",X"EE",X"EE",X"2E",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"CC",X"CC",X"88",
		X"FE",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"10",X"79",X"F0",X"F0",X"F0",X"70",X"50",X"50",X"10",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"01",X"83",X"87",X"1E",X"1E",X"0F",X"0F",X"C0",X"F0",X"F0",X"F0",X"70",X"10",X"10",X"D0",
		X"00",X"08",X"0C",X"0E",X"0F",X"07",X"0F",X"0F",X"00",X"0F",X"0F",X"09",X"C0",X"C0",X"0F",X"0F",
		X"3F",X"FF",X"FF",X"FE",X"FE",X"8F",X"0F",X"0F",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"90",X"F0",
		X"0F",X"03",X"88",X"CC",X"EE",X"FF",X"77",X"7F",X"CF",X"FF",X"FF",X"F7",X"91",X"0E",X"0F",X"0F",
		X"1F",X"1E",X"1E",X"87",X"C3",X"61",X"00",X"00",X"F0",X"F0",X"F0",X"70",X"10",X"00",X"00",X"00",
		X"3F",X"1F",X"8F",X"07",X"07",X"0F",X"0F",X"0E",X"EF",X"FF",X"F3",X"48",X"0C",X"0F",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"40",X"40",X"60",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"30",X"10",X"00",X"00",X"30",X"30",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"F0",X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"70",X"70",X"70",X"70",X"70",X"60",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",
		X"F4",X"F0",X"F0",X"F3",X"F4",X"FB",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FC",X"F2",X"FD",X"E2",X"CC",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F4",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F4",X"F4",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F2",X"F2",X"F2",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",
		X"0C",X"0C",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"0F",X"F0",X"F0",X"F4",X"F4",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",X"08",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"01",X"01",
		X"08",X"08",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",X"08",X"00",X"00",X"00",X"00",X"0F",X"0F",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"F0",X"F0",X"F3",X"F4",X"FB",X"74",X"33",X"0F",X"0E",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F4",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",X"0F",X"0E",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"F4",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"08",X"08",X"0C",X"0F",X"0F",
		X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"00",X"00",X"00",X"08",X"08",X"0C",X"0E",X"0F",
		X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",
		X"F4",X"F0",X"F0",X"F3",X"F4",X"FB",X"74",X"33",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0F",X"0F",X"F4",X"FB",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"0F",X"F2",X"FD",X"E2",X"CC",
		X"30",X"70",X"F0",X"F0",X"0F",X"0F",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"C0",X"C0",X"80",X"00",X"80",X"10",X"30",X"10",X"00",X"00",X"10",X"30",X"10",
		X"C0",X"60",X"C0",X"00",X"00",X"C0",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",X"08",X"C0",X"E0",X"F0",X"F0",X"0F",X"0F",X"01",X"01",
		X"0C",X"0E",X"02",X"02",X"02",X"0E",X"0E",X"00",X"06",X"0F",X"09",X"09",X"09",X"0F",X"0F",X"00",
		X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"80",X"C0",X"3F",X"0F",X"87",X"C3",X"61",X"30",X"10",X"00",
		X"C0",X"80",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"00",X"10",X"30",X"61",X"C3",X"87",X"0F",X"3F",
		X"88",X"88",X"CC",X"FF",X"77",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"77",X"EE",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"FF",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"77",X"33",X"33",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"02",X"02",X"0E",X"0E",X"00",X"00",X"08",X"09",X"09",X"09",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"0F",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"0F",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",X"0F",X"78",X"78",X"78",X"78",X"78",X"78",X"08",X"0F",
		X"E1",X"E1",X"E1",X"E1",X"01",X"01",X"01",X"0F",X"78",X"78",X"78",X"78",X"08",X"08",X"08",X"0F",
		X"E1",X"E1",X"01",X"01",X"01",X"01",X"01",X"0F",X"78",X"78",X"08",X"08",X"08",X"08",X"08",X"0F",
		X"0C",X"0C",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0C",X"0C",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",
		X"F0",X"F0",X"F2",X"F2",X"F2",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E8",X"E4",X"EA",X"C4",X"88",
		X"F4",X"F4",X"F4",X"F4",X"F0",X"F0",X"F0",X"F0",X"80",X"C0",X"E8",X"E8",X"EC",X"E4",X"E4",X"E0",
		X"08",X"08",X"0F",X"0F",X"F2",X"F2",X"F0",X"F0",X"01",X"01",X"0F",X"0F",X"E8",X"E8",X"E0",X"E0",
		X"F0",X"F0",X"F2",X"F2",X"0F",X"0F",X"08",X"08",X"E0",X"E0",X"E0",X"E0",X"0F",X"0F",X"01",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",X"E8",X"E8",X"E8",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F4",X"F4",X"E8",X"E8",X"E8",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"0C",X"0C",X"0F",X"0F",X"F4",X"FB",X"74",X"33",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"30",X"70",X"F0",X"F0",X"0F",X"0F",X"0C",X"0C",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"0F",X"78",X"78",X"78",X"78",X"78",X"78",X"78",
		X"0F",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"78",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0F",X"E1",X"E1",X"E1",X"01",X"01",X"01",X"01",X"0F",X"78",X"78",X"78",X"08",X"08",X"08",X"08",
		X"0F",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",X"01",X"0F",X"78",X"78",X"78",X"78",X"78",X"08",X"08",
		X"00",X"01",X"03",X"07",X"D2",X"F0",X"F0",X"3F",X"A0",X"A0",X"B0",X"F0",X"70",X"70",X"76",X"77",
		X"40",X"40",X"40",X"E0",X"F0",X"F0",X"F0",X"F7",X"20",X"60",X"C0",X"80",X"F0",X"F0",X"F0",X"89",
		X"1F",X"07",X"03",X"88",X"88",X"CC",X"EE",X"66",X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"E6",X"EE",X"EE",X"CC",X"CC",X"CC",X"88",X"CC",X"EE",X"FF",X"77",X"33",X"11",X"00",X"00",
		X"00",X"01",X"03",X"07",X"1F",X"3C",X"F0",X"F0",X"00",X"00",X"A0",X"A0",X"B0",X"F0",X"70",X"70",
		X"00",X"00",X"40",X"40",X"40",X"E0",X"F0",X"F0",X"00",X"00",X"20",X"60",X"C0",X"80",X"F0",X"F0",
		X"F1",X"3F",X"1F",X"07",X"03",X"00",X"88",X"88",X"76",X"77",X"23",X"11",X"00",X"00",X"00",X"00",
		X"F0",X"F7",X"F7",X"E6",X"66",X"33",X"11",X"00",X"F0",X"89",X"88",X"CC",X"66",X"33",X"99",X"CC",
		X"60",X"C0",X"80",X"00",X"F0",X"C0",X"00",X"00",X"0E",X"0F",X"6F",X"FF",X"F0",X"F0",X"F0",X"FF",
		X"00",X"08",X"0E",X"CF",X"F0",X"F0",X"87",X"1E",X"00",X"00",X"10",X"1E",X"F0",X"F0",X"0E",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"0F",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"78",X"F3",X"00",X"00",X"00",X"00",X"00",X"C4",X"FF",X"CC",X"66",X"22",X"22",X"22",X"33",
		X"00",X"70",X"C0",X"80",X"E0",X"08",X"00",X"77",X"0E",X"0F",X"6F",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"00",X"08",X"0E",X"8F",X"FF",X"F0",X"F0",X"C3",X"00",X"00",X"10",X"1E",X"F0",X"C3",X"87",X"2C",
		X"44",X"FF",X"CC",X"66",X"22",X"22",X"22",X"33",X"FF",X"FF",X"EF",X"0F",X"0E",X"00",X"00",X"00",
		X"CF",X"9E",X"1E",X"08",X"00",X"00",X"00",X"00",X"E0",X"F3",X"F7",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E1",X"E7",X"CF",X"0F",X"0C",X"00",X"00",X"00",X"00",X"70",X"10",X"40",X"60",X"20",
		X"80",X"C0",X"60",X"30",X"B0",X"F0",X"E0",X"E0",X"11",X"10",X"30",X"F0",X"F1",X"C3",X"07",X"00",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"00",X"00",X"B0",X"90",X"B0",X"F0",X"70",X"31",X"11",X"00",
		X"E0",X"F3",X"F3",X"F3",X"F0",X"BE",X"CC",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"40",X"40",X"40",X"C0",X"C0",X"08",X"08",X"7F",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"17",
		X"00",X"00",X"00",X"0F",X"0F",X"7F",X"FF",X"FC",X"10",X"10",X"12",X"1E",X"3C",X"F8",X"F0",X"E1",
		X"44",X"FF",X"CC",X"66",X"22",X"22",X"22",X"33",X"17",X"16",X"3C",X"F0",X"F1",X"C3",X"07",X"00",
		X"F0",X"F0",X"E1",X"E7",X"CF",X"0F",X"0C",X"00",X"87",X"3C",X"79",X"48",X"08",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"70",X"10",X"40",X"60",X"20",
		X"1E",X"D2",X"5A",X"70",X"F0",X"F0",X"F0",X"E0",X"F3",X"F3",X"C3",X"87",X"86",X"84",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"00",X"00",X"B0",X"90",X"B0",X"F0",X"70",X"31",X"11",X"00",
		X"E0",X"F3",X"F3",X"F3",X"F0",X"BE",X"CC",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"30",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"A0",X"A0",X"A0",X"E1",X"E1",X"E1",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"48",X"68",X"68",
		X"44",X"FF",X"CC",X"66",X"2A",X"2A",X"2A",X"3F",X"03",X"03",X"07",X"17",X"17",X"17",X"07",X"03",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"3C",X"2C",X"3C",X"9E",X"9E",X"CF",X"CF",X"EF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0A",X"41",X"C1",X"90",X"70",X"10",X"00",X"00",X"01",X"02",X"14",X"04",X"02",X"04",
		X"06",X"0A",X"01",X"00",X"90",X"E0",X"20",X"10",X"06",X"09",X"80",X"80",X"90",X"A0",X"40",X"00",
		X"21",X"C3",X"61",X"30",X"10",X"01",X"02",X"0C",X"38",X"08",X"08",X"06",X"01",X"01",X"00",X"00",
		X"F0",X"00",X"10",X"30",X"E0",X"02",X"0D",X"00",X"00",X"80",X"50",X"A0",X"20",X"20",X"05",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0C",X"06",X"00",X"00",X"00",X"00",X"C0",X"60",X"80",X"41",X"00",
		X"10",X"20",X"60",X"80",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"20",X"C0",X"80",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"24",X"E1",X"41",X"81",X"70",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"0A",X"04",X"38",X"04",X"08",X"00",X"0D",X"02",X"40",X"60",X"90",X"C0",X"20",
		X"21",X"41",X"E1",X"81",X"82",X"04",X"08",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"02",X"0D",X"01",X"01",X"00",X"00",X"C0",X"90",X"40",X"C0",X"00",X"0C",X"03",X"00",
		X"00",X"20",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0D",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"80",X"60",X"00",X"02",X"0C",X"06",X"00",X"00",X"00",X"80",X"00",
		X"00",X"04",X"0A",X"41",X"C1",X"90",X"70",X"10",X"00",X"00",X"01",X"02",X"14",X"04",X"02",X"04",
		X"06",X"0A",X"01",X"00",X"90",X"E0",X"20",X"10",X"06",X"09",X"80",X"80",X"90",X"A0",X"40",X"00",
		X"21",X"C3",X"61",X"30",X"10",X"01",X"02",X"0C",X"38",X"08",X"08",X"06",X"01",X"01",X"00",X"00",
		X"F0",X"00",X"10",X"30",X"E0",X"02",X"0D",X"00",X"00",X"80",X"50",X"A0",X"20",X"20",X"05",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"06",X"00",X"00",X"00",X"00",X"0C",X"06",X"01",X"00",
		X"00",X"00",X"00",X"60",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"B0",X"00",X"00",
		X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"09",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"24",X"E1",X"41",X"81",X"70",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"0A",X"04",X"38",X"04",X"08",X"00",X"0D",X"02",X"40",X"60",X"90",X"C0",X"20",
		X"21",X"41",X"E1",X"81",X"82",X"04",X"08",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"02",X"0D",X"01",X"01",X"00",X"00",X"C0",X"90",X"40",X"C0",X"00",X"0C",X"03",X"00",
		X"CF",X"CF",X"CF",X"8F",X"8F",X"9E",X"1E",X"7F",X"F0",X"F0",X"F0",X"FC",X"FC",X"BC",X"75",X"33",
		X"41",X"E1",X"C3",X"F0",X"F0",X"F0",X"CB",X"CF",X"F8",X"F0",X"F0",X"F0",X"F1",X"F3",X"FF",X"6F",
		X"7C",X"FF",X"FC",X"F6",X"E2",X"22",X"22",X"33",X"33",X"33",X"11",X"11",X"11",X"00",X"00",X"00",
		X"CD",X"CD",X"CC",X"CC",X"CC",X"CC",X"CC",X"44",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",
		X"90",X"F0",X"C2",X"C2",X"C3",X"C3",X"C7",X"CF",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"B0",
		X"00",X"00",X"00",X"00",X"81",X"C1",X"41",X"41",X"70",X"03",X"07",X"0F",X"3E",X"7E",X"7C",X"FC",
		X"CF",X"CF",X"CF",X"8F",X"8F",X"9E",X"1E",X"7F",X"F0",X"F0",X"F0",X"FC",X"FC",X"BC",X"75",X"33",
		X"41",X"E1",X"C3",X"F0",X"F0",X"F0",X"CB",X"CF",X"F8",X"F0",X"F0",X"F0",X"F1",X"F3",X"FF",X"6F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"C0",X"E0",X"F0",X"00",X"00",X"03",X"02",X"02",X"02",X"02",X"03",
		X"00",X"11",X"33",X"77",X"FF",X"BD",X"3C",X"3C",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",
		X"87",X"0E",X"0C",X"08",X"08",X"00",X"00",X"00",X"03",X"06",X"04",X"04",X"06",X"0F",X"00",X"00",
		X"3C",X"3C",X"1E",X"0F",X"07",X"03",X"01",X"00",X"F0",X"F0",X"E1",X"C3",X"0F",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"80",X"80",X"0C",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"03",
		X"00",X"11",X"33",X"70",X"F0",X"96",X"0F",X"0F",X"00",X"EE",X"FF",X"FE",X"F0",X"F0",X"E1",X"0F",
		X"0F",X"0E",X"0C",X"08",X"08",X"00",X"00",X"00",X"03",X"06",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0E",X"0F",X"00",X"00",X"0F",X"06",X"04",X"04",X"06",X"03",
		X"00",X"10",X"30",X"07",X"0F",X"0F",X"0F",X"0F",X"00",X"E0",X"F0",X"E1",X"0F",X"0F",X"0F",X"0F",
		X"7F",X"EE",X"CC",X"88",X"88",X"00",X"00",X"00",X"03",X"02",X"02",X"02",X"02",X"03",X"00",X"00",
		X"0F",X"2F",X"AF",X"FF",X"77",X"33",X"11",X"00",X"0F",X"0F",X"1F",X"3F",X"FF",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"08",X"08",X"CC",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"03",
		X"00",X"01",X"03",X"07",X"0F",X"2F",X"3F",X"3F",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"1F",X"FF",
		X"F8",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"03",X"02",X"03",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3D",X"B5",X"F0",X"70",X"30",X"10",X"00",X"FF",X"FF",X"FE",X"FC",X"F0",X"F0",X"E0",X"00",
		X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"E1",X"C0",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"20",X"30",X"30",X"20",X"0F",X"0F",X"78",X"3C",X"10",X"20",X"E0",X"00",
		X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"01",X"03",X"07",X"0E",X"0C",X"0C",X"0C",X"08",X"09",X"0B",X"03",X"23",X"67",X"FF",X"FF",X"67",
		X"0F",X"0F",X"E1",X"C3",X"90",X"F0",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"20",X"30",X"30",X"20",X"47",X"07",X"70",X"30",X"10",X"30",X"E0",X"00",
		X"08",X"0C",X"0E",X"0F",X"0F",X"87",X"87",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"32",X"22",X"00",X"00",X"11",X"11",X"00",X"0F",X"0F",X"03",X"01",X"01",X"F0",X"F0",X"01",
		X"0E",X"E0",X"E0",X"F0",X"F2",X"F2",X"F0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"B8",X"88",X"F0",X"F0",X"63",X"03",X"10",
		X"08",X"0E",X"0F",X"CF",X"C3",X"C3",X"C3",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"32",X"33",X"11",X"00",X"00",X"03",X"07",X"0F",X"0D",X"81",X"89",X"01",X"01",
		X"0E",X"E0",X"E0",X"F0",X"F2",X"F2",X"F0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"B8",X"88",X"F0",X"F0",X"63",X"03",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"0E",X"0C",X"08",X"08",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"21",
		X"08",X"0C",X"0C",X"0C",X"0E",X"0E",X"8E",X"8F",X"00",X"00",X"01",X"03",X"07",X"0F",X"0E",X"0C",
		X"0C",X"8F",X"88",X"88",X"8F",X"0C",X"07",X"00",X"70",X"71",X"77",X"77",X"FF",X"BB",X"AA",X"AA",
		X"8F",X"FF",X"FF",X"FF",X"EE",X"44",X"44",X"44",X"19",X"FF",X"FF",X"FF",X"99",X"CC",X"66",X"22",
		X"00",X"00",X"08",X"08",X"00",X"07",X"04",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"21",
		X"00",X"00",X"00",X"01",X"03",X"06",X"8E",X"8F",X"00",X"00",X"0C",X"09",X"03",X"06",X"0C",X"08",
		X"88",X"88",X"88",X"88",X"88",X"0F",X"04",X"07",X"70",X"71",X"77",X"77",X"FF",X"BB",X"AA",X"AA",
		X"8F",X"FF",X"FF",X"FF",X"EE",X"44",X"44",X"44",X"19",X"FF",X"FF",X"FF",X"99",X"CC",X"66",X"22",
		X"00",X"00",X"06",X"08",X"0E",X"08",X"06",X"88",X"00",X"11",X"33",X"33",X"11",X"33",X"47",X"CF",
		X"00",X"FF",X"FF",X"FF",X"CF",X"FF",X"C7",X"6F",X"00",X"CC",X"EE",X"88",X"CF",X"EE",X"FF",X"3F",
		X"88",X"88",X"06",X"08",X"0E",X"08",X"06",X"00",X"FF",X"CF",X"47",X"33",X"11",X"33",X"33",X"11",
		X"FF",X"E7",X"4F",X"FF",X"CF",X"FF",X"FF",X"FF",X"0F",X"3F",X"FF",X"EE",X"CF",X"88",X"EE",X"CC",
		X"00",X"01",X"02",X"04",X"0F",X"8C",X"02",X"89",X"00",X"00",X"00",X"00",X"00",X"33",X"47",X"CF",
		X"00",X"77",X"FF",X"FF",X"77",X"FF",X"4F",X"E7",X"00",X"FF",X"FF",X"EE",X"3F",X"FF",X"FF",X"3F",
		X"88",X"89",X"02",X"8C",X"0F",X"04",X"02",X"01",X"FF",X"CF",X"47",X"33",X"00",X"00",X"00",X"00",
		X"FF",X"6F",X"C7",X"FF",X"77",X"FF",X"FF",X"77",X"0F",X"3F",X"FF",X"FF",X"3F",X"EE",X"FF",X"FF",
		X"00",X"07",X"0C",X"8F",X"88",X"88",X"8F",X"0C",X"AA",X"AA",X"BB",X"FF",X"77",X"77",X"71",X"70",
		X"44",X"44",X"44",X"EE",X"FF",X"FF",X"FF",X"8F",X"22",X"66",X"CC",X"99",X"FF",X"FF",X"FF",X"19",
		X"07",X"00",X"00",X"08",X"08",X"0C",X"0E",X"06",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"8E",X"0E",X"0E",X"0C",X"0C",X"0C",X"08",X"0C",X"0E",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"07",X"04",X"0F",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"BB",X"FF",X"77",X"77",X"71",X"70",
		X"44",X"44",X"44",X"EE",X"FF",X"FF",X"FF",X"8F",X"22",X"66",X"CC",X"99",X"FF",X"FF",X"FF",X"19",
		X"0F",X"04",X"07",X"00",X"08",X"08",X"00",X"00",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"8E",X"06",X"03",X"01",X"00",X"00",X"00",X"08",X"0C",X"06",X"03",X"09",X"0C",X"00",X"00",
		X"00",X"00",X"06",X"08",X"0E",X"08",X"06",X"88",X"00",X"11",X"33",X"33",X"11",X"33",X"65",X"CF",
		X"00",X"FF",X"FF",X"FF",X"CF",X"FF",X"4F",X"6F",X"00",X"CC",X"EE",X"88",X"CF",X"EE",X"FF",X"3F",
		X"88",X"88",X"06",X"08",X"0E",X"08",X"06",X"00",X"FF",X"ED",X"47",X"33",X"11",X"33",X"33",X"11",
		X"FF",X"6F",X"4F",X"FF",X"CF",X"FF",X"FF",X"FF",X"0F",X"3F",X"FF",X"EE",X"CF",X"88",X"EE",X"CC",
		X"00",X"01",X"02",X"04",X"0F",X"8C",X"02",X"89",X"00",X"00",X"00",X"00",X"00",X"33",X"47",X"ED",
		X"00",X"77",X"FF",X"FF",X"77",X"FF",X"4F",X"6F",X"00",X"FF",X"FF",X"EE",X"3F",X"FF",X"FF",X"3F",
		X"88",X"89",X"02",X"8C",X"0F",X"04",X"02",X"01",X"FF",X"CF",X"65",X"33",X"00",X"00",X"00",X"00",
		X"FF",X"6F",X"4F",X"FF",X"77",X"FF",X"FF",X"77",X"0F",X"3F",X"FF",X"FF",X"3F",X"EE",X"FF",X"70",
		X"00",X"00",X"00",X"31",X"35",X"3D",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"A0",X"A1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"69",X"69",
		X"0C",X"0C",X"0C",X"E0",X"EE",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"0F",X"0F",X"0F",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"F5",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"A0",X"A1",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"78",
		X"F5",X"3D",X"19",X"00",X"00",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"78",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"62",X"6A",X"6A",X"48",X"08",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"0F",X"0F",
		X"08",X"0C",X"3C",X"34",X"31",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"69",X"69",X"3C",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"35",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"66",X"60",X"60",X"60",X"0F",X"0F",
		X"08",X"0C",X"1E",X"71",X"62",X"44",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"C0",X"00",X"00",X"69",X"69",X"69",X"60",X"60",X"66",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"3D",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"A0",X"A1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"E0",X"EE",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"69",X"69",X"3C",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"62",X"6A",X"6A",X"48",X"08",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"69",X"69",
		X"08",X"0C",X"3D",X"35",X"31",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"0F",X"0F",X"0F",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"35",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"66",X"60",X"60",X"60",X"69",X"69",
		X"08",X"0C",X"1E",X"71",X"62",X"44",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"C0",X"00",X"00",X"0F",X"0F",X"0F",X"60",X"60",X"66",X"00",X"00",
		X"00",X"00",X"00",X"44",X"4C",X"4C",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"31",X"B2",X"F2",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"C0",X"C0",X"40",X"0F",X"0F",
		X"08",X"08",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"0F",X"0F",X"40",X"C8",X"C8",X"C8",X"00",X"00",
		X"00",X"00",X"00",X"26",X"2E",X"2E",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"11",X"91",X"D1",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"C0",X"C0",X"40",X"0F",X"0F",
		X"08",X"08",X"2E",X"2E",X"26",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"D1",X"91",X"11",X"00",X"00",X"0F",X"0F",X"40",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"17",X"1F",X"1F",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"C8",X"C8",X"C8",X"40",X"0F",X"0F",
		X"08",X"08",X"4C",X"4C",X"44",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"F2",X"B2",X"32",X"00",X"00",X"0F",X"0F",X"40",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"1F",X"1F",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"62",X"62",X"62",X"40",X"0F",X"0F",
		X"08",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"C0",X"80",X"00",X"F8",X"F8",X"0F",X"0F",X"41",X"41",X"C0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"88",X"88",X"88",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"F8",X"F8",X"00",X"80",X"C0",X"C0",X"E0",X"E1",X"00",X"80",X"80",X"C0",X"41",X"41",X"0F",X"0F",
		X"08",X"08",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"0F",X"0F",X"40",X"62",X"62",X"62",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"3D",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"81",X"A0",X"A1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"69",X"69",
		X"0C",X"0C",X"0C",X"E0",X"EE",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"0F",X"0F",X"0F",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"F5",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"A0",X"A1",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"78",
		X"F5",X"3D",X"19",X"00",X"00",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"78",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"62",X"6A",X"6A",X"48",X"08",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"0F",X"0F",
		X"08",X"0C",X"3C",X"34",X"31",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"69",X"69",X"3C",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"35",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"66",X"60",X"60",X"60",X"0F",X"0F",
		X"08",X"0C",X"1E",X"71",X"62",X"44",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"69",X"69",X"69",X"60",X"60",X"66",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"3D",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"A0",X"A1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"E0",X"EE",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"69",X"69",X"3C",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"62",X"6A",X"6A",X"48",X"08",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"33",X"30",X"30",X"30",X"69",X"69",
		X"08",X"0C",X"3D",X"35",X"31",X"00",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"0F",X"0F",X"0F",X"30",X"30",X"33",X"00",X"00",
		X"00",X"00",X"00",X"31",X"35",X"35",X"2C",X"0C",X"00",X"00",X"11",X"10",X"30",X"36",X"96",X"F0",
		X"00",X"00",X"00",X"E6",X"80",X"C0",X"C1",X"E1",X"00",X"00",X"66",X"60",X"60",X"60",X"69",X"69",
		X"08",X"0C",X"1E",X"71",X"62",X"44",X"00",X"00",X"F0",X"70",X"30",X"73",X"F7",X"F7",X"70",X"00",
		X"E1",X"E1",X"80",X"80",X"C8",X"80",X"00",X"00",X"0F",X"0F",X"0F",X"60",X"60",X"66",X"00",X"00",
		X"00",X"00",X"00",X"44",X"4C",X"4C",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"31",X"B2",X"F2",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"C0",X"C0",X"40",X"0F",X"0F",
		X"08",X"08",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"0F",X"0F",X"40",X"C8",X"C8",X"C8",X"00",X"00",
		X"00",X"00",X"00",X"26",X"2E",X"2E",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"11",X"91",X"D1",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"C0",X"C0",X"40",X"0F",X"0F",
		X"08",X"08",X"2E",X"2E",X"26",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"D1",X"91",X"11",X"00",X"00",X"0F",X"0F",X"40",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"17",X"1F",X"1F",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"C8",X"C8",X"C8",X"40",X"0F",X"0F",
		X"08",X"08",X"4C",X"4C",X"44",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"F2",X"B2",X"32",X"00",X"00",X"0F",X"0F",X"40",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"1F",X"1F",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"62",X"62",X"62",X"40",X"0F",X"0F",
		X"08",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"C0",X"80",X"00",X"F8",X"F8",X"0F",X"0F",X"41",X"41",X"C0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"88",X"88",X"88",X"08",X"08",X"00",X"00",X"70",X"F0",X"70",X"30",X"70",X"F0",
		X"F8",X"F8",X"00",X"80",X"C0",X"C0",X"E0",X"E1",X"00",X"80",X"80",X"C0",X"41",X"41",X"0F",X"0F",
		X"08",X"08",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"F0",X"70",X"30",X"70",X"F0",X"70",X"00",X"00",
		X"E1",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"0F",X"0F",X"40",X"62",X"62",X"62",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
