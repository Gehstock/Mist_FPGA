`define BUILD_DATE "191004"
`define BUILD_TIME "203008"
