library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity domino_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of domino_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",
		X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",
		X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"FF",X"D5",X"C0",X"F5",X"C0",X"3D",X"C0",X"0F",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"C0",X"0F",X"C0",X"3D",X"C0",X"F5",X"FF",X"D5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"7C",X"00",X"5F",X"00",X"57",X"C0",X"55",X"F0",
		X"55",X"70",X"55",X"70",X"55",X"7C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",
		X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"7C",X"55",X"70",X"55",X"70",
		X"55",X"F0",X"57",X"C0",X"5F",X"00",X"7C",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"FD",X"00",X"D5",X"03",X"D5",X"0F",X"55",
		X"0D",X"55",X"0D",X"55",X"3D",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",
		X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"3D",X"55",X"0D",X"55",X"0D",X"55",
		X"0F",X"55",X"03",X"D5",X"00",X"D5",X"00",X"FD",X"00",X"0F",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FC",X"F5",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"F5",X"7C",X"3D",X"F0",X"0F",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"F0",X"0F",X"7C",X"3D",X"5F",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"5F",X"3F",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"7F",X"00",X"57",X"00",X"57",X"C0",X"55",X"F0",
		X"55",X"70",X"55",X"70",X"55",X"7C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",
		X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"7C",X"55",X"70",X"55",X"70",
		X"55",X"F0",X"57",X"C0",X"57",X"00",X"7F",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"03",X"C0",X"03",X"F0",X"0F",X"70",X"0D",X"70",X"0D",X"7C",X"3D",X"5C",X"35",
		X"5F",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FD",X"7F",X"CD",X"73",X"CD",X"73",X"CF",X"F3",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",
		X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",
		X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"03",X"FF",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"FF",
		X"03",X"FF",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"57",
		X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",
		X"D5",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"FF",X"C0",
		X"FF",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"FF",X"C0",X"00",X"00",
		X"00",X"00",X"C0",X"03",X"C0",X"03",X"F0",X"03",X"70",X"03",X"7C",X"03",X"5C",X"03",X"5F",X"03",
		X"57",X"03",X"57",X"C3",X"55",X"C3",X"55",X"F3",X"55",X"73",X"55",X"7F",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"FD",X"55",X"CD",X"55",X"CF",X"55",X"C3",X"55",X"C3",X"D5",X"C0",X"D5",
		X"C0",X"F5",X"C0",X"35",X"C0",X"3D",X"C0",X"0D",X"C0",X"0F",X"C0",X"03",X"C0",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0D",
		X"00",X"0D",X"00",X"0D",X"00",X"3D",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"F5",X"00",X"D5",
		X"00",X"D5",X"00",X"D5",X"03",X"D5",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"0F",X"55",
		X"0D",X"55",X"3D",X"57",X"35",X"57",X"35",X"5F",X"35",X"5C",X"35",X"5C",X"3F",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"D5",X"57",X"D5",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"D5",X"5F",X"F5",X"5C",X"35",X"5C",X"35",X"7C",X"3D",X"70",X"0D",X"70",X"0D",X"7F",X"FD",
		X"00",X"00",X"05",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"05",X"50",
		X"00",X"00",X"05",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",
		X"00",X"00",X"15",X"50",X"10",X"50",X"00",X"50",X"15",X"50",X"14",X"00",X"14",X"10",X"15",X"50",
		X"00",X"00",X"15",X"50",X"10",X"50",X"00",X"50",X"05",X"40",X"00",X"50",X"10",X"50",X"15",X"50",
		X"00",X"00",X"00",X"50",X"14",X"50",X"14",X"50",X"15",X"54",X"00",X"50",X"00",X"50",X"00",X"50",
		X"00",X"00",X"15",X"50",X"14",X"10",X"14",X"00",X"15",X"50",X"00",X"50",X"10",X"50",X"15",X"50",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"50",X"14",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"05",X"50",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"00",X"14",X"14",X"14",X"15",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"FD",X"70",X"0D",X"F0",X"0F",
		X"C0",X"03",X"C0",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"70",X"00",
		X"70",X"00",X"70",X"00",X"7C",X"00",X"5C",X"00",X"5C",X"00",X"5C",X"00",X"5F",X"00",X"57",X"00",
		X"57",X"00",X"57",X"00",X"57",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"F0",
		X"55",X"70",X"D5",X"7C",X"D5",X"5C",X"F5",X"5C",X"35",X"5C",X"35",X"5C",X"3F",X"FC",X"00",X"00",
		X"06",X"E4",X"0F",X"FC",X"0D",X"DC",X"15",X"55",X"15",X"55",X"0A",X"A8",X"0A",X"28",X"2A",X"2A",
		X"00",X"00",X"05",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"50",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"14",X"00",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"50",X"14",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"54",X"15",X"50",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"00",X"14",X"00",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"14",X"54",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",
		X"00",X"00",X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",
		X"00",X"00",X"01",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"14",X"50",X"14",X"50",X"15",X"50",
		X"00",X"00",X"14",X"10",X"14",X"50",X"15",X"50",X"15",X"00",X"15",X"50",X"14",X"50",X"14",X"50",
		X"00",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"54",X"54",X"55",X"54",X"51",X"14",X"51",X"14",X"50",X"14",X"50",X"14",X"50",X"14",
		X"00",X"00",X"50",X"14",X"54",X"14",X"55",X"14",X"55",X"54",X"51",X"54",X"50",X"54",X"50",X"14",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"00",X"14",X"00",X"14",X"00",
		X"00",X"00",X"55",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"51",X"50",X"51",X"54",X"55",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"50",X"14",X"14",X"14",X"14",X"14",X"14",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"54",X"00",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"15",X"54",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"14",X"04",X"14",X"04",X"14",X"04",X"14",X"14",X"14",X"50",X"15",X"40",X"15",X"00",
		X"00",X"00",X"50",X"14",X"50",X"14",X"50",X"14",X"51",X"14",X"51",X"14",X"55",X"54",X"54",X"54",
		X"00",X"00",X"50",X"14",X"54",X"54",X"15",X"50",X"05",X"40",X"15",X"50",X"54",X"54",X"50",X"14",
		X"00",X"00",X"14",X"14",X"14",X"14",X"15",X"54",X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"15",X"54",X"14",X"14",X"00",X"50",X"01",X"40",X"05",X"00",X"14",X"14",X"15",X"54",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FA",X"FF",X"EA",X"FF",X"AA",X"FE",X"AA",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"56",X"55",X"56",X"55",X"56",X"55",X"AA",X"AA",X"55",X"56",X"55",X"56",X"55",X"56",X"AA",X"AA",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"AA",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"01",X"AA",X"01",X"80",X"01",X"80",X"01",X"80",
		X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",
		X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"AA",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",
		X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"D5",X"55",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"FF",X"FF",
		X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",
		X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"AA",X"A7",X"55",X"57",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"5D",X"D5",X"5D",X"D5",X"7D",X"FD",X"75",X"DD",X"7D",X"F5",X"5D",X"DD",X"7D",X"DD",X"75",
		X"D5",X"FD",X"D5",X"D5",X"D5",X"D5",X"FD",X"FD",X"DD",X"DD",X"F5",X"FD",X"DD",X"DD",X"DD",X"DD",
		X"5D",X"5F",X"7D",X"57",X"75",X"57",X"F7",X"FF",X"D7",X"77",X"F7",X"77",X"77",X"57",X"F7",X"57",
		X"7D",X"55",X"5D",X"55",X"5D",X"55",X"7F",X"F5",X"77",X"75",X"77",X"75",X"75",X"75",X"75",X"75",
		X"7D",X"75",X"5D",X"75",X"5D",X"75",X"7D",X"7D",X"77",X"5D",X"77",X"5D",X"77",X"7D",X"7D",X"75",
		X"75",X"75",X"75",X"75",X"7D",X"7D",X"5D",X"5D",X"5F",X"5D",X"57",X"5D",X"7F",X"7D",X"75",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"80",X"00",
		X"AA",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A8",X"A8",X"08",X"80",X"A8",X"A8",X"80",X"08",X"A8",X"A8",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"A8",X"00",X"80",X"00",X"00",X"00",
		X"AA",X"A0",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"00",X"AA",
		X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"00",X"2A",
		X"40",X"00",X"50",X"00",X"14",X"00",X"05",X"54",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"15",X"40",X"00",X"54",X"00",X"05",
		X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",
		X"15",X"54",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"40",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"80",X"A8",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",
		X"AA",X"80",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"3F",X"30",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"30",X"00",X"F0",X"00",X"F0",X"00",X"C3",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"3C",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"3C",X"00",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"3F",X"00",X"3C",X"00",X"00",X"00",X"10",X"0F",X"14",X"3F",X"00",X"3C",
		X"00",X"0C",X"0F",X"0F",X"3F",X"00",X"3C",X"00",X"00",X"00",X"10",X"0F",X"14",X"3F",X"00",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"02",X"FF",X"02",X"AA",
		X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F8",X"00",X"FA",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"55",X"55",X"55",
		X"55",X"55",X"15",X"55",X"00",X"55",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",
		X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"99",X"99",X"99",
		X"99",X"59",X"99",X"59",X"99",X"59",X"99",X"59",X"99",X"59",X"99",X"59",X"99",X"59",X"99",X"59",
		X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"95",X"99",X"AA",X"9A",X"95",X"A9",X"55",
		X"99",X"59",X"99",X"59",X"99",X"59",X"99",X"69",X"99",X"A5",X"99",X"95",X"9A",X"95",X"AA",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"E9",X"FF",X"A5",X"FE",X"95",X"FE",X"55",X"FA",X"57",
		X"E9",X"5F",X"A5",X"7F",X"95",X"FF",X"97",X"FF",X"97",X"FF",X"AB",X"FA",X"EA",X"A9",X"E5",X"55",
		X"E5",X"55",X"E5",X"55",X"E5",X"55",X"EA",X"55",X"FE",X"55",X"FE",X"55",X"FE",X"57",X"FE",X"FF",
		X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",X"E9",X"FF",X"A9",X"FE",X"BA",X"FE",X"FE",
		X"FA",X"FE",X"FB",X"FE",X"FB",X"FE",X"FB",X"FE",X"FB",X"FE",X"FB",X"FF",X"FB",X"FF",X"FA",X"FF",
		X"FA",X"FF",X"FE",X"BF",X"FE",X"BF",X"FF",X"AF",X"FF",X"EB",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"AA",X"A9",X"55",X"95",X"55",X"55",X"55",X"55",X"FF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"EA",X"FF",X"A9",X"FA",X"95",X"A9",X"55",X"95",X"55",X"55",X"56",X"55",X"5A",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"7A",X"55",X"FA",X"FF",X"FA",X"FF",X"FA",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"F6",X"FF",X"D6",X"D5",X"56",X"55",X"56",X"55",X"56",X"55",X"5A",
		X"A5",X"56",X"AA",X"56",X"AA",X"A6",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"AA",X"BB",X"EA",X"FB",
		X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"F5",X"FF",X"D5",X"AA",X"55",X"FF",X"FF",X"FF",X"FF",
		X"AB",X"FF",X"5A",X"FF",X"5A",X"BF",X"F9",X"BF",X"F9",X"AF",X"F9",X"6F",X"E9",X"6F",X"A5",X"6B",
		X"95",X"59",X"55",X"5A",X"55",X"5E",X"55",X"5E",X"55",X"5E",X"55",X"7E",X"AA",X"BE",X"AA",X"BF",
		X"AA",X"AF",X"AA",X"AD",X"AA",X"AD",X"BF",X"AD",X"BF",X"A9",X"BF",X"A9",X"BF",X"A9",X"AA",X"A9",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"AA",X"AA",X"BF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"BF",X"EA",X"BF",X"BF",X"BE",X"BF",X"BE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"BF",X"FF",X"BF",
		X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"6F",X"FF",X"FB",X"FF",X"FE",X"AA",
		X"FF",X"D7",X"FF",X"5D",X"FD",X"59",X"F6",X"57",X"F5",X"D5",X"D5",X"66",X"6D",X"DD",X"56",X"57",
		X"55",X"97",X"E7",X"5D",X"55",X"59",X"76",X"57",X"59",X"D5",X"95",X"66",X"9D",X"DD",X"96",X"57",
		X"95",X"97",X"A7",X"5D",X"95",X"59",X"B6",X"57",X"99",X"D5",X"95",X"66",X"9D",X"DD",X"96",X"57",
		X"9D",X"97",X"A5",X"5D",X"95",X"59",X"A6",X"55",X"E9",X"D5",X"FA",X"55",X"FE",X"95",X"FF",X"95",
		X"BF",X"A5",X"BF",X"E5",X"AF",X"E5",X"EF",X"E5",X"EF",X"E9",X"EF",X"F9",X"EF",X"F9",X"AF",X"F9",
		X"BF",X"F9",X"FF",X"E9",X"FF",X"E5",X"FF",X"A5",X"FF",X"95",X"FE",X"95",X"EA",X"55",X"A5",X"55",
		X"55",X"9F",X"75",X"57",X"57",X"5D",X"65",X"55",X"55",X"75",X"5D",X"55",X"96",X"5D",X"55",X"55",
		X"95",X"5B",X"56",X"75",X"5D",X"55",X"96",X"75",X"5D",X"56",X"55",X"75",X"75",X"95",X"56",X"56",
		X"95",X"5F",X"56",X"5E",X"5D",X"7F",X"96",X"6E",X"5D",X"FF",X"55",X"EB",X"57",X"EF",X"5F",X"BE",
		X"5E",X"EF",X"7F",X"FE",X"FB",X"BF",X"7F",X"EE",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"97",X"FF",X"65",X"FF",X"55",X"7F",
		X"77",X"5F",X"99",X"D7",X"5D",X"9E",X"75",X"7F",X"D5",X"EF",X"9D",X"FE",X"67",X"EF",X"5E",X"FE",
		X"77",X"EF",X"5F",X"BF",X"7E",X"FE",X"7F",X"FF",X"7B",X"EF",X"7F",X"FE",X"6F",X"EF",X"FE",X"FE",
		X"FE",X"FF",X"EF",X"FB",X"FF",X"BF",X"BF",X"BF",X"EF",X"FE",X"FE",X"EF",X"FF",X"BE",X"BB",X"FF",
		X"EB",X"FF",X"FF",X"BB",X"BF",X"FF",X"EF",X"BE",X"FE",X"FF",X"FF",X"FB",X"55",X"7F",X"55",X"57",
		X"FE",X"FF",X"EF",X"EF",X"FF",X"FF",X"BE",X"EF",X"FF",X"FF",X"FB",X"FB",X"EF",X"BF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FB",X"FF",X"EF",X"BF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"BE",X"FF",
		X"FE",X"FB",X"BF",X"FF",X"FF",X"EE",X"FB",X"FF",X"FF",X"ED",X"EF",X"F5",X"FB",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"B9",X"55",X"FF",X"55",X"EE",X"D5",X"FB",X"D5",X"BF",X"95",
		X"BE",X"55",X"ED",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FE",X"F5",X"EF",X"ED",X"FF",X"FF",X"BE",X"EF",X"FF",X"FF",X"FB",X"FB",X"EF",X"BF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"AA",X"40",X"02",X"40",X"02",X"40",X"02",X"40",
		X"02",X"40",X"02",X"40",X"02",X"40",X"02",X"40",X"02",X"40",X"02",X"40",X"02",X"40",X"02",X"40",
		X"02",X"40",X"02",X"40",X"02",X"40",X"AA",X"40",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"55",X"52",X"AA",X"92",X"00",X"02",X"00",X"02",X"00",X"00",
		X"05",X"50",X"14",X"14",X"11",X"44",X"11",X"04",X"11",X"04",X"11",X"44",X"14",X"14",X"05",X"50",
		X"0F",X"FC",X"03",X"B0",X"0E",X"AC",X"3E",X"FC",X"FE",X"AF",X"FF",X"EF",X"FE",X"AF",X"3F",X"BC",
		X"0F",X"F0",X"3F",X"FC",X"F5",X"5F",X"FD",X"5F",X"7D",X"DD",X"6F",X"F9",X"17",X"D4",X"05",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"A8",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A8",X"A8",X"88",X"88",X"88",X"88",X"88",X"88",X"A8",X"A8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A8",X"00",X"08",X"00",X"A8",X"00",X"80",X"00",X"A8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A8",X"00",X"80",X"00",X"A8",X"00",X"08",X"00",X"A8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A2",X"A2",X"22",X"22",X"82",X"22",X"22",X"22",X"A2",X"A2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A2",X"22",X"22",X"22",X"22",X"22",X"22",X"20",X"22",X"A2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"01",X"55",X"A1",X"AA",X"20",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"F0",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",
		X"FF",X"EA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",
		X"FF",X"EA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"AF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",
		X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",
		X"AB",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FA",X"FF",X"EA",X"FF",X"AA",X"FE",X"AA",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"00",X"30",X"00",X"3C",X"00",X"0C",X"00",X"0F",X"00",X"03",
		X"C0",X"00",X"C0",X"00",X"F0",X"00",X"30",X"00",X"3C",X"00",X"0C",X"00",X"0F",X"00",X"03",X"00",
		X"03",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"30",X"00",X"3C",X"00",X"0C",X"00",X"0F",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"30",X"00",X"3C",X"00",X"0C",X"00",X"0F",X"00",X"03",X"00",
		X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0C",X"00",X"3C",X"00",X"30",X"00",X"F0",
		X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"0C",X"00",X"3C",X"00",X"30",X"00",X"F0",X"00",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"03",X"C0",X"03",X"00",X"0F",X"00",X"0C",X"00",X"3C",X"00",X"30",X"00",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"00",X"0F",X"00",X"0C",X"00",X"3C",X"00",X"30",X"00",X"F0",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"FF",X"FF",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
