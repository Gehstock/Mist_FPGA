`define BUILD_DATE "190303"
`define BUILD_TIME "171430"
