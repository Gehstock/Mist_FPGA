library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ttag_ch_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ttag_ch_bits is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AB",X"AA",X"AA",X"EA",X"AB",X"AA",X"AF",X"FE",X"AA",X"AA",X"AE",X"EE",X"AE",X"EE",X"AF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"3F",X"FC",X"C0",X"03",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"CF",X"F3",X"C0",X"03",X"3F",X"FC",
		X"AA",X"AA",X"AA",X"AE",X"AA",X"AE",X"AF",X"FE",X"AA",X"AA",X"AF",X"EA",X"AE",X"EA",X"AF",X"FE",
		X"AA",X"AA",X"AF",X"EA",X"AA",X"FE",X"AF",X"EA",X"AA",X"AA",X"AB",X"FE",X"AF",X"BA",X"AB",X"FE",
		X"AA",X"AA",X"AF",X"BE",X"AE",X"EA",X"AF",X"FE",X"AA",X"AA",X"AE",X"EE",X"AE",X"EE",X"AF",X"FE",
		X"AF",X"FE",X"AE",X"AA",X"AE",X"AA",X"AF",X"EA",X"AE",X"EA",X"AF",X"FE",X"AA",X"AA",X"AF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"AA",X"FE",X"AF",X"AA",X"AE",X"AA",X"AE",X"AA",
		X"AF",X"EA",X"AE",X"EA",X"AF",X"FE",X"AA",X"AA",X"AE",X"FE",X"AE",X"EE",X"AF",X"EE",X"AA",X"AA",
		X"AE",X"AE",X"AE",X"AE",X"AF",X"FE",X"AA",X"AA",X"AB",X"FE",X"AF",X"BA",X"AB",X"FE",X"AA",X"AA",
		X"AE",X"FE",X"AE",X"EE",X"AF",X"EE",X"AA",X"AA",X"AE",X"EE",X"AE",X"EE",X"AF",X"FE",X"AA",X"AA",
		X"AC",X"00",X"AC",X"00",X"AC",X"FF",X"BC",X"EA",X"B0",X"FA",X"BC",X"3E",X"AF",X"0E",X"AB",X"FE",
		X"00",X"0E",X"00",X"0E",X"FF",X"CE",X"AA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"FE",X"AF",X"0E",X"BC",X"3E",X"B0",X"FA",X"BC",X"EA",X"AC",X"FF",X"AC",X"00",X"AC",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"FF",X"CE",X"00",X"0E",X"00",X"0E",
		X"AF",X"EA",X"AC",X"FF",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"FF",X"AF",X"EA",
		X"AB",X"CE",X"FF",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"3E",X"00",X"FA",X"FF",X"EA",X"AA",X"AA",
		X"AA",X"AA",X"AF",X"EA",X"AC",X"FF",X"AC",X"00",X"AC",X"00",X"AC",X"FF",X"AF",X"EA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"EA",X"00",X"FA",X"00",X"3E",X"FF",X"0E",X"AB",X"CE",X"AA",X"CE",
		X"AC",X"EA",X"AC",X"FA",X"AC",X"3F",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"FF",X"AF",X"EA",
		X"B3",X"BE",X"F3",X"CE",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"FF",X"CE",X"AA",X"FE",
		X"AA",X"AA",X"AA",X"FF",X"AB",X"C0",X"AB",X"00",X"AF",X"00",X"AC",X"03",X"AC",X"3F",X"AC",X"FA",
		X"AA",X"FE",X"FA",X"CE",X"3E",X"CE",X"0F",X"0E",X"0C",X"0E",X"00",X"0E",X"C0",X"CE",X"F3",X"FE",
		X"AC",X"EB",X"AC",X"FF",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"FF",X"AF",X"EA",X"AA",X"AA",
		X"3A",X"CE",X"3F",X"CE",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"FF",X"CE",X"AA",X"FE",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"FF",X"AF",X"03",X"AC",X"00",X"AC",X"00",X"AC",X"FC",
		X"AA",X"AA",X"BF",X"FA",X"F0",X"3E",X"C0",X"0E",X"00",X"0E",X"0F",X"0E",X"3F",X"CE",X"3A",X"CE",
		X"AC",X"EA",X"AC",X"FA",X"AC",X"3F",X"AF",X"00",X"AB",X"00",X"AB",X"C0",X"AA",X"FC",X"AA",X"AF",
		X"AA",X"CE",X"AB",X"CE",X"FF",X"0E",X"00",X"0E",X"00",X"3E",X"00",X"3A",X"00",X"FA",X"FF",X"EA",
		X"AA",X"AF",X"AA",X"FC",X"AB",X"C0",X"AB",X"00",X"AF",X"00",X"AC",X"3F",X"AC",X"FA",X"AC",X"EA",
		X"FF",X"EA",X"00",X"FA",X"00",X"3A",X"00",X"3E",X"00",X"0E",X"FF",X"0E",X"AB",X"CE",X"AA",X"CE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"FE",X"FE",X"9A",X"9A",X"55",X"56",X"75",X"D6",X"55",X"56",X"9A",X"9A",X"FE",X"FE",X"AA",X"AA",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"FF",X"FF",
		X"AF",X"EA",X"AF",X"FE",X"AA",X"AA",X"AF",X"FE",X"AE",X"AE",X"AF",X"FE",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AE",X"EE",X"AE",X"EE",X"AF",X"FE",X"AA",X"AA",X"AF",X"FE",X"AA",X"BE",
		X"AF",X"FF",X"BE",X"AB",X"BA",X"AB",X"BA",X"AB",X"BA",X"AB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AB",X"BF",X"FF",X"BF",X"FF",X"BA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BF",X"EB",X"BF",X"EB",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BA",X"FF",X"BA",X"FF",X"AA",X"AA",
		X"BF",X"FF",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BA",X"AB",X"BE",X"AF",X"BE",X"AF",X"AA",X"AA",
		X"AA",X"EA",X"BF",X"FF",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"BF",X"EA",X"BF",X"EA",X"AA",X"AA",
		X"BA",X"FF",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BF",X"EF",X"BF",X"EF",X"AA",X"AA",
		X"BA",X"FF",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BE",X"AA",X"BB",X"AA",X"BB",X"EA",X"BA",X"FF",X"BA",X"BF",X"BE",X"AA",X"BE",X"AA",X"AA",X"AA",
		X"BF",X"FF",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"FF",X"BF",X"FF",X"BA",X"EA",X"BA",X"EA",X"BA",X"EA",X"BA",X"EA",X"BF",X"EA",X"AA",X"AA",
		X"0F",X"FF",X"3C",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"03",X"3F",X"FF",X"3F",X"FF",X"30",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"C3",X"3F",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"FF",X"30",X"FF",X"00",X"00",
		X"3F",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"03",X"3C",X"0F",X"3C",X"0F",X"00",X"00",
		X"00",X"C0",X"3F",X"FF",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"3F",X"C0",X"3F",X"C0",X"00",X"00",
		X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"CF",X"3F",X"CF",X"00",X"00",
		X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3C",X"00",X"33",X"00",X"33",X"C0",X"30",X"FF",X"30",X"3F",X"3C",X"00",X"3C",X"00",X"00",X"00",
		X"3F",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"FF",X"3F",X"FF",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"3F",X"C0",X"00",X"00",
		X"AA",X"FE",X"AA",X"AE",X"AF",X"FE",X"AA",X"AA",X"AE",X"AA",X"AF",X"FE",X"AE",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AF",X"FE",X"AE",X"AE",X"AF",X"FE",X"AA",X"AA",X"AF",X"FE",X"AA",X"AE",
		X"AF",X"FE",X"AF",X"FE",X"AA",X"AA",X"AA",X"BE",X"AA",X"BE",X"AF",X"FE",X"AF",X"FE",X"AA",X"AA",
		X"AF",X"FE",X"AF",X"FE",X"AF",X"AA",X"AF",X"AA",X"AA",X"AA",X"AF",X"FE",X"AF",X"FE",X"AF",X"BE",
		X"AE",X"EA",X"BF",X"FA",X"AE",X"EA",X"BF",X"FA",X"AE",X"EA",X"AA",X"AA",X"AF",X"AA",X"AF",X"AA",
		X"00",X"00",X"00",X"C3",X"00",X"3C",X"0F",X"33",X"30",X"C3",X"0F",X"C3",X"00",X"3C",X"00",X"00",
		X"9B",X"66",X"9B",X"66",X"9B",X"66",X"9B",X"66",X"9B",X"66",X"9B",X"66",X"9B",X"66",X"9B",X"66",
		X"3F",X"FF",X"3F",X"FF",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"3F",X"33",X"F3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"30",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",X"30",X"0F",X"3F",X"FF",X"3F",X"FC",X"00",X"00",
		X"0F",X"FC",X"3C",X"0F",X"30",X"03",X"30",X"03",X"30",X"03",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"30",X"03",X"30",X"03",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"30",X"00",X"30",X"00",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"03",X"30",X"03",X"3F",X"FF",X"3F",X"FC",X"00",X"00",
		X"3F",X"FF",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"03",X"3F",X"FF",X"3F",X"FF",X"30",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"3F",X"FF",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"00",
		X"3C",X"03",X"0F",X"0F",X"03",X"FC",X"00",X"F0",X"00",X"30",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"00",X"0F",X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"03",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"FF",X"0F",X"00",X"03",X"F0",X"03",X"F0",X"0F",X"00",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"FF",X"00",X"3F",X"03",X"F0",X"3F",X"00",X"30",X"00",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"FF",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"FF",X"30",X"3C",X"30",X"3F",X"30",X"03",X"30",X"03",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"CF",X"30",X"FF",X"30",X"F0",X"30",X"C0",X"30",X"C0",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"30",X"FF",X"30",X"FF",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"3F",X"CF",X"3F",X"CF",X"00",X"00",
		X"00",X"00",X"30",X"00",X"30",X"00",X"3F",X"FF",X"3F",X"FF",X"30",X"00",X"30",X"00",X"00",X"00",
		X"3F",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3F",X"F0",X"00",X"3C",X"00",X"0F",X"00",X"3F",X"00",X"FC",X"3F",X"F0",X"3F",X"C0",X"00",X"00",
		X"3F",X"FF",X"00",X"3C",X"03",X"F0",X"03",X"F0",X"00",X"3C",X"3F",X"FF",X"3F",X"FF",X"00",X"00",
		X"3C",X"0F",X"0F",X"3C",X"03",X"F0",X"00",X"C0",X"03",X"F0",X"0F",X"3C",X"3C",X"0F",X"00",X"00",
		X"3C",X"00",X"0F",X"00",X"03",X"C0",X"00",X"FF",X"03",X"FF",X"0F",X"C0",X"3F",X"00",X"00",X"00",
		X"3C",X"03",X"3F",X"03",X"33",X"C3",X"30",X"C3",X"30",X"F3",X"30",X"3F",X"30",X"0F",X"00",X"00",
		X"BF",X"FF",X"BF",X"FF",X"BA",X"EA",X"BA",X"EA",X"BA",X"EA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"BF",X"BB",X"FB",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BA",X"AF",X"BA",X"AF",X"BA",X"AF",X"BA",X"AF",X"BA",X"AF",X"BF",X"FF",X"BF",X"FE",X"AA",X"AA",
		X"AF",X"FE",X"BE",X"AF",X"BA",X"AB",X"BA",X"AB",X"BA",X"AB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BA",X"AB",X"BA",X"AB",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BA",X"FF",X"BA",X"EB",X"BA",X"EB",X"BA",X"AB",X"BA",X"AB",X"BF",X"FF",X"BF",X"FE",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"BA",X"AB",X"BF",X"FF",X"BF",X"FF",X"BA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"FF",X"AF",X"AA",X"AB",X"FA",X"AB",X"FA",X"AF",X"AA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"FF",X"AA",X"BF",X"AB",X"FA",X"BF",X"AA",X"BA",X"AA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"FF",X"BA",X"AB",X"BA",X"AB",X"BA",X"AB",X"BA",X"AB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"EA",X"BA",X"EA",X"BA",X"EA",X"BA",X"EA",X"BA",X"EA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"FF",X"BA",X"BE",X"BA",X"BF",X"BA",X"AB",X"BA",X"AB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BF",X"EF",X"BA",X"FF",X"BA",X"FA",X"BA",X"EA",X"BA",X"EA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BE",X"FF",X"BE",X"FF",X"BA",X"EB",X"BA",X"EB",X"BA",X"EB",X"BF",X"EF",X"BF",X"EF",X"AA",X"AA",
		X"AA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BF",X"FF",X"BF",X"FF",X"BA",X"AA",X"BA",X"AA",X"AA",X"AA",
		X"BF",X"FF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"BE",X"AA",X"AF",X"AA",X"AB",X"EA",X"AA",X"FF",X"AB",X"FF",X"AF",X"EA",X"BF",X"AA",X"AA",X"AA",
		X"BE",X"AB",X"AF",X"AF",X"AB",X"FE",X"AA",X"FA",X"AA",X"BA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"BF",X"FF",
		X"AA",X"A9",X"9A",X"99",X"A6",X"69",X"A9",X"A9",X"A6",X"69",X"9A",X"99",X"AA",X"A9",X"AA",X"A9",
		X"BA",X"AA",X"BA",X"AA",X"BA",X"EA",X"BA",X"EA",X"BA",X"EA",X"BF",X"FF",X"BF",X"FF",X"AA",X"AA",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"FF",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"AA",X"A9",X"95",X"59",X"9A",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",
		X"BF",X"FF",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"AA",X"AA",X"A5",X"56",X"95",X"55",X"9A",X"A9",X"9A",X"A9",X"9A",X"A9",X"95",X"55",X"A5",X"56",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"95",X"55",X"95",X"55",X"9A",X"A9",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A5",X"A9",X"99",X"69",X"9A",X"69",X"9A",X"59",X"9A",X"99",X"9A",X"95",X"A6",X"A5",
		X"AA",X"AA",X"A5",X"96",X"95",X"55",X"9A",X"69",X"9A",X"69",X"9A",X"A9",X"96",X"A5",X"A6",X"A6",
		X"AA",X"AA",X"AA",X"6A",X"95",X"55",X"95",X"55",X"AA",X"6A",X"AA",X"6A",X"95",X"6A",X"95",X"6A",
		X"AA",X"AA",X"9A",X"56",X"99",X"55",X"99",X"65",X"99",X"A9",X"99",X"A9",X"95",X"A9",X"95",X"A5",
		X"AA",X"AA",X"96",X"96",X"9A",X"55",X"9A",X"69",X"9A",X"69",X"96",X"69",X"A5",X"55",X"A9",X"56",
		X"AA",X"AA",X"96",X"AA",X"95",X"6A",X"9A",X"55",X"9A",X"A5",X"9A",X"AA",X"9A",X"AA",X"96",X"AA",
		X"AA",X"AA",X"A5",X"96",X"95",X"55",X"9A",X"69",X"9A",X"69",X"9A",X"69",X"95",X"55",X"A5",X"96",
		X"AA",X"AA",X"95",X"55",X"95",X"55",X"9A",X"6A",X"9A",X"6A",X"9A",X"6A",X"95",X"6A",X"A5",X"AA",
		X"AA",X"A9",X"A5",X"69",X"96",X"59",X"9A",X"99",X"9A",X"99",X"96",X"59",X"A5",X"69",X"AA",X"A9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
