library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity twotiger_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of twotiger_sp_bits is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"FF",X"EE",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"EE",X"FF",
		X"00",X"55",X"55",X"EE",X"00",X"55",X"55",X"55",X"00",X"55",X"5E",X"F5",X"00",X"6F",X"E1",X"E5",
		X"00",X"EE",X"EF",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"EE",X"FF",X"EE",X"00",X"E5",X"55",X"FF",
		X"00",X"E5",X"5E",X"FF",X"00",X"FF",X"55",X"FE",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"1F",X"55",
		X"00",X"0E",X"EE",X"55",X"00",X"0E",X"00",X"55",X"00",X"EF",X"00",X"5E",X"00",X"EF",X"00",X"5E",
		X"00",X"FF",X"00",X"5E",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"EE",X"FF",X"00",
		X"00",X"5E",X"FF",X"00",X"00",X"5F",X"FF",X"00",X"00",X"6E",X"FF",X"00",X"00",X"F6",X"EF",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"E5",X"EE",X"00",X"F0",X"1E",X"5F",X"00",X"E0",X"F1",X"FF",
		X"00",X"00",X"EE",X"5F",X"00",X"00",X"FE",X"55",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0E",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0E",X"EF",X"00",X"00",X"EF",X"FF",X"00",
		X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"EE",X"00",X"65",X"55",X"FF",
		X"00",X"EF",X"55",X"FF",X"00",X"EE",X"55",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"16",X"FF",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"E0",X"55",X"00",X"0E",X"00",X"55",X"00",X"0E",X"00",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"EF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"5E",X"FF",X"00",X"00",X"6F",X"FF",X"00",X"00",X"FE",X"E5",X"E0",
		X"00",X"E0",X"55",X"FE",X"00",X"00",X"E5",X"FE",X"00",X"00",X"1E",X"FE",X"00",X"00",X"F1",X"E0",
		X"00",X"00",X"EE",X"E0",X"00",X"0E",X"00",X"5E",X"00",X"EF",X"00",X"5E",X"00",X"EF",X"00",X"5E",
		X"00",X"0E",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"5F",X"FF",X"00",X"00",X"6E",X"FF",X"00",X"00",X"6E",X"FF",X"00",X"00",X"EE",X"FF",X"EE",
		X"00",X"E0",X"EF",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"00",X"E5",X"FE",X"00",X"00",X"FE",X"FE",
		X"00",X"00",X"EE",X"E5",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"EE",X"00",X"00",X"F5",X"EF",X"00",
		X"00",X"E6",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"EE",X"EF",X"EE",X"00",X"F0",X"55",X"EF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"F1",X"FF",
		X"00",X"00",X"EE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"EE",X"00",X"00",X"E0",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"0E",X"00",X"00",X"F5",X"EF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"0E",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"E5",X"FE",X"00",X"00",X"1E",X"FE",
		X"00",X"00",X"E1",X"FE",X"00",X"00",X"FE",X"EE",X"00",X"00",X"E0",X"5E",X"00",X"00",X"00",X"5E",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"F5",X"E0",X"00",X"00",X"EF",X"5E",X"00",X"00",X"EE",X"5E",X"00",
		X"00",X"0E",X"EF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"1E",X"E0",
		X"00",X"00",X"EE",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"E0",X"00",X"00",X"EF",X"EE",X"00",X"00",X"EE",X"5E",X"00",X"00",X"0F",X"5E",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"5F",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"0E",X"15",X"00",X"00",X"0E",X"65",X"E0",X"00",X"0E",X"EF",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"E5",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"0F",X"5E",X"00",
		X"00",X"EE",X"5E",X"00",X"00",X"F0",X"EF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5F",X"00",X"00",X"0E",X"5E",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"0E",X"E5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E6",X"E0",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"0E",X"55",X"00",X"00",X"FE",X"55",X"E0",
		X"00",X"00",X"5E",X"E0",X"00",X"00",X"5F",X"E0",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",
		X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"0E",X"E5",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"0E",X"E5",X"00",X"00",X"0E",X"65",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"5E",X"00",X"00",X"EF",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"FF",X"E0",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"0E",X"5E",X"00",X"00",X"EE",X"55",X"00",
		X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"FF",X"E0",
		X"00",X"0E",X"FF",X"E0",X"00",X"EE",X"5F",X"E0",X"00",X"EF",X"5E",X"00",X"00",X"EF",X"55",X"00",
		X"00",X"EE",X"5E",X"00",X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"E0",
		X"00",X"0E",X"FF",X"E0",X"00",X"EF",X"EF",X"E0",X"00",X"EF",X"EF",X"00",X"00",X"0F",X"EF",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"2E",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"EE",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"1E",X"00",
		X"E9",X"00",X"99",X"E0",X"99",X"00",X"99",X"EE",X"99",X"EE",X"EE",X"3E",X"99",X"BE",X"EB",X"9E",
		X"99",X"BB",X"BB",X"E2",X"9E",X"BB",X"BB",X"2E",X"EE",X"BB",X"EB",X"EE",X"0E",X"BB",X"EB",X"EB",
		X"0E",X"BB",X"EB",X"E9",X"0E",X"EE",X"EE",X"E9",X"0E",X"00",X"19",X"EE",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"EE",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"1E",X"00",
		X"E9",X"00",X"99",X"E0",X"9E",X"00",X"BB",X"EF",X"9E",X"EE",X"EE",X"FF",X"9E",X"AA",X"EA",X"EE",
		X"9E",X"AA",X"BE",X"BB",X"9E",X"EE",X"EE",X"BB",X"EE",X"BB",X"BB",X"BB",X"0E",X"BB",X"BB",X"BB",
		X"0E",X"EE",X"BB",X"BB",X"0E",X"F3",X"EE",X"BB",X"0E",X"3F",X"99",X"BB",X"0E",X"EE",X"B9",X"EE",
		X"0E",X"00",X"BB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"F1",X"00",
		X"00",X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"E0",X"00",
		X"EE",X"0E",X"E0",X"00",X"E9",X"EE",X"E0",X"00",X"E9",X"3E",X"FE",X"00",X"E9",X"EE",X"EE",X"00",
		X"E9",X"E1",X"EE",X"E0",X"99",X"11",X"E1",X"EE",X"99",X"E1",X"11",X"3E",X"99",X"EE",X"33",X"EE",
		X"99",X"EE",X"31",X"E2",X"9E",X"EE",X"11",X"2E",X"EE",X"EE",X"1E",X"EE",X"0E",X"11",X"1E",X"E2",
		X"0E",X"11",X"1E",X"E2",X"0E",X"13",X"11",X"E2",X"0E",X"11",X"11",X"EE",X"00",X"11",X"31",X"00",
		X"00",X"1E",X"EE",X"00",X"00",X"1E",X"EE",X"00",X"00",X"1E",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"E0",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"F0",X"00",X"33",X"11",X"00",
		X"EE",X"3E",X"11",X"00",X"E9",X"E3",X"11",X"30",X"E9",X"31",X"FE",X"10",X"E9",X"E1",X"EE",X"00",
		X"E9",X"E1",X"EE",X"E0",X"99",X"EE",X"EE",X"EE",X"99",X"EE",X"EE",X"3E",X"99",X"EE",X"EE",X"EE",
		X"99",X"33",X"EE",X"E2",X"9E",X"11",X"EE",X"2E",X"EE",X"1E",X"EE",X"EE",X"0E",X"1E",X"EE",X"E2",
		X"0E",X"EE",X"EE",X"E2",X"0E",X"EE",X"EE",X"E2",X"0E",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"EE",X"33",X"00",X"EE",X"EE",X"11",X"00",X"EE",X"1E",X"10",X"00",X"EE",X"11",X"00",
		X"00",X"E3",X"E1",X"00",X"00",X"01",X"E1",X"00",X"00",X"11",X"E0",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"AE",X"00",X"00",X"EA",X"AE",X"00",X"00",X"EA",X"AA",X"00",X"00",X"EA",X"AA",X"00",
		X"00",X"AE",X"AA",X"00",X"00",X"AA",X"1A",X"EE",X"00",X"2E",X"1A",X"EE",X"00",X"2E",X"EE",X"AE",
		X"00",X"BE",X"EE",X"BB",X"00",X"EE",X"32",X"1B",X"00",X"EE",X"AA",X"EE",X"00",X"EE",X"AA",X"EB",
		X"00",X"01",X"AA",X"BE",X"00",X"EE",X"EA",X"B9",X"00",X"EB",X"EA",X"B9",X"00",X"BB",X"9E",X"99",
		X"00",X"BB",X"EE",X"EE",X"00",X"B2",X"EA",X"00",X"00",X"B9",X"EA",X"00",X"00",X"99",X"EA",X"00",
		X"00",X"9E",X"EA",X"00",X"00",X"E0",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"3A",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"EA",X"00",X"00",X"AE",X"AA",X"00",X"00",X"E0",X"EE",X"00",X"00",X"0E",X"2E",X"00",
		X"00",X"EE",X"2A",X"00",X"00",X"AE",X"EA",X"00",X"00",X"AE",X"EE",X"00",X"00",X"AA",X"AE",X"00",
		X"00",X"E2",X"AA",X"00",X"00",X"E2",X"EE",X"00",X"00",X"EA",X"EE",X"00",X"00",X"AA",X"AE",X"00",
		X"00",X"AA",X"EA",X"00",X"00",X"EE",X"AE",X"00",X"00",X"2E",X"EE",X"00",X"00",X"12",X"EE",X"00",
		X"00",X"EE",X"12",X"00",X"00",X"EE",X"EE",X"00",X"00",X"AE",X"1E",X"00",X"00",X"AE",X"2E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0A",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"00",X"EF",X"EE",X"E0",X"00",X"BF",X"EE",X"EE",X"00",X"BE",X"EE",X"EE",X"0E",X"EE",X"EA",X"EE",
		X"00",X"AE",X"EE",X"E5",X"00",X"AA",X"EE",X"7E",X"00",X"EE",X"1E",X"BE",X"00",X"BB",X"EE",X"EE",
		X"00",X"BB",X"EE",X"E9",X"00",X"BB",X"99",X"99",X"00",X"EB",X"BB",X"BB",X"00",X"E2",X"92",X"22",
		X"00",X"02",X"20",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"E0",X"00",X"0F",X"01",X"E0",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"E0",X"10",X"E0",X"00",X"00",X"10",X"00",
		X"00",X"10",X"11",X"11",X"00",X"00",X"10",X"00",X"0F",X"E0",X"10",X"E0",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"01",X"E0",X"00",X"0F",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"0E",X"EE",X"00",X"11",X"EE",X"99",X"00",X"01",X"99",X"AA",X"00",X"00",X"99",X"AA",
		X"00",X"F0",X"92",X"EE",X"00",X"EE",X"22",X"00",X"00",X"1E",X"EE",X"E3",X"00",X"11",X"EE",X"EE",
		X"00",X"E1",X"1E",X"E3",X"00",X"EE",X"1E",X"EE",X"00",X"EE",X"3F",X"EE",X"00",X"EE",X"EE",X"EE",
		X"00",X"EE",X"3E",X"EE",X"00",X"FF",X"3F",X"FE",X"00",X"EF",X"3F",X"EE",X"00",X"EE",X"FF",X"EF",
		X"00",X"EE",X"11",X"EF",X"00",X"0E",X"EE",X"EE",X"00",X"EF",X"FE",X"FE",X"00",X"EE",X"11",X"EE",
		X"00",X"13",X"11",X"E3",X"00",X"11",X"EE",X"EE",X"00",X"11",X"EE",X"03",X"00",X"EE",X"22",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"00",X"10",X"00",X"92",X"EE",X"10",X"00",X"AA",X"99",X"11",X"00",X"A1",X"99",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"E1",X"00",X"11",X"11",X"EE",X"01",X"1E",X"1E",X"EE",
		X"01",X"EE",X"EE",X"E0",X"01",X"1E",X"EE",X"30",X"01",X"1E",X"EE",X"30",X"00",X"11",X"EE",X"30",
		X"00",X"11",X"EE",X"E3",X"00",X"EE",X"EE",X"E3",X"0E",X"EE",X"EE",X"33",X"0E",X"EE",X"EE",X"33",
		X"0E",X"EE",X"EE",X"EE",X"00",X"1E",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"00",X"11",X"EE",X"3E",
		X"00",X"11",X"EE",X"31",X"00",X"33",X"E1",X"3E",X"00",X"13",X"E1",X"1E",X"00",X"33",X"11",X"13",
		X"00",X"31",X"11",X"1E",X"00",X"01",X"11",X"EE",X"00",X"11",X"13",X"E1",X"00",X"11",X"13",X"13",
		X"00",X"11",X"10",X"11",X"00",X"EE",X"11",X"00",X"00",X"EE",X"11",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"60",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"F0",X"00",X"06",X"00",X"00",
		X"00",X"26",X"20",X"02",X"00",X"02",X"06",X"00",X"00",X"66",X"66",X"00",X"00",X"0F",X"66",X"06",
		X"0F",X"02",X"F6",X"F0",X"00",X"22",X"F6",X"20",X"00",X"20",X"62",X"00",X"00",X"20",X"62",X"00",
		X"00",X"22",X"22",X"00",X"00",X"02",X"2F",X"02",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"0F",X"F2",X"02",X"20",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"20",X"22",X"00",
		X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"02",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"20",X"06",X"00",X"00",X"22",X"06",X"00",X"00",X"02",X"26",X"06",X"00",X"00",X"26",X"60",
		X"00",X"00",X"2F",X"60",X"00",X"20",X"22",X"00",X"00",X"22",X"22",X"60",X"00",X"00",X"22",X"26",
		X"00",X"02",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",
		X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",
		X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",
		X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"6C",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"4C",
		X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"7F",X"70",
		X"00",X"70",X"00",X"0F",X"00",X"EF",X"00",X"07",X"00",X"70",X"70",X"00",X"F0",X"FF",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"E5",X"00",X"00",X"E6",X"FE",X"00",
		X"00",X"E6",X"FF",X"00",X"00",X"EA",X"FF",X"00",X"00",X"EA",X"FF",X"0E",X"00",X"EF",X"EE",X"EF",
		X"00",X"EE",X"EF",X"FF",X"00",X"66",X"66",X"66",X"00",X"AA",X"EE",X"E2",X"00",X"FF",X"FF",X"EE",
		X"00",X"FF",X"EE",X"BB",X"00",X"FF",X"EE",X"BB",X"00",X"FF",X"EE",X"EE",X"00",X"EE",X"EE",X"00",
		X"0E",X"AA",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E1",X"00",X"00",
		X"00",X"11",X"E0",X"00",X"00",X"EE",X"9E",X"00",X"00",X"0E",X"D9",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"BB",X"E0",X"00",X"00",X"BB",X"EE",
		X"00",X"00",X"BB",X"BE",X"00",X"00",X"EB",X"BB",X"00",X"00",X"EB",X"BB",X"00",X"00",X"EB",X"BB",
		X"00",X"00",X"EB",X"BB",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EE",X"F7",X"0F",X"7F",X"F7",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"EB",X"AA",X"0E",X"00",X"BE",X"AA",X"EB",X"00",X"BE",X"EE",X"BB",X"00",X"BB",X"CC",
		X"EE",X"00",X"EB",X"EF",X"77",X"F7",X"EB",X"EF",X"77",X"10",X"71",X"E7",X"00",X"70",X"00",X"00",
		X"00",X"01",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"07",X"EE",X"9A",X"E0",X"00",X"EE",
		X"BB",X"E7",X"7E",X"BB",X"77",X"E7",X"EE",X"E7",X"77",X"00",X"7E",X"E7",X"00",X"70",X"00",X"06",
		X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"E0",X"00",
		X"0E",X"00",X"2E",X"00",X"0E",X"00",X"21",X"00",X"0E",X"00",X"EE",X"EE",X"0E",X"EE",X"E2",X"2E",
		X"0E",X"22",X"22",X"E1",X"00",X"22",X"22",X"FE",X"E0",X"22",X"E2",X"EE",X"00",X"22",X"E2",X"22",
		X"00",X"EE",X"EE",X"22",X"00",X"00",X"EE",X"EE",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E0",X"00",
		X"E0",X"0E",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"0E",X"2E",X"5E",X"00",X"0E",X"EE",X"EE",X"00",
		X"0E",X"E7",X"2E",X"E0",X"0E",X"77",X"22",X"EE",X"0E",X"E7",X"22",X"6E",X"00",X"26",X"22",X"EE",
		X"00",X"26",X"22",X"E2",X"00",X"26",X"22",X"2E",X"00",X"26",X"E2",X"EE",X"00",X"66",X"E2",X"E2",
		X"0E",X"62",X"22",X"E2",X"0E",X"22",X"26",X"E2",X"0E",X"22",X"77",X"EE",X"0E",X"22",X"26",X"00",
		X"0E",X"6E",X"66",X"00",X"00",X"6E",X"EE",X"00",X"00",X"6E",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"E0",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"DD",X"EE",X"00",X"EE",X"DD",X"DD",X"00",X"EE",X"DD",X"DD",X"00",X"EE",X"EE",X"DD",
		X"00",X"CC",X"CC",X"EE",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CE",X"BC",X"00",X"BB",X"E2",X"EC",
		X"00",X"EE",X"EF",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"ED",X"00",X"00",X"F0",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"0E",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"EE",X"DD",X"EE",X"00",X"EC",X"CC",X"DD",
		X"00",X"EC",X"CE",X"DD",X"00",X"BB",X"CC",X"DE",X"00",X"EE",X"EE",X"DE",X"00",X"00",X"1B",X"CC",
		X"00",X"0E",X"EE",X"CC",X"00",X"0E",X"00",X"CC",X"00",X"ED",X"00",X"CE",X"00",X"ED",X"00",X"CE",
		X"00",X"DD",X"00",X"CE",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"EE",X"DD",X"00",
		X"00",X"CE",X"DD",X"00",X"00",X"CF",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"B6",X"ED",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EC",X"EE",X"00",X"F0",X"2E",X"CD",X"00",X"E0",X"F2",X"DD",
		X"00",X"00",X"EE",X"CD",X"00",X"00",X"DE",X"CC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0E",X"00",X"00",X"0E",X"ED",X"00",X"00",X"0E",X"ED",X"00",X"00",X"EF",X"DD",X"00",
		X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"EE",X"00",X"FC",X"CC",X"DD",
		X"00",X"EB",X"CC",X"DD",X"00",X"EE",X"CC",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"2F",X"DD",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"E0",X"CC",X"00",X"0E",X"00",X"CC",X"00",X"0E",X"00",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"ED",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CE",X"DD",X"00",X"00",X"BB",X"DD",X"00",X"00",X"FE",X"EC",X"E0",
		X"00",X"E0",X"CC",X"DE",X"00",X"00",X"EC",X"DE",X"00",X"00",X"2E",X"DE",X"00",X"00",X"B2",X"E0",
		X"00",X"00",X"EE",X"E0",X"00",X"0E",X"00",X"CE",X"00",X"ED",X"00",X"CE",X"00",X"ED",X"00",X"CE",
		X"00",X"0E",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"ED",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CF",X"DD",X"00",X"00",X"BE",X"DD",X"00",X"00",X"BE",X"DD",X"00",X"00",X"EE",X"DD",X"EE",
		X"00",X"E0",X"EE",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"00",X"EC",X"DE",X"00",X"00",X"FE",X"DE",
		X"00",X"00",X"EE",X"EC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"EE",X"00",X"00",X"BC",X"ED",X"00",
		X"00",X"EB",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0F",X"DD",X"00",
		X"00",X"EE",X"CE",X"EE",X"00",X"F0",X"CC",X"ED",X"00",X"00",X"EE",X"DD",X"00",X"00",X"B2",X"DD",
		X"00",X"00",X"EE",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DE",X"EE",X"00",X"00",X"E0",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"0E",X"00",X"00",X"BC",X"ED",X"00",
		X"00",X"FE",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"FE",X"DD",X"00",X"00",X"0E",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"EC",X"DE",X"00",X"00",X"2E",X"DE",
		X"00",X"00",X"E2",X"DE",X"00",X"00",X"DE",X"EE",X"00",X"00",X"E0",X"CE",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"BC",X"E0",X"00",X"00",X"EB",X"CE",X"00",X"00",X"EE",X"CE",X"00",
		X"00",X"0E",X"ED",X"00",X"00",X"F0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"2E",X"E0",
		X"00",X"00",X"EE",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"BC",X"E0",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"0F",X"CE",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"CD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"0E",X"EC",X"00",
		X"00",X"0E",X"2C",X"00",X"00",X"0E",X"BC",X"E0",X"00",X"0E",X"EB",X"E0",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"EC",X"00",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"0F",X"CE",X"00",
		X"00",X"EE",X"CE",X"00",X"00",X"F0",X"ED",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CD",X"00",X"00",X"0E",X"CE",X"00",X"00",X"0E",X"EC",X"00",
		X"00",X"0E",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EB",X"E0",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"FE",X"CC",X"E0",
		X"00",X"00",X"CE",X"E0",X"00",X"00",X"CD",X"E0",X"00",X"00",X"CD",X"00",X"00",X"00",X"CD",X"00",
		X"00",X"00",X"CD",X"00",X"00",X"00",X"CC",X"00",X"00",X"0E",X"EC",X"00",X"00",X"0E",X"EC",X"00",
		X"00",X"0E",X"EC",X"00",X"00",X"0E",X"BC",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"CE",X"00",X"00",X"EF",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"E0",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"ED",X"00",X"00",X"0E",X"CE",X"00",X"00",X"EE",X"CC",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"E0",X"00",X"00",X"DD",X"E0",
		X"00",X"0E",X"DD",X"E0",X"00",X"EE",X"CD",X"E0",X"00",X"ED",X"CE",X"00",X"00",X"ED",X"CC",X"00",
		X"00",X"EE",X"CE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"E0",
		X"00",X"0E",X"DD",X"E0",X"00",X"ED",X"ED",X"E0",X"00",X"ED",X"ED",X"00",X"00",X"0D",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"2E",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"EE",
		X"00",X"00",X"EE",X"3E",X"00",X"00",X"2E",X"E0",X"00",X"E0",X"22",X"EE",X"00",X"3E",X"22",X"2E",
		X"00",X"E3",X"22",X"2E",X"00",X"EE",X"22",X"E3",X"00",X"E2",X"22",X"3E",X"00",X"22",X"22",X"EE",
		X"00",X"22",X"32",X"EE",X"00",X"22",X"32",X"22",X"00",X"22",X"E2",X"22",X"00",X"3E",X"22",X"22",
		X"00",X"E2",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"E2",X"22",X"22",X"00",X"E2",X"22",X"22",
		X"00",X"EE",X"22",X"22",X"00",X"E3",X"22",X"22",X"00",X"3E",X"22",X"2E",X"00",X"07",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"F5",X"FE",
		X"00",X"00",X"55",X"5F",X"00",X"00",X"55",X"55",X"00",X"00",X"5E",X"55",X"00",X"00",X"EF",X"E5",
		X"00",X"06",X"EF",X"EF",X"00",X"00",X"EE",X"EF",X"00",X"00",X"00",X"FF",X"00",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"F5",X"00",X"EE",X"00",X"55",X"00",X"EE",X"00",X"55",X"00",X"EE",X"00",X"55",
		X"00",X"EE",X"06",X"E5",X"00",X"EE",X"00",X"E5",X"00",X"5E",X"00",X"E5",X"00",X"55",X"00",X"EE",
		X"AE",X"55",X"E6",X"E0",X"AE",X"55",X"00",X"00",X"0D",X"55",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"FC",X"FE",
		X"00",X"00",X"CC",X"CF",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CE",X"CC",X"00",X"00",X"EF",X"EC",
		X"00",X"06",X"EF",X"EF",X"00",X"00",X"EE",X"EF",X"00",X"00",X"00",X"FF",X"00",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"FC",X"00",X"EE",X"00",X"CC",X"00",X"EE",X"00",X"CC",X"00",X"EE",X"00",X"CC",
		X"00",X"EE",X"06",X"EC",X"00",X"EE",X"00",X"EC",X"00",X"BE",X"00",X"EC",X"00",X"CB",X"00",X"EE",
		X"AE",X"CB",X"E6",X"E0",X"AE",X"CC",X"00",X"00",X"0D",X"CC",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"00",X"BE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"55",X"55",X"00",X"0E",X"55",X"5E",X"00",X"0E",X"BB",X"BB",X"E0",X"0E",X"BB",X"BB",X"E0",
		X"0E",X"BB",X"BB",X"E0",X"E9",X"BB",X"BB",X"E0",X"E9",X"BB",X"BB",X"E0",X"E9",X"BB",X"BB",X"E0",
		X"E9",X"BB",X"BB",X"EE",X"7B",X"BB",X"BB",X"BE",X"E7",X"BB",X"BB",X"BE",X"00",X"BB",X"7B",X"7E",
		X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"00",X"30",X"0F",X"00",X"30",X"00",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"03",X"00",X"00",X"F0",X"F0",X"F0",
		X"00",X"01",X"20",X"00",X"00",X"11",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"E6",X"20",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EE",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"10",X"E1",X"00",X"00",X"1E",X"66",X"00",X"00",X"E6",X"E6",X"00",X"00",X"66",X"E6",X"00",
		X"00",X"16",X"66",X"00",X"00",X"66",X"E6",X"00",X"00",X"66",X"BE",X"00",X"00",X"66",X"BE",X"00",
		X"00",X"EE",X"BE",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",
		X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"01",X"20",X"00",X"00",X"11",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"ED",X"20",X"00",
		X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"EE",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"E1",X"00",X"00",X"0E",X"DD",X"00",X"00",X"ED",X"ED",X"00",X"00",X"DD",X"ED",X"00",
		X"00",X"3D",X"DD",X"00",X"00",X"DD",X"ED",X"00",X"00",X"DD",X"BE",X"00",X"00",X"DD",X"BE",X"00",
		X"00",X"EE",X"BE",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"CB",X"00",
		X"00",X"00",X"CB",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"EE",X"FF",X"E0",X"00",X"55",X"FE",X"FE",X"00",X"55",X"E5",X"F5",X"00",X"EE",X"55",X"F5",
		X"00",X"55",X"55",X"E5",X"00",X"55",X"55",X"55",X"00",X"55",X"EE",X"55",X"00",X"FF",X"F1",X"55",
		X"00",X"EE",X"1E",X"55",X"00",X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",
		X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"FF",X"00",
		X"00",X"E5",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"55",X"E5",X"E0",
		X"00",X"55",X"55",X"E0",X"00",X"55",X"55",X"00",X"00",X"FF",X"55",X"E0",X"00",X"EE",X"FF",X"E0",
		X"00",X"FF",X"EE",X"E0",X"00",X"FF",X"00",X"E0",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"EE",X"00",
		X"00",X"E0",X"FF",X"00",X"00",X"E0",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"EE",X"FF",X"00",
		X"00",X"5E",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"FF",X"EE",X"E0",X"00",X"EE",X"55",X"FE",X"00",X"00",X"E5",X"FF",X"00",X"00",X"EF",X"FF",
		X"00",X"0E",X"EE",X"FF",X"00",X"0E",X"0E",X"F5",X"00",X"0E",X"00",X"55",X"00",X"0E",X"00",X"55",
		X"00",X"0E",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"EE",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"E5",X"FF",X"00",X"00",X"5E",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"55",X"E0",
		X"00",X"65",X"55",X"FE",X"00",X"EF",X"55",X"FE",X"00",X"EE",X"E5",X"FE",X"00",X"0E",X"EF",X"EE",
		X"00",X"EF",X"EE",X"5E",X"00",X"EF",X"E0",X"5E",X"00",X"FF",X"E0",X"5E",X"00",X"FF",X"00",X"5E",
		X"00",X"EE",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"00",
		X"00",X"0E",X"EF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"E0",X"FF",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"E5",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"F5",X"FE",X"00",
		X"00",X"EF",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"EF",X"E5",X"00",
		X"00",X"EF",X"E6",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"00",
		X"00",X"0E",X"EF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"F5",X"FF",X"00",
		X"00",X"EF",X"FF",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"FF",X"E0",X"00",X"0E",X"EE",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EF",X"0E",X"00",X"00",X"EE",X"EF",X"00",X"00",X"5E",X"FF",X"00",X"00",X"5E",X"FF",X"00",
		X"00",X"F5",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"0E",X"FF",X"00",
		X"00",X"00",X"FF",X"E0",X"00",X"00",X"EE",X"EE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",
		X"00",X"00",X"EF",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"0E",X"00",X"00",X"EF",X"EF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"F5",X"FF",X"00",X"00",X"EF",X"FF",X"00",
		X"00",X"EE",X"FF",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"0E",X"55",X"00",
		X"00",X"EF",X"55",X"00",X"00",X"EF",X"F5",X"00",X"00",X"EF",X"EE",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5E",X"EE",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"65",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FE",X"00",X"00",X"0E",X"E5",X"00",X"00",X"EF",X"55",X"00",
		X"00",X"EF",X"55",X"00",X"00",X"EF",X"55",X"00",X"00",X"0E",X"E5",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E5",X"EE",X"00",
		X"00",X"E6",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EF",X"5E",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EF",X"0E",X"00",
		X"00",X"E6",X"EF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"FF",X"5E",X"00",X"00",X"EF",X"5E",X"00",X"00",X"EE",X"5E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"0E",X"EF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"EF",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"EF",X"55",X"00",X"00",X"EE",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E6",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"EF",X"5E",X"00",X"00",X"0E",X"EF",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"F0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"5E",X"00",
		X"00",X"0E",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"5E",X"00",X"00",X"EE",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"E0",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"EF",X"EE",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0E",X"FE",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"FE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"E5",X"E0",X"00",X"00",X"E5",X"E0",X"00",X"00",X"E5",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"EE",X"0E",X"00",X"00",X"BB",X"E9",X"F0",X"00",X"BB",X"E9",X"E0",X"00",X"BB",X"E9",X"F0",X"00",
		X"BB",X"E9",X"E1",X"00",X"BB",X"E9",X"EE",X"EE",X"BB",X"EE",X"BB",X"2E",X"BB",X"33",X"BB",X"2E",
		X"EE",X"EE",X"BB",X"EE",X"99",X"BB",X"BB",X"E2",X"99",X"BE",X"BB",X"2B",X"99",X"E9",X"EB",X"BB",
		X"99",X"E9",X"FB",X"99",X"99",X"E9",X"FE",X"9E",X"99",X"E9",X"EE",X"E0",X"EE",X"E9",X"F1",X"00",
		X"00",X"E9",X"9E",X"00",X"00",X"E9",X"E0",X"00",X"00",X"E9",X"F0",X"00",X"00",X"E9",X"E0",X"00",
		X"00",X"E9",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"EE",X"0E",X"00",X"00",X"AA",X"E9",X"F0",X"00",X"AA",X"E9",X"E0",X"00",X"AA",X"E9",X"F0",X"00",
		X"AA",X"E9",X"E0",X"00",X"EE",X"E9",X"E1",X"EE",X"BB",X"E9",X"EA",X"FE",X"BB",X"E9",X"FA",X"EE",
		X"BB",X"E9",X"EB",X"BB",X"BB",X"EE",X"FE",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"EB",X"BB",X"BB",X"BB",X"FE",X"EE",X"BB",X"BB",X"E9",X"EE",X"BB",X"BB",X"E9",X"F1",X"EE",
		X"BB",X"E9",X"BE",X"00",X"EE",X"E9",X"E0",X"00",X"00",X"E9",X"F0",X"00",X"00",X"E9",X"E0",X"00",
		X"00",X"E9",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"EE",X"E2",X"00",X"00",X"AA",X"E2",X"FE",X"00",X"AA",X"EE",X"EE",X"00",X"AA",X"EE",X"FE",X"00",
		X"AA",X"11",X"31",X"00",X"AA",X"EE",X"3E",X"EE",X"A2",X"1E",X"31",X"1E",X"A2",X"11",X"31",X"1E",
		X"EE",X"EE",X"1E",X"EE",X"99",X"EE",X"1E",X"E1",X"99",X"FE",X"E1",X"2F",X"99",X"3E",X"F1",X"2F",
		X"99",X"33",X"11",X"22",X"99",X"31",X"E1",X"2E",X"92",X"1F",X"11",X"E0",X"EE",X"11",X"F1",X"00",
		X"00",X"EE",X"E1",X"00",X"00",X"FE",X"33",X"00",X"00",X"EE",X"FE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"E2",X"FE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"31",X"30",X"00",
		X"EE",X"11",X"30",X"0F",X"AA",X"11",X"FE",X"00",X"AA",X"1E",X"EE",X"00",X"AA",X"33",X"EE",X"00",
		X"AA",X"11",X"EE",X"00",X"A3",X"E1",X"EE",X"EE",X"33",X"EE",X"EE",X"1E",X"A1",X"EE",X"EE",X"1E",
		X"E1",X"EE",X"EE",X"EE",X"93",X"1E",X"EE",X"E1",X"93",X"EE",X"EE",X"2F",X"99",X"EE",X"EE",X"2F",
		X"99",X"EE",X"EE",X"22",X"99",X"EE",X"EE",X"2E",X"92",X"EE",X"EE",X"E0",X"EE",X"EE",X"EE",X"00",
		X"00",X"EE",X"EE",X"10",X"00",X"EE",X"EE",X"10",X"00",X"31",X"EE",X"00",X"00",X"31",X"1E",X"00",
		X"F0",X"33",X"1E",X"00",X"00",X"03",X"13",X"00",X"0F",X"0E",X"01",X"F0",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"BA",X"00",X"00",X"1A",X"3A",X"00",X"00",X"3A",X"AA",X"00",X"00",X"AA",X"EE",X"00",
		X"00",X"AA",X"AE",X"00",X"00",X"EE",X"AE",X"00",X"00",X"EE",X"AA",X"00",X"00",X"A1",X"EA",X"E0",
		X"00",X"AA",X"EE",X"EE",X"00",X"EE",X"2A",X"BE",X"00",X"AA",X"1E",X"1E",X"00",X"AA",X"AE",X"E1",
		X"00",X"AA",X"AE",X"2B",X"00",X"E1",X"AA",X"9B",X"00",X"12",X"AA",X"99",X"00",X"12",X"AA",X"9E",
		X"00",X"22",X"AA",X"E0",X"00",X"22",X"AA",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"AA",X"00",
		X"00",X"EE",X"AE",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"A1",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",
		X"00",X"00",X"EA",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"A0",X"0A",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"0E",X"A0",X"00",X"00",X"0E",X"A0",X"00",X"00",X"0E",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"AA",X"00",
		X"00",X"EE",X"A3",X"00",X"00",X"EE",X"A1",X"00",X"00",X"AA",X"3E",X"00",X"00",X"AA",X"EE",X"00",
		X"0E",X"EE",X"A0",X"00",X"0E",X"AA",X"E0",X"00",X"EA",X"00",X"E0",X"00",X"AE",X"01",X"E0",X"00",
		X"AE",X"02",X"A0",X"00",X"AE",X"00",X"AE",X"00",X"AE",X"0A",X"AE",X"00",X"0A",X"EA",X"EE",X"00",
		X"EA",X"E2",X"AE",X"00",X"EE",X"22",X"EA",X"00",X"EA",X"E2",X"1A",X"00",X"EA",X"EE",X"EA",X"00",
		X"EE",X"EE",X"AA",X"00",X"0E",X"EE",X"AA",X"00",X"00",X"AE",X"3A",X"00",X"00",X"AE",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"E4",X"00",X"00",X"EE",X"EA",X"00",X"00",X"AA",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",
		X"00",X"FE",X"EE",X"00",X"0E",X"EE",X"77",X"EE",X"EA",X"E5",X"EE",X"4E",X"EE",X"55",X"AA",X"EE",
		X"EB",X"55",X"EE",X"E5",X"0E",X"AA",X"77",X"E5",X"00",X"EE",X"77",X"EE",X"00",X"BB",X"EE",X"9B",
		X"00",X"BB",X"EE",X"9B",X"00",X"9B",X"99",X"9B",X"00",X"22",X"99",X"BB",X"00",X"F2",X"99",X"99",
		X"00",X"E2",X"F0",X"2F",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"10",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"99",X"EE",X"00",X"00",X"E9",X"9E",X"00",X"11",X"9E",X"AE",X"00",X"11",X"9E",X"AE",
		X"00",X"11",X"21",X"E0",X"00",X"00",X"E1",X"00",X"00",X"EE",X"E1",X"E0",X"00",X"11",X"11",X"E3",
		X"00",X"11",X"EE",X"E0",X"00",X"EE",X"EE",X"EE",X"00",X"FE",X"EE",X"EE",X"00",X"EE",X"EE",X"22",
		X"00",X"EE",X"E1",X"FF",X"0E",X"F1",X"F1",X"EF",X"0E",X"FE",X"F3",X"E2",X"00",X"EE",X"13",X"F2",
		X"00",X"EE",X"13",X"EE",X"00",X"EE",X"11",X"00",X"00",X"3E",X"11",X"F0",X"00",X"31",X"EE",X"E0",
		X"00",X"3E",X"1E",X"E0",X"00",X"EE",X"EE",X"E0",X"00",X"3E",X"EE",X"0F",X"00",X"EE",X"E2",X"00",
		X"00",X"00",X"2E",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"1E",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"E0",X"00",X"01",X"1A",X"9E",X"11",X"11",X"1E",X"1E",X"11",
		X"11",X"1E",X"11",X"11",X"11",X"31",X"11",X"11",X"11",X"EE",X"EE",X"10",X"11",X"EE",X"EE",X"00",
		X"13",X"EE",X"EE",X"10",X"13",X"EE",X"EE",X"00",X"0E",X"EE",X"EE",X"00",X"0E",X"EE",X"EE",X"00",
		X"0E",X"1E",X"EE",X"1E",X"00",X"EE",X"EE",X"11",X"EE",X"EE",X"EE",X"10",X"11",X"EE",X"EE",X"E0",
		X"EE",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"E0",X"00",X"EE",X"EE",X"E0",X"00",X"EE",X"EE",X"E1",
		X"0E",X"1E",X"EE",X"E1",X"0E",X"1E",X"E3",X"31",X"0E",X"23",X"13",X"11",X"EE",X"2E",X"13",X"11",
		X"EE",X"31",X"13",X"E3",X"EE",X"11",X"33",X"10",X"00",X"11",X"33",X"10",X"00",X"E1",X"33",X"00",
		X"00",X"1E",X"1E",X"00",X"00",X"E1",X"11",X"00",X"00",X"EE",X"1E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"66",X"06",X"F0",X"00",X"22",X"22",X"00",X"66",X"2F",X"22",X"00",
		X"F6",X"00",X"66",X"20",X"00",X"20",X"66",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"F2",X"22",X"22",X"00",X"22",X"22",X"00",
		X"00",X"2F",X"22",X"00",X"00",X"22",X"22",X"20",X"00",X"22",X"22",X"00",X"02",X"22",X"02",X"00",
		X"00",X"22",X"02",X"00",X"06",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"06",X"00",X"02",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"02",X"20",X"00",X"06",X"00",X"20",X"00",
		X"02",X"00",X"20",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"02",X"00",X"20",X"02",X"00",
		X"00",X"22",X"02",X"00",X"00",X"F2",X"02",X"00",X"00",X"72",X"02",X"00",X"00",X"72",X"22",X"00",
		X"00",X"27",X"22",X"60",X"00",X"22",X"22",X"26",X"00",X"22",X"62",X"00",X"00",X"07",X"62",X"02",
		X"00",X"07",X"62",X"00",X"00",X"07",X"22",X"60",X"00",X"77",X"22",X"20",X"00",X"72",X"22",X"20",
		X"00",X"22",X"26",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"08",X"E0",X"00",X"00",X"08",X"E0",X"00",X"00",X"08",X"E0",X"00",X"00",X"08",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"08",X"00",
		X"00",X"0C",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"0C",X"08",X"00",X"00",X"0B",X"08",X"00",
		X"00",X"0C",X"08",X"00",X"00",X"0B",X"08",X"00",X"00",X"0C",X"E8",X"00",X"00",X"0C",X"FE",X"00",
		X"00",X"FE",X"FE",X"00",X"0F",X"EE",X"0F",X"F0",X"00",X"00",X"77",X"00",X"FF",X"FF",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"EF",X"EE",X"00",X"00",X"6E",X"5E",X"00",X"00",X"66",X"A1",X"00",
		X"00",X"66",X"EE",X"00",X"EE",X"AA",X"FF",X"00",X"E6",X"FF",X"FF",X"EE",X"0E",X"FF",X"EE",X"FF",
		X"0E",X"EF",X"FF",X"62",X"00",X"EF",X"66",X"2E",X"00",X"EE",X"EE",X"EF",X"00",X"FF",X"FE",X"BB",
		X"0E",X"FF",X"EE",X"BB",X"0E",X"FF",X"BB",X"BB",X"EF",X"EE",X"FF",X"EE",X"EF",X"55",X"EE",X"00",
		X"FE",X"A1",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"1E",X"00",X"00",X"00",X"1E",X"E0",X"00",X"00",X"EE",X"9E",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"E0",X"00",X"00",X"BB",X"E0",X"00",X"00",X"BB",X"E0",X"00",X"00",X"BB",X"E0",
		X"00",X"00",X"BB",X"EE",X"00",X"00",X"BE",X"FE",X"00",X"00",X"E7",X"FF",X"0F",X"F7",X"70",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"BE",X"E0",
		X"00",X"00",X"E0",X"E0",X"E0",X"00",X"00",X"EE",X"BE",X"00",X"00",X"AE",X"BB",X"00",X"E0",X"AE",
		X"EB",X"00",X"BE",X"FE",X"EB",X"77",X"BB",X"E7",X"F7",X"7F",X"77",X"77",X"00",X"00",X"07",X"00",
		X"00",X"77",X"01",X"77",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"F0",X"0E",X"E0",X"EE",X"00",X"0E",X"E0",
		X"ED",X"00",X"0E",X"EE",X"EE",X"00",X"0E",X"EB",X"00",X"00",X"0E",X"BB",X"AE",X"00",X"EE",X"EE",
		X"BB",X"77",X"E0",X"BB",X"7E",X"00",X"BB",X"77",X"F7",X"0F",X"EE",X"77",X"00",X"00",X"07",X"00",
		X"00",X"07",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"0E",X"F0",X"00",X"2E",X"0E",X"E0",X"00",X"22",X"0E",X"EE",X"00",
		X"22",X"0E",X"E2",X"00",X"22",X"0E",X"EE",X"00",X"22",X"0E",X"EE",X"00",X"22",X"33",X"22",X"F0",
		X"EE",X"EE",X"22",X"EE",X"E2",X"22",X"22",X"ED",X"E2",X"2E",X"22",X"2E",X"E2",X"E2",X"E2",X"2E",
		X"E2",X"EE",X"FE",X"E0",X"E2",X"0E",X"E0",X"00",X"EE",X"0E",X"EE",X"00",X"00",X"0E",X"F1",X"00",
		X"00",X"0E",X"2E",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"EE",X"E2",X"00",X"00",X"EE",X"E2",X"5E",X"00",X"EE",X"EE",X"EE",X"00",X"22",X"EE",X"5E",X"00",
		X"22",X"77",X"27",X"00",X"26",X"E2",X"7E",X"EE",X"E6",X"76",X"26",X"5E",X"E6",X"77",X"26",X"5E",
		X"EE",X"22",X"62",X"6E",X"EE",X"22",X"62",X"E5",X"E6",X"52",X"E2",X"65",X"EE",X"22",X"52",X"65",
		X"EE",X"22",X"52",X"22",X"22",X"26",X"E6",X"6E",X"22",X"65",X"76",X"E0",X"22",X"22",X"77",X"00",
		X"EE",X"66",X"22",X"00",X"EE",X"5E",X"22",X"00",X"00",X"EE",X"5E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"E6",X"5E",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"EE",X"DD",X"E0",X"00",X"CC",X"DE",X"DE",X"00",X"CC",X"EC",X"DC",X"00",X"EE",X"CC",X"DC",
		X"00",X"CC",X"CC",X"EC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"EE",X"CC",X"00",X"BB",X"F2",X"CC",
		X"00",X"EE",X"2E",X"CC",X"00",X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",
		X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"EE",X"DD",X"00",
		X"00",X"EC",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"CC",X"EC",X"E0",
		X"00",X"CC",X"CC",X"E0",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"CC",X"E0",X"00",X"EE",X"BB",X"E0",
		X"00",X"DD",X"EE",X"E0",X"00",X"DD",X"00",X"E0",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"EE",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"E0",X"DD",X"00",X"00",X"FE",X"DD",X"00",X"00",X"EE",X"DD",X"00",
		X"00",X"CE",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"BB",X"EE",X"E0",X"00",X"EE",X"CC",X"DE",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EB",X"DD",
		X"00",X"0E",X"EE",X"DD",X"00",X"0E",X"0E",X"DC",X"00",X"0E",X"00",X"CC",X"00",X"0E",X"00",X"CC",
		X"00",X"0E",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"EE",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"EC",X"DD",X"00",X"00",X"CE",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"CC",X"E0",
		X"00",X"FC",X"CC",X"DE",X"00",X"EB",X"CC",X"DE",X"00",X"EE",X"EC",X"DE",X"00",X"0E",X"EB",X"EE",
		X"00",X"ED",X"EE",X"CE",X"00",X"ED",X"E0",X"CE",X"00",X"DD",X"E0",X"CE",X"00",X"DD",X"00",X"CE",
		X"00",X"EE",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"00",
		X"00",X"0E",X"ED",X"00",X"00",X"FE",X"DD",X"00",X"00",X"E0",X"DD",X"00",X"00",X"BE",X"DD",X"00",
		X"00",X"EC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DE",X"00",
		X"00",X"EB",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"ED",X"EC",X"00",
		X"00",X"ED",X"EB",X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"00",
		X"00",X"0E",X"ED",X"00",X"00",X"F0",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",
		X"00",X"EB",X"DD",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"BB",X"E0",X"00",X"0E",X"EE",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EF",X"0E",X"00",X"00",X"EE",X"ED",X"00",X"00",X"CE",X"DD",X"00",X"00",X"CE",X"DD",X"00",
		X"00",X"FC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"0E",X"DD",X"00",
		X"00",X"00",X"DD",X"E0",X"00",X"00",X"EE",X"EE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",
		X"00",X"00",X"EB",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"0E",X"00",X"00",X"EF",X"ED",X"00",X"00",X"EE",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"EE",X"DD",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"ED",X"CC",X"00",X"00",X"ED",X"BC",X"00",X"00",X"ED",X"EE",X"00",X"00",X"ED",X"00",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"CE",X"EE",X"00",X"00",X"FE",X"DD",X"00",
		X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"ED",X"CC",X"00",
		X"00",X"ED",X"CC",X"00",X"00",X"ED",X"CC",X"00",X"00",X"0E",X"EC",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"EC",X"EE",X"00",
		X"00",X"EB",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",
		X"00",X"0E",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"0E",X"EE",X"00",X"00",X"ED",X"CE",X"00",
		X"00",X"DD",X"CC",X"00",X"00",X"DD",X"CC",X"00",X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EB",X"0E",X"00",
		X"00",X"EB",X"ED",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"DD",X"DE",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"DD",X"CE",X"00",X"00",X"ED",X"CE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"0E",X"ED",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"ED",X"CC",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"CC",X"00",X"00",X"ED",X"CC",X"00",X"00",X"EE",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EB",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"0E",X"DD",X"00",X"00",X"ED",X"DD",X"00",X"00",X"DD",X"DE",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"DD",X"CC",X"00",X"00",X"ED",X"CE",X"00",X"00",X"0E",X"ED",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"ED",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"F0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"CE",X"00",
		X"00",X"0E",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"EE",X"DD",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"DD",X"CE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"E0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"EE",X"DD",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"ED",X"EE",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"0E",X"DE",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"FE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EC",X"E0",X"00",
		X"00",X"EC",X"E0",X"00",X"00",X"EC",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",X"00",X"EE",X"3E",X"00",
		X"00",X"E3",X"3E",X"00",X"00",X"0E",X"E2",X"00",X"00",X"EE",X"22",X"00",X"00",X"E2",X"22",X"EE",
		X"00",X"E2",X"22",X"3E",X"00",X"22",X"22",X"EE",X"00",X"22",X"22",X"EE",X"00",X"22",X"22",X"E2",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"2E",X"22",X"22",X"00",X"EE",X"22",X"22",X"00",X"EE",X"22",X"2E",
		X"00",X"E2",X"22",X"2E",X"00",X"E2",X"22",X"EE",X"00",X"EE",X"22",X"E0",X"00",X"70",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"F5",X"00",X"00",X"EE",X"55",X"00",
		X"00",X"60",X"5E",X"E0",X"00",X"00",X"EF",X"E0",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"5E",
		X"00",X"00",X"FF",X"5E",X"00",X"00",X"EE",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"55",X"00",X"EE",X"00",X"5E",X"00",X"AA",X"00",X"5E",X"00",X"4E",X"06",X"5E",
		X"00",X"44",X"00",X"5E",X"0E",X"44",X"00",X"E0",X"E5",X"44",X"00",X"E0",X"E5",X"EE",X"00",X"00",
		X"55",X"EE",X"00",X"00",X"5E",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"FC",X"00",X"00",X"EE",X"CC",X"00",
		X"00",X"60",X"CE",X"E0",X"00",X"00",X"EF",X"E0",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"CE",
		X"00",X"00",X"FF",X"CE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"EE",X"00",X"CE",X"00",X"AA",X"00",X"CE",X"00",X"4E",X"06",X"CE",
		X"00",X"44",X"00",X"CE",X"0E",X"44",X"00",X"E0",X"EB",X"44",X"00",X"E0",X"EC",X"EE",X"00",X"00",
		X"CC",X"EE",X"00",X"00",X"CE",X"BB",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"00",
		X"E9",X"55",X"55",X"00",X"99",X"E5",X"55",X"00",X"9A",X"BE",X"EB",X"00",X"9A",X"BE",X"EB",X"00",
		X"92",X"BE",X"EB",X"00",X"92",X"BB",X"BE",X"00",X"92",X"BB",X"BE",X"00",X"92",X"BB",X"BE",X"00",
		X"99",X"BB",X"BE",X"00",X"99",X"BB",X"BE",X"00",X"99",X"BB",X"BE",X"70",X"00",X"77",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"F0",X"00",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"E2",X"00",X"00",X"00",X"E2",X"00",X"00",X"02",X"6E",X"00",X"00",X"02",X"6E",X"00",X"00",
		X"01",X"66",X"00",X"00",X"02",X"6E",X"00",X"00",X"02",X"E5",X"00",X"00",X"02",X"E5",X"00",X"00",
		X"00",X"E5",X"1E",X"00",X"00",X"6E",X"61",X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"6E",X"00",X"00",X"66",X"E0",X"00",X"00",X"66",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"E2",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"DE",X"00",X"00",X"03",X"DE",X"00",X"00",
		X"01",X"DD",X"00",X"00",X"01",X"DE",X"00",X"00",X"03",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EC",X"1E",X"00",X"00",X"DE",X"11",X"00",X"00",X"DD",X"11",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DE",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"55",X"5E",X"00",X"00",X"55",X"55",X"E0",X"0E",X"E5",X"55",X"5E",
		X"E5",X"55",X"55",X"5E",X"E5",X"55",X"55",X"5E",X"E6",X"55",X"EF",X"5E",X"0E",X"6F",X"EE",X"5E",
		X"00",X"EE",X"E0",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"55",X"E0",X"00",X"0E",X"5F",X"00",X"00",X"E5",X"EF",X"E0",X"00",X"E5",X"55",X"5E",X"00",
		X"0E",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"EE",X"FE",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"FF",X"0E",X"00",X"00",X"FE",X"0E",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"0E",X"55",X"FE",X"00",
		X"0E",X"E5",X"FE",X"00",X"0E",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"EE",X"00",
		X"00",X"F5",X"55",X"00",X"00",X"F6",X"55",X"00",X"00",X"EE",X"55",X"E0",X"00",X"EF",X"55",X"E0",
		X"00",X"FF",X"FF",X"E0",X"00",X"FF",X"EE",X"E0",X"00",X"FF",X"00",X"5E",X"00",X"FF",X"00",X"5E",
		X"00",X"FF",X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"0E",X"55",X"FE",X"00",
		X"E5",X"55",X"FE",X"00",X"E5",X"55",X"EE",X"00",X"0E",X"55",X"E0",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"FF",X"5E",X"00",X"00",X"EE",X"5E",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"FF",X"0E",X"00",X"00",X"FF",X"0E",X"00",X"00",X"FF",X"0E",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"00",X"E5",X"FE",X"00",X"0E",X"E5",X"FE",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"55",X"E0",X"00",X"00",X"55",X"E0",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"EE",X"00",X"00",X"EF",X"EF",X"00",X"00",X"FE",X"5E",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"65",X"00",X"00",X"FF",X"E5",X"00",X"00",X"FF",X"E5",X"00",X"00",X"FE",X"E5",X"00",
		X"00",X"E0",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"FE",X"00",X"0E",X"EE",X"FE",X"00",X"0E",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"F5",X"EE",X"00",X"00",X"E5",X"55",X"00",X"00",X"EE",X"5E",X"00",X"00",X"EF",X"5E",X"00",
		X"00",X"EF",X"F5",X"00",X"00",X"EF",X"E5",X"00",X"00",X"FF",X"E5",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"00",X"E0",X"FE",X"00",X"00",X"0E",X"FF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"F5",X"E0",X"00",
		X"00",X"EF",X"EE",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"5E",X"00",
		X"00",X"EF",X"55",X"00",X"00",X"EF",X"EF",X"00",X"00",X"EF",X"EE",X"00",X"00",X"EF",X"0E",X"00",
		X"00",X"EE",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"FE",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"5E",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"F5",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EF",X"5E",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"5E",X"FF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"F5",X"FF",X"00",X"00",X"F5",X"FE",X"00",
		X"00",X"EF",X"EE",X"00",X"00",X"EE",X"5E",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"5E",X"00",
		X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"EE",X"5E",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"5E",X"0E",X"00",X"00",X"5E",X"EF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"F5",X"FF",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"E6",X"E0",X"00",X"00",X"FF",X"E0",X"00",X"00",X"FF",X"5E",X"00",
		X"00",X"FF",X"5E",X"00",X"00",X"FF",X"EF",X"00",X"00",X"EE",X"5F",X"00",X"00",X"00",X"5F",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"0E",X"00",X"00",X"55",X"EF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"F5",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"E5",X"FE",X"00",X"00",X"F6",X"E0",X"00",X"00",X"FE",X"00",X"00",X"00",X"F6",X"E0",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"FF",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"65",X"EF",X"00",
		X"00",X"F5",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"E6",X"FF",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"FE",X"E0",X"00",X"00",X"FE",X"E0",X"00",X"00",X"FF",X"E0",X"00",
		X"00",X"FF",X"5E",X"00",X"00",X"FF",X"EE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"EE",X"00",
		X"00",X"65",X"FE",X"00",X"00",X"F5",X"FF",X"00",X"00",X"E6",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"FE",X"FE",X"00",X"00",X"FE",X"EE",X"00",X"00",X"FE",X"E0",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"FE",X"EE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"E6",X"EE",X"00",X"00",X"EF",X"FF",X"00",X"00",X"E6",X"FF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FE",X"EE",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EF",X"FE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"EF",X"EE",X"00",X"00",X"E6",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"E1",X"FF",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"FE",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"EF",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"FE",X"00",
		X"00",X"0F",X"FE",X"00",X"00",X"0F",X"FE",X"00",X"00",X"0F",X"FE",X"00",X"00",X"0E",X"FE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",
		X"BE",X"9E",X"0E",X"00",X"BE",X"99",X"EE",X"00",X"BE",X"E9",X"E9",X"00",X"BB",X"FE",X"E9",X"E0",
		X"EE",X"EB",X"EE",X"BE",X"9E",X"BB",X"BE",X"B9",X"99",X"EE",X"BB",X"B9",X"99",X"99",X"BB",X"9E",
		X"9E",X"99",X"BB",X"E0",X"9E",X"99",X"EB",X"00",X"EE",X"9E",X"EE",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"E0",X"9B",X"00",X"00",X"E0",X"BB",X"00",X"00",X"E0",X"BB",X"00",X"00",
		X"AE",X"B1",X"0E",X"00",X"AE",X"BB",X"EE",X"00",X"EA",X"B1",X"AA",X"00",X"EA",X"BB",X"EE",X"E0",
		X"BE",X"BB",X"EB",X"BE",X"BE",X"EE",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BE",X"EE",X"BB",X"BE",X"BE",X"BE",X"EB",X"E0",X"E0",X"BB",X"0E",X"00",
		X"E0",X"BE",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"9B",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E2",X"00",X"00",X"0F",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"E0",X"FE",X"EE",X"00",X"E0",X"EE",X"3E",X"00",X"E0",X"EF",X"EE",X"00",
		X"2E",X"EE",X"EE",X"00",X"2E",X"EE",X"EE",X"00",X"2E",X"E1",X"EE",X"00",X"22",X"11",X"EE",X"E0",
		X"EE",X"11",X"EE",X"FE",X"2E",X"EF",X"1E",X"FF",X"22",X"EF",X"1E",X"FF",X"92",X"33",X"1E",X"FE",
		X"2E",X"31",X"1E",X"E0",X"2E",X"11",X"EE",X"00",X"EE",X"F1",X"EE",X"00",X"00",X"1E",X"E0",X"00",
		X"00",X"E1",X"EE",X"00",X"00",X"EF",X"3E",X"00",X"0E",X"EF",X"31",X"00",X"FE",X"EF",X"11",X"00",
		X"0E",X"EF",X"EE",X"00",X"0E",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"13",X"00",X"00",X"0F",X"11",X"00",X"00",
		X"00",X"F1",X"00",X"00",X"E0",X"FE",X"EE",X"00",X"E0",X"EE",X"EE",X"F0",X"E0",X"1E",X"EE",X"00",
		X"2E",X"1E",X"EE",X"00",X"31",X"1E",X"EE",X"00",X"33",X"1E",X"E1",X"00",X"22",X"EE",X"E1",X"E0",
		X"11",X"EE",X"E1",X"FE",X"11",X"EE",X"E1",X"FF",X"22",X"EE",X"EE",X"FF",X"31",X"EE",X"EE",X"FE",
		X"31",X"EE",X"EE",X"E0",X"11",X"EE",X"EE",X"00",X"11",X"EE",X"EE",X"00",X"13",X"EE",X"E3",X"0F",
		X"13",X"E3",X"E3",X"00",X"31",X"1E",X"EE",X"F0",X"33",X"1E",X"EE",X"00",X"FE",X"1E",X"EE",X"F0",
		X"0E",X"EE",X"EE",X"00",X"01",X"32",X"33",X"00",X"01",X"22",X"33",X"00",X"00",X"E2",X"13",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"AA",X"EA",X"00",X"0E",X"AA",X"AE",X"00",X"0A",X"AA",X"AE",X"00",X"0A",X"AA",X"AE",X"00",
		X"00",X"AA",X"AE",X"00",X"00",X"AA",X"B3",X"00",X"00",X"A1",X"BE",X"00",X"00",X"AA",X"EE",X"00",
		X"00",X"EE",X"EE",X"E0",X"00",X"EE",X"A3",X"E0",X"00",X"AA",X"E3",X"EE",X"00",X"AA",X"EE",X"EE",
		X"00",X"AA",X"EE",X"2E",X"00",X"AA",X"EE",X"BE",X"00",X"AA",X"E9",X"9E",X"00",X"BB",X"E9",X"E0",
		X"00",X"B9",X"EE",X"00",X"00",X"B9",X"AE",X"00",X"00",X"99",X"AE",X"00",X"00",X"9E",X"AE",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"E3",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"EE",X"AA",X"00",
		X"00",X"AE",X"0A",X"00",X"00",X"2A",X"0A",X"00",X"00",X"EE",X"A1",X"00",X"00",X"0E",X"AA",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"0A",X"A0",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"AA",X"E0",X"00",X"00",X"2A",X"E0",X"00",X"00",X"E0",X"E0",X"00",X"EE",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"EA",X"22",X"00",X"00",X"E0",X"22",X"00",X"00",X"E0",X"E2",X"00",X"00",
		X"0A",X"E3",X"00",X"00",X"00",X"EA",X"00",X"00",X"0A",X"EA",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"E0",X"EE",X"00",X"00",X"E0",X"AE",X"E0",X"00",X"AE",X"3A",X"E0",X"00",X"AE",X"A3",X"E0",X"00",
		X"AA",X"EA",X"E0",X"00",X"AA",X"2A",X"AE",X"00",X"EE",X"EE",X"AE",X"00",X"0E",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"EE",X"AE",X"00",X"00",X"AA",X"CE",X"00",X"00",X"AE",X"CE",X"00",X"00",
		X"AA",X"EE",X"EE",X"00",X"EE",X"5E",X"77",X"00",X"EE",X"5E",X"EE",X"00",X"AA",X"55",X"AA",X"E0",
		X"EE",X"55",X"EE",X"E0",X"BB",X"AA",X"77",X"E0",X"EB",X"EE",X"BB",X"EE",X"EE",X"9B",X"EE",X"BE",
		X"0E",X"BB",X"EE",X"BE",X"00",X"BB",X"99",X"BE",X"00",X"2B",X"99",X"9E",X"00",X"B2",X"B2",X"9E",
		X"00",X"EF",X"FE",X"22",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"99",X"00",X"00",X"0E",X"99",X"00",X"00",X"E9",X"A1",X"00",X"00",X"E2",X"21",X"00",
		X"00",X"1E",X"11",X"00",X"00",X"1E",X"1E",X"F0",X"00",X"EE",X"1E",X"00",X"00",X"E1",X"EE",X"00",
		X"00",X"11",X"EE",X"00",X"F0",X"11",X"E1",X"F0",X"00",X"11",X"11",X"E0",X"0E",X"1F",X"1E",X"E0",
		X"E2",X"1F",X"1E",X"2E",X"22",X"E1",X"11",X"22",X"22",X"11",X"EE",X"22",X"E2",X"33",X"EE",X"2E",
		X"0E",X"31",X"31",X"E0",X"00",X"11",X"31",X"00",X"00",X"F1",X"33",X"00",X"F0",X"11",X"11",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0E",X"E2",X"00",
		X"00",X"0E",X"E3",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"11",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"99",X"00",X"10",X"E2",X"9E",X"00",X"10",X"11",X"E9",X"01",X"13",X"11",X"E1",X"01",X"10",
		X"01",X"EE",X"11",X"10",X"01",X"1E",X"11",X"30",X"0E",X"E1",X"1E",X"00",X"3E",X"E1",X"EE",X"00",
		X"3E",X"E1",X"EE",X"00",X"E1",X"11",X"EE",X"00",X"11",X"E1",X"EE",X"00",X"E1",X"EE",X"EE",X"01",
		X"EE",X"E1",X"E1",X"00",X"EE",X"E1",X"3E",X"00",X"11",X"E1",X"EE",X"00",X"11",X"EE",X"EE",X"00",
		X"E0",X"EE",X"EE",X"11",X"E0",X"EE",X"EE",X"11",X"E0",X"EE",X"EE",X"11",X"EE",X"EE",X"EE",X"11",
		X"EE",X"EE",X"33",X"31",X"EE",X"EE",X"3E",X"11",X"12",X"EE",X"33",X"10",X"E1",X"3E",X"33",X"30",
		X"E1",X"13",X"31",X"00",X"E1",X"33",X"31",X"00",X"EE",X"33",X"11",X"00",X"EE",X"11",X"1E",X"00",
		X"EE",X"11",X"EE",X"00",X"00",X"11",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",
		X"00",X"F6",X"22",X"00",X"00",X"22",X"00",X"00",X"06",X"FF",X"00",X"00",X"00",X"02",X"66",X"00",
		X"00",X"22",X"60",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"20",X"00",X"06",X"20",X"22",X"00",
		X"06",X"20",X"2F",X"00",X"00",X"20",X"2F",X"60",X"00",X"20",X"FF",X"00",X"00",X"F2",X"F2",X"06",
		X"F2",X"F2",X"F2",X"02",X"02",X"F2",X"22",X"02",X"00",X"26",X"22",X"00",X"0F",X"26",X"2F",X"00",
		X"00",X"26",X"2F",X"00",X"00",X"22",X"2F",X"00",X"00",X"62",X"22",X"60",X"60",X"62",X"02",X"22",
		X"00",X"62",X"02",X"02",X"00",X"22",X"F2",X"00",X"00",X"22",X"F2",X"00",X"00",X"22",X"02",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"20",X"00",X"00",X"06",X"26",X"60",X"00",X"22",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"20",X"00",X"00",X"20",X"20",X"02",X"00",
		X"00",X"60",X"02",X"00",X"00",X"20",X"06",X"00",X"00",X"26",X"20",X"66",X"00",X"02",X"60",X"06",
		X"00",X"07",X"00",X"02",X"00",X"07",X"02",X"02",X"00",X"27",X"22",X"00",X"00",X"26",X"22",X"00",
		X"60",X"26",X"26",X"00",X"00",X"27",X"66",X"00",X"00",X"27",X"62",X"00",X"00",X"27",X"27",X"00",
		X"00",X"27",X"22",X"00",X"00",X"27",X"72",X"00",X"00",X"27",X"72",X"00",X"00",X"27",X"72",X"60",
		X"00",X"27",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"86",X"00",
		X"00",X"00",X"C4",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"64",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"FF",X"00",X"00",X"70",X"FF",X"00",
		X"00",X"EF",X"F0",X"00",X"0F",X"7F",X"7F",X"00",X"00",X"00",X"0F",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"6E",X"E0",X"00",
		X"00",X"66",X"00",X"00",X"EE",X"AA",X"E0",X"00",X"66",X"FF",X"FE",X"00",X"66",X"FF",X"EE",X"E0",
		X"66",X"FF",X"FF",X"EE",X"E6",X"FF",X"66",X"FF",X"EA",X"FF",X"EE",X"FF",X"EA",X"FF",X"EB",X"BB",
		X"AA",X"FF",X"BA",X"BD",X"FF",X"FE",X"AA",X"BE",X"FF",X"EE",X"AA",X"E0",X"FF",X"EE",X"EE",X"00",
		X"EE",X"1E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"ED",X"00",X"00",
		X"00",X"ED",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EB",X"BB",X"00",X"00",X"0E",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"EE",X"F0",X"00",X"60",X"7E",X"7F",X"F0",X"7F",X"F7",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"0F",X"00",X"EC",X"00",X"E0",X"00",X"EC",X"0F",
		X"EE",X"00",X"EC",X"F0",X"BB",X"77",X"EC",X"97",X"77",X"70",X"7E",X"00",X"F0",X"00",X"77",X"70",
		X"00",X"00",X"10",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"EE",X"00",
		X"00",X"00",X"EA",X"00",X"00",X"00",X"AA",X"00",X"EE",X"00",X"AE",X"00",X"ED",X"00",X"AF",X"EE",
		X"DB",X"00",X"AC",X"EB",X"EB",X"00",X"AA",X"BB",X"EB",X"00",X"AE",X"EE",X"EE",X"77",X"EE",X"EE",
		X"EE",X"77",X"BB",X"BB",X"7E",X"00",X"BB",X"B7",X"77",X"70",X"E7",X"70",X"F0",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"E2",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"E0",X"2E",X"E0",X"00",X"20",X"22",X"E0",X"00",X"2E",X"E2",X"EE",X"00",X"22",X"FE",X"E2",X"00",
		X"EE",X"E2",X"EE",X"00",X"2E",X"22",X"2E",X"00",X"2E",X"EE",X"22",X"00",X"2E",X"22",X"22",X"00",
		X"2E",X"22",X"EE",X"00",X"E0",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E2",X"00",X"00",X"05",X"66",X"00",X"00",
		X"00",X"55",X"00",X"00",X"E0",X"5E",X"EE",X"00",X"E0",X"EE",X"7E",X"00",X"E0",X"E5",X"EE",X"00",
		X"6E",X"EE",X"EE",X"00",X"6E",X"22",X"EE",X"00",X"2E",X"62",X"EE",X"00",X"22",X"22",X"EE",X"E0",
		X"EE",X"22",X"EE",X"5E",X"2E",X"22",X"26",X"55",X"22",X"2E",X"26",X"55",X"E2",X"22",X"2E",X"5E",
		X"6E",X"2E",X"2E",X"E0",X"6E",X"22",X"2E",X"00",X"EE",X"52",X"22",X"00",X"E0",X"26",X"22",X"00",
		X"E0",X"22",X"EE",X"00",X"E0",X"E5",X"2E",X"00",X"0E",X"E5",X"27",X"00",X"5E",X"E5",X"77",X"00",
		X"0E",X"E5",X"EE",X"00",X"0E",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"CC",X"E0",X"0E",X"EC",X"CC",X"CE",
		X"EC",X"CC",X"CC",X"CE",X"EC",X"CC",X"CC",X"CE",X"EB",X"CC",X"EB",X"CE",X"0E",X"BB",X"EE",X"CE",
		X"00",X"EE",X"E0",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"CC",X"E0",X"00",X"0E",X"CD",X"00",X"00",X"EC",X"ED",X"E0",X"00",X"EC",X"CC",X"CE",X"00",
		X"0E",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"CC",X"00",X"00",X"EE",X"BE",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"0E",X"00",X"00",X"DE",X"0E",X"00",X"00",X"DE",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"0E",X"CC",X"DE",X"00",
		X"0E",X"EC",X"DE",X"00",X"0E",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"EE",X"00",
		X"00",X"BC",X"CC",X"00",X"00",X"BB",X"CC",X"00",X"00",X"EE",X"CC",X"E0",X"00",X"ED",X"CC",X"E0",
		X"00",X"DD",X"BB",X"E0",X"00",X"DD",X"EE",X"E0",X"00",X"DD",X"00",X"CE",X"00",X"DD",X"00",X"CE",
		X"00",X"DD",X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"0E",X"CC",X"DE",X"00",
		X"EC",X"CC",X"DE",X"00",X"EC",X"CC",X"EE",X"00",X"0E",X"CC",X"E0",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"BB",X"CE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"DD",X"BB",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"0E",X"00",X"00",X"DD",X"0E",X"00",X"00",X"DD",X"0E",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"00",X"EC",X"DE",X"00",X"0E",X"EC",X"DE",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"BC",X"EE",X"00",X"00",X"EB",X"ED",X"00",X"00",X"DE",X"CE",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"BC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DE",X"EC",X"00",
		X"00",X"E0",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"DE",X"00",X"0E",X"EE",X"DE",X"00",X"0E",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"EE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"BC",X"EE",X"00",X"00",X"EC",X"CC",X"00",X"00",X"EE",X"CE",X"00",X"00",X"ED",X"CE",X"00",
		X"00",X"ED",X"BC",X"00",X"00",X"ED",X"EC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"00",X"E0",X"DE",X"00",X"00",X"0E",X"DD",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"BC",X"E0",X"00",
		X"00",X"EB",X"EE",X"00",X"00",X"0E",X"EC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"ED",X"CC",X"00",X"00",X"ED",X"EB",X"00",X"00",X"ED",X"EE",X"00",X"00",X"ED",X"0E",X"00",
		X"00",X"EE",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"DE",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"CE",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"BC",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"ED",X"CE",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"CD",X"00",X"00",X"DD",X"CD",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"CE",X"DD",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DE",X"00",
		X"00",X"EB",X"EE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"ED",X"00",X"00",X"DD",X"ED",X"00",X"00",X"DD",X"ED",X"00",X"00",X"EE",X"CE",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CE",X"0E",X"00",X"00",X"CE",X"ED",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DD",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"EB",X"E0",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"CE",X"00",
		X"00",X"DD",X"CE",X"00",X"00",X"DD",X"ED",X"00",X"00",X"EE",X"CD",X"00",X"00",X"00",X"CD",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"0E",X"00",X"00",X"CC",X"ED",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"EC",X"DE",X"00",X"00",X"DB",X"E0",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"E0",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"ED",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"BC",X"ED",X"00",
		X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"DE",X"E0",X"00",X"00",X"DE",X"E0",X"00",X"00",X"DD",X"E0",X"00",
		X"00",X"DD",X"CE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"BC",X"EE",X"00",
		X"00",X"BC",X"DE",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"DE",X"DE",X"00",X"00",X"DE",X"EE",X"00",X"00",X"DE",X"E0",X"00",
		X"00",X"DD",X"E0",X"00",X"00",X"DE",X"EE",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DE",X"DD",X"00",X"00",X"DE",X"EE",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EB",X"FE",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"EF",X"DD",X"00",X"00",X"E2",X"DD",X"00",X"00",X"DE",X"DD",X"00",
		X"00",X"DE",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"EF",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"DE",X"00",X"00",X"0E",X"DE",X"00",
		X"00",X"0F",X"DE",X"00",X"00",X"0F",X"DE",X"00",X"00",X"0F",X"DE",X"00",X"00",X"0E",X"DE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"EE",X"2E",X"00",X"00",X"E2",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"EE",X"00",X"22",X"22",X"E3",
		X"00",X"22",X"22",X"EE",X"0E",X"22",X"22",X"EE",X"E3",X"22",X"22",X"2E",X"E3",X"22",X"22",X"2E",
		X"EE",X"22",X"22",X"2E",X"00",X"22",X"22",X"2E",X"00",X"22",X"22",X"33",X"00",X"22",X"22",X"2E",
		X"00",X"E3",X"E3",X"EE",X"00",X"3E",X"EE",X"E0",X"00",X"3E",X"EE",X"E0",X"00",X"E2",X"EE",X"E0",
		X"00",X"22",X"22",X"3E",X"00",X"22",X"22",X"EE",X"00",X"22",X"22",X"00",X"00",X"77",X"07",X"00",
		X"70",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FF",X"55",X"00",X"00",X"EF",X"EE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"E5",X"E0",
		X"00",X"00",X"E5",X"E0",X"00",X"EE",X"EE",X"E0",X"00",X"AE",X"EE",X"00",X"00",X"AA",X"00",X"00",
		X"0E",X"4A",X"00",X"00",X"0E",X"EA",X"00",X"00",X"E0",X"4A",X"00",X"00",X"5E",X"EE",X"00",X"00",
		X"55",X"EE",X"60",X"00",X"55",X"EE",X"00",X"00",X"E5",X"5E",X"00",X"00",X"0E",X"55",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"EE",X"0E",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FF",X"CC",X"00",X"00",X"EF",X"EE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"EC",X"E0",
		X"00",X"00",X"EC",X"E0",X"00",X"EE",X"EE",X"E0",X"00",X"AE",X"EE",X"00",X"00",X"AA",X"00",X"00",
		X"0E",X"4A",X"00",X"00",X"0E",X"EA",X"00",X"00",X"E0",X"4A",X"00",X"00",X"BE",X"EE",X"00",X"00",
		X"CB",X"EE",X"60",X"00",X"CC",X"EE",X"00",X"00",X"EC",X"BE",X"00",X"00",X"0E",X"CB",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"EE",X"0E",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",
		X"E5",X"55",X"55",X"00",X"9E",X"55",X"55",X"00",X"9E",X"BB",X"BB",X"00",X"AE",X"BB",X"BB",X"00",
		X"AE",X"BB",X"BB",X"00",X"A9",X"EB",X"BB",X"00",X"2A",X"EB",X"BB",X"00",X"2A",X"EB",X"BB",X"00",
		X"2A",X"EB",X"BB",X"00",X"2A",X"EA",X"AB",X"00",X"2A",X"EA",X"AB",X"00",X"22",X"BA",X"7B",X"00",
		X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"30",X"30",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"30",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"32",X"00",X"00",
		X"01",X"02",X"00",X"00",X"01",X"22",X"00",X"00",X"30",X"2E",X"00",X"00",X"10",X"25",X"00",X"00",
		X"10",X"55",X"00",X"00",X"20",X"25",X"00",X"00",X"20",X"52",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"22",X"55",X"00",X"00",
		X"23",X"55",X"00",X"00",X"21",X"55",X"E0",X"00",X"01",X"E5",X"6E",X"00",X"00",X"6E",X"6E",X"00",
		X"0E",X"6E",X"E0",X"00",X"0E",X"66",X"00",X"00",X"0E",X"66",X"00",X"00",X"00",X"6E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"32",X"00",X"00",
		X"01",X"02",X"00",X"00",X"01",X"22",X"00",X"00",X"30",X"2E",X"00",X"00",X"10",X"2C",X"00",X"00",
		X"10",X"CC",X"00",X"00",X"00",X"2C",X"00",X"00",X"00",X"C2",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"03",X"CC",X"00",X"00",X"01",X"CC",X"E0",X"00",X"01",X"EC",X"DE",X"00",X"00",X"DE",X"DE",X"00",
		X"0E",X"DE",X"E0",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DE",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",
		X"0E",X"EF",X"0E",X"00",X"0E",X"EF",X"EF",X"00",X"0E",X"EF",X"EE",X"00",X"EE",X"5E",X"5E",X"00",
		X"5F",X"55",X"55",X"00",X"5E",X"55",X"55",X"00",X"5E",X"55",X"FF",X"00",X"6F",X"FF",X"EE",X"00",
		X"EE",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"EF",X"00",X"00",
		X"0F",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"5E",X"55",X"0E",X"00",
		X"5E",X"55",X"EF",X"00",X"E6",X"55",X"FF",X"00",X"0E",X"FF",X"5E",X"00",X"0F",X"EE",X"55",X"00",
		X"0E",X"E0",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",
		X"0E",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"55",X"EE",X"00",X"00",
		X"55",X"EF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"EF",X"EF",X"00",X"00",X"EE",X"5E",X"E0",X"00",
		X"0E",X"55",X"5E",X"00",X"00",X"55",X"55",X"00",X"00",X"EE",X"55",X"00",X"00",X"FE",X"55",X"00",
		X"0F",X"FF",X"65",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"FE",X"E5",X"00",X"00",X"E0",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"E5",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"5F",X"0E",X"00",X"E6",X"55",X"EE",X"00",
		X"0E",X"55",X"EF",X"00",X"0F",X"55",X"FF",X"00",X"0E",X"FE",X"FF",X"00",X"0E",X"EE",X"EE",X"00",
		X"F0",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E5",X"5E",X"00",X"00",X"55",X"55",X"00",X"00",
		X"E5",X"5F",X"00",X"00",X"E6",X"5F",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"55",X"EE",X"00",
		X"00",X"55",X"FF",X"00",X"0E",X"55",X"FF",X"00",X"F0",X"EE",X"FF",X"00",X"00",X"FE",X"EF",X"00",
		X"00",X"F6",X"55",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"5E",X"E0",X"00",X"00",X"55",X"5E",X"00",X"00",X"E5",X"5F",X"00",X"00",
		X"E5",X"5F",X"00",X"00",X"0E",X"5E",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"55",X"0E",X"00",
		X"00",X"55",X"EF",X"00",X"0F",X"55",X"EF",X"00",X"0F",X"E1",X"FF",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"FE",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"55",X"00",X"00",X"FE",X"55",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"0E",X"5E",X"E0",X"00",X"0E",X"55",X"E0",X"00",
		X"00",X"5E",X"E0",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"E5",X"EE",X"00",X"00",X"F1",X"EE",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"FE",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"E6",X"5E",X"E0",X"00",X"EE",X"55",X"E0",X"00",
		X"0E",X"5E",X"E0",X"00",X"00",X"5E",X"E0",X"00",X"00",X"EF",X"00",X"00",X"0E",X"5E",X"00",X"00",
		X"0E",X"55",X"00",X"00",X"F0",X"55",X"EE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"EF",X"FF",X"00",
		X"00",X"EE",X"FF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FE",X"55",X"00",
		X"00",X"E0",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"E0",X"00",X"00",X"E5",X"FE",X"00",
		X"00",X"55",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"0F",X"5E",X"E0",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",X"0E",X"00",X"00",X"EF",X"EF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"E0",X"00",X"00",X"E5",X"FE",X"00",
		X"00",X"55",X"FE",X"00",X"0F",X"5E",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"EF",X"E0",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"FE",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"5E",X"FE",X"00",
		X"00",X"55",X"FE",X"00",X"0E",X"55",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"00",X"5E",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E1",X"00",X"00",
		X"00",X"FE",X"E0",X"00",X"00",X"EE",X"FE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"5E",X"EE",X"00",X"00",X"55",X"FE",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"E1",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E0",X"FE",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"5E",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"0F",X"5E",X"00",X"00",X"0F",X"5E",X"E0",X"00",
		X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"5E",X"FF",X"00",X"00",X"5E",X"FE",X"00",
		X"00",X"5E",X"EE",X"00",X"00",X"E5",X"E0",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"FE",X"00",X"00",X"5E",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"E5",X"FE",X"00",X"00",X"1E",X"E0",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FE",X"00",X"00",X"E5",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"99",X"99",X"00",X"EE",X"99",X"99",X"00",X"BB",X"EE",X"99",X"00",
		X"BB",X"BB",X"99",X"00",X"EB",X"BB",X"EE",X"E0",X"EB",X"EE",X"BB",X"E0",X"EB",X"99",X"BB",X"00",
		X"BB",X"99",X"BB",X"00",X"EE",X"99",X"BE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"99",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"BB",X"AA",X"00",X"EE",X"BB",X"AA",X"00",X"AA",X"BB",X"EE",X"00",
		X"AA",X"BB",X"BB",X"00",X"EE",X"EE",X"BB",X"E0",X"BB",X"BB",X"BB",X"E0",X"BB",X"BB",X"BB",X"E0",
		X"BE",X"BB",X"BB",X"E0",X"EF",X"EE",X"BB",X"00",X"0E",X"1E",X"BB",X"00",X"00",X"BB",X"EE",X"00",
		X"00",X"1E",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"3F",X"00",X"00",
		X"00",X"3F",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",
		X"03",X"22",X"F0",X"00",X"EE",X"EF",X"00",X"00",X"3E",X"EF",X"30",X"00",X"EE",X"EE",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"F2",X"00",X"2E",X"EE",X"EE",X"00",
		X"2E",X"33",X"E2",X"00",X"EE",X"F1",X"EE",X"E0",X"EE",X"FF",X"E2",X"E0",X"EE",X"3F",X"E2",X"00",
		X"2E",X"11",X"E2",X"00",X"E1",X"11",X"2E",X"00",X"E1",X"13",X"EE",X"00",X"EE",X"13",X"00",X"00",
		X"E1",X"EE",X"EE",X"00",X"E1",X"FE",X"3E",X"00",X"E1",X"FE",X"1E",X"00",X"11",X"EE",X"1E",X"00",
		X"1E",X"E2",X"EE",X"00",X"EE",X"22",X"03",X"00",X"00",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"1E",X"00",X"00",X"03",X"22",X"00",X"00",
		X"03",X"22",X"11",X"00",X"EE",X"EF",X"11",X"00",X"3E",X"EF",X"11",X"00",X"E1",X"EE",X"10",X"00",
		X"11",X"EE",X"1E",X"00",X"1E",X"EE",X"13",X"00",X"EE",X"EE",X"12",X"00",X"3E",X"EE",X"3E",X"00",
		X"13",X"EE",X"13",X"00",X"11",X"EE",X"1E",X"E0",X"EE",X"EE",X"13",X"E0",X"1E",X"EE",X"11",X"00",
		X"2E",X"EE",X"E1",X"00",X"1E",X"EE",X"2E",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"33",X"00",
		X"3E",X"EE",X"13",X"00",X"EE",X"EE",X"33",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"00",
		X"EE",X"E2",X"EE",X"00",X"EE",X"22",X"03",X"00",X"10",X"22",X"00",X"00",X"11",X"2E",X"00",X"00",
		X"31",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2B",X"EA",X"00",X"00",X"2B",X"AE",X"00",X"00",X"00",X"AA",X"00",X"00",X"A2",X"AA",X"00",X"00",
		X"AA",X"AA",X"EE",X"00",X"EE",X"A1",X"AA",X"00",X"EE",X"33",X"3A",X"00",X"0E",X"A3",X"BA",X"00",
		X"0E",X"A3",X"EA",X"00",X"0E",X"AA",X"EE",X"00",X"0E",X"AA",X"EE",X"00",X"0E",X"AA",X"3E",X"00",
		X"0E",X"AA",X"EE",X"00",X"EE",X"A3",X"BB",X"00",X"EE",X"A3",X"9B",X"00",X"0E",X"39",X"99",X"00",
		X"EE",X"99",X"99",X"00",X"EB",X"99",X"EE",X"00",X"EB",X"99",X"00",X"00",X"E9",X"EE",X"00",X"00",
		X"E9",X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AE",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"A1",X"00",X"00",X"00",X"AE",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AE",X"00",X"00",
		X"00",X"AE",X"00",X"00",X"0A",X"0A",X"00",X"00",X"AA",X"0A",X"00",X"00",X"AE",X"EE",X"00",X"00",
		X"E0",X"0E",X"00",X"00",X"0E",X"AA",X"00",X"00",X"0E",X"EA",X"00",X"00",X"AE",X"EA",X"00",X"00",
		X"AE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"AE",X"AA",X"00",X"00",X"A1",X"AE",X"00",X"00",
		X"EA",X"AA",X"00",X"00",X"2A",X"EE",X"00",X"00",X"EE",X"AE",X"00",X"00",X"3E",X"AA",X"00",X"00",
		X"EE",X"AA",X"00",X"00",X"E2",X"E3",X"00",X"00",X"2A",X"AE",X"00",X"00",X"AE",X"E1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"77",X"00",X"AE",X"EE",X"77",X"00",X"AA",X"55",X"AA",X"00",
		X"AA",X"5E",X"EE",X"00",X"EE",X"EE",X"77",X"00",X"BB",X"EE",X"BB",X"00",X"BB",X"BE",X"EE",X"00",
		X"EB",X"BB",X"EE",X"00",X"EE",X"9B",X"99",X"E0",X"0E",X"B9",X"9B",X"E0",X"00",X"B9",X"2B",X"E0",
		X"00",X"FE",X"E0",X"20",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"F1",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"1A",X"00",
		X"00",X"22",X"12",X"00",X"EE",X"EE",X"EE",X"00",X"E1",X"E2",X"EE",X"00",X"EE",X"1E",X"EE",X"00",
		X"0E",X"11",X"1E",X"00",X"00",X"31",X"11",X"00",X"0E",X"33",X"E1",X"00",X"E2",X"13",X"E1",X"00",
		X"2E",X"13",X"EE",X"00",X"2F",X"11",X"EE",X"E0",X"2E",X"11",X"EE",X"E0",X"22",X"11",X"EE",X"00",
		X"EE",X"11",X"EE",X"00",X"00",X"1E",X"1E",X"00",X"0F",X"E1",X"33",X"00",X"0E",X"11",X"E1",X"00",
		X"0E",X"E1",X"EE",X"00",X"0E",X"EE",X"EE",X"00",X"0E",X"2E",X"EE",X"00",X"3E",X"E2",X"EE",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"22",X"E0",X"00",X"00",X"22",X"E0",X"00",X"00",X"E2",X"E0",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E0",X"21",X"00",X"11",X"2E",X"01",X"00",X"1A",X"99",X"11",X"00",X"1A",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"1E",X"00",X"3E",X"E1",X"EE",X"00",X"E1",X"EE",X"EE",X"00",
		X"3E",X"11",X"EE",X"00",X"11",X"EE",X"EE",X"00",X"11",X"EE",X"33",X"00",X"E1",X"EE",X"11",X"00",
		X"E1",X"EE",X"11",X"01",X"EE",X"EE",X"EE",X"10",X"EE",X"11",X"EE",X"00",X"3E",X"E1",X"EE",X"00",
		X"1E",X"E1",X"11",X"00",X"11",X"1E",X"EE",X"10",X"00",X"EE",X"E3",X"10",X"EE",X"1E",X"E3",X"10",
		X"E1",X"EE",X"E3",X"30",X"E1",X"EE",X"E3",X"00",X"31",X"EE",X"EE",X"00",X"13",X"31",X"EE",X"00",
		X"11",X"1E",X"11",X"00",X"12",X"11",X"11",X"00",X"11",X"11",X"EE",X"00",X"11",X"11",X"E0",X"00",
		X"EE",X"11",X"E1",X"00",X"EE",X"1E",X"03",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"02",X"00",X"6F",X"00",
		X"02",X"20",X"02",X"00",X"00",X"F0",X"F0",X"00",X"00",X"F0",X"20",X"00",X"62",X"F0",X"02",X"00",
		X"F0",X"FF",X"02",X"00",X"02",X"2F",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"26",X"00",X"00",
		X"00",X"26",X"00",X"20",X"60",X"26",X"00",X"20",X"FF",X"22",X"02",X"00",X"F2",X"22",X"22",X"00",
		X"22",X"22",X"22",X"00",X"02",X"22",X"20",X"00",X"02",X"22",X"00",X"00",X"00",X"22",X"00",X"20",
		X"00",X"22",X"00",X"20",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"62",X"02",X"00",X"00",X"00",X"62",X"60",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"02",X"00",X"60",X"22",X"00",X"00",X"20",X"62",X"60",X"00",
		X"00",X"62",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"62",X"02",X"00",X"62",X"62",X"60",X"20",X"20",X"26",X"60",X"00",X"00",X"26",X"22",X"60",
		X"00",X"22",X"22",X"60",X"00",X"22",X"20",X"60",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"70",X"20",X"00",X"00",X"72",X"20",X"00",X"00",X"72",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"4C",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"E7",X"F7",X"00",
		X"00",X"F7",X"F7",X"00",X"77",X"00",X"77",X"00",X"00",X"00",X"F0",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E0",X"00",X"00",X"E6",X"FE",X"00",X"00",X"06",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"0E",X"AE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"6E",X"FF",X"EE",X"00",
		X"66",X"FE",X"FF",X"E0",X"66",X"FE",X"66",X"FE",X"AA",X"FF",X"6B",X"FF",X"FF",X"FF",X"BF",X"BE",
		X"FF",X"FF",X"BB",X"E0",X"FF",X"EE",X"BB",X"00",X"FF",X"EE",X"EE",X"00",X"EE",X"EE",X"E0",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"9E",X"00",X"00",
		X"0E",X"9E",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"BB",X"EE",X"00",X"00",X"EB",X"BB",X"00",
		X"00",X"0E",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"77",X"00",X"77",X"F7",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"0E",X"AA",X"00",X"00",X"EB",X"EE",X"00",X"00",X"0E",X"EF",X"00",
		X"00",X"00",X"CC",X"00",X"E7",X"7F",X"CC",X"F7",X"70",X"07",X"EE",X"07",X"00",X"00",X"77",X"00",
		X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"CC",X"00",X"E0",X"00",X"EC",X"00",X"E0",X"00",X"EC",X"EE",
		X"E0",X"00",X"CC",X"CC",X"EE",X"00",X"CC",X"EE",X"BE",X"00",X"EE",X"E0",X"BE",X"07",X"BB",X"E0",
		X"BB",X"07",X"BB",X"CC",X"EE",X"7F",X"EE",X"77",X"70",X"07",X"77",X"07",X"10",X"10",X"07",X"06",
		X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"22",X"EE",X"00",X"00",X"22",X"E2",X"00",X"EE",X"EE",X"22",X"00",
		X"22",X"22",X"22",X"00",X"22",X"22",X"EE",X"00",X"22",X"EE",X"EE",X"00",X"22",X"22",X"E2",X"00",
		X"EE",X"22",X"EE",X"00",X"00",X"22",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"66",X"00",X"00",
		X"02",X"62",X"50",X"00",X"26",X"E5",X"00",X"00",X"66",X"E5",X"60",X"00",X"EE",X"EE",X"00",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"26",X"EE",X"00",X"EE",X"66",X"52",X"00",X"2E",X"22",X"EE",X"00",
		X"2E",X"2E",X"E2",X"00",X"EE",X"EE",X"EE",X"E0",X"EE",X"EE",X"E2",X"E0",X"EE",X"EE",X"E2",X"00",
		X"2E",X"EE",X"E2",X"00",X"E2",X"E2",X"2E",X"00",X"E2",X"22",X"EE",X"00",X"EE",X"22",X"00",X"00",
		X"E6",X"66",X"EE",X"00",X"E6",X"5E",X"2E",X"00",X"E6",X"5E",X"7E",X"00",X"22",X"EE",X"6E",X"00",
		X"2E",X"E6",X"EE",X"00",X"EE",X"22",X"06",X"00",X"00",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",
		X"0E",X"ED",X"0E",X"00",X"0E",X"ED",X"ED",X"00",X"0E",X"ED",X"EE",X"00",X"EE",X"CE",X"CE",X"00",
		X"CF",X"CC",X"CC",X"00",X"CE",X"CC",X"CC",X"00",X"CE",X"CC",X"BB",X"00",X"BB",X"BB",X"EE",X"00",
		X"EE",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"ED",X"00",X"00",
		X"0F",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"CE",X"CC",X"0E",X"00",
		X"CE",X"CC",X"ED",X"00",X"EB",X"CC",X"DD",X"00",X"0E",X"BB",X"CD",X"00",X"0F",X"EE",X"CC",X"00",
		X"0E",X"E0",X"CC",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",
		X"0E",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"CC",X"EE",X"00",X"00",
		X"CC",X"ED",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EB",X"ED",X"00",X"00",X"EE",X"CE",X"E0",X"00",
		X"0E",X"CC",X"CE",X"00",X"00",X"CC",X"CC",X"00",X"00",X"EE",X"CC",X"00",X"00",X"DE",X"CC",X"00",
		X"0F",X"DD",X"CC",X"00",X"00",X"DD",X"BE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"DE",X"EC",X"00",X"00",X"E0",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"EC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"CD",X"0E",X"00",X"EB",X"CC",X"EE",X"00",
		X"0E",X"CC",X"ED",X"00",X"0F",X"CC",X"DD",X"00",X"0E",X"BE",X"DD",X"00",X"0E",X"EE",X"EE",X"00",
		X"F0",X"DD",X"CC",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EC",X"CE",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"EC",X"CD",X"00",X"00",X"EB",X"CD",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"CC",X"EE",X"00",
		X"00",X"CC",X"DD",X"00",X"0E",X"CC",X"DD",X"00",X"F0",X"EE",X"DD",X"00",X"00",X"DE",X"ED",X"00",
		X"00",X"DB",X"CC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"CE",X"E0",X"00",X"00",X"CC",X"CE",X"00",X"00",X"EC",X"CD",X"00",X"00",
		X"EC",X"CD",X"00",X"00",X"0E",X"CE",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"CC",X"0E",X"00",
		X"00",X"CC",X"ED",X"00",X"0F",X"CC",X"ED",X"00",X"0F",X"E2",X"DD",X"00",X"00",X"DE",X"DD",X"00",
		X"00",X"DE",X"ED",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DE",X"CC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"0E",X"CE",X"E0",X"00",X"0E",X"CC",X"E0",X"00",
		X"00",X"CE",X"E0",X"00",X"00",X"CD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"EE",X"00",X"00",X"D2",X"EE",X"00",X"00",X"DE",X"DD",X"00",
		X"00",X"DE",X"ED",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"EB",X"CE",X"E0",X"00",X"EE",X"CC",X"E0",X"00",
		X"0E",X"CE",X"E0",X"00",X"00",X"CE",X"E0",X"00",X"00",X"ED",X"00",X"00",X"0E",X"CE",X"00",X"00",
		X"0E",X"CC",X"00",X"00",X"F0",X"CC",X"EE",X"00",X"00",X"EE",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"EE",X"DD",X"00",X"00",X"DD",X"ED",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DE",X"CC",X"00",
		X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"E0",X"00",X"00",X"EC",X"DE",X"00",
		X"00",X"CC",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"0F",X"CE",X"E0",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"E2",X"0E",X"00",X"00",X"EF",X"ED",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"E0",X"00",X"00",X"EC",X"DE",X"00",
		X"00",X"CC",X"DE",X"00",X"0F",X"CE",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EF",X"E0",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"DE",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"CE",X"DE",X"00",
		X"00",X"CC",X"DE",X"00",X"0E",X"CC",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"00",X"CE",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"DE",X"E0",X"00",X"00",X"EE",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CE",X"EE",X"00",X"00",X"CC",X"DE",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E0",X"DE",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"CE",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"0F",X"CE",X"00",X"00",X"0F",X"CE",X"E0",X"00",
		X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CE",X"DD",X"00",X"00",X"CE",X"DE",X"00",
		X"00",X"CE",X"EE",X"00",X"00",X"EC",X"E0",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CE",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"EC",X"DE",X"00",X"00",X"2E",X"E0",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DE",X"00",X"00",X"EC",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E2",X"EE",X"00",X"EE",X"22",X"2E",X"00",X"E3",X"22",X"22",X"00",X"EE",X"22",X"22",X"00",
		X"0E",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"0E",X"22",X"2E",X"E0",X"0E",X"23",X"22",X"E0",
		X"0E",X"2E",X"22",X"00",X"EE",X"2E",X"22",X"00",X"E2",X"EE",X"22",X"00",X"33",X"EE",X"22",X"00",
		X"EE",X"22",X"22",X"00",X"EE",X"22",X"22",X"EE",X"E2",X"22",X"22",X"3E",X"E2",X"22",X"22",X"3E",
		X"EE",X"22",X"22",X"EE",X"0E",X"22",X"32",X"00",X"0E",X"22",X"32",X"00",X"0E",X"22",X"EE",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"0E",X"22",X"22",X"00",X"70",X"07",X"77",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"5F",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"E5",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",
		X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"60",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"E0",X"00",X"EF",X"00",X"E4",X"00",X"FF",X"00",X"E5",X"E0",X"EF",X"00",X"E5",X"E0",X"0E",X"00",
		X"5E",X"E0",X"00",X"00",X"55",X"E0",X"00",X"00",X"E5",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"E5",X"E4",X"60",X"00",X"55",X"5E",X"00",X"00",X"55",X"5E",X"00",X"00",X"55",X"5E",X"00",X"00",
		X"E5",X"E0",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"CF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FC",X"00",X"00",X"EC",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"60",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"E0",X"00",X"EF",X"00",X"E4",X"00",X"FF",X"00",X"EC",X"E0",X"EF",X"00",X"EC",X"E0",X"0E",X"00",
		X"CE",X"E0",X"00",X"00",X"CB",X"E0",X"00",X"00",X"EC",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"EC",X"E4",X"60",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"CE",X"00",X"00",
		X"EC",X"E0",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",
		X"55",X"55",X"E0",X"00",X"55",X"55",X"5E",X"00",X"5B",X"BB",X"BB",X"00",X"5B",X"BB",X"BB",X"00",
		X"5B",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"00",
		X"E5",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"70",X"E5",X"BB",X"BB",X"07",X"75",X"BB",X"BB",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"0F",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"F0",X"03",X"03",X"00",X"00",X"F0",X"F0",X"00",
		X"00",X"30",X"00",X"00",X"03",X"22",X"00",X"00",X"21",X"00",X"00",X"00",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"BE",X"00",X"00",X"10",X"BE",X"00",X"00",
		X"11",X"BE",X"00",X"00",X"31",X"BE",X"00",X"00",X"13",X"EF",X"00",X"00",X"31",X"5F",X"00",X"00",
		X"E1",X"5E",X"00",X"00",X"66",X"E5",X"00",X"00",X"66",X"E5",X"00",X"00",X"E6",X"E5",X"00",X"00",
		X"0E",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"30",X"00",X"00",X"03",X"22",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"00",
		X"00",X"BE",X"00",X"00",X"30",X"BE",X"00",X"00",X"13",X"EF",X"00",X"00",X"33",X"CF",X"00",X"00",
		X"E3",X"CE",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"ED",X"EC",X"00",X"00",
		X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
