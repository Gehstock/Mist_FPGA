library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"60",X"CB",X"BE",X"CB",X"86",X"CB",X"6E",X"28",X"02",X"3E",X"02",X"DD",X"77",X"02",X"DD",X"36",
		X"03",X"0A",X"DD",X"36",X"04",X"00",X"3E",X"00",X"CD",X"A0",X"1B",X"CD",X"21",X"40",X"C3",X"44",
		X"40",X"21",X"53",X"41",X"CD",X"39",X"1D",X"CD",X"39",X"1D",X"CD",X"39",X"1D",X"DD",X"7E",X"02",
		X"FE",X"02",X"20",X"03",X"21",X"98",X"41",X"CD",X"39",X"1D",X"21",X"B1",X"41",X"CD",X"39",X"1D",
		X"CD",X"39",X"41",X"C9",X"EF",X"DD",X"E5",X"CD",X"73",X"3B",X"DD",X"E1",X"CD",X"53",X"1B",X"DD",
		X"35",X"01",X"20",X"17",X"DD",X"36",X"01",X"14",X"DD",X"7E",X"00",X"D6",X"01",X"27",X"DD",X"77",
		X"00",X"CD",X"39",X"41",X"DD",X"7E",X"00",X"A7",X"CA",X"1F",X"41",X"DD",X"35",X"03",X"20",X"07",
		X"DD",X"36",X"03",X"0A",X"DD",X"34",X"04",X"3A",X"04",X"60",X"A7",X"20",X"13",X"21",X"53",X"41",
		X"DD",X"CB",X"04",X"46",X"20",X"05",X"CD",X"39",X"1D",X"18",X"03",X"CD",X"46",X"41",X"18",X"B4",
		X"21",X"7F",X"41",X"DD",X"7E",X"02",X"FE",X"02",X"20",X"03",X"21",X"98",X"41",X"DD",X"CB",X"04",
		X"46",X"20",X"05",X"CD",X"39",X"1D",X"18",X"03",X"CD",X"46",X"41",X"21",X"00",X"90",X"DD",X"7E",
		X"02",X"FE",X"02",X"28",X"1B",X"CB",X"6E",X"C2",X"44",X"40",X"21",X"00",X"60",X"CB",X"A6",X"CB",
		X"96",X"21",X"17",X"60",X"11",X"0C",X"60",X"AF",X"32",X"2A",X"60",X"01",X"1A",X"60",X"18",X"19",
		X"CB",X"76",X"C2",X"44",X"40",X"21",X"00",X"60",X"CB",X"9E",X"CB",X"8E",X"21",X"18",X"60",X"11",
		X"0F",X"60",X"AF",X"32",X"2B",X"60",X"01",X"21",X"60",X"AF",X"12",X"13",X"12",X"13",X"12",X"E5",
		X"C5",X"E1",X"01",X"01",X"07",X"D7",X"3A",X"02",X"90",X"07",X"07",X"E6",X"03",X"5F",X"16",X"00",
		X"21",X"44",X"06",X"19",X"7E",X"E1",X"3C",X"77",X"3A",X"04",X"60",X"3D",X"32",X"04",X"60",X"3A",
		X"5B",X"6B",X"3D",X"32",X"5B",X"6B",X"3A",X"91",X"6E",X"3D",X"32",X"91",X"6E",X"DD",X"E1",X"CD",
		X"7C",X"1B",X"21",X"00",X"60",X"CB",X"FE",X"CB",X"C6",X"21",X"DB",X"61",X"36",X"00",X"21",X"0B",
		X"60",X"36",X"00",X"CD",X"21",X"40",X"DD",X"E1",X"C9",X"DD",X"E5",X"06",X"02",X"21",X"D9",X"D2",
		X"CD",X"95",X"1E",X"DD",X"E1",X"C9",X"5E",X"23",X"56",X"23",X"46",X"3E",X"24",X"EB",X"77",X"23",
		X"10",X"FC",X"C9",X"25",X"D1",X"0D",X"19",X"1E",X"1D",X"24",X"16",X"18",X"1B",X"0E",X"24",X"0C",
		X"18",X"12",X"17",X"66",X"D1",X"13",X"1D",X"18",X"24",X"0C",X"18",X"17",X"1D",X"12",X"17",X"1E",
		X"0E",X"24",X"1D",X"18",X"24",X"19",X"15",X"0A",X"22",X"CE",X"D1",X"03",X"0A",X"17",X"0D",X"25",
		X"D2",X"16",X"19",X"1E",X"1C",X"11",X"24",X"24",X"01",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",
		X"24",X"24",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"25",X"D2",X"16",X"19",X"1E",X"1C",X"11",X"24",
		X"24",X"02",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"24",X"0B",X"1E",X"1D",X"1D",X"18",
		X"17",X"D4",X"D2",X"04",X"1D",X"12",X"16",X"0E",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"62",
		X"00",X"42",X"00",X"42",X"05",X"42",X"02",X"42",X"02",X"42",X"00",X"42",X"02",X"42",X"00",X"42",
		X"00",X"42",X"02",X"42",X"02",X"42",X"02",X"42",X"02",X"42",X"02",X"42",X"02",X"42",X"02",X"42",
		X"0C",X"42",X"0C",X"42",X"0C",X"42",X"0C",X"42",X"0C",X"42",X"0C",X"42",X"0C",X"42",X"0C",X"42",
		X"01",X"00",X"02",X"00",X"10",X"06",X"00",X"10",X"20",X"30",X"60",X"70",X"02",X"40",X"50",X"FD",
		X"21",X"00",X"6C",X"DD",X"21",X"06",X"6C",X"FD",X"36",X"02",X"00",X"01",X"00",X"18",X"21",X"3C",
		X"43",X"DD",X"7E",X"00",X"E6",X"03",X"20",X"07",X"DD",X"36",X"00",X"00",X"C3",X"17",X"43",X"E5",
		X"DD",X"CB",X"00",X"56",X"28",X"15",X"DD",X"36",X"00",X"00",X"CF",X"23",X"36",X"00",X"FD",X"7E",
		X"02",X"A7",X"C2",X"16",X"43",X"CD",X"9C",X"43",X"C3",X"16",X"43",X"FD",X"34",X"02",X"CB",X"47",
		X"28",X"1B",X"DD",X"CB",X"00",X"86",X"DD",X"CB",X"00",X"CE",X"CF",X"71",X"23",X"36",X"80",X"FD",
		X"7E",X"02",X"FE",X"01",X"C2",X"16",X"43",X"CD",X"9C",X"43",X"C3",X"16",X"43",X"C5",X"DD",X"E5",
		X"CF",X"E5",X"DD",X"E1",X"79",X"FE",X"10",X"38",X"08",X"FD",X"7E",X"02",X"FE",X"01",X"C2",X"13",
		X"43",X"DD",X"CB",X"01",X"76",X"28",X"09",X"DD",X"35",X"02",X"20",X"0F",X"DD",X"CB",X"01",X"B6",
		X"EB",X"CF",X"FD",X"E5",X"01",X"99",X"42",X"C5",X"E9",X"FD",X"E1",X"FD",X"7E",X"02",X"FE",X"01",
		X"C2",X"13",X"43",X"DD",X"CB",X"01",X"7E",X"CA",X"13",X"43",X"DD",X"6E",X"00",X"26",X"00",X"29",
		X"11",X"D0",X"41",X"19",X"CF",X"7E",X"47",X"23",X"7E",X"23",X"E5",X"21",X"00",X"B0",X"FE",X"40",
		X"38",X"05",X"D6",X"40",X"21",X"00",X"C0",X"87",X"C6",X"80",X"4F",X"FE",X"E0",X"28",X"1E",X"DD",
		X"7E",X"03",X"E6",X"0F",X"81",X"77",X"DD",X"7E",X"03",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"5F",
		X"DD",X"7E",X"04",X"E6",X"03",X"07",X"07",X"07",X"07",X"83",X"77",X"18",X"11",X"DD",X"CB",X"04",
		X"7E",X"28",X"0B",X"DD",X"CB",X"04",X"BE",X"DD",X"7E",X"03",X"E6",X"07",X"81",X"77",X"DD",X"7E",
		X"05",X"2F",X"E6",X"0F",X"81",X"C6",X"10",X"77",X"E1",X"11",X"03",X"00",X"DD",X"19",X"10",X"A8",
		X"C3",X"13",X"43",X"DD",X"E1",X"C1",X"E1",X"11",X"04",X"00",X"19",X"DD",X"23",X"0C",X"79",X"FE",
		X"10",X"20",X"0A",X"FD",X"7E",X"02",X"FD",X"77",X"05",X"FD",X"36",X"02",X"00",X"05",X"C2",X"21",
		X"42",X"FD",X"7E",X"02",X"FD",X"86",X"05",X"C0",X"CD",X"9C",X"43",X"C9",X"1E",X"6C",X"DA",X"45",
		X"2A",X"6C",X"63",X"46",X"32",X"6C",X"37",X"47",X"49",X"6C",X"A0",X"49",X"56",X"6C",X"E1",X"49",
		X"68",X"6C",X"22",X"46",X"73",X"6C",X"E1",X"49",X"85",X"6C",X"22",X"46",X"90",X"6C",X"22",X"46",
		X"9B",X"6C",X"09",X"48",X"AC",X"6C",X"05",X"48",X"BA",X"6C",X"2D",X"49",X"CC",X"6C",X"F1",X"48",
		X"DA",X"6C",X"7E",X"46",X"F1",X"6C",X"B2",X"48",X"FE",X"6C",X"E1",X"49",X"10",X"6D",X"4E",X"4A",
		X"2D",X"6D",X"4E",X"4A",X"4A",X"6D",X"4E",X"4A",X"67",X"6D",X"4E",X"4A",X"84",X"6D",X"4E",X"4A",
		X"A1",X"6D",X"4E",X"4A",X"BE",X"6D",X"4E",X"4A",X"DB",X"6D",X"4E",X"4A",X"3E",X"9F",X"32",X"00",
		X"B0",X"32",X"00",X"C0",X"C6",X"20",X"30",X"F6",X"C9",X"DD",X"36",X"01",X"00",X"DD",X"5E",X"00",
		X"16",X"00",X"21",X"06",X"6C",X"19",X"36",X"00",X"3A",X"02",X"6C",X"FE",X"01",X"C0",X"CD",X"9C",
		X"43",X"C9",X"00",X"00",X"F8",X"03",X"BF",X"03",X"89",X"03",X"56",X"03",X"26",X"03",X"FA",X"02",
		X"CE",X"02",X"A6",X"02",X"80",X"02",X"5C",X"02",X"3A",X"02",X"1A",X"02",X"FC",X"01",X"DF",X"01",
		X"C4",X"01",X"AB",X"01",X"93",X"01",X"7D",X"01",X"67",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",
		X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E2",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",
		X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",
		X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4B",X"00",
		X"47",X"00",X"43",X"00",X"3F",X"00",X"3C",X"00",X"39",X"00",X"D5",X"21",X"00",X"00",X"78",X"A7",
		X"28",X"0A",X"CB",X"3F",X"30",X"01",X"19",X"EB",X"29",X"EB",X"18",X"F3",X"D1",X"79",X"CB",X"3A",
		X"CB",X"1B",X"A7",X"C8",X"CB",X"27",X"30",X"F6",X"19",X"18",X"F3",X"FD",X"E5",X"FD",X"21",X"00",
		X"00",X"11",X"00",X"01",X"78",X"B1",X"28",X"18",X"AF",X"ED",X"42",X"38",X"04",X"FD",X"19",X"18",
		X"F7",X"09",X"CB",X"38",X"CB",X"19",X"78",X"B1",X"28",X"06",X"CB",X"3A",X"CB",X"1B",X"30",X"E8",
		X"FD",X"E5",X"D1",X"FD",X"E1",X"C9",X"DD",X"CB",X"01",X"EE",X"DD",X"6E",X"00",X"26",X"00",X"29",
		X"11",X"92",X"44",X"19",X"CF",X"4E",X"23",X"06",X"00",X"DD",X"E5",X"D1",X"13",X"13",X"13",X"ED",
		X"B0",X"C9",X"C2",X"44",X"CC",X"44",X"71",X"45",X"F7",X"44",X"E7",X"44",X"00",X"45",X"61",X"45",
		X"09",X"45",X"12",X"45",X"1B",X"45",X"86",X"45",X"2A",X"45",X"45",X"45",X"D2",X"44",X"3A",X"45",
		X"51",X"45",X"92",X"45",X"9B",X"45",X"A4",X"45",X"AD",X"45",X"B6",X"45",X"BF",X"45",X"C8",X"45",
		X"D1",X"45",X"09",X"00",X"00",X"0F",X"F0",X"60",X"50",X"EE",X"81",X"04",X"05",X"00",X"00",X"0F",
		X"F6",X"FE",X"14",X"40",X"00",X"0A",X"48",X"00",X"0A",X"06",X"0E",X"0C",X"20",X"11",X"09",X"00",
		X"11",X"0F",X"80",X"01",X"81",X"01",X"08",X"0F",X"AD",X"01",X"0F",X"00",X"01",X"0F",X"00",X"F0",
		X"1C",X"1C",X"5E",X"05",X"04",X"03",X"50",X"08",X"60",X"00",X"0F",X"57",X"01",X"0F",X"36",X"F0",
		X"08",X"80",X"03",X"0F",X"18",X"08",X"77",X"50",X"01",X"08",X"FF",X"03",X"0F",X"07",X"07",X"00",
		X"A0",X"01",X"08",X"00",X"00",X"0F",X"07",X"00",X"A0",X"00",X"01",X"0E",X"00",X"03",X"0F",X"01",
		X"03",X"0F",X"F0",X"67",X"00",X"AA",X"00",X"03",X"02",X"04",X"0F",X"A0",X"03",X"0F",X"30",X"03",
		X"0F",X"F0",X"00",X"10",X"03",X"40",X"06",X"06",X"FF",X"00",X"0A",X"10",X"00",X"0C",X"01",X"00",
		X"0C",X"FF",X"01",X"40",X"02",X"0B",X"00",X"00",X"0C",X"01",X"00",X"0C",X"88",X"02",X"88",X"02",
		X"02",X"0F",X"80",X"03",X"0F",X"00",X"00",X"0F",X"00",X"F0",X"06",X"1C",X"1D",X"BB",X"18",X"03",
		X"50",X"0F",X"01",X"03",X"00",X"00",X"03",X"00",X"00",X"F0",X"07",X"1C",X"1D",X"0E",X"0E",X"03",
		X"50",X"14",X"01",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"03",X"C0",X"00",X"00",X"00",
		X"00",X"07",X"C0",X"00",X"00",X"00",X"0B",X"50",X"00",X"0F",X"60",X"00",X"0F",X"F0",X"03",X"03",
		X"04",X"02",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"4C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"73",X"4D",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"4D",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"4E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"4E",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"4F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"B1",
		X"4F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"4F",X"DD",X"CB",X"01",X"6E",X"20",X"04",
		X"CD",X"76",X"44",X"C9",X"DD",X"7E",X"07",X"DD",X"BE",X"08",X"38",X"0F",X"28",X"0D",X"DD",X"7E",
		X"03",X"DD",X"86",X"09",X"30",X"10",X"DD",X"34",X"04",X"18",X"0B",X"DD",X"7E",X"03",X"DD",X"96",
		X"0A",X"30",X"03",X"DD",X"35",X"04",X"DD",X"77",X"03",X"DD",X"35",X"07",X"DD",X"7E",X"06",X"DD",
		X"96",X"0B",X"DD",X"77",X"06",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"05",X"20",X"03",X"CD",X"A9",
		X"43",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"76",X"44",X"C9",X"DD",X"7E",X"06",X"DD",
		X"BE",X"07",X"38",X"0F",X"28",X"0D",X"DD",X"7E",X"03",X"DD",X"86",X"08",X"30",X"10",X"DD",X"34",
		X"04",X"18",X"0B",X"DD",X"7E",X"03",X"DD",X"96",X"09",X"30",X"03",X"DD",X"35",X"04",X"DD",X"77",
		X"03",X"DD",X"CB",X"01",X"F6",X"DD",X"7E",X"0A",X"DD",X"77",X"02",X"DD",X"35",X"06",X"C0",X"CD",
		X"A9",X"43",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"76",X"44",X"C9",X"DD",X"7E",X"06",
		X"DD",X"86",X"03",X"DD",X"77",X"03",X"DD",X"A6",X"07",X"C0",X"CD",X"A9",X"43",X"C9",X"DD",X"CB",
		X"01",X"6E",X"20",X"08",X"CD",X"76",X"44",X"DD",X"CB",X"01",X"A6",X"C9",X"DD",X"7E",X"0C",X"A7",
		X"20",X"04",X"CD",X"A9",X"43",X"C9",X"DD",X"7E",X"09",X"A7",X"20",X"43",X"DD",X"CB",X"01",X"66",
		X"20",X"1D",X"DD",X"CB",X"01",X"E6",X"DD",X"7E",X"12",X"DD",X"77",X"03",X"DD",X"7E",X"13",X"DD",
		X"77",X"04",X"DD",X"7E",X"14",X"DD",X"77",X"06",X"DD",X"7E",X"15",X"DD",X"77",X"07",X"C9",X"DD",
		X"7E",X"03",X"DD",X"96",X"16",X"30",X"03",X"DD",X"35",X"04",X"DD",X"77",X"03",X"DD",X"7E",X"06",
		X"DD",X"96",X"16",X"30",X"03",X"DD",X"35",X"07",X"DD",X"77",X"06",X"DD",X"35",X"0C",X"C9",X"DD",
		X"7E",X"0F",X"DD",X"BE",X"0D",X"20",X"08",X"DD",X"36",X"0F",X"00",X"DD",X"35",X"09",X"C9",X"DD",
		X"7E",X"0F",X"DD",X"BE",X"0E",X"38",X"20",X"28",X"1E",X"DD",X"7E",X"03",X"DD",X"96",X"0B",X"30",
		X"03",X"DD",X"35",X"04",X"DD",X"77",X"03",X"DD",X"7E",X"06",X"DD",X"96",X"11",X"30",X"03",X"DD",
		X"35",X"07",X"DD",X"77",X"06",X"18",X"1C",X"DD",X"7E",X"03",X"DD",X"86",X"0A",X"30",X"03",X"DD",
		X"34",X"04",X"DD",X"77",X"03",X"DD",X"7E",X"06",X"DD",X"86",X"10",X"30",X"03",X"DD",X"34",X"07",
		X"DD",X"77",X"06",X"DD",X"34",X"0F",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"08",X"CD",X"76",X"44",
		X"DD",X"CB",X"01",X"A6",X"C9",X"DD",X"CB",X"01",X"66",X"20",X"33",X"DD",X"7E",X"16",X"C6",X"02",
		X"DD",X"77",X"16",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"0B",X"DD",X"77",X"11",X"DD",X"77",X"14",
		X"DD",X"7E",X"15",X"C6",X"03",X"DD",X"77",X"15",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"08",X"DD",
		X"77",X"0E",X"E6",X"0F",X"FE",X"0F",X"20",X"38",X"DD",X"CB",X"01",X"E6",X"18",X"32",X"DD",X"7E",
		X"0B",X"E6",X"0F",X"20",X"04",X"CD",X"A9",X"43",X"C9",X"DD",X"7E",X"16",X"D6",X"07",X"DD",X"77",
		X"16",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"0B",X"DD",X"77",X"11",X"DD",X"77",X"14",X"DD",X"7E",
		X"15",X"D6",X"0A",X"DD",X"77",X"15",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"08",X"DD",X"77",X"0E",
		X"DD",X"7E",X"03",X"DD",X"CB",X"01",X"5E",X"20",X"0B",X"C6",X"1A",X"DD",X"77",X"03",X"DD",X"CB",
		X"01",X"DE",X"18",X"09",X"D6",X"18",X"DD",X"77",X"03",X"DD",X"CB",X"01",X"9E",X"DD",X"7E",X"06",
		X"C6",X"04",X"38",X"05",X"DD",X"77",X"06",X"18",X"0A",X"DD",X"7E",X"06",X"D6",X"04",X"38",X"ED",
		X"DD",X"77",X"06",X"DD",X"7E",X"09",X"C6",X"01",X"30",X"02",X"3E",X"00",X"DD",X"77",X"09",X"DD",
		X"7E",X"0F",X"C6",X"04",X"30",X"03",X"DD",X"34",X"10",X"DD",X"77",X"0F",X"DD",X"CB",X"01",X"F6",
		X"DD",X"36",X"02",X"02",X"C9",X"CD",X"A9",X"43",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",
		X"76",X"44",X"C9",X"DD",X"7E",X"05",X"FE",X"00",X"20",X"04",X"CD",X"A9",X"43",X"C9",X"DD",X"7E",
		X"0C",X"FE",X"00",X"20",X"08",X"30",X"06",X"DD",X"36",X"0C",X"00",X"18",X"6D",X"DD",X"6E",X"03",
		X"DD",X"66",X"04",X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"19",X"DD",X"75",X"03",X"DD",X"74",X"04",
		X"DD",X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"19",X"DD",X"75",X"06",
		X"DD",X"74",X"07",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"DD",X"4E",X"0A",X"06",X"00",X"CB",X"79",
		X"28",X"01",X"05",X"09",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"5E",X"0D",X"DD",X"56",X"0E",
		X"EB",X"AF",X"ED",X"52",X"F2",X"7E",X"48",X"11",X"00",X"00",X"EB",X"AF",X"ED",X"52",X"DD",X"5E",
		X"0C",X"16",X"00",X"AF",X"ED",X"52",X"28",X"09",X"FA",X"91",X"48",X"79",X"ED",X"44",X"DD",X"77",
		X"0A",X"DD",X"7E",X"0C",X"DD",X"96",X"0F",X"DD",X"77",X"0C",X"DD",X"7E",X"09",X"DD",X"96",X"10",
		X"DD",X"77",X"09",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"05",X"DD",X"77",
		X"08",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"05",X"CD",X"76",X"44",X"18",X"29",X"DD",X"7E",X"09",
		X"A7",X"20",X"04",X"CD",X"A9",X"43",X"C9",X"DD",X"7E",X"03",X"DD",X"86",X"0A",X"30",X"03",X"DD",
		X"34",X"04",X"DD",X"77",X"03",X"DD",X"7E",X"06",X"DD",X"86",X"0B",X"30",X"03",X"DD",X"34",X"07",
		X"DD",X"77",X"06",X"DD",X"35",X"09",X"DD",X"CB",X"01",X"F6",X"DD",X"7E",X"0C",X"DD",X"77",X"02",
		X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"05",X"CD",X"76",X"44",X"18",X"26",X"DD",X"6E",X"03",X"DD",
		X"66",X"04",X"DD",X"5E",X"09",X"DD",X"56",X"0A",X"19",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",
		X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"0B",X"DD",X"56",X"0C",X"19",X"DD",X"75",X"06",X"DD",
		X"74",X"07",X"DD",X"CB",X"01",X"F6",X"DD",X"7E",X"0D",X"DD",X"77",X"02",X"C9",X"DD",X"CB",X"01",
		X"6E",X"20",X"04",X"CD",X"76",X"44",X"C9",X"DD",X"7E",X"0A",X"DD",X"BE",X"0B",X"30",X"20",X"28",
		X"1E",X"DD",X"7E",X"03",X"DD",X"86",X"0E",X"30",X"03",X"DD",X"34",X"04",X"DD",X"77",X"03",X"DD",
		X"7E",X"06",X"DD",X"86",X"0F",X"30",X"03",X"DD",X"34",X"07",X"DD",X"77",X"06",X"18",X"1C",X"DD",
		X"7E",X"03",X"DD",X"96",X"10",X"30",X"03",X"DD",X"35",X"04",X"DD",X"77",X"03",X"DD",X"7E",X"06",
		X"DD",X"86",X"11",X"30",X"03",X"DD",X"34",X"07",X"DD",X"77",X"06",X"DD",X"7E",X"09",X"DD",X"96",
		X"0C",X"DD",X"77",X"09",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"05",X"DD",
		X"77",X"08",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"DD",X"BE",X"0D",X"C0",X"CD",X"A9",X"43",X"C9",
		X"DD",X"CB",X"01",X"6E",X"20",X"0C",X"DD",X"36",X"0B",X"04",X"DD",X"36",X"0C",X"01",X"CD",X"76",
		X"44",X"C9",X"DD",X"7E",X"09",X"A7",X"20",X"0D",X"DD",X"35",X"0C",X"DD",X"7E",X"0C",X"A7",X"20",
		X"ED",X"CD",X"A9",X"43",X"C9",X"DD",X"35",X"09",X"DD",X"7E",X"05",X"A7",X"C8",X"DD",X"7E",X"0A",
		X"DD",X"96",X"0B",X"DD",X"77",X"0A",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"05",X"DD",X"77",X"08",
		X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"76",X"44",X"C9",X"DD",X"7E",X"09",X"DD",X"BE",
		X"0B",X"30",X"1E",X"DD",X"7E",X"0C",X"DD",X"86",X"03",X"30",X"03",X"DD",X"34",X"04",X"DD",X"77",
		X"03",X"DD",X"7E",X"06",X"DD",X"86",X"0D",X"30",X"03",X"DD",X"34",X"07",X"DD",X"77",X"06",X"18",
		X"1C",X"DD",X"7E",X"03",X"DD",X"96",X"0E",X"30",X"03",X"DD",X"35",X"04",X"DD",X"77",X"03",X"DD",
		X"7E",X"06",X"DD",X"96",X"0F",X"30",X"03",X"DD",X"35",X"07",X"DD",X"77",X"06",X"DD",X"7E",X"0A",
		X"DD",X"96",X"10",X"DD",X"77",X"0A",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"05",X"DD",X"77",X"08",
		X"DD",X"34",X"09",X"DD",X"7E",X"09",X"DD",X"BE",X"11",X"C0",X"CD",X"A9",X"43",X"C9",X"DD",X"CB",
		X"01",X"6E",X"20",X"44",X"DD",X"CB",X"01",X"EE",X"DD",X"E5",X"06",X"1A",X"DD",X"36",X"03",X"00",
		X"DD",X"23",X"10",X"F8",X"DD",X"E1",X"CD",X"76",X"44",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"7E",
		X"DD",X"77",X"0B",X"23",X"7E",X"DD",X"77",X"0C",X"23",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"DD",
		X"7E",X"0C",X"E6",X"0F",X"DD",X"CB",X"01",X"8E",X"DD",X"CB",X"01",X"96",X"DD",X"CB",X"01",X"9E",
		X"DD",X"CB",X"01",X"A6",X"DD",X"77",X"14",X"C9",X"DD",X"CB",X"01",X"66",X"28",X"41",X"DD",X"CB",
		X"01",X"4E",X"28",X"22",X"DD",X"7E",X"11",X"DD",X"BE",X"13",X"30",X"30",X"DD",X"7E",X"1A",X"DD",
		X"96",X"1C",X"30",X"02",X"3E",X"00",X"DD",X"77",X"1A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"DD",X"77",X"08",X"18",X"16",X"DD",X"7E",X"13",X"DD",X"BE",X"11",X"38",X"0E",X"DD",X"36",
		X"08",X"00",X"DD",X"CB",X"01",X"A6",X"DD",X"36",X"11",X"00",X"18",X"03",X"DD",X"35",X"11",X"DD",
		X"7E",X"10",X"FE",X"00",X"28",X"38",X"DD",X"CB",X"01",X"56",X"28",X"22",X"DD",X"7E",X"10",X"DD",
		X"BE",X"12",X"30",X"26",X"DD",X"7E",X"19",X"DD",X"96",X"1B",X"30",X"02",X"3E",X"00",X"DD",X"77",
		X"19",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"05",X"18",X"0C",X"DD",X"7E",
		X"12",X"DD",X"BE",X"10",X"38",X"04",X"DD",X"36",X"05",X"00",X"DD",X"35",X"10",X"C9",X"DD",X"6E",
		X"09",X"DD",X"66",X"0A",X"7E",X"DD",X"77",X"0B",X"23",X"7E",X"DD",X"77",X"0C",X"23",X"DD",X"75",
		X"09",X"DD",X"74",X"0A",X"DD",X"CB",X"0C",X"7E",X"28",X"3D",X"DD",X"7E",X"0C",X"E6",X"F0",X"FE",
		X"F0",X"20",X"04",X"CD",X"A9",X"43",X"C9",X"FE",X"90",X"20",X"13",X"DD",X"7E",X"0B",X"DD",X"77",
		X"0D",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"C9",X"FE",X"A0",
		X"C0",X"DD",X"7E",X"0D",X"FE",X"00",X"C8",X"DD",X"7E",X"0E",X"DD",X"77",X"09",X"DD",X"7E",X"0F",
		X"DD",X"77",X"0A",X"DD",X"35",X"0D",X"C9",X"DD",X"CB",X"0C",X"76",X"28",X"08",X"DD",X"CB",X"01",
		X"DE",X"DD",X"CB",X"01",X"E6",X"DD",X"7E",X"0C",X"E6",X"3F",X"CB",X"27",X"E6",X"FF",X"28",X"18",
		X"4F",X"06",X"00",X"21",X"C2",X"43",X"09",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"04",
		X"DD",X"7E",X"14",X"DD",X"77",X"05",X"18",X"04",X"DD",X"36",X"05",X"00",X"DD",X"7E",X"0B",X"E6",
		X"0F",X"21",X"D4",X"4C",X"4F",X"06",X"00",X"09",X"7E",X"DD",X"77",X"15",X"DD",X"7E",X"00",X"21",
		X"06",X"6C",X"4F",X"06",X"00",X"09",X"7E",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",
		X"DF",X"4C",X"4F",X"06",X"00",X"09",X"4E",X"DD",X"71",X"17",X"23",X"46",X"DD",X"70",X"18",X"DD",
		X"5E",X"15",X"16",X"00",X"CD",X"2A",X"44",X"DD",X"75",X"10",X"CB",X"3D",X"DD",X"75",X"12",X"DD",
		X"7E",X"0B",X"E6",X"40",X"20",X"06",X"DD",X"CB",X"01",X"D6",X"18",X"06",X"DD",X"CB",X"01",X"96",
		X"18",X"2E",X"DD",X"7E",X"05",X"6F",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"DD",X"77",
		X"19",X"26",X"00",X"DD",X"4E",X"12",X"06",X"00",X"CD",X"4B",X"44",X"CB",X"22",X"CB",X"22",X"CB",
		X"22",X"CB",X"22",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"7A",X"83",X"DD",X"77",X"1B",
		X"DD",X"CB",X"01",X"5E",X"C8",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"7E",X"DD",X"77",X"0B",X"23",
		X"7E",X"DD",X"77",X"0C",X"23",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"DD",X"7E",X"0C",X"E6",X"3F",
		X"CB",X"27",X"4F",X"06",X"00",X"21",X"C2",X"43",X"09",X"7E",X"DD",X"77",X"06",X"23",X"7E",X"DD",
		X"77",X"07",X"DD",X"7E",X"14",X"DD",X"77",X"08",X"DD",X"7E",X"0B",X"E6",X"0F",X"21",X"D4",X"4C",
		X"4F",X"06",X"00",X"09",X"7E",X"DD",X"77",X"16",X"DD",X"4E",X"17",X"DD",X"46",X"18",X"DD",X"5E",
		X"16",X"16",X"00",X"CD",X"2A",X"44",X"DD",X"75",X"11",X"CB",X"3D",X"DD",X"75",X"13",X"DD",X"7E",
		X"0B",X"E6",X"40",X"20",X"06",X"DD",X"CB",X"01",X"CE",X"18",X"06",X"DD",X"CB",X"01",X"8E",X"18",
		X"2E",X"DD",X"7E",X"08",X"6F",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"DD",X"77",X"1A",
		X"26",X"00",X"DD",X"4E",X"13",X"06",X"00",X"CD",X"4B",X"44",X"CB",X"22",X"CB",X"22",X"CB",X"22",
		X"CB",X"22",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"7A",X"83",X"DD",X"77",X"1C",X"DD",
		X"CB",X"01",X"9E",X"C9",X"04",X"06",X"08",X"0C",X"10",X"18",X"20",X"30",X"40",X"60",X"80",X"80",
		X"01",X"70",X"01",X"60",X"01",X"50",X"01",X"40",X"01",X"30",X"01",X"20",X"01",X"10",X"01",X"00",
		X"01",X"F0",X"00",X"E0",X"00",X"D0",X"00",X"C0",X"00",X"B0",X"00",X"A0",X"00",X"90",X"00",X"00",
		X"8C",X"FF",X"90",X"02",X"63",X"05",X"14",X"02",X"23",X"02",X"23",X"04",X"61",X"04",X"12",X"02",
		X"60",X"02",X"10",X"05",X"54",X"07",X"23",X"02",X"10",X"02",X"12",X"02",X"14",X"02",X"65",X"05",
		X"15",X"02",X"21",X"02",X"25",X"04",X"68",X"02",X"17",X"02",X"65",X"02",X"15",X"04",X"54",X"07",
		X"23",X"02",X"14",X"02",X"10",X"02",X"12",X"02",X"14",X"02",X"65",X"05",X"15",X"02",X"21",X"02",
		X"25",X"02",X"68",X"04",X"17",X"02",X"27",X"02",X"65",X"02",X"15",X"02",X"63",X"05",X"14",X"02",
		X"25",X"02",X"23",X"02",X"60",X"05",X"10",X"02",X"1C",X"02",X"20",X"02",X"63",X"05",X"12",X"02",
		X"23",X"02",X"23",X"04",X"65",X"04",X"10",X"02",X"67",X"02",X"0F",X"07",X"68",X"07",X"10",X"01",
		X"00",X"00",X"A0",X"00",X"8A",X"FF",X"90",X"05",X"63",X"05",X"20",X"05",X"60",X"05",X"1C",X"05",
		X"63",X"05",X"20",X"05",X"60",X"05",X"1C",X"05",X"65",X"05",X"21",X"05",X"60",X"05",X"1C",X"05",
		X"65",X"05",X"21",X"05",X"60",X"05",X"1C",X"05",X"67",X"05",X"23",X"05",X"60",X"05",X"1C",X"05",
		X"67",X"05",X"23",X"05",X"60",X"05",X"1C",X"03",X"65",X"03",X"21",X"03",X"60",X"03",X"1C",X"05",
		X"63",X"05",X"20",X"05",X"60",X"05",X"1C",X"05",X"60",X"05",X"1C",X"00",X"A0",X"00",X"8C",X"FF",
		X"90",X"04",X"63",X"06",X"14",X"02",X"23",X"02",X"25",X"04",X"63",X"06",X"14",X"04",X"21",X"04",
		X"60",X"04",X"10",X"04",X"61",X"04",X"12",X"06",X"63",X"06",X"14",X"04",X"5E",X"04",X"0F",X"04",
		X"60",X"04",X"10",X"06",X"61",X"06",X"12",X"04",X"60",X"04",X"10",X"04",X"61",X"04",X"12",X"06",
		X"63",X"06",X"14",X"04",X"63",X"06",X"14",X"02",X"23",X"02",X"25",X"04",X"63",X"06",X"14",X"04",
		X"21",X"04",X"60",X"04",X"10",X"04",X"61",X"04",X"12",X"06",X"63",X"06",X"14",X"06",X"5E",X"06",
		X"0F",X"06",X"63",X"06",X"0F",X"04",X"60",X"04",X"10",X"07",X"5C",X"07",X"10",X"00",X"A0",X"00",
		X"8C",X"FF",X"90",X"04",X"60",X"06",X"14",X"02",X"1C",X"02",X"17",X"04",X"60",X"06",X"14",X"02",
		X"1C",X"02",X"17",X"04",X"61",X"06",X"15",X"02",X"1E",X"02",X"17",X"04",X"63",X"06",X"17",X"02",
		X"20",X"02",X"17",X"04",X"63",X"06",X"17",X"02",X"20",X"02",X"17",X"04",X"61",X"06",X"15",X"02",
		X"1E",X"02",X"17",X"04",X"60",X"06",X"14",X"02",X"1C",X"02",X"17",X"04",X"5E",X"06",X"12",X"02",
		X"1B",X"02",X"17",X"04",X"5C",X"06",X"10",X"02",X"17",X"02",X"14",X"04",X"5C",X"06",X"10",X"02",
		X"17",X"02",X"14",X"04",X"5E",X"06",X"12",X"02",X"1B",X"02",X"17",X"04",X"60",X"06",X"14",X"02",
		X"1C",X"02",X"17",X"04",X"60",X"06",X"14",X"02",X"1C",X"02",X"17",X"04",X"60",X"05",X"14",X"02",
		X"1C",X"02",X"5E",X"02",X"12",X"04",X"5E",X"06",X"12",X"02",X"1B",X"02",X"17",X"04",X"5E",X"04",
		X"0B",X"02",X"5B",X"02",X"17",X"02",X"57",X"02",X"12",X"00",X"A0",X"00",X"89",X"FF",X"90",X"03",
		X"5C",X"05",X"04",X"03",X"1E",X"03",X"60",X"03",X"04",X"05",X"60",X"05",X"08",X"03",X"5E",X"03",
		X"08",X"03",X"5C",X"05",X"0B",X"03",X"00",X"03",X"5C",X"05",X"04",X"03",X"1E",X"03",X"5E",X"03",
		X"04",X"03",X"60",X"05",X"08",X"03",X"00",X"03",X"60",X"03",X"08",X"03",X"5E",X"05",X"0B",X"03",
		X"1C",X"03",X"59",X"05",X"01",X"03",X"1B",X"03",X"5C",X"03",X"01",X"05",X"5C",X"05",X"04",X"03",
		X"5B",X"03",X"04",X"03",X"59",X"05",X"08",X"03",X"00",X"03",X"59",X"05",X"01",X"03",X"1B",X"03",
		X"5B",X"03",X"01",X"03",X"5C",X"05",X"04",X"03",X"00",X"03",X"5C",X"03",X"04",X"03",X"5E",X"05",
		X"08",X"03",X"1C",X"03",X"5E",X"05",X"06",X"03",X"20",X"03",X"61",X"03",X"06",X"05",X"61",X"05",
		X"09",X"03",X"60",X"03",X"09",X"03",X"5E",X"05",X"0D",X"03",X"00",X"03",X"5E",X"05",X"06",X"03",
		X"20",X"03",X"60",X"03",X"06",X"03",X"61",X"05",X"09",X"03",X"00",X"03",X"61",X"03",X"09",X"03",
		X"60",X"05",X"0D",X"03",X"21",X"03",X"63",X"04",X"0B",X"03",X"00",X"03",X"63",X"04",X"0B",X"03",
		X"00",X"03",X"63",X"04",X"0B",X"05",X"00",X"05",X"63",X"06",X"0B",X"03",X"23",X"03",X"61",X"05",
		X"09",X"03",X"21",X"03",X"60",X"05",X"08",X"03",X"20",X"03",X"5E",X"05",X"06",X"03",X"1E",X"00",
		X"A0",X"00",X"8C",X"05",X"50",X"05",X"14",X"02",X"50",X"02",X"14",X"04",X"50",X"04",X"14",X"04",
		X"5C",X"04",X"20",X"04",X"5B",X"04",X"1E",X"04",X"59",X"04",X"1C",X"04",X"57",X"04",X"1B",X"04",
		X"55",X"04",X"19",X"05",X"54",X"05",X"17",X"02",X"55",X"02",X"19",X"04",X"54",X"04",X"17",X"04",
		X"52",X"04",X"15",X"04",X"50",X"04",X"14",X"04",X"52",X"04",X"15",X"05",X"54",X"05",X"17",X"FF",
		X"FF",X"00",X"8C",X"04",X"5C",X"04",X"0B",X"02",X"68",X"02",X"14",X"02",X"67",X"02",X"10",X"04",
		X"65",X"04",X"10",X"04",X"63",X"04",X"0F",X"04",X"61",X"04",X"0D",X"04",X"60",X"04",X"0B",X"04",
		X"5E",X"04",X"09",X"04",X"00",X"04",X"5C",X"04",X"08",X"02",X"57",X"02",X"01",X"02",X"59",X"02",
		X"03",X"02",X"5B",X"02",X"04",X"02",X"5C",X"02",X"06",X"02",X"5E",X"02",X"08",X"02",X"60",X"02",
		X"08",X"04",X"1C",X"04",X"00",X"06",X"5C",X"06",X"04",X"FF",X"FF",X"00",X"8C",X"02",X"5C",X"02",
		X"17",X"02",X"63",X"02",X"10",X"02",X"60",X"02",X"17",X"02",X"5C",X"02",X"10",X"02",X"5E",X"04",
		X"12",X"02",X"1B",X"04",X"57",X"04",X"0F",X"02",X"5E",X"04",X"17",X"02",X"21",X"02",X"65",X"04",
		X"14",X"02",X"23",X"02",X"61",X"04",X"12",X"02",X"1B",X"04",X"60",X"04",X"10",X"04",X"60",X"04",
		X"10",X"04",X"63",X"04",X"14",X"04",X"68",X"04",X"17",X"FF",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"4C",X"50",X"86",X"50",X"F2",X"50",X"48",X"51",X"0E",X"52",X"8E",X"52",X"04",X"01",X"00",X"07",
		X"01",X"01",X"00",X"00",X"02",X"05",X"00",X"02",X"1F",X"11",X"3B",X"21",X"01",X"02",X"00",X"03",
		X"0A",X"12",X"27",X"21",X"3F",X"11",X"A6",X"13",X"00",X"00",X"A8",X"14",X"00",X"01",X"03",X"51",
		X"A6",X"13",X"00",X"01",X"1F",X"40",X"A8",X"14",X"00",X"00",X"0F",X"15",X"00",X"04",X"10",X"12",
		X"2B",X"11",X"3C",X"60",X"58",X"60",X"05",X"03",X"00",X"0C",X"01",X"04",X"00",X"01",X"3D",X"30",
		X"03",X"09",X"00",X"02",X"3A",X"12",X"3D",X"31",X"03",X"0C",X"00",X"03",X"19",X"23",X"2B",X"30",
		X"3F",X"12",X"02",X"08",X"00",X"03",X"23",X"13",X"2B",X"21",X"2C",X"35",X"01",X"03",X"00",X"02",
		X"2B",X"22",X"38",X"21",X"A6",X"13",X"00",X"01",X"01",X"34",X"A6",X"13",X"00",X"00",X"85",X"09",
		X"12",X"02",X"1C",X"50",X"3C",X"41",X"85",X"0C",X"12",X"01",X"23",X"50",X"85",X"09",X"12",X"03",
		X"02",X"21",X"1B",X"52",X"3E",X"41",X"A8",X"14",X"00",X"01",X"10",X"20",X"A8",X"14",X"00",X"02",
		X"00",X"51",X"1C",X"40",X"0F",X"15",X"00",X"05",X"10",X"12",X"2B",X"11",X"3C",X"60",X"40",X"12",
		X"5A",X"60",X"06",X"03",X"00",X"05",X"04",X"0D",X"00",X"03",X"23",X"75",X"24",X"12",X"3C",X"13",
		X"04",X"0F",X"00",X"06",X"10",X"13",X"16",X"74",X"22",X"70",X"24",X"12",X"2E",X"71",X"38",X"13",
		X"04",X"0F",X"00",X"05",X"00",X"21",X"16",X"75",X"22",X"71",X"24",X"50",X"2E",X"74",X"85",X"0E",
		X"11",X"04",X"18",X"22",X"1A",X"70",X"26",X"71",X"34",X"21",X"04",X"0F",X"00",X"05",X"16",X"70",
		X"1F",X"13",X"22",X"74",X"2E",X"75",X"3C",X"13",X"0F",X"15",X"00",X"06",X"02",X"23",X"14",X"12",
		X"2C",X"12",X"3E",X"60",X"42",X"11",X"5C",X"60",X"01",X"03",X"00",X"12",X"03",X"0A",X"00",X"01",
		X"3E",X"41",X"03",X"0C",X"00",X"04",X"0A",X"13",X"1A",X"40",X"29",X"12",X"38",X"41",X"03",X"0A",
		X"00",X"04",X"0B",X"11",X"1E",X"40",X"28",X"13",X"38",X"40",X"03",X"0B",X"00",X"04",X"08",X"12",
		X"1C",X"41",X"29",X"13",X"3A",X"40",X"02",X"06",X"00",X"06",X"08",X"13",X"1C",X"23",X"22",X"21",
		X"2E",X"21",X"39",X"12",X"3F",X"23",X"03",X"0A",X"00",X"05",X"0E",X"23",X"1C",X"21",X"26",X"23",
		X"30",X"13",X"3D",X"21",X"02",X"05",X"00",X"03",X"0E",X"21",X"1F",X"23",X"30",X"23",X"A6",X"13",
		X"00",X"02",X"04",X"41",X"1E",X"51",X"A6",X"13",X"00",X"00",X"A8",X"14",X"00",X"02",X"04",X"50",
		X"1F",X"41",X"A8",X"14",X"00",X"01",X"10",X"52",X"03",X"0C",X"00",X"04",X"08",X"12",X"14",X"52",
		X"28",X"41",X"3F",X"50",X"A6",X"13",X"00",X"01",X"18",X"52",X"A6",X"13",X"00",X"01",X"18",X"52",
		X"04",X"0E",X"00",X"03",X"1A",X"74",X"26",X"71",X"3F",X"21",X"85",X"0E",X"10",X"03",X"1A",X"71",
		X"26",X"74",X"3C",X"31",X"04",X"0F",X"00",X"06",X"16",X"74",X"20",X"12",X"22",X"75",X"2E",X"70",
		X"3C",X"12",X"3F",X"31",X"04",X"0D",X"00",X"03",X"20",X"12",X"22",X"70",X"3F",X"13",X"0F",X"15",
		X"00",X"06",X"00",X"31",X"14",X"12",X"28",X"12",X"34",X"12",X"3C",X"60",X"58",X"60",X"00",X"03",
		X"00",X"0C",X"A6",X"13",X"00",X"01",X"1B",X"52",X"85",X"0C",X"11",X"02",X"1F",X"50",X"34",X"52",
		X"85",X"0B",X"12",X"04",X"00",X"21",X"20",X"51",X"2C",X"52",X"3C",X"52",X"85",X"0C",X"12",X"03",
		X"10",X"22",X"1C",X"51",X"3E",X"51",X"85",X"0A",X"11",X"03",X"0A",X"21",X"18",X"50",X"34",X"50",
		X"A8",X"14",X"00",X"02",X"06",X"50",X"12",X"52",X"85",X"06",X"10",X"03",X"1A",X"21",X"34",X"41",
		X"3A",X"40",X"85",X"0C",X"11",X"03",X"12",X"40",X"1A",X"41",X"3A",X"23",X"85",X"0C",X"10",X"03",
		X"16",X"40",X"1E",X"41",X"3E",X"20",X"85",X"07",X"12",X"03",X"06",X"20",X"1C",X"40",X"32",X"41",
		X"A8",X"14",X"00",X"03",X"06",X"21",X"12",X"41",X"18",X"40",X"A8",X"14",X"00",X"00",X"0F",X"15",
		X"00",X"06",X"0E",X"12",X"20",X"11",X"2A",X"12",X"3C",X"60",X"48",X"11",X"58",X"60",X"02",X"03",
		X"00",X"15",X"A6",X"13",X"00",X"00",X"04",X"0E",X"00",X"06",X"0E",X"31",X"1A",X"71",X"1E",X"12",
		X"26",X"70",X"32",X"13",X"36",X"31",X"85",X"0F",X"12",X"06",X"12",X"23",X"16",X"74",X"22",X"71",
		X"23",X"34",X"2E",X"70",X"3E",X"30",X"85",X"0F",X"11",X"05",X"16",X"70",X"17",X"21",X"22",X"71",
		X"2A",X"30",X"2E",X"74",X"04",X"0E",X"00",X"06",X"0E",X"31",X"1A",X"70",X"1E",X"13",X"26",X"71",
		X"36",X"22",X"3C",X"12",X"A6",X"13",X"00",X"02",X"06",X"41",X"1A",X"21",X"A6",X"13",X"00",X"02",
		X"0A",X"41",X"0B",X"34",X"A6",X"13",X"00",X"01",X"06",X"40",X"A6",X"13",X"00",X"02",X"02",X"31",
		X"08",X"41",X"85",X"0B",X"11",X"05",X"0C",X"22",X"0E",X"31",X"1E",X"40",X"26",X"41",X"3E",X"35",
		X"A6",X"13",X"00",X"03",X"06",X"41",X"0E",X"34",X"1F",X"22",X"A6",X"13",X"00",X"03",X"02",X"41",
		X"0A",X"40",X"14",X"35",X"A6",X"13",X"00",X"02",X"06",X"41",X"1C",X"35",X"A6",X"13",X"00",X"01",
		X"06",X"40",X"A8",X"14",X"00",X"02",X"12",X"21",X"18",X"31",X"85",X"0C",X"12",X"04",X"0C",X"21",
		X"20",X"22",X"2E",X"21",X"3C",X"21",X"A6",X"13",X"00",X"01",X"0A",X"41",X"A6",X"13",X"00",X"02",
		X"08",X"41",X"12",X"31",X"85",X"08",X"12",X"03",X"0C",X"20",X"28",X"22",X"32",X"31",X"85",X"0A",
		X"12",X"01",X"2E",X"31",X"03",X"16",X"00",X"02",X"22",X"12",X"36",X"12",X"0F",X"15",X"00",X"05",
		X"0A",X"12",X"26",X"12",X"3A",X"12",X"3C",X"60",X"58",X"60",X"98",X"53",X"A1",X"53",X"A6",X"53",
		X"AC",X"53",X"B1",X"53",X"B7",X"53",X"BC",X"53",X"C1",X"53",X"C6",X"53",X"CB",X"53",X"D0",X"53",
		X"D5",X"53",X"DC",X"53",X"E4",X"53",X"ED",X"53",X"F7",X"53",X"02",X"54",X"0D",X"54",X"19",X"54",
		X"24",X"54",X"32",X"54",X"40",X"54",X"66",X"54",X"08",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"04",X"03",X"03",X"03",X"03",X"05",X"03",X"02",X"03",X"03",X"02",X"04",X"04",X"03",X"04",
		X"03",X"05",X"02",X"04",X"03",X"04",X"02",X"04",X"04",X"03",X"05",X"03",X"04",X"04",X"05",X"04",
		X"05",X"04",X"05",X"03",X"06",X"04",X"04",X"06",X"05",X"06",X"05",X"04",X"05",X"03",X"07",X"04",
		X"04",X"05",X"07",X"05",X"06",X"06",X"05",X"01",X"02",X"07",X"01",X"06",X"07",X"02",X"02",X"07",
		X"01",X"02",X"07",X"01",X"08",X"03",X"0F",X"10",X"12",X"10",X"11",X"01",X"02",X"09",X"02",X"0F",
		X"10",X"12",X"10",X"12",X"10",X"11",X"02",X"0A",X"01",X"0F",X"10",X"12",X"10",X"12",X"10",X"12",
		X"10",X"11",X"0A",X"0E",X"0C",X"0B",X"0B",X"0D",X"0E",X"0D",X"0C",X"0B",X"0C",X"0B",X"0E",X"0B",
		X"0D",X"0C",X"0E",X"0C",X"0B",X"0D",X"0E",X"0B",X"0E",X"0A",X"0E",X"0C",X"0A",X"0C",X"0C",X"0E",
		X"0D",X"0B",X"0A",X"0D",X"FF",X"09",X"13",X"09",X"02",X"09",X"03",X"06",X"00",X"00",X"00",X"00",
		X"0A",X"0C",X"FF",X"0D",X"17",X"09",X"02",X"03",X"09",X"06",X"0C",X"0A",X"00",X"00",X"00",X"00",
		X"25",X"02",X"0F",X"14",X"15",X"16",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"0B",X"0F",X"14",X"15",X"16",X"16",X"16",X"16",X"14",X"15",
		X"14",X"0F",X"A0",X"54",X"A9",X"54",X"B2",X"54",X"BF",X"54",X"D4",X"54",X"E9",X"54",X"FE",X"54",
		X"13",X"55",X"28",X"55",X"39",X"55",X"4E",X"55",X"5B",X"55",X"68",X"55",X"75",X"55",X"7E",X"55",
		X"87",X"55",X"94",X"55",X"A1",X"55",X"AE",X"55",X"B7",X"55",X"C0",X"55",X"CD",X"55",X"DA",X"55",
		X"A0",X"00",X"E1",X"55",X"04",X"00",X"00",X"00",X"00",X"A4",X"00",X"F1",X"55",X"04",X"01",X"01",
		X"01",X"01",X"A8",X"00",X"01",X"56",X"08",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"B0",
		X"00",X"21",X"56",X"10",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"C0",X"00",X"61",X"56",X"10",X"01",X"01",X"01",X"02",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"02",X"01",X"01",X"01",X"D2",X"00",X"A1",X"56",X"10",X"01",X"01",
		X"01",X"02",X"11",X"12",X"21",X"21",X"21",X"21",X"12",X"11",X"02",X"01",X"01",X"01",X"E6",X"00",
		X"E1",X"56",X"10",X"01",X"01",X"02",X"12",X"21",X"22",X"31",X"31",X"31",X"31",X"22",X"21",X"12",
		X"02",X"01",X"01",X"00",X"01",X"21",X"57",X"10",X"01",X"01",X"02",X"12",X"22",X"32",X"41",X"41",
		X"32",X"32",X"32",X"31",X"22",X"12",X"02",X"01",X"1A",X"01",X"61",X"57",X"0C",X"01",X"01",X"01",
		X"02",X"11",X"12",X"22",X"32",X"42",X"52",X"62",X"71",X"40",X"01",X"C1",X"57",X"10",X"01",X"02",
		X"12",X"22",X"33",X"52",X"62",X"72",X"72",X"62",X"52",X"33",X"22",X"12",X"02",X"01",X"60",X"01",
		X"01",X"58",X"08",X"10",X"50",X"54",X"18",X"18",X"54",X"50",X"10",X"78",X"01",X"21",X"58",X"08",
		X"10",X"30",X"22",X"22",X"12",X"22",X"21",X"20",X"87",X"01",X"41",X"58",X"08",X"10",X"20",X"21",
		X"12",X"12",X"21",X"20",X"10",X"93",X"01",X"61",X"58",X"04",X"40",X"33",X"33",X"40",X"A1",X"01",
		X"71",X"58",X"04",X"20",X"31",X"31",X"20",X"AB",X"01",X"81",X"58",X"08",X"01",X"01",X"02",X"11",
		X"12",X"21",X"22",X"31",X"B6",X"01",X"A1",X"58",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"D6",X"01",X"C1",X"58",X"08",X"31",X"22",X"21",X"12",X"11",X"02",X"01",X"01",X"A0",X"00",
		X"E1",X"58",X"04",X"00",X"00",X"00",X"00",X"20",X"01",X"F1",X"58",X"04",X"02",X"02",X"02",X"02",
		X"AB",X"01",X"01",X"59",X"08",X"41",X"41",X"42",X"51",X"52",X"61",X"62",X"71",X"AB",X"01",X"21",
		X"59",X"08",X"81",X"81",X"82",X"91",X"92",X"A1",X"A2",X"B1",X"A4",X"00",X"41",X"59",X"02",X"C1",
		X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"06",X"07",
		X"07",X"07",X"07",X"06",X"06",X"05",X"05",X"04",X"04",X"03",X"03",X"02",X"02",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",X"03",X"03",
		X"03",X"03",X"04",X"04",X"04",X"04",X"05",X"05",X"05",X"05",X"06",X"06",X"06",X"06",X"07",X"07",
		X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",X"05",X"05",X"05",X"05",X"04",X"04",X"04",X"04",
		X"03",X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"06",X"07",
		X"08",X"09",X"09",X"0A",X"0B",X"0B",X"0C",X"0C",X"0C",X"0D",X"0D",X"0E",X"0E",X"0E",X"0E",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0D",X"0D",X"0D",X"0C",X"0C",X"0B",X"0B",X"0A",X"0A",
		X"09",X"08",X"08",X"07",X"06",X"05",X"04",X"03",X"03",X"02",X"02",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"03",X"03",X"04",X"05",X"06",X"07",X"08",X"09",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"15",X"16",X"16",X"16",
		X"17",X"17",X"17",X"16",X"16",X"15",X"15",X"14",X"13",X"12",X"11",X"10",X"0F",X"0E",X"0D",X"0C",
		X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"03",X"02",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"09",X"0A",X"0C",X"0D",X"0F",
		X"10",X"12",X"13",X"14",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1D",X"1E",X"1E",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1E",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"14",X"13",
		X"12",X"10",X"0F",X"0D",X"0C",X"0A",X"09",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"03",X"05",X"06",X"08",X"0A",X"0C",X"0E",X"10",X"12",
		X"14",X"16",X"18",X"1A",X"1C",X"1E",X"20",X"22",X"24",X"26",X"27",X"27",X"26",X"24",X"23",X"22",
		X"21",X"1F",X"1E",X"1C",X"1B",X"1B",X"1B",X"1C",X"1E",X"20",X"22",X"21",X"20",X"1F",X"1E",X"1C",
		X"1A",X"18",X"16",X"14",X"12",X"10",X"0E",X"0C",X"0A",X"08",X"06",X"04",X"02",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"02",X"03",X"04",X"05",X"06",X"07",X"08",
		X"09",X"0A",X"0C",X"0D",X"0E",X"0F",X"11",X"12",X"13",X"15",X"17",X"18",X"19",X"1B",X"1C",X"1E",
		X"1F",X"21",X"23",X"25",X"27",X"29",X"2B",X"2E",X"31",X"32",X"35",X"38",X"3C",X"40",X"40",X"40",
		X"40",X"3F",X"3F",X"3F",X"3F",X"3E",X"3A",X"37",X"34",X"31",X"2F",X"2C",X"2A",X"28",X"26",X"24",
		X"22",X"20",X"1F",X"1D",X"1C",X"1A",X"19",X"17",X"16",X"14",X"13",X"11",X"10",X"0F",X"0D",X"0C",
		X"0B",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"03",X"02",X"02",X"02",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"01",X"02",X"03",X"05",X"06",X"08",X"0A",X"0C",X"0E",X"10",X"14",X"16",X"19",
		X"1C",X"1E",X"21",X"24",X"27",X"2A",X"2D",X"30",X"32",X"35",X"38",X"3B",X"3E",X"40",X"42",X"43",
		X"43",X"43",X"43",X"43",X"41",X"3F",X"3C",X"39",X"36",X"34",X"31",X"2E",X"2B",X"28",X"25",X"23",
		X"20",X"1D",X"1A",X"18",X"15",X"12",X"0F",X"0D",X"0B",X"09",X"07",X"05",X"03",X"02",X"01",X"01",
		X"00",X"01",X"01",X"02",X"04",X"08",X"10",X"1A",X"22",X"2B",X"33",X"3A",X"40",X"43",X"45",X"46",
		X"48",X"48",X"47",X"46",X"44",X"41",X"3B",X"33",X"2B",X"24",X"1D",X"15",X"0C",X"06",X"03",X"02",
		X"01",X"01",X"02",X"04",X"07",X"0A",X"0E",X"11",X"14",X"17",X"1A",X"1E",X"20",X"20",X"1D",X"1A",
		X"17",X"14",X"12",X"12",X"15",X"17",X"19",X"1A",X"19",X"17",X"13",X"10",X"0C",X"09",X"05",X"02",
		X"01",X"01",X"01",X"03",X"05",X"07",X"09",X"0B",X"0D",X"0F",X"11",X"13",X"13",X"12",X"11",X"12",
		X"13",X"15",X"17",X"18",X"18",X"16",X"14",X"12",X"0F",X"0D",X"0B",X"09",X"06",X"04",X"03",X"02",
		X"01",X"01",X"04",X"0B",X"17",X"22",X"2A",X"2E",X"30",X"30",X"2F",X"2C",X"26",X"1E",X"11",X"07",
		X"02",X"01",X"02",X"04",X"08",X"11",X"1A",X"1E",X"20",X"20",X"1F",X"1C",X"16",X"0D",X"05",X"02",
		X"01",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",
		X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",
		X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",
		X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",
		X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",
		X"3F",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",
		X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",
		X"5F",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"0E",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"F5",X"C5",X"D5",X"E5",X"4F",X"E6",X"F0",X"FE",X"50",X"30",X"13",X"0F",X"0F",X"0F",X"5F",X"16",
		X"00",X"21",X"73",X"59",X"19",X"5E",X"23",X"56",X"EB",X"11",X"6E",X"59",X"D5",X"E9",X"E1",X"D1",
		X"C1",X"F1",X"C9",X"7D",X"59",X"8B",X"59",X"D6",X"59",X"E9",X"59",X"4D",X"5A",X"21",X"00",X"6F",
		X"36",X"00",X"11",X"01",X"6F",X"01",X"7D",X"00",X"ED",X"B0",X"C9",X"21",X"0C",X"6F",X"11",X"E4",
		X"5A",X"CD",X"B7",X"5A",X"3A",X"06",X"6F",X"FE",X"38",X"30",X"24",X"E6",X"FC",X"0F",X"5F",X"16",
		X"00",X"21",X"85",X"5A",X"19",X"CD",X"58",X"5A",X"21",X"07",X"6F",X"7E",X"2B",X"FE",X"02",X"28",
		X"0B",X"47",X"7E",X"E6",X"03",X"20",X"03",X"78",X"A7",X"C0",X"34",X"C9",X"36",X"00",X"C9",X"CD",
		X"93",X"5B",X"3A",X"06",X"6F",X"FE",X"38",X"20",X"05",X"CD",X"AF",X"5A",X"20",X"F4",X"CD",X"59",
		X"5D",X"AF",X"32",X"06",X"6F",X"C9",X"11",X"E4",X"5A",X"CB",X"41",X"20",X"05",X"21",X"58",X"6F",
		X"18",X"03",X"21",X"5D",X"6F",X"CD",X"B7",X"5A",X"C9",X"CB",X"41",X"28",X"2E",X"21",X"0C",X"6F",
		X"11",X"5D",X"6F",X"CD",X"B7",X"5A",X"21",X"11",X"6F",X"11",X"5D",X"6F",X"CD",X"B7",X"5A",X"21",
		X"13",X"6F",X"11",X"E4",X"5A",X"CD",X"D4",X"5A",X"21",X"5B",X"6F",X"CD",X"E5",X"5A",X"21",X"03",
		X"6F",X"CD",X"FA",X"5A",X"21",X"59",X"6F",X"CD",X"8B",X"5B",X"C9",X"21",X"0C",X"6F",X"11",X"58",
		X"6F",X"CD",X"B7",X"5A",X"21",X"11",X"6F",X"11",X"58",X"6F",X"CD",X"B7",X"5A",X"21",X"13",X"6F",
		X"11",X"E4",X"5A",X"CD",X"D4",X"5A",X"21",X"56",X"6F",X"CD",X"E5",X"5A",X"21",X"00",X"6F",X"CD",
		X"FA",X"5A",X"21",X"54",X"6F",X"CD",X"8B",X"5B",X"AF",X"32",X"06",X"6F",X"C9",X"3A",X"06",X"6F",
		X"FE",X"38",X"C0",X"3C",X"32",X"06",X"6F",X"C9",X"AF",X"32",X"07",X"6F",X"5E",X"23",X"56",X"EB",
		X"5E",X"23",X"56",X"7A",X"B3",X"C8",X"23",X"1A",X"A6",X"23",X"BE",X"20",X"04",X"23",X"23",X"18",
		X"EF",X"47",X"3E",X"01",X"32",X"07",X"6F",X"78",X"23",X"BE",X"20",X"03",X"23",X"18",X"E1",X"3E",
		X"02",X"32",X"07",X"6F",X"C9",X"A1",X"5A",X"A8",X"5A",X"A1",X"5A",X"A8",X"5A",X"A1",X"5A",X"A8",
		X"5A",X"A1",X"5A",X"A8",X"5A",X"A1",X"5A",X"A8",X"5A",X"A1",X"5A",X"A8",X"5A",X"A1",X"5A",X"A8",
		X"5A",X"00",X"90",X"7F",X"1B",X"1F",X"00",X"00",X"00",X"90",X"7F",X"1F",X"1B",X"00",X"00",X"3A",
		X"00",X"90",X"E6",X"1F",X"FE",X"1E",X"C9",X"06",X"03",X"37",X"3F",X"1A",X"8E",X"27",X"38",X"08",
		X"FE",X"60",X"38",X"06",X"D6",X"60",X"18",X"02",X"C6",X"40",X"77",X"1B",X"2B",X"10",X"EB",X"3F",
		X"CD",X"D5",X"5A",X"C9",X"AF",X"06",X"02",X"1A",X"8E",X"27",X"77",X"1B",X"2B",X"10",X"F8",X"C9",
		X"00",X"00",X"00",X"00",X"01",X"11",X"0F",X"5B",X"CD",X"69",X"5B",X"CB",X"21",X"06",X"00",X"21",
		X"15",X"6F",X"09",X"11",X"E4",X"5A",X"CD",X"D4",X"5A",X"C9",X"11",X"3C",X"5B",X"CD",X"69",X"5B",
		X"CB",X"21",X"06",X"00",X"21",X"35",X"6F",X"09",X"11",X"E4",X"5A",X"CD",X"D4",X"5A",X"C9",X"01",
		X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"06",X"00",
		X"00",X"07",X"00",X"00",X"08",X"00",X"00",X"09",X"00",X"00",X"10",X"00",X"00",X"12",X"00",X"00",
		X"14",X"00",X"00",X"16",X"00",X"00",X"18",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"50",X"00",X"01",X"00",X"00",X"01",X"30",X"00",X"01",X"60",X"00",X"02",X"00",X"00",X"02",X"50",
		X"00",X"03",X"00",X"00",X"03",X"50",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"06",X"00",X"00",
		X"08",X"00",X"00",X"10",X"00",X"00",X"15",X"00",X"00",X"01",X"00",X"0F",X"C5",X"D5",X"E5",X"06",
		X"03",X"1A",X"BE",X"20",X"06",X"13",X"23",X"10",X"F8",X"18",X"0C",X"30",X"0A",X"E1",X"D1",X"13",
		X"13",X"13",X"C1",X"0C",X"10",X"E6",X"C9",X"E1",X"D1",X"C1",X"C9",X"AF",X"06",X"05",X"77",X"23",
		X"10",X"FC",X"C9",X"21",X"00",X"D0",X"11",X"5E",X"6F",X"01",X"04",X"08",X"C5",X"E5",X"7E",X"12",
		X"36",X"00",X"13",X"23",X"10",X"F8",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",X"20",X"ED",X"21",
		X"80",X"D0",X"36",X"24",X"11",X"81",X"D0",X"01",X"FF",X"02",X"ED",X"B0",X"21",X"80",X"D4",X"01",
		X"00",X"03",X"36",X"00",X"23",X"0B",X"78",X"B1",X"20",X"F8",X"0E",X"40",X"11",X"20",X"00",X"21",
		X"00",X"70",X"06",X"20",X"36",X"00",X"19",X"10",X"FB",X"0D",X"20",X"F3",X"21",X"71",X"5C",X"0E",
		X"25",X"CD",X"15",X"5C",X"0D",X"20",X"FA",X"11",X"AF",X"D0",X"21",X"08",X"6F",X"CD",X"22",X"5C",
		X"11",X"EF",X"D0",X"21",X"0D",X"6F",X"CD",X"22",X"5C",X"11",X"2F",X"D1",X"21",X"12",X"6F",X"CD",
		X"40",X"5C",X"11",X"6A",X"D1",X"21",X"14",X"6F",X"CD",X"2E",X"5C",X"11",X"78",X"D1",X"21",X"34",
		X"6F",X"CD",X"2E",X"5C",X"C9",X"5E",X"23",X"56",X"23",X"46",X"23",X"7E",X"12",X"13",X"23",X"10",
		X"FA",X"C9",X"CD",X"40",X"5C",X"13",X"CD",X"44",X"5C",X"13",X"CD",X"44",X"5C",X"C9",X"06",X"10",
		X"C5",X"D5",X"CD",X"40",X"5C",X"D1",X"EB",X"01",X"20",X"00",X"09",X"EB",X"C1",X"10",X"F1",X"C9",
		X"06",X"04",X"18",X"02",X"06",X"02",X"AF",X"ED",X"6F",X"28",X"13",X"CB",X"FF",X"F5",X"D5",X"E5",
		X"E6",X"0F",X"5F",X"16",X"00",X"21",X"4F",X"5D",X"19",X"7E",X"E1",X"D1",X"12",X"F1",X"13",X"CB",
		X"40",X"28",X"05",X"ED",X"6F",X"23",X"18",X"06",X"CB",X"48",X"28",X"02",X"CB",X"FF",X"10",X"D7",
		X"C9",X"A6",X"D0",X"05",X"1D",X"18",X"1D",X"0A",X"15",X"B3",X"D0",X"07",X"11",X"24",X"24",X"16",
		X"24",X"24",X"1C",X"E6",X"D0",X"07",X"12",X"17",X"24",X"19",X"15",X"0A",X"22",X"F3",X"D0",X"07",
		X"11",X"24",X"24",X"16",X"24",X"24",X"1C",X"26",X"D1",X"05",X"1D",X"12",X"16",X"0E",X"1C",X"65",
		X"D1",X"04",X"01",X"16",X"12",X"17",X"72",X"D1",X"05",X"02",X"14",X"19",X"1D",X"1C",X"85",X"D1",
		X"01",X"02",X"92",X"D1",X"02",X"05",X"14",X"A5",X"D1",X"01",X"03",X"B1",X"D1",X"03",X"01",X"00",
		X"14",X"C5",X"D1",X"01",X"04",X"D1",X"D1",X"03",X"01",X"03",X"14",X"E5",X"D1",X"01",X"05",X"F1",
		X"D1",X"03",X"01",X"06",X"14",X"05",X"D2",X"01",X"06",X"11",X"D2",X"03",X"02",X"00",X"14",X"25",
		X"D2",X"01",X"07",X"31",X"D2",X"03",X"02",X"05",X"14",X"45",X"D2",X"01",X"08",X"51",X"D2",X"03",
		X"03",X"00",X"14",X"65",X"D2",X"01",X"09",X"71",X"D2",X"03",X"03",X"05",X"14",X"84",X"D2",X"02",
		X"01",X"00",X"91",X"D2",X"03",X"04",X"00",X"14",X"A4",X"D2",X"02",X"01",X"02",X"B1",X"D2",X"03",
		X"05",X"00",X"14",X"C4",X"D2",X"02",X"01",X"04",X"D1",X"D2",X"03",X"06",X"00",X"14",X"E4",X"D2",
		X"02",X"01",X"06",X"F1",X"D2",X"03",X"08",X"00",X"14",X"04",X"D3",X"02",X"01",X"08",X"10",X"D3",
		X"04",X"01",X"00",X"00",X"14",X"24",X"D3",X"02",X"02",X"00",X"30",X"D3",X"04",X"01",X"05",X"00",
		X"14",X"44",X"D3",X"04",X"18",X"1F",X"0E",X"1B",X"50",X"D3",X"04",X"18",X"1F",X"0E",X"1B",X"00",
		X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"21",X"80",X"D0",X"36",X"24",X"11",X"81",
		X"D0",X"01",X"FF",X"02",X"ED",X"B0",X"21",X"5E",X"6F",X"11",X"00",X"D0",X"01",X"08",X"04",X"C5",
		X"06",X"00",X"ED",X"B0",X"EB",X"01",X"18",X"00",X"09",X"EB",X"C1",X"10",X"F2",X"C9",X"C7",X"C7",
		X"21",X"00",X"B0",X"36",X"9F",X"36",X"BF",X"36",X"DF",X"36",X"FF",X"21",X"00",X"C0",X"36",X"9F",
		X"36",X"BF",X"36",X"DF",X"36",X"FF",X"21",X"80",X"D0",X"36",X"24",X"23",X"7C",X"FE",X"E0",X"38",
		X"F8",X"21",X"00",X"D0",X"36",X"00",X"11",X"01",X"D0",X"01",X"7F",X"00",X"ED",X"B0",X"0E",X"40",
		X"11",X"20",X"00",X"21",X"00",X"70",X"06",X"20",X"36",X"00",X"19",X"10",X"FB",X"0D",X"20",X"F3",
		X"DD",X"21",X"ED",X"D1",X"DD",X"36",X"00",X"1B",X"DD",X"36",X"01",X"18",X"DD",X"36",X"02",X"16",
		X"21",X"00",X"00",X"11",X"00",X"00",X"AF",X"06",X"10",X"86",X"2C",X"20",X"FC",X"24",X"10",X"F9",
		X"BB",X"28",X"10",X"16",X"FF",X"7B",X"C6",X"01",X"DD",X"77",X"04",X"01",X"00",X"00",X"0B",X"78",
		X"B1",X"20",X"FB",X"1C",X"7B",X"FE",X"06",X"38",X"DD",X"CB",X"7A",X"C2",X"00",X"00",X"DD",X"36",
		X"04",X"18",X"DD",X"36",X"05",X"14",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"DD",X"36",
		X"00",X"1B",X"DD",X"36",X"01",X"0A",X"DD",X"36",X"02",X"16",X"DD",X"36",X"04",X"24",X"DD",X"36",
		X"05",X"24",X"1E",X"FF",X"21",X"00",X"60",X"16",X"10",X"7B",X"0E",X"10",X"06",X"10",X"C6",X"2F",
		X"77",X"23",X"10",X"FA",X"3D",X"0D",X"20",X"F4",X"3D",X"15",X"20",X"EE",X"21",X"00",X"60",X"16",
		X"10",X"7B",X"0E",X"10",X"06",X"10",X"C6",X"2F",X"BE",X"20",X"23",X"23",X"10",X"F8",X"3D",X"0D",
		X"20",X"F2",X"3D",X"15",X"20",X"EC",X"7B",X"D6",X"0F",X"5F",X"30",X"C8",X"DD",X"36",X"04",X"18",
		X"DD",X"36",X"05",X"14",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"18",X"15",X"7C",X"E6",
		X"0C",X"0F",X"0F",X"C6",X"01",X"DD",X"77",X"04",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",
		X"C3",X"00",X"00",X"DD",X"36",X"00",X"1C",X"DD",X"36",X"01",X"18",X"DD",X"36",X"02",X"1E",X"DD",
		X"36",X"03",X"17",X"DD",X"36",X"04",X"0D",X"DD",X"36",X"05",X"24",X"CD",X"E0",X"5E",X"3E",X"03",
		X"21",X"81",X"D0",X"11",X"81",X"D4",X"06",X"1D",X"36",X"4D",X"12",X"13",X"23",X"10",X"F9",X"36",
		X"4F",X"12",X"21",X"A1",X"D0",X"11",X"A1",X"D4",X"01",X"17",X"1D",X"C5",X"36",X"4C",X"12",X"23",
		X"13",X"10",X"F9",X"36",X"4E",X"12",X"23",X"23",X"23",X"13",X"13",X"13",X"C1",X"0D",X"20",X"EB",
		X"18",X"FE",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"DD",X"21",X"00",X"6C",X"16",X"02",X"21",X"00",X"B0",X"18",X"03",X"21",X"00",X"C0",X"06",X"04",
		X"3E",X"9F",X"77",X"C6",X"20",X"10",X"FB",X"15",X"28",X"02",X"18",X"EF",X"21",X"00",X"B0",X"0E",
		X"00",X"11",X"EC",X"5F",X"06",X"03",X"1A",X"77",X"13",X"1A",X"13",X"DD",X"77",X"00",X"DD",X"36",
		X"01",X"00",X"CD",X"A0",X"5F",X"28",X"05",X"CD",X"CD",X"5F",X"18",X"F6",X"1A",X"77",X"13",X"10",
		X"E5",X"CD",X"C6",X"5F",X"06",X"02",X"36",X"E3",X"36",X"F0",X"DD",X"36",X"00",X"C0",X"DD",X"36",
		X"01",X"00",X"CD",X"A0",X"5F",X"28",X"05",X"CD",X"CD",X"5F",X"18",X"F6",X"36",X"E7",X"10",X"EA",
		X"36",X"FF",X"CD",X"C6",X"5F",X"11",X"F5",X"5F",X"06",X"06",X"36",X"F0",X"1A",X"13",X"77",X"CD",
		X"C6",X"5F",X"10",X"F8",X"36",X"FF",X"CD",X"C6",X"5F",X"11",X"EC",X"5F",X"06",X"03",X"1A",X"77",
		X"DD",X"77",X"00",X"13",X"1A",X"77",X"13",X"36",X"0F",X"CD",X"94",X"5F",X"28",X"05",X"CD",X"BF",
		X"5F",X"18",X"F6",X"13",X"10",X"E8",X"CD",X"C6",X"5F",X"36",X"E4",X"DD",X"36",X"00",X"F0",X"CD",
		X"94",X"5F",X"28",X"05",X"CD",X"BF",X"5F",X"18",X"F6",X"79",X"FE",X"00",X"C0",X"0C",X"21",X"00",
		X"C0",X"C3",X"01",X"5F",X"DD",X"34",X"00",X"DD",X"7E",X"00",X"77",X"E6",X"0F",X"FE",X"0F",X"C9",
		X"DD",X"34",X"00",X"DD",X"7E",X"00",X"E6",X"0F",X"FE",X"0F",X"20",X"0B",X"DD",X"34",X"01",X"DD",
		X"7E",X"00",X"D6",X"0F",X"DD",X"77",X"00",X"DD",X"7E",X"01",X"E6",X"3F",X"FE",X"3F",X"C9",X"D9",
		X"08",X"11",X"89",X"1D",X"18",X"14",X"D9",X"08",X"11",X"24",X"76",X"18",X"0D",X"DD",X"7E",X"00",
		X"77",X"DD",X"7E",X"01",X"77",X"D9",X"08",X"11",X"7B",X"00",X"DD",X"CB",X"00",X"46",X"1B",X"7A",
		X"FE",X"00",X"20",X"F6",X"7B",X"FE",X"00",X"20",X"F1",X"D9",X"08",X"C9",X"90",X"80",X"9F",X"B0",
		X"A0",X"BF",X"D0",X"C0",X"DF",X"E0",X"E1",X"E2",X"E4",X"E5",X"E6",X"C7",X"C7",X"C7",X"C7",X"C7");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
