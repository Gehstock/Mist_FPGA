library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bagman_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bagman_tile_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"E6",X"E4",X"00",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"00",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"42",X"A5",X"A5",X"A5",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"0C",X"1A",X"18",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"04",X"04",X"00",X"09",X"08",X"18",X"3A",X"48",X"90",X"90",X"00",X"C0",X"00",X"00",X"48",
		X"3A",X"18",X"08",X"09",X"00",X"04",X"04",X"02",X"48",X"00",X"00",X"C0",X"00",X"90",X"90",X"48",
		X"08",X"08",X"04",X"00",X"09",X"08",X"18",X"3A",X"20",X"40",X"98",X"04",X"C0",X"00",X"00",X"48",
		X"3A",X"18",X"08",X"09",X"00",X"04",X"08",X"08",X"48",X"00",X"00",X"C0",X"04",X"98",X"40",X"20",
		X"00",X"00",X"01",X"03",X"0F",X"60",X"81",X"08",X"00",X"00",X"80",X"C0",X"F0",X"06",X"81",X"10",
		X"68",X"89",X"00",X"60",X"81",X"00",X"00",X"00",X"16",X"91",X"00",X"06",X"81",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"CF",X"20",X"01",X"08",X"00",X"00",X"80",X"C0",X"F3",X"04",X"80",X"10",
		X"28",X"49",X"80",X"20",X"21",X"10",X"00",X"00",X"14",X"92",X"01",X"04",X"84",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"19",X"05",X"0C",X"1C",X"00",X"00",X"00",X"C0",X"1C",X"20",X"00",X"A0",
		X"1E",X"1C",X"0C",X"05",X"19",X"00",X"00",X"00",X"00",X"A0",X"00",X"20",X"1C",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"05",X"0C",X"0C",X"00",X"00",X"00",X"98",X"20",X"20",X"00",X"A0",
		X"1E",X"1C",X"0C",X"05",X"09",X"08",X"00",X"00",X"00",X"A0",X"00",X"20",X"20",X"98",X"00",X"00",
		X"00",X"00",X"00",X"13",X"17",X"0F",X"01",X"18",X"00",X"00",X"00",X"90",X"D0",X"E0",X"00",X"30",
		X"22",X"20",X"0A",X"10",X"10",X"10",X"00",X"00",X"88",X"08",X"A0",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"03",X"37",X"0F",X"01",X"18",X"00",X"00",X"00",X"80",X"D8",X"E0",X"00",X"30",
		X"22",X"00",X"0A",X"20",X"20",X"00",X"00",X"00",X"88",X"00",X"A0",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"E4",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"01",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"C8",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"03",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"04",X"08",X"04",X"05",X"03",X"E7",X"27",X"00",X"88",X"48",X"24",X"7C",X"7E",X"7F",X"3F",
		X"3F",X"27",X"E7",X"03",X"05",X"04",X"08",X"04",X"80",X"3F",X"7E",X"7C",X"7C",X"24",X"48",X"88",
		X"00",X"00",X"00",X"08",X"15",X"03",X"E7",X"27",X"00",X"10",X"23",X"24",X"7C",X"7E",X"7F",X"3F",
		X"3F",X"27",X"E7",X"03",X"15",X"08",X"00",X"00",X"80",X"3F",X"7F",X"7E",X"7C",X"24",X"23",X"10",
		X"04",X"04",X"07",X"01",X"41",X"B7",X"0F",X"1F",X"40",X"40",X"C0",X"00",X"04",X"DA",X"E0",X"F0",
		X"81",X"5C",X"3E",X"1E",X"DE",X"3E",X"0E",X"06",X"02",X"74",X"F8",X"F0",X"F6",X"F8",X"E0",X"C0",
		X"04",X"04",X"07",X"11",X"21",X"17",X"0F",X"1F",X"40",X"40",X"C0",X"10",X"08",X"D0",X"E0",X"F0",
		X"01",X"1C",X"7E",X"9E",X"1E",X"3E",X"4E",X"46",X"00",X"70",X"FC",X"F2",X"F0",X"F8",X"E4",X"C4",
		X"00",X"00",X"03",X"01",X"01",X"38",X"CC",X"07",X"00",X"40",X"44",X"24",X"12",X"FC",X"FF",X"FF",
		X"01",X"07",X"CC",X"38",X"01",X"01",X"03",X"00",X"FF",X"FF",X"FF",X"FC",X"12",X"24",X"44",X"40",
		X"00",X"00",X"06",X"02",X"01",X"00",X"7C",X"87",X"00",X"04",X"0D",X"11",X"12",X"FC",X"FF",X"FF",
		X"01",X"87",X"7C",X"00",X"01",X"02",X"06",X"00",X"FF",X"FF",X"FF",X"FC",X"12",X"11",X"0D",X"04",
		X"04",X"04",X"08",X"08",X"0C",X"06",X"42",X"73",X"40",X"40",X"20",X"20",X"60",X"C0",X"84",X"9C",
		X"0F",X"CF",X"2F",X"1F",X"0F",X"6F",X"17",X"07",X"E0",X"E6",X"E8",X"F0",X"E0",X"EC",X"D0",X"C0",
		X"02",X"04",X"04",X"04",X"04",X"46",X"62",X"13",X"80",X"40",X"40",X"40",X"40",X"C4",X"8C",X"90",
		X"0F",X"0F",X"0F",X"3F",X"4F",X"CF",X"17",X"67",X"E0",X"E0",X"E0",X"F8",X"E4",X"E6",X"D0",X"CC",
		X"00",X"00",X"00",X"02",X"03",X"18",X"24",X"32",X"00",X"00",X"00",X"00",X"80",X"E4",X"F8",X"B0",
		X"2B",X"15",X"25",X"19",X"0A",X"0E",X"00",X"00",X"3C",X"70",X"78",X"64",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"1A",X"00",X"00",X"00",X"00",X"00",X"C8",X"04",X"00",
		X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"05",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"6E",X"77",X"3B",X"DF",X"EF",X"7F",X"9F",X"B0",X"76",X"6E",X"FC",X"FB",X"F7",X"FE",X"FD",
		X"BF",X"7F",X"EF",X"DF",X"3B",X"76",X"6E",X"0D",X"F9",X"FE",X"F7",X"FB",X"DC",X"EE",X"76",X"B0",
		X"00",X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"00",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"03",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",X"10",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"03",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",X"10",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"03",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",X"10",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1F",X"03",X"21",X"35",X"11",X"00",X"F0",X"E0",X"80",X"00",X"80",X"C0",X"80",
		X"1D",X"11",X"35",X"21",X"03",X"1F",X"0F",X"03",X"90",X"80",X"C0",X"80",X"00",X"80",X"E0",X"F0",
		X"00",X"FF",X"0F",X"07",X"03",X"21",X"35",X"11",X"00",X"00",X"C0",X"C0",X"00",X"80",X"C0",X"80",
		X"1D",X"11",X"35",X"21",X"03",X"07",X"0F",X"FF",X"90",X"80",X"C0",X"80",X"00",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"07",X"07",X"01",X"1B",X"1C",X"00",X"1E",X"F0",X"C0",X"80",X"80",X"E0",X"30",
		X"1E",X"1C",X"1B",X"01",X"07",X"07",X"00",X"00",X"18",X"30",X"E0",X"80",X"80",X"C0",X"F0",X"1E",
		X"00",X"07",X"3F",X"0F",X"07",X"01",X"1B",X"1C",X"00",X"F8",X"E0",X"C0",X"80",X"80",X"E0",X"30",
		X"1E",X"1C",X"1B",X"01",X"07",X"0F",X"3F",X"07",X"18",X"30",X"E0",X"80",X"80",X"C0",X"E0",X"F8",
		X"00",X"0F",X"10",X"10",X"0F",X"00",X"0F",X"10",X"00",X"F8",X"04",X"04",X"F8",X"00",X"F8",X"04",
		X"10",X"0F",X"00",X"0F",X"10",X"10",X"10",X"0C",X"04",X"F8",X"00",X"04",X"84",X"44",X"24",X"1C",
		X"00",X"0F",X"10",X"10",X"0F",X"00",X"0F",X"10",X"00",X"F8",X"04",X"04",X"F8",X"00",X"F8",X"04",
		X"10",X"0F",X"00",X"00",X"08",X"06",X"01",X"00",X"04",X"F8",X"00",X"10",X"FC",X"10",X"90",X"70",
		X"00",X"0F",X"10",X"10",X"0F",X"00",X"0F",X"10",X"00",X"F8",X"04",X"04",X"F8",X"00",X"F8",X"04",
		X"10",X"0F",X"00",X"0F",X"10",X"10",X"10",X"0F",X"04",X"F8",X"00",X"78",X"84",X"84",X"84",X"78",
		X"1F",X"10",X"1F",X"00",X"1F",X"10",X"1F",X"00",X"FC",X"04",X"FC",X"00",X"FC",X"04",X"FC",X"00",
		X"0C",X"11",X"11",X"0F",X"00",X"00",X"1F",X"10",X"F8",X"04",X"04",X"F8",X"00",X"04",X"FC",X"04",
		X"1F",X"10",X"1F",X"00",X"1F",X"10",X"1F",X"00",X"FC",X"04",X"FC",X"00",X"FC",X"04",X"FC",X"00",
		X"1F",X"10",X"1C",X"00",X"1F",X"10",X"10",X"1C",X"04",X"C4",X"3C",X"00",X"7C",X"84",X"84",X"1C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"22",
		X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"02",X"10",X"02",X"12",X"12",X"12",
		X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"10",X"02",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"08",X"40",X"48",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"08",X"40",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",
		X"00",X"00",X"00",X"05",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"F4",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"04",X"04",X"00",X"01",X"C0",X"00",X"10",X"00",X"08",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",
		X"00",X"02",X"00",X"04",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"04",X"00",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"13",X"3F",X"3F",X"00",X"00",X"00",X"00",X"22",X"77",X"DD",X"DD",
		X"3F",X"3F",X"13",X"03",X"00",X"00",X"00",X"00",X"DD",X"DD",X"77",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"09",X"1F",X"1F",X"00",X"00",X"02",X"17",X"BD",X"ED",X"ED",X"ED",
		X"1F",X"19",X"09",X"07",X"00",X"00",X"00",X"00",X"EF",X"FA",X"90",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"77",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"DD",X"DD",X"77",X"22",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"E8",X"BC",X"B6",X"B7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B7",X"F6",X"5C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"03",X"03",X"0F",X"0F",X"00",X"00",X"C0",X"E0",X"C0",X"C0",X"F0",X"F0",
		X"03",X"07",X"0C",X"07",X"03",X"07",X"0C",X"07",X"C0",X"E0",X"30",X"E0",X"C0",X"E0",X"30",X"E0",
		X"00",X"00",X"00",X"03",X"07",X"09",X"09",X"0F",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"C0",X"F0",
		X"0F",X"03",X"03",X"06",X"03",X"01",X"03",X"01",X"F0",X"E0",X"F0",X"18",X"F0",X"F8",X"0C",X"F8",
		X"03",X"07",X"0C",X"07",X"03",X"07",X"0C",X"07",X"C0",X"E0",X"30",X"E0",X"C0",X"E0",X"30",X"E0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"06",X"03",X"07",X"0C",X"07",X"03",X"01",X"F0",X"18",X"F0",X"E0",X"30",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"0A",X"EA",X"20",X"02",X"3E",X"C8",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"C8",X"3E",X"02",X"20",X"EA",
		X"A8",X"A8",X"00",X"F0",X"4C",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"4C",X"F0",X"00",X"A8",X"00",X"00",X"FE",X"FE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0A",X"EA",X"27",X"06",X"3E",X"EA",X"1A",X"FE",
		X"1F",X"31",X"75",X"00",X"00",X"00",X"00",X"00",X"26",X"64",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"64",
		X"1F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"26",X"FE",X"1A",X"EA",X"3E",X"06",X"27",X"EA",
		X"A8",X"A8",X"80",X"F0",X"FE",X"DF",X"FC",X"7A",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",
		X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"9E",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"9E",
		X"10",X"7A",X"FC",X"DF",X"FE",X"F0",X"80",X"A8",X"F0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0A",X"EA",X"27",X"06",X"3E",X"FE",X"FE",X"FE",
		X"0F",X"1F",X"3F",X"7D",X"44",X"54",X"47",X"7C",X"FE",X"FE",X"FE",X"8E",X"AC",X"88",X"F8",X"00",
		X"00",X"7C",X"47",X"54",X"44",X"7D",X"3F",X"1F",X"00",X"00",X"F8",X"88",X"AC",X"8E",X"FE",X"FE",
		X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"3E",X"06",X"27",X"EA",
		X"A8",X"A8",X"80",X"F8",X"FE",X"FF",X"F8",X"FA",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",
		X"E0",X"6B",X"23",X"3E",X"1C",X"00",X"00",X"00",X"C0",X"E0",X"30",X"1E",X"0A",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"23",X"6B",X"00",X"00",X"00",X"0E",X"0A",X"1E",X"30",X"E0",
		X"E0",X"FA",X"F8",X"FF",X"FE",X"F8",X"80",X"A8",X"C0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"50",X"48",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"67",X"37",X"37",X"10",X"17",X"1C",X"07",
		X"00",X"04",X"04",X"04",X"04",X"14",X"24",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"CC",X"D8",X"D8",X"10",X"D0",X"70",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1B",X"08",X"2B",X"30",X"71",X"30",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"20",X"20",X"60",X"60",X"60",X"00",
		X"60",X"B0",X"20",X"A8",X"18",X"1C",X"18",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"07",X"07",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"90",X"C8",X"C4",
		X"07",X"05",X"07",X"07",X"01",X"03",X"01",X"00",X"E3",X"E7",X"F7",X"F7",X"F0",X"FF",X"FC",X"07",
		X"00",X"00",X"00",X"01",X"01",X"13",X"27",X"47",X"00",X"40",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",
		X"8F",X"CF",X"DF",X"DF",X"1F",X"FF",X"7F",X"C0",X"C0",X"40",X"C0",X"C0",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"03",X"7C",X"DB",X"A8",X"DB",X"F0",X"F1",X"70",X"E0",
		X"03",X"01",X"01",X"03",X"06",X"06",X"06",X"00",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"B6",X"2A",X"B7",X"1F",X"1E",X"1D",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"00",
		X"00",X"F8",X"FC",X"DE",X"FF",X"FF",X"7F",X"77",X"00",X"00",X"00",X"00",X"00",X"90",X"C8",X"C4",
		X"7F",X"7F",X"6F",X"7F",X"7F",X"1F",X"0F",X"00",X"E3",X"E7",X"F7",X"F7",X"F0",X"FF",X"FC",X"07",
		X"00",X"00",X"00",X"00",X"01",X"13",X"27",X"47",X"00",X"3E",X"7E",X"F6",X"FE",X"FE",X"FC",X"DC",
		X"8F",X"CF",X"DF",X"DF",X"1F",X"FF",X"7F",X"C0",X"FC",X"FC",X"EC",X"FC",X"FC",X"F0",X"E0",X"00",
		X"01",X"03",X"0F",X"1F",X"1D",X"1F",X"0F",X"07",X"FC",X"3B",X"E8",X"DB",X"F8",X"F1",X"70",X"E0",
		X"03",X"03",X"06",X"0C",X"38",X"38",X"38",X"00",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"B9",X"2F",X"B7",X"3F",X"1F",X"1D",X"0F",X"00",X"80",X"E0",X"F0",X"70",X"F0",X"E0",X"C0",
		X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"60",X"38",X"38",X"38",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"02",X"03",X"00",X"00",X"00",X"3F",X"3F",X"21",X"21",X"E3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"01",X"01",X"01",X"01",X"00",X"00",X"1B",X"F2",X"FD",X"11",X"11",X"FD",X"01",X"0D",X"CD",X"41",
		X"03",X"03",X"02",X"02",X"03",X"00",X"03",X"00",X"03",X"01",X"01",X"3F",X"FF",X"00",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"05",
		X"FD",X"FF",X"FC",X"FC",X"FC",X"CC",X"84",X"84",X"C0",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",
		X"12",X"1E",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"41",X"CD",X"DD",X"3D",X"FD",X"FD",X"FF",X"FD",
		X"00",X"03",X"00",X"03",X"03",X"00",X"00",X"03",X"00",X"FF",X"C0",X"00",X"FF",X"3F",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"19",X"11",X"31",X"21",X"21",X"40",X"40",
		X"CC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"FD",X"3D",X"1D",X"4D",X"61",X"7F",X"FF",
		X"02",X"82",X"82",X"43",X"40",X"40",X"23",X"22",X"3F",X"03",X"03",X"FF",X"00",X"3F",X"E0",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"4F",X"47",X"47",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"01",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F0",X"F0",X"C0",
		X"22",X"23",X"20",X"23",X"22",X"23",X"22",X"23",X"3F",X"FF",X"00",X"00",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"23",X"21",X"30",X"10",X"18",X"08",X"0C",
		X"FF",X"FF",X"FF",X"7C",X"7C",X"7C",X"7C",X"3C",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"7F",X"7F",
		X"FF",X"FC",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"0D",X"1D",X"3D",X"FD",X"FD",
		X"20",X"23",X"43",X"42",X"42",X"C3",X"80",X"02",X"00",X"03",X"01",X"01",X"3F",X"FF",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"24",X"24",X"DC",X"FC",X"3C",X"3C",X"1F",X"05",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"0E",X"FD",X"FF",X"FD",X"FD",X"3D",X"7D",X"8D",X"00",
		X"02",X"02",X"02",X"03",X"00",X"00",X"00",X"00",X"21",X"21",X"3F",X"FF",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"02",X"02",X"02",X"02",X"03",X"FF",X"3F",X"00",X"21",X"21",X"21",X"3F",X"FF",
		X"00",X"3F",X"48",X"48",X"48",X"48",X"48",X"3F",X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",
		X"00",X"7F",X"04",X"08",X"10",X"20",X"40",X"7F",X"00",X"41",X"49",X"49",X"49",X"49",X"49",X"7F",
		X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"31",X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",
		X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",
		X"3F",X"40",X"40",X"41",X"42",X"42",X"42",X"42",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"F8",X"04",X"02",X"82",X"82",X"42",X"42",X"42",
		X"42",X"42",X"42",X"41",X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",X"80",X"43",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"01",X"FE",X"00",X"00",X"42",X"82",X"82",X"82",X"02",X"04",X"04",X"08",
		X"08",X"06",X"01",X"00",X"00",X"38",X"44",X"43",X"00",X"00",X"C0",X"3F",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"03",X"FC",X"00",X"00",X"00",X"FF",X"30",X"40",X"80",X"00",X"00",X"1C",X"22",X"C2",
		X"40",X"40",X"40",X"40",X"40",X"27",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"C2",X"22",X"1C",X"00",
		X"00",X"00",X"1F",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"C0",X"38",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"FC",X"00",X"00",X"01",X"00",X"00",X"FC",X"02",X"02",X"02",X"02",X"F2",
		X"20",X"27",X"18",X"00",X"00",X"01",X"31",X"4E",X"00",X"F0",X"20",X"40",X"80",X"00",X"01",X"02",
		X"06",X"18",X"10",X"20",X"40",X"80",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",
		X"40",X"40",X"40",X"40",X"40",X"33",X"0C",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"F2",X"02",X"02",X"02",X"02",X"F2",X"0C",X"00",
		X"00",X"00",X"01",X"0E",X"10",X"20",X"40",X"41",X"00",X"00",X"FC",X"03",X"00",X"00",X"00",X"FE",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"F2",X"02",X"02",X"02",X"02",
		X"42",X"44",X"44",X"44",X"44",X"44",X"48",X"48",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"07",X"88",X"88",X"88",X"88",X"88",X"04",X"03",X"FA",X"06",X"00",X"00",X"00",X"00",X"06",X"FA",
		X"48",X"47",X"40",X"40",X"20",X"10",X"0F",X"00",X"3C",X"C0",X"00",X"00",X"1F",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"82",X"62",X"1C",X"00",
		X"00",X"00",X"0E",X"11",X"21",X"41",X"41",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"7F",X"00",X"00",X"00",X"00",X"7F",X"80",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"E3",X"1C",X"22",X"C2",X"02",X"02",X"02",X"02",X"C2",X"22",
		X"41",X"41",X"41",X"41",X"21",X"12",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"06",X"08",X"10",X"20",X"20",X"00",X"00",X"FC",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0C",X"06",X"02",X"02",X"02",
		X"41",X"42",X"44",X"44",X"44",X"44",X"44",X"42",X"FC",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"22",X"12",X"12",X"12",X"12",X"12",X"22",
		X"41",X"20",X"20",X"10",X"08",X"04",X"03",X"00",X"03",X"FC",X"00",X"00",X"00",X"07",X"F8",X"00",
		X"FC",X"03",X"00",X"00",X"00",X"FF",X"00",X"00",X"62",X"82",X"02",X"02",X"02",X"84",X"78",X"00",
		X"00",X"00",X"00",X"03",X"04",X"08",X"08",X"10",X"00",X"00",X"FC",X"02",X"01",X"01",X"01",X"00",
		X"00",X"00",X"03",X"1C",X"20",X"40",X"80",X"07",X"00",X"00",X"80",X"78",X"04",X"02",X"02",X"82",
		X"10",X"21",X"22",X"22",X"22",X"42",X"44",X"44",X"E0",X"10",X"0C",X"04",X"02",X"02",X"02",X"04",
		X"08",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"62",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"44",X"43",X"40",X"40",X"20",X"10",X"0F",X"00",X"18",X"E0",X"00",X"00",X"01",X"3E",X"C0",X"00",
		X"18",X"07",X"00",X"00",X"FC",X"03",X"00",X"00",X"22",X"C2",X"02",X"02",X"02",X"E2",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"08",X"08",X"08",X"04",X"04",
		X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"01",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"02",X"01",X"00",X"F1",X"F2",X"05",X"92",X"8C",X"44",X"42",X"C2",X"31",X"08",
		X"04",X"08",X"10",X"20",X"20",X"43",X"4C",X"30",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"3F",
		X"F0",X"E0",X"00",X"01",X"06",X"18",X"00",X"00",X"07",X"19",X"60",X"82",X"02",X"05",X"14",X"28",
		X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"40",X"7F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"11",X"10",X"10",X"01",X"03",X"03",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"10",X"20",X"20",X"40",X"5F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"9F",X"9F",X"00",X"00",X"00",X"00",X"80",X"40",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"05",X"12",X"0C",X"04",X"02",X"02",X"F9",X"F8",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F9",X"20",X"02",X"02",X"05",X"14",X"28",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"83",X"8F",X"47",X"42",X"C2",X"31",X"08",X"C0",X"C0",X"C0",X"E0",X"20",X"43",X"4C",X"30",
		X"07",X"19",X"60",X"82",X"03",X"07",X"03",X"03",X"80",X"80",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"07",X"07",X"0F",X"0F",X"3F",X"FF",X"FC",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FF",X"3F",X"0F",X"0F",X"07",X"03",X"03",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"F0",X"FC",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"7F",X"7F",X"FC",X"F8",X"E0",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"07",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"07",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"07",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"07",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"07",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"FF",X"FF",
		X"FF",X"FF",X"07",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"01",X"C1",X"28",X"C8",X"2C",X"00",X"40",X"90",X"24",X"48",X"98",X"23",X"FF",
		X"3E",X"3E",X"2C",X"C8",X"28",X"C0",X"00",X"00",X"7F",X"7F",X"FC",X"00",X"88",X"00",X"00",X"00",
		X"00",X"60",X"00",X"20",X"38",X"20",X"0C",X"80",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"06",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",X"00",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"FF",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"06",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"00",
		X"00",X"00",X"02",X"FF",X"00",X"00",X"02",X"01",X"80",X"80",X"00",X"FF",X"80",X"80",X"40",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"70",X"F8",X"7C",X"3E",X"7C",X"F8",X"70",
		X"00",X"40",X"9C",X"9E",X"5F",X"1E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
