`define BUILD_DATE "190715"
`define BUILD_TIME "162500"
