-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity OMEGA_ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of OMEGA_ROM_PGM_0 is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"AF",x"32",x"01",x"70",x"C3",x"69",x"00",x"FF", -- 0x0000
    x"77",x"3C",x"23",x"77",x"3C",x"19",x"C9",x"FF", -- 0x0008
    x"77",x"23",x"10",x"FC",x"C9",x"FF",x"FF",x"FF", -- 0x0010
    x"77",x"23",x"10",x"FC",x"0D",x"20",x"F9",x"C9", -- 0x0018
    x"85",x"6F",x"3E",x"00",x"8C",x"67",x"7E",x"C9", -- 0x0020
    x"87",x"E1",x"5F",x"16",x"00",x"19",x"5E",x"23", -- 0x0028
    x"56",x"EB",x"E9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
    x"E5",x"26",x"40",x"3A",x"A0",x"40",x"6F",x"CB", -- 0x0038
    x"7E",x"28",x"0E",x"72",x"2C",x"73",x"2C",x"7D", -- 0x0040
    x"FE",x"C0",x"30",x"02",x"3E",x"C0",x"32",x"A0", -- 0x0048
    x"40",x"E1",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"94", -- 0x0060
    x"08",x"21",x"00",x"40",x"11",x"01",x"40",x"01", -- 0x0068
    x"00",x"04",x"36",x"00",x"ED",x"B0",x"31",x"00", -- 0x0070
    x"44",x"21",x"C0",x"40",x"06",x"40",x"3E",x"FF", -- 0x0078
    x"D7",x"32",x"00",x"78",x"3A",x"00",x"78",x"AF", -- 0x0080
    x"32",x"01",x"70",x"32",x"00",x"68",x"32",x"01", -- 0x0088
    x"68",x"32",x"02",x"68",x"32",x"04",x"60",x"32", -- 0x0090
    x"05",x"60",x"32",x"06",x"60",x"32",x"07",x"60", -- 0x0098
    x"3E",x"01",x"32",x"06",x"70",x"32",x"07",x"70", -- 0x00A0
    x"21",x"C0",x"C0",x"22",x"A0",x"40",x"32",x"04", -- 0x00A8
    x"70",x"21",x"00",x"50",x"22",x"0B",x"40",x"3E", -- 0x00B0
    x"20",x"32",x"08",x"40",x"3A",x"00",x"70",x"47", -- 0x00B8
    x"E6",x"01",x"3E",x"10",x"28",x"02",x"3E",x"20", -- 0x00C0
    x"32",x"17",x"40",x"78",x"0F",x"0F",x"E6",x"01", -- 0x00C8
    x"3E",x"05",x"20",x"02",x"3E",x"03",x"32",x"07", -- 0x00D0
    x"40",x"78",x"0F",x"0F",x"0F",x"E6",x"01",x"32", -- 0x00D8
    x"0F",x"40",x"3A",x"00",x"68",x"07",x"07",x"E6", -- 0x00E0
    x"03",x"32",x"00",x"40",x"21",x"00",x"00",x"2B", -- 0x00E8
    x"3A",x"00",x"78",x"7D",x"B4",x"21",x"00",x"58", -- 0x00F0
    x"01",x"00",x"01",x"16",x"00",x"72",x"23",x"0B", -- 0x00F8
    x"78",x"B1",x"20",x"F9",x"16",x"5D",x"21",x"00", -- 0x0100
    x"50",x"01",x"00",x"04",x"72",x"3A",x"00",x"78", -- 0x0108
    x"23",x"0B",x"78",x"B1",x"20",x"F6",x"3E",x"01", -- 0x0110
    x"32",x"01",x"70",x"26",x"40",x"3A",x"A1",x"40", -- 0x0118
    x"6F",x"7E",x"87",x"30",x"05",x"CD",x"5E",x"01", -- 0x0120
    x"18",x"F1",x"E6",x"0F",x"4F",x"06",x"00",x"36", -- 0x0128
    x"FF",x"23",x"5E",x"36",x"FF",x"2C",x"7D",x"FE", -- 0x0130
    x"C0",x"30",x"02",x"3E",x"C0",x"32",x"A1",x"40", -- 0x0138
    x"7B",x"21",x"4E",x"01",x"09",x"5E",x"23",x"56", -- 0x0140
    x"21",x"1B",x"01",x"E5",x"EB",x"E9",x"F0",x"02", -- 0x0148
    x"24",x"03",x"35",x"03",x"AD",x"03",x"4E",x"04", -- 0x0150
    x"6A",x"04",x"B1",x"04",x"BC",x"07",x"3A",x"5F", -- 0x0158
    x"42",x"47",x"E6",x"0F",x"CA",x"82",x"01",x"21", -- 0x0160
    x"81",x"42",x"CB",x"46",x"C0",x"E6",x"03",x"CA", -- 0x0168
    x"A6",x"02",x"FE",x"01",x"28",x"53",x"FE",x"02", -- 0x0170
    x"28",x"76",x"3A",x"00",x"41",x"A7",x"C8",x"C3", -- 0x0178
    x"F0",x"02",x"11",x"E0",x"FF",x"21",x"E0",x"50", -- 0x0180
    x"3A",x"0E",x"40",x"A7",x"28",x"22",x"36",x"02", -- 0x0188
    x"CD",x"BA",x"01",x"21",x"40",x"53",x"CD",x"B8", -- 0x0190
    x"01",x"3A",x"0D",x"40",x"A7",x"21",x"40",x"53", -- 0x0198
    x"28",x"03",x"21",x"E0",x"50",x"CB",x"60",x"C8", -- 0x01A0
    x"3A",x"06",x"40",x"0F",x"D0",x"C3",x"C1",x"01", -- 0x01A8
    x"21",x"E0",x"50",x"CD",x"C1",x"01",x"18",x"DB", -- 0x01B0
    x"36",x"01",x"19",x"36",x"25",x"19",x"36",x"20", -- 0x01B8
    x"C9",x"3E",x"10",x"77",x"19",x"77",x"19",x"77", -- 0x01C0
    x"C9",x"21",x"7D",x"53",x"11",x"4F",x"41",x"06", -- 0x01C8
    x"02",x"CD",x"3E",x"02",x"01",x"E2",x"FF",x"09", -- 0x01D0
    x"7B",x"FE",x"3F",x"28",x"09",x"FE",x"2F",x"28", -- 0x01D8
    x"0A",x"FE",x"1F",x"20",x"EA",x"C9",x"21",x"3D", -- 0x01E0
    x"52",x"18",x"E4",x"21",x"FD",x"50",x"18",x"DF", -- 0x01E8
    x"21",x"68",x"50",x"11",x"50",x"41",x"06",x"03", -- 0x01F0
    x"CD",x"17",x"02",x"01",x"1D",x"00",x"09",x"7B", -- 0x01F8
    x"FE",x"80",x"28",x"09",x"FE",x"B0",x"28",x"0A", -- 0x0200
    x"FE",x"E0",x"C8",x"18",x"E9",x"21",x"88",x"51", -- 0x0208
    x"18",x"E4",x"21",x"A8",x"52",x"18",x"DF",x"1A", -- 0x0210
    x"F5",x"13",x"1A",x"4F",x"F1",x"CB",x"4F",x"28", -- 0x0218
    x"10",x"79",x"CB",x"4F",x"28",x"07",x"36",x"C8", -- 0x0220
    x"23",x"13",x"10",x"EB",x"C9",x"36",x"C9",x"18", -- 0x0228
    x"F7",x"79",x"CB",x"4F",x"28",x"04",x"36",x"CA", -- 0x0230
    x"18",x"EE",x"36",x"10",x"18",x"EA",x"E5",x"D5", -- 0x0238
    x"1A",x"CB",x"4F",x"28",x"25",x"CB",x"57",x"20", -- 0x0240
    x"28",x"CB",x"5F",x"20",x"2B",x"1D",x"1A",x"CB", -- 0x0248
    x"4F",x"28",x"30",x"CB",x"57",x"20",x"30",x"CB", -- 0x0250
    x"5F",x"20",x"36",x"36",x"C8",x"2D",x"1D",x"10", -- 0x0258
    x"DF",x"D1",x"E1",x"2D",x"2D",x"7B",x"D6",x"04", -- 0x0260
    x"5F",x"C9",x"36",x"10",x"2D",x"36",x"10",x"18", -- 0x0268
    x"F0",x"CD",x"9E",x"02",x"36",x"5E",x"18",x"F4", -- 0x0270
    x"D6",x"10",x"12",x"E6",x"70",x"20",x"F5",x"1A", -- 0x0278
    x"CB",x"9F",x"12",x"36",x"CA",x"18",x"E5",x"CD", -- 0x0280
    x"9E",x"02",x"36",x"C8",x"2D",x"36",x"5F",x"18", -- 0x0288
    x"D0",x"D6",x"10",x"12",x"E6",x"70",x"20",x"F2", -- 0x0290
    x"1A",x"CB",x"9F",x"12",x"18",x"CE",x"CB",x"97", -- 0x0298
    x"CB",x"DF",x"F6",x"70",x"12",x"C9",x"3A",x"BA", -- 0x02A0
    x"40",x"0F",x"D0",x"78",x"E6",x"08",x"21",x"D8", -- 0x02A8
    x"02",x"28",x"03",x"21",x"E4",x"02",x"06",x"06", -- 0x02B0
    x"11",x"20",x"00",x"DD",x"21",x"AC",x"51",x"7E", -- 0x02B8
    x"DD",x"77",x"00",x"23",x"DD",x"19",x"10",x"F7", -- 0x02C0
    x"06",x"06",x"DD",x"21",x"AD",x"51",x"7E",x"DD", -- 0x02C8
    x"77",x"00",x"23",x"DD",x"19",x"10",x"F7",x"C9", -- 0x02D0
    x"10",x"10",x"10",x"10",x"10",x"10",x"30",x"31", -- 0x02D8
    x"32",x"33",x"34",x"35",x"10",x"10",x"10",x"10", -- 0x02E0
    x"10",x"10",x"4F",x"4E",x"36",x"37",x"4D",x"4C", -- 0x02E8
    x"21",x"A5",x"51",x"11",x"1F",x"00",x"06",x"06", -- 0x02F0
    x"DD",x"21",x"04",x"41",x"3A",x"5F",x"42",x"E6", -- 0x02F8
    x"10",x"28",x"15",x"FD",x"21",x"0A",x"41",x"DD", -- 0x0300
    x"7E",x"00",x"77",x"23",x"FD",x"7E",x"00",x"77", -- 0x0308
    x"19",x"DD",x"23",x"FD",x"23",x"10",x"F0",x"C9", -- 0x0310
    x"FD",x"21",x"1E",x"03",x"18",x"E9",x"4F",x"4E", -- 0x0318
    x"32",x"33",x"4D",x"4C",x"21",x"A5",x"51",x"11", -- 0x0320
    x"1F",x"00",x"06",x"06",x"3E",x"10",x"77",x"23", -- 0x0328
    x"77",x"19",x"10",x"FA",x"C9",x"FE",x"06",x"30", -- 0x0330
    x"4A",x"A7",x"28",x"39",x"3D",x"28",x"22",x"3D", -- 0x0338
    x"87",x"87",x"87",x"87",x"2F",x"E6",x"30",x"C6", -- 0x0340
    x"C0",x"21",x"D8",x"51",x"CD",x"9A",x"03",x"21", -- 0x0348
    x"DA",x"51",x"CD",x"9A",x"03",x"21",x"18",x"52", -- 0x0350
    x"CD",x"9A",x"03",x"21",x"1A",x"52",x"C3",x"9A", -- 0x0358
    x"03",x"21",x"D8",x"51",x"11",x"1C",x"00",x"0E", -- 0x0360
    x"04",x"06",x"04",x"36",x"10",x"23",x"10",x"FB", -- 0x0368
    x"19",x"0D",x"20",x"F5",x"C9",x"CD",x"61",x"03", -- 0x0370
    x"3E",x"58",x"32",x"0D",x"42",x"21",x"F9",x"51", -- 0x0378
    x"C3",x"9A",x"03",x"FE",x"06",x"47",x"3E",x"58", -- 0x0380
    x"28",x"09",x"78",x"FE",x"07",x"3E",x"60",x"28", -- 0x0388
    x"02",x"3E",x"54",x"21",x"F9",x"51",x"18",x"02", -- 0x0390
    x"3E",x"10",x"D5",x"11",x"1F",x"00",x"CF",x"CF", -- 0x0398
    x"D1",x"C9",x"3E",x"10",x"D5",x"11",x"DF",x"FF", -- 0x03A0
    x"CF",x"C6",x"FC",x"18",x"F2",x"A7",x"28",x"48", -- 0x03A8
    x"4F",x"CD",x"03",x"04",x"87",x"81",x"4F",x"06", -- 0x03B0
    x"00",x"21",x"12",x"04",x"09",x"A7",x"06",x"03", -- 0x03B8
    x"1A",x"8E",x"27",x"12",x"13",x"23",x"10",x"F8", -- 0x03C0
    x"D5",x"3A",x"0D",x"40",x"0F",x"30",x"02",x"3E", -- 0x03C8
    x"01",x"CD",x"6A",x"04",x"D1",x"1B",x"21",x"AA", -- 0x03D0
    x"40",x"06",x"03",x"1A",x"BE",x"D8",x"20",x"05", -- 0x03D8
    x"1B",x"2B",x"10",x"F7",x"C9",x"CD",x"03",x"04", -- 0x03E0
    x"21",x"A8",x"40",x"06",x"03",x"1A",x"77",x"13", -- 0x03E8
    x"23",x"10",x"FA",x"3E",x"02",x"C3",x"6A",x"04", -- 0x03F0
    x"CD",x"03",x"04",x"21",x"AB",x"40",x"A7",x"06", -- 0x03F8
    x"03",x"18",x"BD",x"F5",x"3A",x"0D",x"40",x"11", -- 0x0400
    x"A2",x"40",x"0F",x"30",x"03",x"11",x"A5",x"40", -- 0x0408
    x"F1",x"C9",x"00",x"00",x"00",x"20",x"00",x"00", -- 0x0410
    x"40",x"00",x"00",x"60",x"00",x"00",x"80",x"00", -- 0x0418
    x"00",x"00",x"01",x"00",x"20",x"01",x"00",x"40", -- 0x0420
    x"01",x"00",x"60",x"01",x"00",x"00",x"02",x"00", -- 0x0428
    x"00",x"02",x"00",x"00",x"02",x"00",x"00",x"02", -- 0x0430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0440
    x"00",x"04",x"00",x"00",x"04",x"00",x"F5",x"21", -- 0x0448
    x"A2",x"40",x"A7",x"28",x"09",x"21",x"A5",x"40", -- 0x0450
    x"3D",x"28",x"03",x"21",x"A8",x"40",x"36",x"00", -- 0x0458
    x"23",x"36",x"00",x"23",x"36",x"00",x"F1",x"C3", -- 0x0460
    x"6A",x"04",x"21",x"A4",x"40",x"DD",x"21",x"81", -- 0x0468
    x"53",x"A7",x"28",x"11",x"21",x"A7",x"40",x"DD", -- 0x0470
    x"21",x"21",x"51",x"3D",x"28",x"07",x"21",x"AA", -- 0x0478
    x"40",x"DD",x"21",x"41",x"52",x"11",x"E0",x"FF", -- 0x0480
    x"06",x"03",x"0E",x"04",x"7E",x"0F",x"0F",x"0F", -- 0x0488
    x"0F",x"CD",x"9C",x"04",x"7E",x"CD",x"9C",x"04", -- 0x0490
    x"2B",x"10",x"F1",x"C9",x"E6",x"0F",x"28",x"08", -- 0x0498
    x"0E",x"00",x"DD",x"77",x"00",x"DD",x"19",x"C9", -- 0x04A0
    x"79",x"A7",x"28",x"F6",x"3E",x"10",x"0D",x"18", -- 0x04A8
    x"F1",x"87",x"F5",x"21",x"1E",x"05",x"E6",x"7F", -- 0x04B0
    x"5F",x"16",x"00",x"19",x"5E",x"23",x"56",x"EB", -- 0x04B8
    x"5E",x"23",x"56",x"23",x"EB",x"01",x"E0",x"FF", -- 0x04C0
    x"F1",x"38",x"0E",x"FA",x"E3",x"04",x"1A",x"FE", -- 0x04C8
    x"3F",x"C8",x"D6",x"30",x"77",x"13",x"09",x"18", -- 0x04D0
    x"F5",x"1A",x"FE",x"3F",x"C8",x"36",x"10",x"13", -- 0x04D8
    x"09",x"18",x"F6",x"22",x"B5",x"40",x"ED",x"53", -- 0x04E0
    x"B3",x"40",x"EB",x"7B",x"E6",x"1F",x"47",x"87", -- 0x04E8
    x"C6",x"20",x"6F",x"26",x"40",x"22",x"B1",x"40", -- 0x04F0
    x"CB",x"3B",x"CB",x"3B",x"7A",x"E6",x"03",x"0F", -- 0x04F8
    x"0F",x"B3",x"E6",x"F8",x"4F",x"21",x"00",x"50", -- 0x0500
    x"78",x"85",x"6F",x"11",x"20",x"00",x"43",x"36", -- 0x0508
    x"10",x"19",x"10",x"FB",x"2A",x"B1",x"40",x"71", -- 0x0510
    x"3E",x"01",x"32",x"B0",x"40",x"C9",x"6E",x"05", -- 0x0518
    x"7B",x"05",x"8F",x"05",x"9C",x"05",x"A9",x"05", -- 0x0520
    x"B6",x"05",x"D4",x"05",x"E4",x"05",x"ED",x"05", -- 0x0528
    x"FB",x"05",x"07",x"06",x"0F",x"06",x"16",x"06", -- 0x0530
    x"24",x"06",x"3E",x"06",x"4E",x"06",x"5E",x"06", -- 0x0538
    x"6E",x"06",x"7F",x"06",x"82",x"06",x"85",x"06", -- 0x0540
    x"88",x"06",x"8B",x"06",x"9C",x"06",x"A6",x"06", -- 0x0548
    x"B8",x"06",x"CD",x"06",x"E7",x"06",x"FA",x"06", -- 0x0550
    x"0D",x"07",x"20",x"07",x"33",x"07",x"46",x"07", -- 0x0558
    x"54",x"07",x"62",x"07",x"70",x"07",x"7E",x"07", -- 0x0560
    x"8C",x"07",x"9B",x"07",x"B5",x"07",x"96",x"52", -- 0x0568
    x"47",x"41",x"4D",x"45",x"40",x"40",x"4F",x"56", -- 0x0570
    x"45",x"52",x"3F",x"F1",x"52",x"50",x"55",x"53", -- 0x0578
    x"48",x"40",x"53",x"54",x"41",x"52",x"54",x"40", -- 0x0580
    x"42",x"55",x"54",x"54",x"4F",x"4E",x"3F",x"94", -- 0x0588
    x"52",x"50",x"4C",x"41",x"59",x"45",x"52",x"40", -- 0x0590
    x"4F",x"4E",x"45",x"3F",x"94",x"52",x"50",x"4C", -- 0x0598
    x"41",x"59",x"45",x"52",x"40",x"54",x"57",x"4F", -- 0x05A0
    x"3F",x"80",x"52",x"48",x"49",x"47",x"48",x"40", -- 0x05A8
    x"53",x"43",x"4F",x"52",x"45",x"3F",x"9F",x"53", -- 0x05B0
    x"40",x"43",x"52",x"45",x"44",x"49",x"54",x"40", -- 0x05B8
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x05C0
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x05C8
    x"40",x"40",x"40",x"3F",x"D1",x"52",x"49",x"4E", -- 0x05D0
    x"53",x"45",x"52",x"54",x"40",x"40",x"43",x"4F", -- 0x05D8
    x"49",x"4E",x"53",x"3F",x"1E",x"51",x"40",x"40", -- 0x05E0
    x"40",x"40",x"40",x"40",x"3F",x"5F",x"52",x"43", -- 0x05E8
    x"48",x"41",x"4E",x"43",x"45",x"40",x"54",x"49", -- 0x05F0
    x"4D",x"45",x"3F",x"94",x"52",x"46",x"49",x"52", -- 0x05F8
    x"45",x"40",x"40",x"55",x"46",x"4F",x"3F",x"4D", -- 0x0600
    x"52",x"40",x"40",x"40",x"40",x"40",x"3F",x"26", -- 0x0608
    x"52",x"50",x"4C",x"41",x"59",x"3F",x"89",x"52", -- 0x0610
    x"5B",x"40",x"40",x"4F",x"4D",x"45",x"47",x"41", -- 0x0618
    x"40",x"40",x"5B",x"3F",x"4F",x"53",x"5B",x"40", -- 0x0620
    x"53",x"43",x"4F",x"52",x"45",x"40",x"41",x"44", -- 0x0628
    x"56",x"41",x"4E",x"43",x"45",x"40",x"54",x"41", -- 0x0630
    x"42",x"4C",x"45",x"40",x"5B",x"3F",x"92",x"52", -- 0x0638
    x"34",x"30",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0640
    x"40",x"40",x"40",x"38",x"30",x"3F",x"95",x"52", -- 0x0648
    x"38",x"30",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0650
    x"40",x"40",x"31",x"36",x"30",x"3F",x"98",x"52", -- 0x0658
    x"32",x"30",x"30",x"40",x"40",x"40",x"40",x"40", -- 0x0660
    x"40",x"40",x"34",x"30",x"30",x"3F",x"BC",x"52", -- 0x0668
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0670
    x"40",x"40",x"40",x"40",x"40",x"40",x"3F",x"D5", -- 0x0678
    x"52",x"3F",x"D5",x"52",x"3F",x"D5",x"52",x"3F", -- 0x0680
    x"D5",x"52",x"3F",x"78",x"53",x"42",x"4F",x"4E", -- 0x0688
    x"55",x"53",x"40",x"42",x"45",x"45",x"54",x"4C", -- 0x0690
    x"45",x"40",x"40",x"3F",x"58",x"51",x"30",x"30", -- 0x0698
    x"30",x"40",x"50",x"54",x"53",x"3F",x"D4",x"52", -- 0x06A0
    x"4F",x"4E",x"45",x"40",x"50",x"4C",x"41",x"59", -- 0x06A8
    x"45",x"52",x"40",x"4F",x"4E",x"4C",x"59",x"3F", -- 0x06B0
    x"F4",x"52",x"4F",x"4E",x"45",x"40",x"4F",x"52", -- 0x06B8
    x"40",x"54",x"57",x"4F",x"40",x"50",x"4C",x"41", -- 0x06C0
    x"59",x"45",x"52",x"53",x"3F",x"4D",x"53",x"5B", -- 0x06C8
    x"40",x"53",x"43",x"4F",x"52",x"45",x"40",x"52", -- 0x06D0
    x"41",x"4E",x"4B",x"49",x"4E",x"47",x"40",x"54", -- 0x06D8
    x"41",x"42",x"4C",x"45",x"40",x"5B",x"3F",x"F0", -- 0x06E0
    x"52",x"31",x"53",x"54",x"40",x"40",x"40",x"40", -- 0x06E8
    x"40",x"40",x"40",x"40",x"40",x"40",x"50",x"54", -- 0x06F0
    x"53",x"3F",x"F2",x"52",x"32",x"4E",x"44",x"40", -- 0x06F8
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0700
    x"40",x"50",x"54",x"53",x"3F",x"F4",x"52",x"33", -- 0x0708
    x"52",x"44",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0710
    x"40",x"40",x"40",x"40",x"50",x"54",x"53",x"3F", -- 0x0718
    x"F6",x"52",x"34",x"54",x"48",x"40",x"40",x"40", -- 0x0720
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"50", -- 0x0728
    x"54",x"53",x"3F",x"F8",x"52",x"35",x"54",x"48", -- 0x0730
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0738
    x"40",x"40",x"50",x"54",x"53",x"3F",x"8F",x"52", -- 0x0740
    x"31",x"53",x"54",x"40",x"40",x"41",x"54",x"54", -- 0x0748
    x"41",x"43",x"4B",x"3F",x"8F",x"52",x"32",x"4E", -- 0x0750
    x"44",x"40",x"40",x"41",x"54",x"54",x"41",x"43", -- 0x0758
    x"4B",x"3F",x"8F",x"52",x"33",x"52",x"44",x"40", -- 0x0760
    x"40",x"41",x"54",x"54",x"41",x"43",x"4B",x"3F", -- 0x0768
    x"8F",x"52",x"34",x"54",x"48",x"40",x"40",x"41", -- 0x0770
    x"54",x"54",x"41",x"43",x"4B",x"3F",x"8F",x"52", -- 0x0778
    x"4E",x"45",x"58",x"54",x"40",x"41",x"54",x"54", -- 0x0780
    x"41",x"43",x"4B",x"3F",x"AF",x"52",x"4C",x"41", -- 0x0788
    x"53",x"54",x"40",x"41",x"54",x"54",x"41",x"43", -- 0x0790
    x"4B",x"40",x"3F",x"4F",x"53",x"43",x"48",x"41", -- 0x0798
    x"4C",x"4C",x"45",x"4E",x"47",x"45",x"40",x"4E", -- 0x07A0
    x"45",x"58",x"54",x"40",x"50",x"41",x"54",x"54", -- 0x07A8
    x"45",x"52",x"4E",x"40",x"3F",x"2D",x"52",x"47", -- 0x07B0
    x"4F",x"4F",x"44",x"3F",x"A7",x"CA",x"CB",x"07", -- 0x07B8
    x"3D",x"CA",x"EE",x"07",x"3D",x"CA",x"49",x"08", -- 0x07C0
    x"C3",x"2C",x"08",x"21",x"9F",x"53",x"11",x"E0", -- 0x07C8
    x"FF",x"3A",x"10",x"41",x"FE",x"15",x"38",x"02", -- 0x07D0
    x"3E",x"14",x"47",x"A7",x"28",x"06",x"36",x"CE", -- 0x07D8
    x"19",x"3D",x"20",x"F7",x"3E",x"15",x"90",x"47", -- 0x07E0
    x"36",x"10",x"19",x"10",x"FB",x"C9",x"3E",x"05", -- 0x07E8
    x"CD",x"B1",x"04",x"3A",x"02",x"40",x"FE",x"63", -- 0x07F0
    x"38",x"02",x"3E",x"63",x"CD",x"12",x"08",x"47", -- 0x07F8
    x"E6",x"F0",x"28",x"07",x"0F",x"0F",x"0F",x"0F", -- 0x0800
    x"32",x"9F",x"52",x"78",x"E6",x"0F",x"32",x"7F", -- 0x0808
    x"52",x"C9",x"47",x"E6",x"0F",x"C6",x"00",x"27", -- 0x0810
    x"4F",x"78",x"E6",x"F0",x"28",x"0B",x"0F",x"0F", -- 0x0818
    x"0F",x"0F",x"47",x"AF",x"C6",x"16",x"27",x"10", -- 0x0820
    x"FB",x"81",x"27",x"C9",x"3A",x"1D",x"41",x"47", -- 0x0828
    x"4F",x"21",x"7F",x"50",x"11",x"20",x"00",x"A7", -- 0x0830
    x"28",x"05",x"36",x"CC",x"19",x"10",x"FB",x"3E", -- 0x0838
    x"06",x"91",x"47",x"36",x"10",x"19",x"10",x"FB", -- 0x0840
    x"C9",x"DD",x"21",x"CE",x"43",x"FD",x"21",x"38", -- 0x0848
    x"52",x"0E",x"05",x"06",x"03",x"11",x"E0",x"FF", -- 0x0850
    x"26",x"04",x"DD",x"7E",x"00",x"0F",x"0F",x"0F", -- 0x0858
    x"0F",x"CD",x"77",x"08",x"DD",x"7E",x"00",x"CD", -- 0x0860
    x"77",x"08",x"DD",x"2B",x"10",x"EC",x"11",x"BE", -- 0x0868
    x"00",x"FD",x"19",x"0D",x"20",x"DD",x"C9",x"E6", -- 0x0870
    x"0F",x"6F",x"7C",x"A7",x"20",x"06",x"FD",x"75", -- 0x0878
    x"00",x"FD",x"19",x"C9",x"7D",x"A7",x"20",x"04", -- 0x0880
    x"25",x"FD",x"19",x"C9",x"26",x"00",x"FD",x"75", -- 0x0888
    x"00",x"FD",x"19",x"C9",x"F5",x"C5",x"D5",x"E5", -- 0x0890
    x"DD",x"E5",x"FD",x"E5",x"AF",x"32",x"01",x"70", -- 0x0898
    x"21",x"20",x"40",x"11",x"00",x"58",x"01",x"80", -- 0x08A0
    x"00",x"ED",x"B0",x"3A",x"00",x"78",x"3A",x"15", -- 0x08A8
    x"40",x"32",x"16",x"40",x"3A",x"13",x"40",x"32", -- 0x08B0
    x"15",x"40",x"2A",x"10",x"40",x"22",x"13",x"40", -- 0x08B8
    x"21",x"12",x"40",x"3A",x"00",x"70",x"77",x"2B", -- 0x08C0
    x"3A",x"00",x"68",x"77",x"2B",x"3A",x"00",x"60", -- 0x08C8
    x"77",x"21",x"5F",x"42",x"35",x"CD",x"1A",x"09", -- 0x08D0
    x"CD",x"3D",x"09",x"CD",x"86",x"09",x"CD",x"B8", -- 0x08D8
    x"09",x"3A",x"06",x"40",x"0F",x"38",x"10",x"AF", -- 0x08E0
    x"32",x"C0",x"58",x"32",x"A0",x"58",x"32",x"B0", -- 0x08E8
    x"58",x"32",x"D0",x"58",x"32",x"E0",x"58",x"CD", -- 0x08F0
    x"CC",x"2A",x"21",x"0C",x"09",x"E5",x"3A",x"05", -- 0x08F8
    x"40",x"EF",x"FF",x"09",x"C1",x"0A",x"05",x"0F", -- 0x0900
    x"80",x"11",x"A7",x"11",x"FD",x"E1",x"DD",x"E1", -- 0x0908
    x"E1",x"D1",x"C1",x"3E",x"01",x"32",x"01",x"70", -- 0x0910
    x"F1",x"C9",x"21",x"10",x"40",x"7E",x"23",x"23", -- 0x0918
    x"23",x"B6",x"23",x"23",x"2F",x"A6",x"23",x"A6", -- 0x0920
    x"E6",x"03",x"C8",x"CB",x"47",x"C4",x"38",x"09", -- 0x0928
    x"CB",x"4F",x"C8",x"21",x"81",x"58",x"34",x"C9", -- 0x0930
    x"21",x"85",x"58",x"34",x"C9",x"21",x"84",x"58", -- 0x0938
    x"7E",x"A7",x"20",x"3A",x"23",x"B6",x"C8",x"35", -- 0x0940
    x"2B",x"36",x"0F",x"3A",x"00",x"40",x"CB",x"47", -- 0x0948
    x"28",x"1C",x"21",x"02",x"40",x"7E",x"FE",x"63", -- 0x0950
    x"C8",x"30",x"10",x"34",x"21",x"90",x"58",x"CB", -- 0x0958
    x"CE",x"3A",x"06",x"40",x"0F",x"D8",x"11",x"01", -- 0x0960
    x"07",x"FF",x"C9",x"36",x"63",x"C9",x"21",x"01", -- 0x0968
    x"40",x"CB",x"46",x"28",x"06",x"36",x"00",x"23", -- 0x0970
    x"C3",x"55",x"09",x"36",x"01",x"C9",x"0F",x"0F", -- 0x0978
    x"0F",x"32",x"03",x"60",x"35",x"C9",x"21",x"80", -- 0x0980
    x"58",x"7E",x"A7",x"20",x"6A",x"23",x"B6",x"C8", -- 0x0988
    x"35",x"2B",x"36",x"0F",x"21",x"02",x"40",x"34", -- 0x0990
    x"34",x"34",x"3A",x"00",x"40",x"CB",x"4F",x"20", -- 0x0998
    x"02",x"34",x"34",x"7E",x"FE",x"63",x"C8",x"30", -- 0x09A0
    x"4B",x"21",x"90",x"58",x"CB",x"CE",x"3A",x"06", -- 0x09A8
    x"40",x"0F",x"D8",x"11",x"01",x"07",x"FF",x"C9", -- 0x09B0
    x"21",x"03",x"40",x"5E",x"16",x"06",x"1A",x"1C", -- 0x09B8
    x"73",x"23",x"86",x"3D",x"77",x"3A",x"B0",x"40", -- 0x09C0
    x"0F",x"D0",x"2A",x"B1",x"40",x"7E",x"E6",x"07", -- 0x09C8
    x"20",x"1B",x"EB",x"2A",x"B3",x"40",x"7E",x"FE", -- 0x09D0
    x"3F",x"28",x"11",x"23",x"22",x"B3",x"40",x"D6", -- 0x09D8
    x"30",x"2A",x"B5",x"40",x"77",x"01",x"E0",x"FF", -- 0x09E0
    x"09",x"22",x"B5",x"40",x"EB",x"35",x"C0",x"AF", -- 0x09E8
    x"32",x"B0",x"40",x"C9",x"36",x"63",x"C9",x"0F", -- 0x09F0
    x"0F",x"0F",x"32",x"04",x"68",x"35",x"C9",x"2A", -- 0x09F8
    x"0B",x"40",x"06",x"20",x"3E",x"10",x"D7",x"22", -- 0x0A00
    x"0B",x"40",x"21",x"08",x"40",x"35",x"C0",x"2D", -- 0x0A08
    x"2D",x"36",x"00",x"2D",x"36",x"01",x"AF",x"32", -- 0x0A10
    x"0A",x"40",x"21",x"41",x"0A",x"CD",x"30",x"0A", -- 0x0A18
    x"11",x"04",x"06",x"FF",x"11",x"00",x"05",x"FF", -- 0x0A20
    x"1E",x"02",x"FF",x"AF",x"32",x"80",x"42",x"C9", -- 0x0A28
    x"11",x"21",x"40",x"06",x"20",x"7E",x"12",x"23", -- 0x0A30
    x"1C",x"EB",x"36",x"00",x"EB",x"1C",x"10",x"F5", -- 0x0A38
    x"C9",x"00",x"05",x"00",x"00",x"00",x"01",x"06", -- 0x0A40
    x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x0A48
    x"00",x"00",x"00",x"00",x"05",x"05",x"05",x"05", -- 0x0A50
    x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06", -- 0x0A58
    x"06",x"00",x"05",x"00",x"00",x"01",x"01",x"06", -- 0x0A60
    x"03",x"03",x"04",x"04",x"04",x"04",x"00",x"00", -- 0x0A68
    x"00",x"06",x"06",x"06",x"00",x"00",x"00",x"05", -- 0x0A70
    x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06", -- 0x0A78
    x"06",x"00",x"05",x"02",x"02",x"02",x"02",x"06", -- 0x0A80
    x"02",x"00",x"00",x"02",x"01",x"01",x"01",x"01", -- 0x0A88
    x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06", -- 0x0A90
    x"06",x"06",x"06",x"06",x"06",x"00",x"06",x"06", -- 0x0A98
    x"06",x"00",x"05",x"00",x"00",x"00",x"00",x"06", -- 0x0AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA8
    x"00",x"05",x"05",x"02",x"02",x"06",x"06",x"07", -- 0x0AB0
    x"07",x"04",x"04",x"00",x"00",x"00",x"06",x"06", -- 0x0AB8
    x"06",x"21",x"E9",x"0E",x"E5",x"3A",x"80",x"42", -- 0x0AC0
    x"EF",x"E9",x"0A",x"34",x"0B",x"6F",x"0B",x"90", -- 0x0AC8
    x"0B",x"C2",x"0B",x"D6",x"0B",x"F3",x"0B",x"34", -- 0x0AD0
    x"0C",x"5D",x"0C",x"5E",x"0C",x"5F",x"0C",x"79", -- 0x0AD8
    x"0C",x"F9",x"0C",x"49",x"0D",x"64",x"0D",x"65", -- 0x0AE0
    x"0D",x"AF",x"32",x"C0",x"58",x"32",x"A0",x"58", -- 0x0AE8
    x"32",x"B0",x"58",x"32",x"D0",x"58",x"32",x"E0", -- 0x0AF0
    x"58",x"21",x"20",x"40",x"11",x"21",x"40",x"01", -- 0x0AF8
    x"7F",x"00",x"36",x"00",x"ED",x"B0",x"21",x"00", -- 0x0B00
    x"41",x"11",x"01",x"41",x"01",x"FF",x"01",x"36", -- 0x0B08
    x"00",x"ED",x"B0",x"21",x"A0",x"42",x"11",x"A1", -- 0x0B10
    x"42",x"01",x"FF",x"00",x"36",x"00",x"ED",x"B0", -- 0x0B18
    x"21",x"02",x"50",x"22",x"0B",x"40",x"21",x"09", -- 0x0B20
    x"40",x"36",x"20",x"21",x"80",x"42",x"34",x"AF", -- 0x0B28
    x"32",x"06",x"40",x"C9",x"2A",x"0B",x"40",x"06", -- 0x0B30
    x"1E",x"3E",x"10",x"D7",x"11",x"02",x"00",x"19", -- 0x0B38
    x"22",x"0B",x"40",x"21",x"09",x"40",x"35",x"C0", -- 0x0B40
    x"21",x"81",x"0A",x"CD",x"30",x"0A",x"3E",x"01", -- 0x0B48
    x"32",x"06",x"70",x"32",x"07",x"70",x"21",x"80", -- 0x0B50
    x"42",x"34",x"2C",x"36",x"01",x"2C",x"36",x"0B", -- 0x0B58
    x"2C",x"36",x"1E",x"11",x"01",x"07",x"FF",x"11", -- 0x0B60
    x"11",x"06",x"FF",x"1E",x"07",x"FF",x"C9",x"21", -- 0x0B68
    x"83",x"42",x"35",x"C0",x"36",x"1E",x"2D",x"5E", -- 0x0B70
    x"34",x"16",x"06",x"FF",x"7B",x"FE",x"0E",x"C0", -- 0x0B78
    x"2D",x"2D",x"34",x"21",x"1C",x"0C",x"22",x"84", -- 0x0B80
    x"42",x"21",x"60",x"40",x"22",x"86",x"42",x"C9", -- 0x0B88
    x"21",x"83",x"42",x"35",x"C0",x"36",x"1E",x"2D", -- 0x0B90
    x"5E",x"34",x"16",x"06",x"FF",x"2A",x"84",x"42", -- 0x0B98
    x"ED",x"5B",x"86",x"42",x"01",x"08",x"00",x"ED", -- 0x0BA0
    x"B0",x"22",x"84",x"42",x"ED",x"53",x"86",x"42", -- 0x0BA8
    x"3A",x"82",x"42",x"FE",x"12",x"C0",x"21",x"80", -- 0x0BB0
    x"42",x"34",x"2C",x"2C",x"36",x"0C",x"2C",x"36", -- 0x0BB8
    x"1E",x"C9",x"21",x"83",x"42",x"35",x"C0",x"36", -- 0x0BC0
    x"0F",x"11",x"0E",x"06",x"FF",x"1C",x"FF",x"1C", -- 0x0BC8
    x"FF",x"2D",x"2D",x"2D",x"34",x"C9",x"21",x"83", -- 0x0BD0
    x"42",x"35",x"C0",x"36",x"0F",x"11",x"8E",x"06", -- 0x0BD8
    x"FF",x"1C",x"FF",x"1C",x"FF",x"2D",x"35",x"28", -- 0x0BE0
    x"04",x"2D",x"2D",x"35",x"C9",x"36",x"14",x"2D", -- 0x0BE8
    x"2D",x"34",x"C9",x"21",x"82",x"42",x"35",x"C0", -- 0x0BF0
    x"36",x"96",x"11",x"8D",x"06",x"FF",x"21",x"60", -- 0x0BF8
    x"40",x"11",x"61",x"40",x"01",x"1F",x"00",x"36", -- 0x0C00
    x"00",x"ED",x"B0",x"3A",x"00",x"40",x"C6",x"12", -- 0x0C08
    x"5F",x"16",x"06",x"FF",x"1E",x"06",x"FF",x"21", -- 0x0C10
    x"80",x"42",x"34",x"C9",x"34",x"EB",x"07",x"8B", -- 0x0C18
    x"8B",x"22",x"07",x"8B",x"34",x"EB",x"03",x"A3", -- 0x0C20
    x"8B",x"22",x"03",x"A3",x"34",x"EB",x"01",x"BB", -- 0x0C28
    x"8B",x"22",x"01",x"BB",x"21",x"82",x"42",x"35", -- 0x0C30
    x"C0",x"21",x"A1",x"0A",x"CD",x"30",x"0A",x"11", -- 0x0C38
    x"92",x"06",x"FF",x"1E",x"86",x"FF",x"1E",x"1A", -- 0x0C40
    x"06",x"06",x"FF",x"1C",x"10",x"FC",x"11",x"02", -- 0x0C48
    x"07",x"FF",x"21",x"80",x"42",x"34",x"34",x"34", -- 0x0C50
    x"2C",x"2C",x"36",x"DC",x"C9",x"C9",x"C9",x"3A", -- 0x0C58
    x"5F",x"42",x"0F",x"D8",x"21",x"82",x"42",x"35", -- 0x0C60
    x"C0",x"3E",x"20",x"32",x"09",x"40",x"21",x"02", -- 0x0C68
    x"50",x"22",x"0B",x"40",x"21",x"80",x"42",x"34", -- 0x0C70
    x"C9",x"2A",x"0B",x"40",x"06",x"1D",x"3E",x"10", -- 0x0C78
    x"D7",x"11",x"03",x"00",x"19",x"22",x"0B",x"40", -- 0x0C80
    x"21",x"09",x"40",x"35",x"C0",x"21",x"41",x"0A", -- 0x0C88
    x"CD",x"30",x"0A",x"21",x"E8",x"0C",x"22",x"07", -- 0x0C90
    x"42",x"AF",x"32",x"5F",x"42",x"3E",x"01",x"32", -- 0x0C98
    x"06",x"70",x"32",x"07",x"70",x"AF",x"32",x"0D", -- 0x0CA0
    x"40",x"21",x"92",x"10",x"11",x"00",x"41",x"01", -- 0x0CA8
    x"E0",x"00",x"ED",x"B0",x"21",x"66",x"0D",x"11", -- 0x0CB0
    x"50",x"41",x"01",x"90",x"00",x"ED",x"B0",x"3E", -- 0x0CB8
    x"01",x"32",x"00",x"41",x"3E",x"0B",x"32",x"1A", -- 0x0CC0
    x"41",x"21",x"01",x"00",x"22",x"00",x"42",x"3E", -- 0x0CC8
    x"18",x"32",x"02",x"42",x"3E",x"67",x"32",x"52", -- 0x0CD0
    x"40",x"32",x"54",x"40",x"11",x"00",x"02",x"FF", -- 0x0CD8
    x"21",x"80",x"42",x"34",x"2C",x"36",x"00",x"C9", -- 0x0CE0
    x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08", -- 0x0CE8
    x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08", -- 0x0CF0
    x"FF",x"CD",x"1C",x"15",x"CD",x"85",x"1C",x"CD", -- 0x0CF8
    x"AB",x"1C",x"CD",x"7B",x"18",x"CD",x"8E",x"18", -- 0x0D00
    x"3A",x"16",x"41",x"A7",x"CC",x"E0",x"1C",x"CD", -- 0x0D08
    x"1F",x"18",x"CD",x"13",x"19",x"CD",x"6D",x"0E", -- 0x0D10
    x"CD",x"65",x"1A",x"3A",x"8B",x"42",x"A7",x"CC", -- 0x0D18
    x"E0",x"1B",x"CD",x"41",x"1B",x"3A",x"1A",x"41", -- 0x0D20
    x"A7",x"28",x"07",x"3A",x"11",x"41",x"A7",x"28", -- 0x0D28
    x"01",x"C9",x"21",x"80",x"42",x"34",x"2C",x"2C", -- 0x0D30
    x"36",x"B4",x"AF",x"32",x"90",x"42",x"CD",x"00", -- 0x0D38
    x"12",x"11",x"00",x"06",x"FF",x"1E",x"02",x"FF", -- 0x0D40
    x"C9",x"CD",x"AB",x"1C",x"CD",x"7B",x"18",x"CD", -- 0x0D48
    x"8E",x"18",x"CD",x"C1",x"15",x"3A",x"5F",x"42", -- 0x0D50
    x"0F",x"D8",x"21",x"82",x"42",x"35",x"C0",x"2D", -- 0x0D58
    x"2D",x"36",x"00",x"C9",x"C9",x"C9",x"03",x"03", -- 0x0D60
    x"03",x"03",x"01",x"01",x"03",x"03",x"03",x"03", -- 0x0D68
    x"01",x"01",x"00",x"00",x"00",x"00",x"01",x"01", -- 0x0D70
    x"00",x"00",x"00",x"03",x"01",x"00",x"00",x"00", -- 0x0D78
    x"03",x"03",x"00",x"00",x"00",x"03",x"03",x"00", -- 0x0D80
    x"00",x"00",x"03",x"03",x"03",x"03",x"01",x"01", -- 0x0D88
    x"03",x"03",x"03",x"03",x"01",x"01",x"03",x"03", -- 0x0D90
    x"00",x"00",x"03",x"03",x"03",x"03",x"00",x"00", -- 0x0D98
    x"03",x"03",x"03",x"03",x"00",x"00",x"03",x"03", -- 0x0DA0
    x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03", -- 0x0DA8
    x"03",x"03",x"03",x"03",x"03",x"03",x"00",x"00", -- 0x0DB0
    x"03",x"03",x"03",x"03",x"00",x"00",x"03",x"03", -- 0x0DB8
    x"03",x"03",x"00",x"00",x"03",x"03",x"03",x"00", -- 0x0DC0
    x"00",x"00",x"00",x"00",x"03",x"00",x"03",x"03", -- 0x0DC8
    x"00",x"00",x"03",x"00",x"03",x"03",x"00",x"00", -- 0x0DD0
    x"03",x"00",x"03",x"03",x"00",x"00",x"03",x"00", -- 0x0DD8
    x"03",x"03",x"00",x"00",x"03",x"00",x"03",x"03", -- 0x0DE0
    x"00",x"00",x"03",x"03",x"03",x"03",x"03",x"03", -- 0x0DE8
    x"03",x"03",x"03",x"03",x"03",x"03",x"3A",x"16", -- 0x0DF0
    x"41",x"A7",x"C8",x"3A",x"88",x"42",x"EF",x"05", -- 0x0DF8
    x"0E",x"1B",x"0E",x"3E",x"0E",x"ED",x"5F",x"0F", -- 0x0E00
    x"3E",x"68",x"38",x"02",x"3E",x"B8",x"21",x"88", -- 0x0E08
    x"42",x"34",x"2C",x"77",x"2C",x"36",x"28",x"2C", -- 0x0E10
    x"36",x"01",x"C9",x"21",x"02",x"42",x"3A",x"89", -- 0x0E18
    x"42",x"BE",x"28",x"11",x"38",x"03",x"34",x"18", -- 0x0E20
    x"01",x"35",x"7E",x"2F",x"C6",x"80",x"32",x"58", -- 0x0E28
    x"40",x"32",x"5A",x"40",x"C9",x"21",x"88",x"42", -- 0x0E30
    x"34",x"AF",x"32",x"8B",x"42",x"C9",x"21",x"64", -- 0x0E38
    x"42",x"CB",x"46",x"C8",x"2C",x"3A",x"02",x"42", -- 0x0E40
    x"C6",x"08",x"96",x"D8",x"FE",x"10",x"D0",x"2C", -- 0x0E48
    x"2C",x"7E",x"FE",x"B8",x"D8",x"21",x"02",x"42", -- 0x0E50
    x"35",x"7E",x"2F",x"C6",x"80",x"32",x"58",x"40", -- 0x0E58
    x"32",x"5A",x"40",x"21",x"8A",x"42",x"35",x"C0", -- 0x0E60
    x"2D",x"2D",x"36",x"00",x"C9",x"3A",x"7C",x"42", -- 0x0E68
    x"0F",x"D8",x"DD",x"21",x"A0",x"42",x"11",x"20", -- 0x0E70
    x"00",x"06",x"08",x"D9",x"CD",x"85",x"0E",x"D9", -- 0x0E78
    x"DD",x"19",x"10",x"F7",x"C9",x"DD",x"CB",x"00", -- 0x0E80
    x"46",x"C8",x"DD",x"CB",x"08",x"46",x"C8",x"DD", -- 0x0E88
    x"CB",x"09",x"46",x"C0",x"DD",x"7E",x"0B",x"FE", -- 0x0E90
    x"80",x"D0",x"DD",x"7E",x"03",x"FE",x"60",x"D8", -- 0x0E98
    x"FE",x"C0",x"D0",x"DD",x"4E",x"06",x"DD",x"46", -- 0x0EA0
    x"08",x"3A",x"02",x"42",x"05",x"28",x"09",x"B9", -- 0x0EA8
    x"D8",x"4F",x"DD",x"7E",x"04",x"91",x"18",x"05", -- 0x0EB0
    x"B9",x"D0",x"DD",x"96",x"04",x"D8",x"47",x"3E", -- 0x0EB8
    x"E0",x"DD",x"96",x"03",x"DD",x"CB",x"19",x"46", -- 0x0EC0
    x"20",x"13",x"DD",x"4E",x"16",x"0D",x"28",x"0D", -- 0x0EC8
    x"0F",x"0F",x"0F",x"E6",x"1F",x"B8",x"C0",x"3E", -- 0x0ED0
    x"01",x"32",x"7C",x"42",x"C9",x"0F",x"0F",x"E6", -- 0x0ED8
    x"3F",x"B8",x"C0",x"3E",x"01",x"32",x"7C",x"42", -- 0x0EE0
    x"C9",x"3A",x"02",x"40",x"A7",x"C8",x"21",x"05", -- 0x0EE8
    x"40",x"34",x"AF",x"32",x"0A",x"40",x"32",x"81", -- 0x0EF0
    x"42",x"21",x"96",x"10",x"11",x"04",x"41",x"01", -- 0x0EF8
    x"0C",x"00",x"ED",x"B0",x"C9",x"21",x"E8",x"0F", -- 0x0F00
    x"E5",x"3A",x"0A",x"40",x"EF",x"13",x"0F",x"49", -- 0x0F08
    x"0F",x"DA",x"0F",x"AF",x"32",x"00",x"41",x"11", -- 0x0F10
    x"00",x"01",x"FF",x"21",x"61",x"0A",x"CD",x"30", -- 0x0F18
    x"0A",x"21",x"60",x"40",x"06",x"40",x"AF",x"D7", -- 0x0F20
    x"21",x"60",x"42",x"D7",x"06",x"40",x"D7",x"21", -- 0x0F28
    x"20",x"41",x"06",x"C0",x"D7",x"32",x"B0",x"40", -- 0x0F30
    x"32",x"06",x"40",x"21",x"02",x"50",x"22",x"0B", -- 0x0F38
    x"40",x"21",x"09",x"40",x"36",x"10",x"2C",x"34", -- 0x0F40
    x"C9",x"2A",x"0B",x"40",x"06",x"1D",x"3E",x"10", -- 0x0F48
    x"D7",x"11",x"03",x"00",x"19",x"06",x"1D",x"D7", -- 0x0F50
    x"19",x"22",x"0B",x"40",x"21",x"09",x"40",x"35", -- 0x0F58
    x"C0",x"2C",x"34",x"3E",x"01",x"32",x"06",x"70", -- 0x0F60
    x"32",x"07",x"70",x"AF",x"32",x"0D",x"40",x"11", -- 0x0F68
    x"01",x"07",x"FF",x"11",x"01",x"06",x"FF",x"1E", -- 0x0F70
    x"16",x"FF",x"1C",x"FF",x"3A",x"17",x"40",x"47", -- 0x0F78
    x"E6",x"0F",x"32",x"78",x"51",x"78",x"E6",x"F0", -- 0x0F80
    x"C8",x"0F",x"0F",x"0F",x"0F",x"32",x"98",x"51", -- 0x0F88
    x"C9",x"3A",x"00",x"42",x"0F",x"D0",x"DD",x"21", -- 0x0F90
    x"A0",x"42",x"11",x"20",x"00",x"06",x"08",x"D9", -- 0x0F98
    x"CD",x"A9",x"0F",x"D9",x"DD",x"19",x"10",x"F7", -- 0x0FA0
    x"C9",x"DD",x"CB",x"00",x"46",x"C8",x"DD",x"7E", -- 0x0FA8
    x"03",x"C6",x"39",x"D6",x"05",x"38",x"10",x"D6", -- 0x0FB0
    x"0C",x"D0",x"3A",x"02",x"42",x"DD",x"96",x"04", -- 0x0FB8
    x"C6",x"0A",x"FE",x"15",x"D0",x"18",x"0B",x"3A", -- 0x0FC0
    x"02",x"42",x"DD",x"96",x"04",x"C6",x"07",x"FE", -- 0x0FC8
    x"0F",x"D0",x"3E",x"01",x"32",x"04",x"42",x"C3", -- 0x0FD0
    x"9C",x"1A",x"3A",x"02",x"40",x"A7",x"C8",x"3D", -- 0x0FD8
    x"11",x"18",x"06",x"28",x"01",x"1C",x"FF",x"C9", -- 0x0FE0
    x"3A",x"11",x"40",x"CB",x"47",x"C2",x"7C",x"10", -- 0x0FE8
    x"CB",x"4F",x"C8",x"3A",x"02",x"40",x"FE",x"02", -- 0x0FF0
    x"D8",x"D6",x"02",x"32",x"02",x"40",x"21",x"00", -- 0x0FF8
    x"01",x"22",x"0D",x"40",x"AF",x"32",x"0A",x"40", -- 0x1000
    x"3E",x"03",x"32",x"05",x"40",x"3E",x"01",x"32", -- 0x1008
    x"06",x"40",x"11",x"04",x"06",x"FF",x"21",x"92", -- 0x1010
    x"10",x"11",x"00",x"41",x"01",x"E0",x"00",x"ED", -- 0x1018
    x"B0",x"21",x"92",x"10",x"11",x"E0",x"41",x"01", -- 0x1020
    x"20",x"00",x"ED",x"B0",x"DD",x"21",x"20",x"41", -- 0x1028
    x"21",x"10",x"42",x"0E",x"30",x"06",x"04",x"CB", -- 0x1030
    x"26",x"CB",x"26",x"DD",x"CB",x"00",x"46",x"28", -- 0x1038
    x"02",x"CB",x"C6",x"DD",x"CB",x"00",x"4E",x"28", -- 0x1040
    x"02",x"CB",x"CE",x"DD",x"23",x"10",x"E8",x"23", -- 0x1048
    x"0D",x"20",x"E2",x"3E",x"01",x"32",x"00",x"41", -- 0x1050
    x"32",x"E0",x"41",x"3A",x"07",x"40",x"32",x"1D", -- 0x1058
    x"41",x"32",x"FD",x"41",x"AF",x"32",x"52",x"40", -- 0x1060
    x"32",x"54",x"40",x"21",x"A0",x"58",x"CB",x"C6", -- 0x1068
    x"11",x"00",x"04",x"FF",x"3A",x"0E",x"40",x"0F", -- 0x1070
    x"D0",x"1C",x"FF",x"C9",x"3A",x"02",x"40",x"A7", -- 0x1078
    x"28",x"0A",x"3D",x"32",x"02",x"40",x"21",x"00", -- 0x1080
    x"00",x"C3",x"01",x"10",x"3E",x"01",x"32",x"05", -- 0x1088
    x"40",x"C9",x"00",x"80",x"00",x"06",x"6C",x"64", -- 0x1090
    x"64",x"64",x"64",x"65",x"30",x"31",x"32",x"33", -- 0x1098
    x"34",x"35",x"00",x"2E",x"00",x"00",x"00",x"00", -- 0x10A0
    x"00",x"1C",x"20",x"24",x"60",x"30",x"00",x"03", -- 0x10A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10D8
    x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x10E0
    x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00", -- 0x10E8
    x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"01", -- 0x10F0
    x"01",x"00",x"00",x"00",x"01",x"01",x"00",x"00", -- 0x10F8
    x"00",x"01",x"01",x"00",x"00",x"00",x"01",x"01", -- 0x1100
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1108
    x"01",x"01",x"01",x"01",x"00",x"00",x"01",x"01", -- 0x1110
    x"01",x"01",x"00",x"00",x"01",x"01",x"01",x"01", -- 0x1118
    x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1120
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1128
    x"01",x"01",x"00",x"00",x"01",x"01",x"01",x"01", -- 0x1130
    x"00",x"00",x"01",x"01",x"01",x"01",x"00",x"00", -- 0x1138
    x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x1140
    x"01",x"00",x"01",x"01",x"00",x"00",x"01",x"00", -- 0x1148
    x"01",x"01",x"00",x"00",x"01",x"00",x"01",x"01", -- 0x1150
    x"00",x"00",x"01",x"00",x"01",x"01",x"00",x"00", -- 0x1158
    x"01",x"00",x"01",x"01",x"00",x"00",x"01",x"01", -- 0x1160
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1168
    x"01",x"01",x"21",x"09",x"40",x"35",x"C0",x"36", -- 0x1170
    x"00",x"11",x"60",x"06",x"FF",x"2C",x"34",x"C9", -- 0x1178
    x"CD",x"85",x"1C",x"CD",x"AB",x"1C",x"CD",x"7B", -- 0x1180
    x"18",x"CD",x"8E",x"18",x"CD",x"1C",x"15",x"3A", -- 0x1188
    x"0A",x"40",x"EF",x"CE",x"11",x"0F",x"12",x"28", -- 0x1190
    x"12",x"A6",x"12",x"B7",x"12",x"F1",x"12",x"A0", -- 0x1198
    x"13",x"D1",x"13",x"6C",x"15",x"AB",x"15",x"CD", -- 0x11A0
    x"85",x"1C",x"CD",x"AB",x"1C",x"CD",x"7B",x"18", -- 0x11A8
    x"CD",x"8E",x"18",x"CD",x"1C",x"15",x"3A",x"0A", -- 0x11B0
    x"40",x"EF",x"CE",x"11",x"0F",x"12",x"69",x"12", -- 0x11B8
    x"A6",x"12",x"B7",x"12",x"F1",x"12",x"13",x"14", -- 0x11C0
    x"35",x"14",x"6C",x"15",x"AB",x"15",x"AF",x"32", -- 0x11C8
    x"B0",x"58",x"32",x"D0",x"58",x"32",x"E0",x"58", -- 0x11D0
    x"AF",x"32",x"81",x"42",x"21",x"00",x"42",x"06", -- 0x11D8
    x"10",x"D7",x"21",x"60",x"42",x"D7",x"06",x"40", -- 0x11E0
    x"D7",x"CD",x"00",x"12",x"21",x"89",x"1B",x"22", -- 0x11E8
    x"07",x"42",x"21",x"0A",x"40",x"34",x"2D",x"36", -- 0x11F0
    x"20",x"21",x"00",x"50",x"22",x"0B",x"40",x"C9", -- 0x11F8
    x"21",x"60",x"40",x"06",x"40",x"AF",x"D7",x"AF", -- 0x1200
    x"32",x"52",x"40",x"32",x"54",x"40",x"C9",x"2A", -- 0x1208
    x"0B",x"40",x"06",x"20",x"3E",x"10",x"D7",x"22", -- 0x1210
    x"0B",x"40",x"21",x"09",x"40",x"35",x"C0",x"2C", -- 0x1218
    x"34",x"21",x"41",x"0A",x"CD",x"30",x"0A",x"C9", -- 0x1220
    x"AF",x"32",x"5F",x"42",x"3E",x"01",x"32",x"06", -- 0x1228
    x"70",x"32",x"07",x"70",x"AF",x"32",x"0D",x"40", -- 0x1230
    x"21",x"0A",x"40",x"34",x"2D",x"36",x"00",x"3A", -- 0x1238
    x"0E",x"40",x"0F",x"38",x"1E",x"11",x"00",x"05", -- 0x1240
    x"FF",x"1E",x"02",x"FF",x"14",x"FF",x"1E",x"04", -- 0x1248
    x"FF",x"3A",x"14",x"41",x"A7",x"C2",x"5B",x"12", -- 0x1250
    x"1E",x"60",x"FF",x"11",x"03",x"07",x"FF",x"1E", -- 0x1258
    x"00",x"FF",x"C9",x"11",x"01",x"05",x"FF",x"18", -- 0x1260
    x"DC",x"AF",x"32",x"5F",x"42",x"3A",x"0F",x"40", -- 0x1268
    x"0F",x"30",x"07",x"AF",x"32",x"06",x"70",x"32", -- 0x1270
    x"07",x"70",x"3E",x"01",x"32",x"0D",x"40",x"21", -- 0x1278
    x"0A",x"40",x"34",x"2D",x"36",x"00",x"11",x"00", -- 0x1280
    x"05",x"FF",x"1C",x"FF",x"1C",x"FF",x"11",x"03", -- 0x1288
    x"06",x"FF",x"1C",x"FF",x"3A",x"14",x"41",x"A7", -- 0x1290
    x"C2",x"9E",x"12",x"1E",x"60",x"FF",x"11",x"03", -- 0x1298
    x"07",x"FF",x"1E",x"00",x"FF",x"C9",x"21",x"09", -- 0x12A0
    x"40",x"35",x"C0",x"36",x"14",x"2C",x"34",x"11", -- 0x12A8
    x"82",x"06",x"FF",x"1E",x"A0",x"FF",x"C9",x"21", -- 0x12B0
    x"09",x"40",x"35",x"C0",x"36",x"0A",x"2C",x"34", -- 0x12B8
    x"21",x"60",x"42",x"06",x"20",x"AF",x"D7",x"21", -- 0x12C0
    x"01",x"00",x"22",x"00",x"42",x"3E",x"18",x"32", -- 0x12C8
    x"02",x"42",x"AF",x"32",x"52",x"40",x"32",x"54", -- 0x12D0
    x"40",x"3A",x"07",x"40",x"A7",x"20",x"05",x"3E", -- 0x12D8
    x"02",x"32",x"1D",x"41",x"21",x"1D",x"41",x"35", -- 0x12E0
    x"11",x"03",x"07",x"FF",x"11",x"00",x"02",x"FF", -- 0x12E8
    x"C9",x"CD",x"4D",x"13",x"CD",x"76",x"17",x"CD", -- 0x12F0
    x"54",x"15",x"CD",x"AF",x"17",x"CD",x"C5",x"17", -- 0x12F8
    x"CD",x"1F",x"18",x"CD",x"13",x"19",x"CD",x"91", -- 0x1300
    x"0F",x"CD",x"DC",x"18",x"CD",x"65",x"1A",x"CD", -- 0x1308
    x"0A",x"1B",x"CD",x"A2",x"1B",x"CD",x"E0",x"1B", -- 0x1310
    x"CD",x"5E",x"1C",x"CD",x"41",x"1B",x"3A",x"1A", -- 0x1318
    x"41",x"A7",x"28",x"43",x"3A",x"11",x"41",x"A7", -- 0x1320
    x"28",x"4E",x"21",x"00",x"42",x"CB",x"46",x"C0", -- 0x1328
    x"23",x"CB",x"46",x"C0",x"3A",x"7C",x"42",x"0F", -- 0x1330
    x"D8",x"3A",x"60",x"42",x"47",x"3A",x"64",x"42", -- 0x1338
    x"4F",x"3A",x"68",x"42",x"B0",x"B1",x"0F",x"D8", -- 0x1340
    x"21",x"0A",x"40",x"34",x"C9",x"21",x"A0",x"42", -- 0x1348
    x"11",x"20",x"00",x"06",x"08",x"AF",x"B6",x"19", -- 0x1350
    x"10",x"FC",x"0F",x"21",x"C0",x"58",x"CB",x"D6", -- 0x1358
    x"D8",x"21",x"C0",x"58",x"CB",x"96",x"C9",x"3A", -- 0x1360
    x"01",x"42",x"0F",x"D8",x"AF",x"32",x"1D",x"41", -- 0x1368
    x"32",x"00",x"42",x"21",x"0A",x"40",x"34",x"C9", -- 0x1370
    x"21",x"00",x"42",x"CB",x"46",x"20",x"06",x"2C", -- 0x1378
    x"CB",x"46",x"C0",x"18",x"AF",x"AF",x"21",x"60", -- 0x1380
    x"42",x"06",x"20",x"D7",x"21",x"80",x"40",x"06", -- 0x1388
    x"20",x"D7",x"21",x"B7",x"40",x"36",x"00",x"23", -- 0x1390
    x"36",x"32",x"3E",x"08",x"32",x"0A",x"40",x"C9", -- 0x1398
    x"3A",x"1D",x"41",x"A7",x"20",x"14",x"11",x"00", -- 0x13A0
    x"06",x"FF",x"1E",x"02",x"FF",x"21",x"0A",x"40", -- 0x13A8
    x"36",x"09",x"2B",x"36",x"B4",x"AF",x"32",x"90", -- 0x13B0
    x"42",x"C9",x"3A",x"0E",x"40",x"0F",x"38",x"09", -- 0x13B8
    x"21",x"0A",x"40",x"36",x"04",x"2B",x"36",x"64", -- 0x13C0
    x"C9",x"21",x"0A",x"40",x"34",x"2D",x"36",x"64", -- 0x13C8
    x"C9",x"21",x"09",x"40",x"35",x"C0",x"3A",x"1D", -- 0x13D0
    x"41",x"A7",x"20",x"0C",x"3A",x"0E",x"40",x"0F", -- 0x13D8
    x"38",x"15",x"3E",x"01",x"32",x"05",x"40",x"C9", -- 0x13E0
    x"3A",x"FD",x"41",x"A7",x"20",x"15",x"21",x"0A", -- 0x13E8
    x"40",x"36",x"04",x"2B",x"36",x"01",x"C9",x"3A", -- 0x13F0
    x"FD",x"41",x"A7",x"20",x"06",x"3E",x"01",x"32", -- 0x13F8
    x"05",x"40",x"C9",x"CD",x"6B",x"14",x"CD",x"AC", -- 0x1400
    x"14",x"AF",x"32",x"0A",x"40",x"3E",x"04",x"32", -- 0x1408
    x"05",x"40",x"C9",x"3A",x"1D",x"41",x"A7",x"20", -- 0x1410
    x"14",x"11",x"00",x"06",x"FF",x"1E",x"03",x"FF", -- 0x1418
    x"21",x"0A",x"40",x"36",x"09",x"2B",x"36",x"B4", -- 0x1420
    x"AF",x"32",x"90",x"42",x"C9",x"21",x"0A",x"40", -- 0x1428
    x"34",x"2D",x"36",x"64",x"C9",x"21",x"09",x"40", -- 0x1430
    x"35",x"C0",x"3A",x"1D",x"41",x"A7",x"20",x"0C", -- 0x1438
    x"3A",x"FD",x"41",x"A7",x"20",x"15",x"3E",x"01", -- 0x1440
    x"32",x"05",x"40",x"C9",x"3A",x"FD",x"41",x"A7", -- 0x1448
    x"20",x"09",x"21",x"0A",x"40",x"36",x"04",x"2B", -- 0x1450
    x"36",x"01",x"C9",x"CD",x"6B",x"14",x"CD",x"AC", -- 0x1458
    x"14",x"AF",x"32",x"0A",x"40",x"3E",x"03",x"32", -- 0x1460
    x"05",x"40",x"C9",x"AF",x"21",x"A0",x"42",x"11", -- 0x1468
    x"20",x"00",x"06",x"08",x"CB",x"46",x"28",x"01", -- 0x1470
    x"3C",x"19",x"10",x"F8",x"47",x"21",x"12",x"41", -- 0x1478
    x"7E",x"90",x"77",x"21",x"96",x"10",x"11",x"04", -- 0x1480
    x"41",x"01",x"0C",x"00",x"ED",x"B0",x"3A",x"12", -- 0x1488
    x"41",x"A7",x"C8",x"47",x"16",x"00",x"DD",x"21", -- 0x1490
    x"2A",x"20",x"21",x"04",x"41",x"DD",x"5E",x"00", -- 0x1498
    x"19",x"DD",x"7E",x"01",x"77",x"1E",x"05",x"DD", -- 0x14A0
    x"19",x"10",x"EF",x"C9",x"21",x"00",x"41",x"DD", -- 0x14A8
    x"21",x"E0",x"41",x"06",x"20",x"DD",x"7E",x"00", -- 0x14B0
    x"4E",x"DD",x"71",x"00",x"77",x"DD",x"23",x"23", -- 0x14B8
    x"10",x"F3",x"DD",x"21",x"20",x"41",x"FD",x"21", -- 0x14C0
    x"10",x"42",x"06",x"30",x"FD",x"4E",x"00",x"3E", -- 0x14C8
    x"03",x"A1",x"6F",x"CB",x"09",x"CB",x"09",x"3E", -- 0x14D0
    x"03",x"A1",x"67",x"CB",x"09",x"CB",x"09",x"3E", -- 0x14D8
    x"03",x"A1",x"5F",x"CB",x"09",x"CB",x"09",x"3E", -- 0x14E0
    x"03",x"A1",x"57",x"FD",x"23",x"0E",x"04",x"CB", -- 0x14E8
    x"27",x"CB",x"27",x"DD",x"CB",x"00",x"4E",x"28", -- 0x14F0
    x"02",x"CB",x"CF",x"DD",x"CB",x"00",x"46",x"28", -- 0x14F8
    x"02",x"CB",x"C7",x"DD",x"23",x"0D",x"20",x"E7", -- 0x1500
    x"DD",x"72",x"FC",x"DD",x"73",x"FD",x"DD",x"74", -- 0x1508
    x"FE",x"DD",x"75",x"FF",x"FD",x"77",x"FF",x"05", -- 0x1510
    x"C2",x"CC",x"14",x"C9",x"3A",x"00",x"42",x"0F", -- 0x1518
    x"D0",x"3A",x"5F",x"42",x"E6",x"0F",x"C0",x"3A", -- 0x1520
    x"0D",x"42",x"16",x"02",x"FE",x"58",x"28",x"09", -- 0x1528
    x"FE",x"60",x"28",x"0E",x"FE",x"54",x"28",x"13", -- 0x1530
    x"C9",x"3E",x"60",x"32",x"0D",x"42",x"1E",x"07", -- 0x1538
    x"FF",x"C9",x"3E",x"54",x"32",x"0D",x"42",x"1E", -- 0x1540
    x"08",x"FF",x"C9",x"3E",x"58",x"32",x"0D",x"42", -- 0x1548
    x"1E",x"06",x"FF",x"C9",x"3A",x"1C",x"41",x"0F", -- 0x1550
    x"D0",x"3E",x"01",x"32",x"13",x"41",x"3A",x"5F", -- 0x1558
    x"42",x"E6",x"10",x"11",x"08",x"06",x"28",x"02", -- 0x1560
    x"1E",x"88",x"FF",x"C9",x"3A",x"16",x"41",x"A7", -- 0x1568
    x"CC",x"E0",x"1C",x"3A",x"B7",x"40",x"EF",x"68", -- 0x1570
    x"26",x"BC",x"26",x"F8",x"26",x"03",x"27",x"0F", -- 0x1578
    x"27",x"2B",x"27",x"78",x"27",x"79",x"27",x"AF", -- 0x1580
    x"27",x"E0",x"27",x"0D",x"28",x"84",x"28",x"A9", -- 0x1588
    x"28",x"B7",x"28",x"D2",x"28",x"DF",x"28",x"01", -- 0x1590
    x"29",x"10",x"29",x"79",x"29",x"93",x"29",x"B6", -- 0x1598
    x"29",x"C5",x"29",x"DF",x"29",x"F1",x"29",x"0A", -- 0x15A0
    x"2A",x"53",x"2A",x"CD",x"C1",x"15",x"3A",x"5F", -- 0x15A8
    x"42",x"0F",x"D8",x"21",x"09",x"40",x"35",x"C0", -- 0x15B0
    x"36",x"0A",x"2C",x"36",x"07",x"CD",x"23",x"17", -- 0x15B8
    x"C9",x"CD",x"D2",x"15",x"3A",x"90",x"42",x"EF", -- 0x15C0
    x"0B",x"16",x"32",x"16",x"8A",x"16",x"D9",x"16", -- 0x15C8
    x"F6",x"16",x"3A",x"5F",x"42",x"E6",x"07",x"C0", -- 0x15D0
    x"21",x"9B",x"42",x"7E",x"3C",x"FE",x"06",x"20", -- 0x15D8
    x"01",x"AF",x"77",x"21",x"1D",x"17",x"4F",x"06", -- 0x15E0
    x"00",x"09",x"7E",x"32",x"31",x"40",x"32",x"33", -- 0x15E8
    x"40",x"32",x"35",x"40",x"C9",x"21",x"4C",x"50", -- 0x15F0
    x"22",x"92",x"42",x"22",x"96",x"42",x"21",x"5E", -- 0x15F8
    x"50",x"22",x"94",x"42",x"21",x"AC",x"53",x"22", -- 0x1600
    x"98",x"42",x"C9",x"CD",x"00",x"12",x"CD",x"F5", -- 0x1608
    x"15",x"21",x"90",x"42",x"34",x"2C",x"36",x"32", -- 0x1610
    x"21",x"9A",x"42",x"36",x"07",x"2C",x"36",x"00", -- 0x1618
    x"2C",x"36",x"00",x"21",x"A0",x"58",x"CB",x"CE", -- 0x1620
    x"21",x"C0",x"58",x"CB",x"96",x"AF",x"32",x"B0", -- 0x1628
    x"58",x"C9",x"21",x"91",x"42",x"35",x"C0",x"36", -- 0x1630
    x"01",x"2D",x"34",x"21",x"39",x"40",x"D9",x"06", -- 0x1638
    x"00",x"3A",x"9C",x"42",x"4F",x"21",x"85",x"16", -- 0x1640
    x"09",x"7E",x"D9",x"06",x"13",x"77",x"2C",x"2C", -- 0x1648
    x"10",x"FB",x"3E",x"01",x"32",x"81",x"42",x"AF", -- 0x1650
    x"06",x"18",x"21",x"30",x"40",x"77",x"2C",x"2C", -- 0x1658
    x"10",x"FB",x"21",x"4C",x"50",x"0E",x"1C",x"06", -- 0x1660
    x"13",x"36",x"10",x"23",x"10",x"FB",x"11",x"0D", -- 0x1668
    x"00",x"19",x"0D",x"20",x"F2",x"11",x"00",x"06", -- 0x1670
    x"FF",x"3A",x"0D",x"40",x"1E",x"02",x"0F",x"D2", -- 0x1678
    x"38",x"00",x"1C",x"FF",x"C9",x"06",x"02",x"03", -- 0x1680
    x"07",x"00",x"21",x"91",x"42",x"35",x"C0",x"36", -- 0x1688
    x"03",x"06",x"13",x"3E",x"C8",x"2A",x"96",x"42", -- 0x1690
    x"ED",x"5B",x"98",x"42",x"77",x"12",x"13",x"23", -- 0x1698
    x"10",x"FA",x"06",x"28",x"2A",x"92",x"42",x"11", -- 0x16A0
    x"20",x"00",x"77",x"19",x"10",x"FC",x"2A",x"94", -- 0x16A8
    x"42",x"06",x"1C",x"77",x"19",x"10",x"FC",x"21", -- 0x16B0
    x"92",x"42",x"34",x"2C",x"2C",x"35",x"2A",x"96", -- 0x16B8
    x"42",x"19",x"22",x"96",x"42",x"2A",x"98",x"42", -- 0x16C0
    x"11",x"E0",x"FF",x"19",x"22",x"98",x"42",x"21", -- 0x16C8
    x"9A",x"42",x"35",x"C0",x"21",x"90",x"42",x"34", -- 0x16D0
    x"C9",x"CD",x"F5",x"15",x"21",x"90",x"42",x"36", -- 0x16D8
    x"01",x"2C",x"36",x"0A",x"21",x"9A",x"42",x"36", -- 0x16E0
    x"07",x"2C",x"2C",x"34",x"7E",x"FE",x"05",x"C0", -- 0x16E8
    x"3E",x"04",x"32",x"90",x"42",x"C9",x"3A",x"5F", -- 0x16F0
    x"42",x"E6",x"07",x"C0",x"3A",x"9B",x"42",x"2E", -- 0x16F8
    x"13",x"11",x"39",x"40",x"06",x"00",x"D6",x"01", -- 0x1700
    x"30",x"02",x"3E",x"05",x"4F",x"E5",x"F5",x"21", -- 0x1708
    x"1D",x"17",x"09",x"7E",x"12",x"1C",x"1C",x"F1", -- 0x1710
    x"E1",x"2D",x"20",x"EA",x"C9",x"00",x"03",x"02", -- 0x1718
    x"06",x"07",x"04",x"11",x"FD",x"FF",x"DD",x"21", -- 0x1720
    x"A4",x"40",x"3A",x"0D",x"40",x"0F",x"30",x"04", -- 0x1728
    x"DD",x"21",x"A7",x"40",x"FD",x"21",x"CE",x"43", -- 0x1730
    x"06",x"05",x"FD",x"7E",x"00",x"DD",x"BE",x"00", -- 0x1738
    x"20",x"0F",x"FD",x"7E",x"FF",x"DD",x"BE",x"FF", -- 0x1740
    x"20",x"07",x"FD",x"7E",x"FE",x"DD",x"BE",x"FE", -- 0x1748
    x"C8",x"30",x"04",x"FD",x"19",x"10",x"E3",x"3E", -- 0x1750
    x"05",x"90",x"C8",x"21",x"CE",x"43",x"11",x"D1", -- 0x1758
    x"43",x"47",x"87",x"80",x"06",x"00",x"4F",x"ED", -- 0x1760
    x"B8",x"2C",x"EB",x"DD",x"E5",x"E1",x"2D",x"2D", -- 0x1768
    x"01",x"03",x"00",x"ED",x"B0",x"C9",x"3A",x"1E", -- 0x1770
    x"41",x"0F",x"D8",x"21",x"A4",x"40",x"3A",x"0D", -- 0x1778
    x"40",x"0F",x"30",x"03",x"21",x"A7",x"40",x"3A", -- 0x1780
    x"17",x"40",x"47",x"7E",x"E6",x"0F",x"07",x"07", -- 0x1788
    x"07",x"07",x"4F",x"2D",x"7E",x"E6",x"F0",x"0F", -- 0x1790
    x"0F",x"0F",x"0F",x"B1",x"B8",x"D8",x"21",x"90", -- 0x1798
    x"58",x"CB",x"C6",x"21",x"1D",x"41",x"34",x"11", -- 0x17A0
    x"03",x"07",x"FF",x"2C",x"36",x"01",x"C9",x"3A", -- 0x17A8
    x"16",x"41",x"A7",x"C0",x"21",x"1C",x"41",x"7E", -- 0x17B0
    x"0F",x"D2",x"E0",x"1C",x"11",x"88",x"06",x"FF", -- 0x17B8
    x"36",x"00",x"C3",x"E0",x"1C",x"21",x"00",x"42", -- 0x17C0
    x"CB",x"46",x"28",x"3A",x"2C",x"2C",x"3A",x"0F", -- 0x17C8
    x"40",x"0F",x"30",x"06",x"3A",x"0D",x"40",x"0F", -- 0x17D0
    x"38",x"3F",x"3A",x"10",x"40",x"47",x"CB",x"5F", -- 0x17D8
    x"28",x"07",x"7E",x"FE",x"17",x"38",x"02",x"35", -- 0x17E0
    x"35",x"CB",x"50",x"28",x"07",x"7E",x"FE",x"E9", -- 0x17E8
    x"30",x"02",x"34",x"34",x"7E",x"2F",x"C6",x"80", -- 0x17F0
    x"0E",x"06",x"21",x"50",x"40",x"06",x"04",x"77", -- 0x17F8
    x"2C",x"71",x"2C",x"10",x"FA",x"C9",x"2C",x"CB", -- 0x1800
    x"46",x"20",x"05",x"2C",x"36",x"00",x"18",x"E4", -- 0x1808
    x"2C",x"7E",x"2F",x"C6",x"80",x"0E",x"07",x"18", -- 0x1810
    x"E1",x"3A",x"11",x"40",x"47",x"18",x"BE",x"21", -- 0x1818
    x"7C",x"42",x"CB",x"46",x"23",x"23",x"23",x"28", -- 0x1820
    x"0C",x"7E",x"D6",x"05",x"77",x"FE",x"34",x"30", -- 0x1828
    x"16",x"AF",x"32",x"7C",x"42",x"36",x"C7",x"2D", -- 0x1830
    x"2D",x"3A",x"00",x"42",x"0F",x"30",x"06",x"3A", -- 0x1838
    x"02",x"42",x"77",x"18",x"02",x"36",x"00",x"DD", -- 0x1840
    x"21",x"9D",x"40",x"FD",x"21",x"7D",x"42",x"3A", -- 0x1848
    x"0F",x"40",x"0F",x"30",x"17",x"3A",x"0D",x"40", -- 0x1850
    x"0F",x"30",x"11",x"FD",x"7E",x"02",x"2F",x"C6", -- 0x1858
    x"FC",x"DD",x"77",x"02",x"FD",x"7E",x"00",x"2F", -- 0x1860
    x"DD",x"77",x"00",x"C9",x"FD",x"7E",x"02",x"3D", -- 0x1868
    x"DD",x"77",x"02",x"FD",x"7E",x"00",x"2F",x"DD", -- 0x1870
    x"77",x"00",x"C9",x"DD",x"21",x"A0",x"42",x"11", -- 0x1878
    x"20",x"00",x"06",x"08",x"D9",x"CD",x"1D",x"1D", -- 0x1880
    x"D9",x"DD",x"19",x"10",x"F7",x"C9",x"DD",x"21", -- 0x1888
    x"A0",x"42",x"FD",x"21",x"60",x"40",x"01",x"08", -- 0x1890
    x"08",x"DD",x"CB",x"00",x"46",x"28",x"27",x"DD", -- 0x1898
    x"7E",x"16",x"FD",x"77",x"02",x"DD",x"7E",x"03", -- 0x18A0
    x"91",x"FD",x"77",x"03",x"DD",x"7E",x"04",x"2F", -- 0x18A8
    x"91",x"FD",x"77",x"00",x"DD",x"7E",x"12",x"FD", -- 0x18B0
    x"77",x"01",x"11",x"20",x"00",x"DD",x"19",x"1E", -- 0x18B8
    x"04",x"FD",x"19",x"10",x"D4",x"C9",x"DD",x"CB", -- 0x18C0
    x"01",x"46",x"28",x"06",x"FD",x"36",x"02",x"07", -- 0x18C8
    x"18",x"CD",x"FD",x"36",x"03",x"F8",x"FD",x"36", -- 0x18D0
    x"00",x"F8",x"18",x"DE",x"3A",x"00",x"42",x"0F", -- 0x18D8
    x"D0",x"3A",x"7C",x"42",x"0F",x"D8",x"3A",x"0F", -- 0x18E0
    x"40",x"0F",x"30",x"06",x"3A",x"0D",x"40",x"0F", -- 0x18E8
    x"38",x"17",x"3A",x"13",x"40",x"2F",x"47",x"3A", -- 0x18F0
    x"10",x"40",x"A0",x"E6",x"10",x"C8",x"3E",x"01", -- 0x18F8
    x"32",x"7C",x"42",x"21",x"C0",x"58",x"CB",x"C6", -- 0x1900
    x"C9",x"3A",x"14",x"40",x"2F",x"47",x"3A",x"11", -- 0x1908
    x"40",x"18",x"E7",x"CD",x"89",x"19",x"CD",x"DC", -- 0x1910
    x"19",x"CD",x"FB",x"19",x"CD",x"3E",x"1A",x"C3", -- 0x1918
    x"22",x"19",x"06",x"08",x"21",x"60",x"42",x"CB", -- 0x1920
    x"46",x"20",x"07",x"2C",x"2C",x"2C",x"2C",x"10", -- 0x1928
    x"F6",x"C9",x"2C",x"2C",x"2C",x"7E",x"C6",x"20", -- 0x1930
    x"D6",x"10",x"30",x"F2",x"2D",x"2D",x"7E",x"C6", -- 0x1938
    x"E0",x"D6",x"20",x"30",x"05",x"11",x"20",x"41", -- 0x1940
    x"18",x"14",x"D6",x"30",x"D6",x"20",x"30",x"05", -- 0x1948
    x"11",x"30",x"41",x"18",x"09",x"D6",x"30",x"D6", -- 0x1950
    x"20",x"30",x"D1",x"11",x"40",x"41",x"C6",x"20", -- 0x1958
    x"E6",x"F8",x"1F",x"83",x"5F",x"2C",x"2C",x"7E", -- 0x1960
    x"D6",x"E0",x"E6",x"0C",x"1F",x"1F",x"83",x"5F", -- 0x1968
    x"1A",x"CB",x"4F",x"28",x"B9",x"4F",x"7D",x"FE", -- 0x1970
    x"7C",x"79",x"30",x"03",x"CB",x"D7",x"12",x"0E", -- 0x1978
    x"04",x"AF",x"77",x"2D",x"0D",x"20",x"FB",x"18", -- 0x1980
    x"A2",x"DD",x"21",x"60",x"42",x"11",x"04",x"00", -- 0x1988
    x"06",x"04",x"CD",x"9A",x"19",x"DD",x"19",x"10", -- 0x1990
    x"F9",x"C9",x"DD",x"CB",x"00",x"46",x"28",x"2B", -- 0x1998
    x"DD",x"CB",x"02",x"4E",x"28",x"18",x"DD",x"34", -- 0x19A0
    x"01",x"DD",x"CB",x"02",x"46",x"28",x"0F",x"DD", -- 0x19A8
    x"35",x"01",x"DD",x"35",x"01",x"DD",x"7E",x"01", -- 0x19B0
    x"C6",x"10",x"D6",x"21",x"38",x"0D",x"DD",x"7E", -- 0x19B8
    x"03",x"C6",x"02",x"DD",x"77",x"03",x"FE",x"DF", -- 0x19C0
    x"30",x"01",x"C9",x"DD",x"36",x"00",x"00",x"DD", -- 0x19C8
    x"36",x"01",x"00",x"DD",x"36",x"02",x"00",x"DD", -- 0x19D0
    x"36",x"03",x"00",x"C9",x"DD",x"21",x"68",x"42", -- 0x19D8
    x"DD",x"CB",x"00",x"46",x"28",x"E5",x"3A",x"10", -- 0x19E0
    x"41",x"FE",x"05",x"30",x"03",x"AF",x"18",x"02", -- 0x19E8
    x"3E",x"02",x"DD",x"86",x"03",x"DD",x"77",x"03", -- 0x19F0
    x"C3",x"C6",x"19",x"DD",x"21",x"60",x"42",x"11", -- 0x19F8
    x"04",x"00",x"06",x"03",x"CD",x"0C",x"1A",x"DD", -- 0x1A00
    x"19",x"10",x"F9",x"C9",x"DD",x"CB",x"00",x"46", -- 0x1A08
    x"C8",x"DD",x"7E",x"03",x"C6",x"37",x"D6",x"05", -- 0x1A10
    x"38",x"17",x"D6",x"09",x"D0",x"3A",x"02",x"42", -- 0x1A18
    x"DD",x"96",x"01",x"C6",x"06",x"D6",x"0D",x"D0", -- 0x1A20
    x"CD",x"CB",x"19",x"3E",x"01",x"32",x"04",x"42", -- 0x1A28
    x"C9",x"3A",x"02",x"42",x"DD",x"96",x"01",x"C6", -- 0x1A30
    x"02",x"D6",x"05",x"D0",x"18",x"EA",x"21",x"81", -- 0x1A38
    x"40",x"11",x"61",x"42",x"06",x"03",x"1A",x"2F", -- 0x1A40
    x"77",x"2C",x"2C",x"1C",x"1C",x"1A",x"77",x"3A", -- 0x1A48
    x"0F",x"40",x"0F",x"30",x"09",x"3A",x"0D",x"40", -- 0x1A50
    x"0F",x"30",x"03",x"7E",x"2F",x"77",x"2C",x"2C", -- 0x1A58
    x"1C",x"1C",x"10",x"E2",x"C9",x"3A",x"7C",x"42", -- 0x1A60
    x"0F",x"D0",x"DD",x"21",x"A0",x"42",x"11",x"20", -- 0x1A68
    x"00",x"06",x"08",x"D9",x"CD",x"7D",x"1A",x"D9", -- 0x1A70
    x"DD",x"19",x"10",x"F7",x"C9",x"DD",x"CB",x"00", -- 0x1A78
    x"46",x"C8",x"3A",x"7F",x"42",x"6F",x"3A",x"7D", -- 0x1A80
    x"42",x"67",x"DD",x"7E",x"03",x"95",x"C6",x"02", -- 0x1A88
    x"FE",x"06",x"D0",x"DD",x"7E",x"04",x"94",x"C6", -- 0x1A90
    x"05",x"FE",x"0C",x"D0",x"DD",x"36",x"00",x"00", -- 0x1A98
    x"DD",x"36",x"01",x"01",x"DD",x"36",x"02",x"00", -- 0x1AA0
    x"3A",x"06",x"40",x"0F",x"30",x"34",x"DD",x"CB", -- 0x1AA8
    x"19",x"46",x"28",x"07",x"21",x"B0",x"58",x"CB", -- 0x1AB0
    x"D6",x"18",x"05",x"21",x"B0",x"58",x"CB",x"DE", -- 0x1AB8
    x"16",x"03",x"DD",x"7E",x"16",x"FE",x"07",x"28", -- 0x1AC0
    x"06",x"FE",x"03",x"28",x"06",x"18",x"08",x"1E", -- 0x1AC8
    x"02",x"18",x"06",x"1E",x"04",x"18",x"02",x"1E", -- 0x1AD0
    x"09",x"DD",x"7E",x"19",x"0F",x"30",x"02",x"CB", -- 0x1AD8
    x"23",x"FF",x"AF",x"32",x"7C",x"42",x"21",x"11", -- 0x1AE0
    x"41",x"35",x"DD",x"7E",x"18",x"DD",x"36",x"18", -- 0x1AE8
    x"00",x"3D",x"28",x"04",x"3D",x"28",x"0C",x"C9", -- 0x1AF0
    x"DD",x"7E",x"17",x"C6",x"20",x"6F",x"26",x"41", -- 0x1AF8
    x"CB",x"BE",x"C9",x"DD",x"7E",x"17",x"C6",x"50", -- 0x1B00
    x"18",x"F3",x"21",x"04",x"42",x"CB",x"46",x"28", -- 0x1B08
    x"18",x"36",x"00",x"21",x"00",x"01",x"22",x"00", -- 0x1B10
    x"42",x"21",x"0A",x"04",x"22",x"05",x"42",x"11", -- 0x1B18
    x"03",x"02",x"FF",x"21",x"C0",x"58",x"CB",x"CE", -- 0x1B20
    x"C9",x"3A",x"01",x"42",x"0F",x"D0",x"21",x"05", -- 0x1B28
    x"42",x"35",x"C0",x"36",x"0A",x"23",x"16",x"02", -- 0x1B30
    x"5E",x"FF",x"35",x"C0",x"AF",x"32",x"01",x"42", -- 0x1B38
    x"C9",x"3A",x"12",x"41",x"FE",x"2E",x"C8",x"3A", -- 0x1B40
    x"00",x"42",x"0F",x"D0",x"3A",x"16",x"41",x"A7", -- 0x1B48
    x"C8",x"3A",x"5F",x"42",x"E6",x"07",x"C0",x"3A", -- 0x1B50
    x"5F",x"42",x"A7",x"20",x"0E",x"2A",x"07",x"42", -- 0x1B58
    x"23",x"7E",x"3C",x"20",x"03",x"21",x"89",x"1B", -- 0x1B60
    x"22",x"07",x"42",x"2A",x"07",x"42",x"46",x"21", -- 0x1B68
    x"A0",x"42",x"11",x"1F",x"00",x"7E",x"23",x"B6", -- 0x1B70
    x"0F",x"30",x"04",x"19",x"10",x"F7",x"C9",x"23", -- 0x1B78
    x"36",x"00",x"2B",x"36",x"00",x"2B",x"36",x"01", -- 0x1B80
    x"C9",x"08",x"08",x"04",x"04",x"04",x"05",x"05", -- 0x1B88
    x"05",x"06",x"06",x"06",x"07",x"07",x"07",x"08", -- 0x1B90
    x"08",x"08",x"08",x"08",x"08",x"04",x"04",x"04", -- 0x1B98
    x"04",x"FF",x"3A",x"10",x"41",x"FE",x"04",x"D8", -- 0x1BA0
    x"3A",x"11",x"41",x"FE",x"0F",x"D8",x"3A",x"00", -- 0x1BA8
    x"42",x"0F",x"D0",x"21",x"B8",x"42",x"11",x"20", -- 0x1BB0
    x"00",x"06",x"08",x"CB",x"46",x"20",x"04",x"19", -- 0x1BB8
    x"10",x"F9",x"C9",x"7D",x"D6",x"15",x"6F",x"3A", -- 0x1BC0
    x"60",x"42",x"0F",x"D8",x"7E",x"2C",x"46",x"FE", -- 0x1BC8
    x"B0",x"D0",x"FE",x"60",x"D8",x"21",x"60",x"42", -- 0x1BD0
    x"36",x"01",x"2C",x"70",x"2C",x"2C",x"77",x"C9", -- 0x1BD8
    x"3A",x"00",x"42",x"0F",x"D0",x"3A",x"10",x"41", -- 0x1BE0
    x"A7",x"C8",x"3A",x"11",x"41",x"FE",x"0F",x"D8", -- 0x1BE8
    x"3A",x"02",x"42",x"4F",x"26",x"FF",x"2E",x"00", -- 0x1BF0
    x"DD",x"21",x"A0",x"42",x"11",x"20",x"00",x"06", -- 0x1BF8
    x"08",x"DD",x"CB",x"00",x"46",x"28",x"12",x"DD", -- 0x1C00
    x"7E",x"04",x"B9",x"30",x"06",x"79",x"DD",x"96", -- 0x1C08
    x"04",x"18",x"01",x"91",x"BC",x"30",x"02",x"67", -- 0x1C10
    x"68",x"DD",x"19",x"10",x"E4",x"7D",x"A7",x"C8", -- 0x1C18
    x"3E",x"08",x"95",x"21",x"A0",x"42",x"A7",x"28", -- 0x1C20
    x"04",x"3D",x"19",x"18",x"F9",x"2C",x"2C",x"2C", -- 0x1C28
    x"DD",x"21",x"64",x"42",x"DD",x"CB",x"00",x"46", -- 0x1C30
    x"C0",x"7E",x"FE",x"60",x"D8",x"47",x"3A",x"10", -- 0x1C38
    x"41",x"0E",x"A8",x"A7",x"28",x"07",x"0E",x"B0", -- 0x1C40
    x"3D",x"28",x"02",x"0E",x"B8",x"78",x"B9",x"D0", -- 0x1C48
    x"DD",x"36",x"00",x"01",x"7E",x"DD",x"77",x"03", -- 0x1C50
    x"2C",x"7E",x"DD",x"77",x"01",x"C9",x"3A",x"00", -- 0x1C58
    x"42",x"0F",x"D0",x"3A",x"11",x"41",x"FE",x"0F", -- 0x1C60
    x"D8",x"3A",x"00",x"41",x"0F",x"D0",x"3A",x"10", -- 0x1C68
    x"41",x"FE",x"02",x"D8",x"21",x"68",x"42",x"CB", -- 0x1C70
    x"46",x"C0",x"34",x"2C",x"3A",x"01",x"41",x"77", -- 0x1C78
    x"2C",x"2C",x"36",x"38",x"C9",x"21",x"DF",x"41", -- 0x1C80
    x"1E",x"06",x"0E",x"06",x"06",x"18",x"CB",x"4E", -- 0x1C88
    x"20",x"0C",x"7D",x"93",x"6F",x"10",x"F7",x"7D", -- 0x1C90
    x"C6",x"8F",x"6F",x"0D",x"20",x"EE",x"3E",x"40", -- 0x1C98
    x"41",x"0E",x"04",x"04",x"81",x"10",x"FD",x"32", -- 0x1CA0
    x"1B",x"41",x"C9",x"3A",x"00",x"41",x"A7",x"C8", -- 0x1CA8
    x"3A",x"5F",x"42",x"E6",x"01",x"C8",x"21",x"02", -- 0x1CB0
    x"41",x"7E",x"2D",x"0F",x"38",x"12",x"7E",x"FE", -- 0x1CB8
    x"27",x"38",x"15",x"3D",x"77",x"2F",x"C6",x"80", -- 0x1CC0
    x"21",x"2A",x"40",x"77",x"2C",x"2C",x"77",x"C9", -- 0x1CC8
    x"7E",x"FE",x"D9",x"30",x"07",x"3C",x"18",x"EC", -- 0x1CD0
    x"2C",x"36",x"01",x"C9",x"2C",x"36",x"00",x"C9", -- 0x1CD8
    x"3A",x"58",x"40",x"A7",x"20",x"0E",x"3E",x"30", -- 0x1CE0
    x"32",x"58",x"40",x"32",x"5A",x"40",x"21",x"20", -- 0x1CE8
    x"41",x"C3",x"14",x"1D",x"21",x"58",x"40",x"34", -- 0x1CF0
    x"23",x"23",x"34",x"7E",x"FE",x"80",x"21",x"30", -- 0x1CF8
    x"41",x"CA",x"14",x"1D",x"FE",x"D0",x"21",x"40", -- 0x1D00
    x"41",x"CA",x"14",x"1D",x"A7",x"C0",x"21",x"16", -- 0x1D08
    x"41",x"36",x"30",x"C9",x"06",x"10",x"3E",x"02", -- 0x1D10
    x"77",x"23",x"10",x"FC",x"C9",x"DD",x"CB",x"01", -- 0x1D18
    x"46",x"C2",x"61",x"1D",x"DD",x"CB",x"00",x"46", -- 0x1D20
    x"C8",x"DD",x"7E",x"02",x"EF",x"BD",x"1F",x"76", -- 0x1D28
    x"21",x"A5",x"21",x"B7",x"21",x"C1",x"21",x"EE", -- 0x1D30
    x"21",x"12",x"22",x"1C",x"22",x"2B",x"22",x"A9", -- 0x1D38
    x"23",x"B3",x"23",x"C1",x"23",x"CB",x"23",x"FA", -- 0x1D40
    x"23",x"04",x"24",x"0E",x"24",x"18",x"24",x"25", -- 0x1D48
    x"24",x"28",x"24",x"32",x"24",x"41",x"24",x"F2", -- 0x1D50
    x"25",x"FC",x"25",x"0A",x"26",x"14",x"26",x"43", -- 0x1D58
    x"26",x"DD",x"7E",x"02",x"EF",x"69",x"1D",x"79", -- 0x1D60
    x"1D",x"DD",x"36",x"10",x"04",x"DD",x"36",x"11", -- 0x1D68
    x"04",x"DD",x"36",x"12",x"1C",x"DD",x"34",x"02", -- 0x1D70
    x"C9",x"DD",x"35",x"10",x"C0",x"DD",x"36",x"10", -- 0x1D78
    x"04",x"DD",x"34",x"12",x"DD",x"35",x"11",x"C0", -- 0x1D80
    x"DD",x"36",x"01",x"00",x"C9",x"DD",x"7E",x"16", -- 0x1D88
    x"FE",x"01",x"F5",x"CC",x"AC",x"1D",x"F1",x"28", -- 0x1D90
    x"13",x"DD",x"CB",x"19",x"46",x"20",x"0D",x"DD", -- 0x1D98
    x"7E",x"16",x"FE",x"03",x"28",x"06",x"3A",x"5F", -- 0x1DA0
    x"42",x"0F",x"3F",x"D0",x"DD",x"7E",x"04",x"DD", -- 0x1DA8
    x"BE",x"06",x"28",x"4A",x"DD",x"7E",x"03",x"DD", -- 0x1DB0
    x"BE",x"05",x"28",x"58",x"DD",x"CB",x"09",x"46", -- 0x1DB8
    x"28",x"1E",x"DD",x"7E",x"07",x"DD",x"86",x"03", -- 0x1DC0
    x"DD",x"77",x"03",x"DD",x"7E",x"0B",x"DD",x"86", -- 0x1DC8
    x"0A",x"DD",x"77",x"0A",x"D0",x"DD",x"7E",x"08", -- 0x1DD0
    x"DD",x"86",x"04",x"DD",x"77",x"04",x"A7",x"C9", -- 0x1DD8
    x"DD",x"7E",x"08",x"DD",x"86",x"04",x"DD",x"77", -- 0x1DE0
    x"04",x"DD",x"7E",x"0B",x"DD",x"86",x"0A",x"DD", -- 0x1DE8
    x"77",x"0A",x"D0",x"DD",x"7E",x"07",x"DD",x"86", -- 0x1DF0
    x"03",x"DD",x"77",x"03",x"A7",x"C9",x"DD",x"7E", -- 0x1DF8
    x"03",x"DD",x"BE",x"05",x"28",x"0C",x"30",x"05", -- 0x1E00
    x"DD",x"34",x"03",x"A7",x"C9",x"DD",x"35",x"03", -- 0x1E08
    x"A7",x"C9",x"37",x"C9",x"DD",x"7E",x"04",x"DD", -- 0x1E10
    x"BE",x"06",x"30",x"05",x"DD",x"34",x"04",x"A7", -- 0x1E18
    x"C9",x"DD",x"35",x"04",x"A7",x"C9",x"DD",x"35", -- 0x1E20
    x"0E",x"C0",x"DD",x"6E",x"0C",x"DD",x"66",x"0D", -- 0x1E28
    x"7E",x"FE",x"FF",x"20",x"06",x"23",x"5E",x"23", -- 0x1E30
    x"56",x"EB",x"7E",x"DD",x"77",x"12",x"23",x"7E", -- 0x1E38
    x"DD",x"77",x"0E",x"23",x"DD",x"75",x"0C",x"DD", -- 0x1E40
    x"74",x"0D",x"C9",x"8E",x"0A",x"8F",x"0A",x"90", -- 0x1E48
    x"0A",x"91",x"0A",x"92",x"0A",x"F1",x"05",x"F0", -- 0x1E50
    x"05",x"EF",x"05",x"EE",x"05",x"ED",x"05",x"FF", -- 0x1E58
    x"79",x"1E",x"0E",x"0A",x"0F",x"0A",x"10",x"0A", -- 0x1E60
    x"11",x"0A",x"12",x"0A",x"71",x"05",x"70",x"05", -- 0x1E68
    x"6F",x"05",x"6E",x"05",x"6D",x"05",x"FF",x"79", -- 0x1E70
    x"1E",x"E9",x"05",x"EA",x"05",x"EB",x"05",x"EC", -- 0x1E78
    x"05",x"FF",x"79",x"1E",x"6E",x"05",x"6F",x"05", -- 0x1E80
    x"6E",x"05",x"6D",x"05",x"E9",x"05",x"EA",x"05", -- 0x1E88
    x"EB",x"05",x"EC",x"05",x"ED",x"05",x"EE",x"05", -- 0x1E90
    x"EF",x"05",x"EE",x"05",x"ED",x"05",x"FF",x"79", -- 0x1E98
    x"1E",x"E4",x"03",x"E5",x"03",x"E6",x"03",x"E7", -- 0x1EA0
    x"03",x"E8",x"03",x"A7",x"03",x"A6",x"03",x"A5", -- 0x1EA8
    x"03",x"A4",x"03",x"FF",x"B6",x"1E",x"20",x"05", -- 0x1EB0
    x"21",x"05",x"22",x"05",x"23",x"05",x"FF",x"B6", -- 0x1EB8
    x"1E",x"25",x"05",x"26",x"05",x"25",x"05",x"24", -- 0x1EC0
    x"05",x"20",x"05",x"21",x"05",x"22",x"05",x"23", -- 0x1EC8
    x"05",x"A4",x"05",x"A5",x"05",x"A6",x"05",x"A5", -- 0x1ED0
    x"05",x"A4",x"05",x"FF",x"B6",x"1E",x"2D",x"03", -- 0x1ED8
    x"2E",x"03",x"2F",x"03",x"30",x"03",x"31",x"03", -- 0x1EE0
    x"70",x"03",x"6F",x"03",x"6E",x"03",x"6D",x"03", -- 0x1EE8
    x"FF",x"79",x"1E",x"DD",x"E5",x"E1",x"3E",x"07", -- 0x1EF0
    x"85",x"6F",x"DD",x"36",x"0A",x"00",x"DD",x"7E", -- 0x1EF8
    x"05",x"DD",x"BE",x"03",x"28",x"04",x"38",x"1E", -- 0x1F00
    x"18",x"56",x"DD",x"7E",x"06",x"DD",x"BE",x"04", -- 0x1F08
    x"28",x"0E",x"38",x"06",x"36",x"00",x"2C",x"36", -- 0x1F10
    x"01",x"C9",x"36",x"00",x"2C",x"36",x"FF",x"C9", -- 0x1F18
    x"36",x"00",x"2C",x"36",x"00",x"C9",x"DD",x"7E", -- 0x1F20
    x"06",x"DD",x"BE",x"04",x"28",x"2C",x"38",x"15", -- 0x1F28
    x"36",x"FF",x"2C",x"36",x"01",x"DD",x"7E",x"03", -- 0x1F30
    x"DD",x"96",x"05",x"47",x"DD",x"7E",x"06",x"DD", -- 0x1F38
    x"96",x"04",x"4F",x"18",x"55",x"36",x"FF",x"2C", -- 0x1F40
    x"36",x"FF",x"DD",x"7E",x"03",x"DD",x"96",x"05", -- 0x1F48
    x"47",x"DD",x"7E",x"04",x"DD",x"96",x"06",x"4F", -- 0x1F50
    x"18",x"40",x"36",x"FF",x"2C",x"36",x"00",x"C9", -- 0x1F58
    x"DD",x"7E",x"06",x"DD",x"BE",x"04",x"28",x"2C", -- 0x1F60
    x"38",x"15",x"36",x"01",x"2C",x"36",x"01",x"DD", -- 0x1F68
    x"7E",x"05",x"DD",x"96",x"03",x"47",x"DD",x"7E", -- 0x1F70
    x"06",x"DD",x"96",x"04",x"4F",x"18",x"1B",x"36", -- 0x1F78
    x"01",x"2C",x"36",x"FF",x"DD",x"7E",x"05",x"DD", -- 0x1F80
    x"96",x"03",x"47",x"DD",x"7E",x"04",x"DD",x"96", -- 0x1F88
    x"06",x"4F",x"18",x"06",x"36",x"01",x"2C",x"36", -- 0x1F90
    x"00",x"C9",x"79",x"B8",x"28",x"16",x"38",x"0B", -- 0x1F98
    x"DD",x"36",x"09",x"00",x"CD",x"4F",x"26",x"DD", -- 0x1FA0
    x"77",x"0B",x"C9",x"DD",x"36",x"09",x"01",x"78", -- 0x1FA8
    x"41",x"4F",x"18",x"F0",x"DD",x"36",x"09",x"01", -- 0x1FB0
    x"DD",x"36",x"0B",x"FF",x"C9",x"DD",x"36",x"18", -- 0x1FB8
    x"00",x"DD",x"36",x"19",x"00",x"21",x"0E",x"21", -- 0x1FC0
    x"DD",x"75",x"13",x"DD",x"74",x"14",x"DD",x"36", -- 0x1FC8
    x"10",x"30",x"DD",x"36",x"0E",x"01",x"21",x"12", -- 0x1FD0
    x"41",x"7E",x"34",x"47",x"87",x"87",x"80",x"5F", -- 0x1FD8
    x"16",x"00",x"21",x"28",x"20",x"19",x"3E",x"30", -- 0x1FE0
    x"86",x"DD",x"77",x"03",x"23",x"3A",x"01",x"41", -- 0x1FE8
    x"86",x"DD",x"77",x"04",x"23",x"5E",x"23",x"46", -- 0x1FF0
    x"23",x"7E",x"DD",x"77",x"16",x"21",x"04",x"41", -- 0x1FF8
    x"19",x"70",x"DD",x"36",x"12",x"0B",x"3A",x"01", -- 0x2000
    x"41",x"FE",x"80",x"30",x"11",x"DD",x"36",x"15", -- 0x2008
    x"00",x"21",x"4B",x"1E",x"DD",x"75",x"0C",x"DD", -- 0x2010
    x"74",x"0D",x"DD",x"34",x"02",x"C9",x"DD",x"36", -- 0x2018
    x"15",x"01",x"21",x"62",x"1E",x"C3",x"14",x"20", -- 0x2020
    x"F1",x"EF",x"00",x"66",x"07",x"F1",x"12",x"05", -- 0x2028
    x"66",x"07",x"F3",x"EB",x"00",x"6D",x"07",x"F3", -- 0x2030
    x"16",x"05",x"67",x"07",x"F3",x"EE",x"00",x"68", -- 0x2038
    x"07",x"F3",x"13",x"05",x"68",x"07",x"F5",x"EA", -- 0x2040
    x"00",x"6E",x"07",x"F5",x"17",x"05",x"69",x"07", -- 0x2048
    x"F5",x"EF",x"00",x"6A",x"07",x"F5",x"12",x"05", -- 0x2050
    x"6A",x"07",x"F7",x"EB",x"00",x"6F",x"07",x"F7", -- 0x2058
    x"16",x"05",x"6B",x"03",x"F7",x"EE",x"00",x"10", -- 0x2060
    x"03",x"F7",x"13",x"05",x"10",x"03",x"F1",x"F2", -- 0x2068
    x"01",x"6C",x"03",x"F1",x"0F",x"04",x"65",x"03", -- 0x2070
    x"F1",x"F7",x"01",x"66",x"03",x"F1",x"0A",x"04", -- 0x2078
    x"66",x"03",x"F3",x"F3",x"01",x"6D",x"03",x"F3", -- 0x2080
    x"0E",x"04",x"67",x"03",x"F3",x"F6",x"01",x"68", -- 0x2088
    x"03",x"F3",x"0B",x"04",x"68",x"03",x"F5",x"F2", -- 0x2090
    x"01",x"6E",x"03",x"F5",x"0F",x"04",x"69",x"03", -- 0x2098
    x"F5",x"F7",x"01",x"6A",x"03",x"F5",x"0A",x"04", -- 0x20A0
    x"6A",x"03",x"F7",x"F3",x"01",x"6F",x"03",x"F7", -- 0x20A8
    x"0E",x"04",x"6B",x"03",x"F7",x"F6",x"01",x"10", -- 0x20B0
    x"03",x"F7",x"0B",x"04",x"10",x"03",x"F1",x"FA", -- 0x20B8
    x"02",x"6C",x"03",x"F1",x"07",x"03",x"65",x"03", -- 0x20C0
    x"F1",x"FF",x"02",x"66",x"03",x"F1",x"02",x"03", -- 0x20C8
    x"66",x"03",x"F3",x"FB",x"02",x"6D",x"03",x"F3", -- 0x20D0
    x"06",x"03",x"67",x"03",x"F3",x"FE",x"02",x"68", -- 0x20D8
    x"03",x"F3",x"03",x"03",x"68",x"01",x"F5",x"FA", -- 0x20E0
    x"02",x"6E",x"01",x"F5",x"07",x"03",x"69",x"01", -- 0x20E8
    x"F5",x"FF",x"02",x"6A",x"01",x"F5",x"02",x"03", -- 0x20F0
    x"6A",x"01",x"F7",x"FB",x"02",x"6F",x"01",x"F7", -- 0x20F8
    x"06",x"03",x"6B",x"01",x"F7",x"FE",x"02",x"10", -- 0x2100
    x"01",x"F7",x"03",x"03",x"10",x"01",x"FF",x"00", -- 0x2108
    x"FF",x"00",x"FF",x"00",x"FF",x"01",x"FF",x"00", -- 0x2110
    x"FF",x"00",x"FF",x"01",x"FF",x"00",x"FF",x"01", -- 0x2118
    x"FF",x"00",x"00",x"01",x"FF",x"00",x"FF",x"01", -- 0x2120
    x"00",x"01",x"FF",x"00",x"00",x"01",x"FF",x"01", -- 0x2128
    x"00",x"01",x"FF",x"01",x"00",x"01",x"00",x"01", -- 0x2130
    x"FF",x"01",x"00",x"01",x"00",x"01",x"00",x"01", -- 0x2138
    x"00",x"01",x"00",x"01",x"00",x"01",x"01",x"01", -- 0x2140
    x"00",x"01",x"00",x"01",x"01",x"01",x"00",x"01", -- 0x2148
    x"01",x"01",x"00",x"01",x"01",x"00",x"00",x"01", -- 0x2150
    x"01",x"01",x"01",x"00",x"00",x"01",x"01",x"00", -- 0x2158
    x"01",x"01",x"01",x"00",x"01",x"01",x"01",x"00", -- 0x2160
    x"01",x"00",x"01",x"01",x"01",x"00",x"01",x"00", -- 0x2168
    x"01",x"00",x"01",x"00",x"01",x"00",x"DD",x"35", -- 0x2170
    x"10",x"28",x"27",x"DD",x"6E",x"13",x"DD",x"66", -- 0x2178
    x"14",x"DD",x"7E",x"03",x"86",x"DD",x"77",x"03", -- 0x2180
    x"23",x"7E",x"23",x"DD",x"75",x"13",x"DD",x"74", -- 0x2188
    x"14",x"DD",x"CB",x"15",x"46",x"28",x"02",x"ED", -- 0x2190
    x"44",x"DD",x"86",x"04",x"DD",x"77",x"04",x"C3", -- 0x2198
    x"26",x"1E",x"DD",x"34",x"02",x"3A",x"1B",x"41", -- 0x21A0
    x"DD",x"77",x"05",x"DD",x"7E",x"04",x"DD",x"77", -- 0x21A8
    x"06",x"CD",x"F3",x"1E",x"DD",x"34",x"02",x"CD", -- 0x21B0
    x"26",x"1E",x"CD",x"8D",x"1D",x"D0",x"DD",x"34", -- 0x21B8
    x"02",x"3A",x"1C",x"41",x"0F",x"3E",x"01",x"30", -- 0x21C0
    x"1F",x"3E",x"03",x"18",x"1B",x"3A",x"04",x"40", -- 0x21C8
    x"47",x"3A",x"10",x"41",x"A7",x"28",x"07",x"3D", -- 0x21D0
    x"28",x"0A",x"3E",x"01",x"18",x"0A",x"3E",x"03", -- 0x21D8
    x"A0",x"3C",x"18",x"04",x"3E",x"01",x"A0",x"3C", -- 0x21E0
    x"DD",x"77",x"10",x"DD",x"34",x"02",x"3A",x"04", -- 0x21E8
    x"40",x"47",x"E6",x"70",x"FE",x"60",x"38",x"02", -- 0x21F0
    x"D6",x"20",x"C6",x"58",x"DD",x"77",x"05",x"78", -- 0x21F8
    x"FE",x"D0",x"38",x"02",x"D6",x"80",x"C6",x"18", -- 0x2200
    x"DD",x"77",x"06",x"CD",x"F3",x"1E",x"DD",x"34", -- 0x2208
    x"02",x"C9",x"CD",x"26",x"1E",x"CD",x"8D",x"1D", -- 0x2210
    x"D0",x"DD",x"34",x"02",x"DD",x"35",x"10",x"28", -- 0x2218
    x"07",x"DD",x"35",x"02",x"DD",x"35",x"02",x"C9", -- 0x2220
    x"DD",x"34",x"02",x"DD",x"36",x"02",x"04",x"3A", -- 0x2228
    x"00",x"42",x"0F",x"D0",x"3A",x"16",x"41",x"A7", -- 0x2230
    x"C8",x"ED",x"5F",x"E6",x"03",x"28",x"13",x"3D", -- 0x2238
    x"28",x"44",x"3D",x"28",x"72",x"3A",x"02",x"42", -- 0x2240
    x"FE",x"58",x"38",x"6B",x"FE",x"A8",x"38",x"02", -- 0x2248
    x"18",x"34",x"21",x"20",x"41",x"CD",x"11",x"23", -- 0x2250
    x"DA",x"E8",x"22",x"21",x"2C",x"41",x"CD",x"2D", -- 0x2258
    x"23",x"DA",x"E8",x"22",x"21",x"30",x"41",x"CD", -- 0x2260
    x"11",x"23",x"DA",x"E8",x"22",x"21",x"3C",x"41", -- 0x2268
    x"CD",x"2D",x"23",x"38",x"73",x"21",x"40",x"41", -- 0x2270
    x"CD",x"11",x"23",x"38",x"6B",x"21",x"4C",x"41", -- 0x2278
    x"CD",x"2D",x"23",x"38",x"63",x"C9",x"21",x"3C", -- 0x2280
    x"41",x"CD",x"2D",x"23",x"38",x"5A",x"21",x"30", -- 0x2288
    x"41",x"CD",x"11",x"23",x"38",x"52",x"21",x"4C", -- 0x2290
    x"41",x"CD",x"2D",x"23",x"38",x"4A",x"21",x"40", -- 0x2298
    x"41",x"CD",x"11",x"23",x"38",x"42",x"21",x"20", -- 0x22A0
    x"41",x"CD",x"11",x"23",x"38",x"3A",x"21",x"2C", -- 0x22A8
    x"41",x"CD",x"2D",x"23",x"38",x"32",x"C9",x"21", -- 0x22B0
    x"40",x"41",x"CD",x"11",x"23",x"38",x"29",x"21", -- 0x22B8
    x"4C",x"41",x"CD",x"2D",x"23",x"38",x"21",x"21", -- 0x22C0
    x"20",x"41",x"CD",x"11",x"23",x"38",x"19",x"21", -- 0x22C8
    x"2C",x"41",x"CD",x"2D",x"23",x"38",x"11",x"21", -- 0x22D0
    x"30",x"41",x"CD",x"11",x"23",x"38",x"09",x"21", -- 0x22D8
    x"3C",x"41",x"CD",x"2D",x"23",x"38",x"01",x"C9", -- 0x22E0
    x"CB",x"FE",x"7D",x"D6",x"20",x"DD",x"77",x"17", -- 0x22E8
    x"DD",x"36",x"18",x"01",x"87",x"5F",x"16",x"00", -- 0x22F0
    x"21",x"49",x"23",x"19",x"7E",x"D6",x"10",x"DD", -- 0x22F8
    x"77",x"05",x"23",x"7E",x"DD",x"77",x"06",x"CD", -- 0x2300
    x"F3",x"1E",x"DD",x"36",x"02",x"09",x"C3",x"A9", -- 0x2308
    x"23",x"11",x"0F",x"04",x"4A",x"42",x"CB",x"4E", -- 0x2310
    x"20",x"0D",x"7D",x"82",x"6F",x"10",x"F7",x"7D", -- 0x2318
    x"93",x"6F",x"0D",x"20",x"F0",x"A7",x"C9",x"A7", -- 0x2320
    x"CB",x"7E",x"C0",x"37",x"C9",x"11",x"11",x"04", -- 0x2328
    x"4A",x"42",x"CB",x"4E",x"20",x"0D",x"7D",x"92", -- 0x2330
    x"6F",x"10",x"F7",x"7D",x"83",x"6F",x"0D",x"20", -- 0x2338
    x"F0",x"A7",x"C9",x"A7",x"CB",x"7E",x"C0",x"37", -- 0x2340
    x"C9",x"E0",x"24",x"E4",x"24",x"E8",x"24",x"EC", -- 0x2348
    x"24",x"E0",x"2C",x"E4",x"2C",x"E8",x"2C",x"EC", -- 0x2350
    x"2C",x"E0",x"34",x"E4",x"34",x"E8",x"34",x"EC", -- 0x2358
    x"34",x"E0",x"3C",x"E4",x"3C",x"E8",x"3C",x"EC", -- 0x2360
    x"3C",x"E0",x"74",x"E4",x"74",x"E8",x"74",x"EC", -- 0x2368
    x"74",x"E0",x"7C",x"E4",x"7C",x"E8",x"7C",x"EC", -- 0x2370
    x"7C",x"E0",x"84",x"E4",x"84",x"E8",x"84",x"EC", -- 0x2378
    x"84",x"E0",x"8C",x"E4",x"8C",x"E8",x"8C",x"EC", -- 0x2380
    x"8C",x"E0",x"C4",x"E4",x"C4",x"E8",x"C4",x"EC", -- 0x2388
    x"C4",x"E0",x"CC",x"E4",x"CC",x"E8",x"CC",x"EC", -- 0x2390
    x"CC",x"E0",x"D4",x"E4",x"D4",x"E8",x"D4",x"EC", -- 0x2398
    x"D4",x"E0",x"DC",x"E4",x"DC",x"E8",x"DC",x"EC", -- 0x23A0
    x"DC",x"CD",x"26",x"1E",x"CD",x"8D",x"1D",x"D0", -- 0x23A8
    x"DD",x"34",x"02",x"DD",x"7E",x"05",x"C6",x"10", -- 0x23B0
    x"DD",x"77",x"05",x"CD",x"F3",x"1E",x"DD",x"34", -- 0x23B8
    x"02",x"CD",x"26",x"1E",x"CD",x"8D",x"1D",x"D0", -- 0x23C0
    x"DD",x"34",x"02",x"21",x"B0",x"58",x"CB",x"CE", -- 0x23C8
    x"21",x"A1",x"1E",x"DD",x"75",x"0C",x"DD",x"74", -- 0x23D0
    x"0D",x"DD",x"36",x"0E",x"01",x"DD",x"36",x"10", -- 0x23D8
    x"0F",x"DD",x"36",x"18",x"00",x"DD",x"36",x"19", -- 0x23E0
    x"01",x"DD",x"7E",x"17",x"C6",x"20",x"6F",x"26", -- 0x23E8
    x"41",x"36",x"00",x"21",x"16",x"41",x"35",x"DD", -- 0x23F0
    x"34",x"02",x"CD",x"26",x"1E",x"DD",x"35",x"10", -- 0x23F8
    x"C0",x"DD",x"34",x"02",x"DD",x"36",x"05",x"B8", -- 0x2400
    x"CD",x"F3",x"1E",x"DD",x"34",x"02",x"CD",x"26", -- 0x2408
    x"1E",x"CD",x"8D",x"1D",x"D0",x"DD",x"34",x"02", -- 0x2410
    x"3A",x"04",x"40",x"E6",x"03",x"3E",x"01",x"DD", -- 0x2418
    x"77",x"10",x"DD",x"34",x"02",x"CD",x"EE",x"21", -- 0x2420
    x"CD",x"26",x"1E",x"CD",x"8D",x"1D",x"D0",x"DD", -- 0x2428
    x"34",x"02",x"DD",x"35",x"10",x"28",x"07",x"DD", -- 0x2430
    x"35",x"02",x"DD",x"35",x"02",x"C9",x"DD",x"34", -- 0x2438
    x"02",x"3A",x"04",x"40",x"E6",x"03",x"21",x"50", -- 0x2440
    x"41",x"3D",x"28",x"09",x"21",x"80",x"41",x"3D", -- 0x2448
    x"28",x"03",x"21",x"B0",x"41",x"CD",x"7D",x"24", -- 0x2450
    x"DD",x"36",x"02",x"10",x"D0",x"DD",x"6E",x"17", -- 0x2458
    x"26",x"00",x"29",x"EB",x"21",x"D2",x"24",x"19", -- 0x2460
    x"7E",x"C6",x"10",x"DD",x"77",x"05",x"23",x"7E", -- 0x2468
    x"DD",x"77",x"06",x"CD",x"F3",x"1E",x"DD",x"36", -- 0x2470
    x"02",x"15",x"C3",x"F2",x"25",x"08",x"3E",x"01", -- 0x2478
    x"08",x"16",x"06",x"ED",x"5F",x"E6",x"07",x"4F", -- 0x2480
    x"87",x"47",x"87",x"80",x"85",x"6F",x"1E",x"08", -- 0x2488
    x"7B",x"91",x"47",x"7E",x"CB",x"46",x"20",x"24", -- 0x2490
    x"7D",x"C6",x"06",x"6F",x"1D",x"10",x"F4",x"7B", -- 0x2498
    x"A7",x"28",x"0A",x"7D",x"D6",x"30",x"6F",x"43", -- 0x24A0
    x"08",x"AF",x"08",x"18",x"E6",x"08",x"A7",x"28", -- 0x24A8
    x"04",x"7D",x"D6",x"30",x"6F",x"08",x"2C",x"15", -- 0x24B0
    x"20",x"D4",x"A7",x"C9",x"CB",x"4E",x"20",x"D8", -- 0x24B8
    x"A7",x"CB",x"7E",x"C0",x"CB",x"FE",x"7D",x"D6", -- 0x24C0
    x"50",x"DD",x"77",x"17",x"DD",x"36",x"18",x"02", -- 0x24C8
    x"37",x"C9",x"44",x"1C",x"48",x"1C",x"4C",x"1C", -- 0x24D0
    x"50",x"1C",x"54",x"1C",x"58",x"1C",x"44",x"24", -- 0x24D8
    x"48",x"24",x"4C",x"24",x"50",x"24",x"54",x"24", -- 0x24E0
    x"58",x"24",x"44",x"2C",x"48",x"2C",x"4C",x"2C", -- 0x24E8
    x"50",x"2C",x"54",x"2C",x"58",x"2C",x"44",x"34", -- 0x24F0
    x"48",x"34",x"4C",x"34",x"50",x"34",x"54",x"34", -- 0x24F8
    x"58",x"34",x"44",x"3C",x"48",x"3C",x"4C",x"3C", -- 0x2500
    x"50",x"3C",x"54",x"3C",x"58",x"3C",x"44",x"44", -- 0x2508
    x"48",x"44",x"4C",x"44",x"50",x"44",x"54",x"44", -- 0x2510
    x"58",x"44",x"44",x"4C",x"48",x"4C",x"4C",x"4C", -- 0x2518
    x"50",x"4C",x"54",x"4C",x"58",x"4C",x"44",x"54", -- 0x2520
    x"48",x"54",x"4C",x"54",x"50",x"54",x"54",x"54", -- 0x2528
    x"58",x"54",x"44",x"64",x"48",x"64",x"4C",x"64", -- 0x2530
    x"50",x"64",x"54",x"64",x"58",x"64",x"44",x"6C", -- 0x2538
    x"48",x"6C",x"4C",x"6C",x"50",x"6C",x"54",x"6C", -- 0x2540
    x"58",x"6C",x"44",x"74",x"48",x"74",x"4C",x"74", -- 0x2548
    x"50",x"74",x"54",x"74",x"58",x"74",x"44",x"7C", -- 0x2550
    x"48",x"7C",x"4C",x"7C",x"50",x"7C",x"54",x"7C", -- 0x2558
    x"58",x"7C",x"44",x"84",x"48",x"84",x"4C",x"84", -- 0x2560
    x"50",x"84",x"54",x"84",x"58",x"84",x"44",x"8C", -- 0x2568
    x"48",x"8C",x"4C",x"8C",x"50",x"8C",x"54",x"8C", -- 0x2570
    x"58",x"8C",x"44",x"94",x"48",x"94",x"4C",x"94", -- 0x2578
    x"50",x"94",x"54",x"94",x"58",x"94",x"44",x"9C", -- 0x2580
    x"48",x"9C",x"4C",x"9C",x"50",x"9C",x"54",x"9C", -- 0x2588
    x"58",x"9C",x"44",x"AC",x"48",x"AC",x"4C",x"AC", -- 0x2590
    x"50",x"AC",x"54",x"AC",x"58",x"AC",x"44",x"B4", -- 0x2598
    x"48",x"B4",x"4C",x"B4",x"50",x"B4",x"54",x"B4", -- 0x25A0
    x"58",x"B4",x"44",x"BC",x"48",x"BC",x"4C",x"BC", -- 0x25A8
    x"50",x"BC",x"54",x"BC",x"58",x"BC",x"44",x"C4", -- 0x25B0
    x"48",x"C4",x"4C",x"C4",x"50",x"C4",x"54",x"C4", -- 0x25B8
    x"58",x"C4",x"44",x"CC",x"48",x"CC",x"4C",x"CC", -- 0x25C0
    x"50",x"CC",x"54",x"CC",x"58",x"CC",x"44",x"D4", -- 0x25C8
    x"48",x"D4",x"4C",x"D4",x"50",x"D4",x"54",x"D4", -- 0x25D0
    x"58",x"D4",x"44",x"DC",x"48",x"DC",x"4C",x"DC", -- 0x25D8
    x"50",x"DC",x"54",x"DC",x"58",x"DC",x"44",x"E4", -- 0x25E0
    x"48",x"E4",x"4C",x"E4",x"50",x"E4",x"54",x"E4", -- 0x25E8
    x"58",x"E4",x"CD",x"26",x"1E",x"CD",x"8D",x"1D", -- 0x25F0
    x"D0",x"DD",x"34",x"02",x"DD",x"7E",x"05",x"D6", -- 0x25F8
    x"10",x"DD",x"77",x"05",x"CD",x"F3",x"1E",x"DD", -- 0x2600
    x"34",x"02",x"CD",x"26",x"1E",x"CD",x"8D",x"1D", -- 0x2608
    x"D0",x"DD",x"34",x"02",x"21",x"B0",x"58",x"CB", -- 0x2610
    x"C6",x"21",x"DE",x"1E",x"DD",x"75",x"0C",x"DD", -- 0x2618
    x"74",x"0D",x"DD",x"36",x"0E",x"01",x"DD",x"7E", -- 0x2620
    x"17",x"C6",x"50",x"6F",x"26",x"41",x"36",x"03", -- 0x2628
    x"DD",x"36",x"18",x"00",x"DD",x"36",x"19",x"00", -- 0x2630
    x"21",x"1A",x"41",x"35",x"DD",x"36",x"10",x"0F", -- 0x2638
    x"DD",x"34",x"02",x"CD",x"26",x"1E",x"DD",x"35", -- 0x2640
    x"10",x"C0",x"DD",x"36",x"02",x"02",x"C9",x"AF", -- 0x2648
    x"67",x"68",x"57",x"59",x"06",x"08",x"CB",x"FF", -- 0x2650
    x"07",x"29",x"A7",x"ED",x"52",x"38",x"03",x"10", -- 0x2658
    x"F5",x"C9",x"19",x"CB",x"87",x"10",x"EF",x"C9", -- 0x2660
    x"AF",x"32",x"B0",x"58",x"32",x"D0",x"58",x"32", -- 0x2668
    x"E0",x"58",x"21",x"B8",x"40",x"35",x"C0",x"2D", -- 0x2670
    x"3A",x"1C",x"41",x"47",x"0F",x"38",x"13",x"3A", -- 0x2678
    x"1A",x"41",x"FE",x"2C",x"30",x"34",x"78",x"A7", -- 0x2680
    x"20",x"30",x"3E",x"01",x"32",x"1C",x"41",x"36", -- 0x2688
    x"02",x"C9",x"AF",x"32",x"1C",x"41",x"11",x"88", -- 0x2690
    x"06",x"FF",x"36",x"07",x"26",x"40",x"2E",x"AE", -- 0x2698
    x"36",x"20",x"2E",x"BF",x"36",x"12",x"3A",x"09", -- 0x26A0
    x"42",x"3C",x"32",x"09",x"42",x"FE",x"7F",x"C0", -- 0x26A8
    x"AF",x"32",x"09",x"42",x"26",x"40",x"2E",x"A1", -- 0x26B0
    x"34",x"C9",x"34",x"C9",x"21",x"10",x"41",x"34", -- 0x26B8
    x"21",x"14",x"41",x"34",x"11",x"00",x"07",x"FF", -- 0x26C0
    x"21",x"96",x"10",x"11",x"04",x"41",x"01",x"0C", -- 0x26C8
    x"00",x"ED",x"B0",x"21",x"11",x"41",x"36",x"2E", -- 0x26D0
    x"23",x"36",x"00",x"21",x"89",x"1B",x"22",x"07", -- 0x26D8
    x"42",x"21",x"B7",x"40",x"36",x"15",x"3A",x"15", -- 0x26E0
    x"41",x"0F",x"D8",x"36",x"13",x"3A",x"13",x"41", -- 0x26E8
    x"0F",x"D0",x"3E",x"01",x"32",x"15",x"41",x"C9", -- 0x26F0
    x"21",x"B7",x"40",x"34",x"2C",x"36",x"01",x"23", -- 0x26F8
    x"36",x"01",x"C9",x"21",x"B9",x"40",x"35",x"C0", -- 0x2700
    x"36",x"01",x"21",x"B7",x"40",x"34",x"C9",x"21", -- 0x2708
    x"B9",x"40",x"35",x"C0",x"36",x"10",x"21",x"20", -- 0x2710
    x"41",x"3A",x"15",x"41",x"0F",x"3E",x"00",x"38", -- 0x2718
    x"02",x"3E",x"02",x"06",x"30",x"D7",x"21",x"B7", -- 0x2720
    x"40",x"34",x"C9",x"21",x"B9",x"40",x"35",x"C0", -- 0x2728
    x"2D",x"36",x"00",x"3E",x"30",x"32",x"16",x"41", -- 0x2730
    x"21",x"10",x"41",x"34",x"21",x"14",x"41",x"34", -- 0x2738
    x"11",x"00",x"07",x"FF",x"11",x"08",x"06",x"3A", -- 0x2740
    x"15",x"41",x"0F",x"D4",x"38",x"00",x"21",x"72", -- 0x2748
    x"27",x"11",x"04",x"41",x"01",x"06",x"00",x"ED", -- 0x2750
    x"B0",x"21",x"11",x"41",x"36",x"18",x"2C",x"36", -- 0x2758
    x"16",x"21",x"B7",x"40",x"36",x"15",x"3A",x"15", -- 0x2760
    x"41",x"0F",x"D8",x"36",x"13",x"C9",x"2D",x"36", -- 0x2768
    x"03",x"C9",x"10",x"68",x"64",x"64",x"68",x"10", -- 0x2770
    x"C9",x"21",x"00",x"41",x"36",x"00",x"2C",x"34", -- 0x2778
    x"7E",x"47",x"2F",x"C6",x"80",x"32",x"2A",x"40", -- 0x2780
    x"32",x"2C",x"40",x"78",x"FE",x"FF",x"C0",x"36", -- 0x2788
    x"80",x"21",x"B7",x"40",x"34",x"16",x"01",x"FF", -- 0x2790
    x"23",x"36",x"19",x"3A",x"09",x"42",x"3C",x"32", -- 0x2798
    x"09",x"42",x"FE",x"7F",x"C0",x"AF",x"32",x"09", -- 0x27A0
    x"42",x"3E",x"01",x"32",x"0A",x"40",x"C9",x"21", -- 0x27A8
    x"B8",x"40",x"35",x"C0",x"3E",x"F7",x"32",x"BB", -- 0x27B0
    x"40",x"2F",x"32",x"38",x"40",x"32",x"3A",x"40", -- 0x27B8
    x"21",x"B7",x"40",x"34",x"21",x"A0",x"58",x"CB", -- 0x27C0
    x"D6",x"11",x"09",x"06",x"FF",x"3A",x"09",x"42", -- 0x27C8
    x"3C",x"32",x"09",x"42",x"FE",x"7F",x"C0",x"AF", -- 0x27D0
    x"32",x"09",x"42",x"21",x"1A",x"41",x"34",x"C9", -- 0x27D8
    x"21",x"BA",x"40",x"36",x"01",x"2C",x"35",x"7E", -- 0x27E0
    x"47",x"2F",x"C6",x"80",x"32",x"38",x"40",x"32", -- 0x27E8
    x"3A",x"40",x"78",x"FE",x"80",x"C0",x"11",x"89", -- 0x27F0
    x"06",x"FF",x"E5",x"21",x"A0",x"58",x"CB",x"96", -- 0x27F8
    x"E1",x"16",x"40",x"23",x"1E",x"BF",x"36",x"00", -- 0x2800
    x"21",x"B7",x"40",x"34",x"C9",x"CD",x"C5",x"17", -- 0x2808
    x"CD",x"1F",x"18",x"CD",x"DC",x"18",x"21",x"BC", -- 0x2810
    x"40",x"7E",x"2D",x"0F",x"38",x"08",x"35",x"7E", -- 0x2818
    x"FE",x"27",x"38",x"13",x"18",x"06",x"34",x"7E", -- 0x2820
    x"FE",x"D9",x"30",x"0B",x"2F",x"C6",x"80",x"32", -- 0x2828
    x"38",x"40",x"32",x"3A",x"40",x"18",x"02",x"2C", -- 0x2830
    x"34",x"CD",x"6A",x"28",x"38",x"13",x"3A",x"BC", -- 0x2838
    x"40",x"FE",x"0A",x"C0",x"AF",x"32",x"9D",x"40", -- 0x2840
    x"11",x"89",x"06",x"FF",x"21",x"B7",x"40",x"34", -- 0x2848
    x"C9",x"21",x"E0",x"58",x"CB",x"C6",x"AF",x"32", -- 0x2850
    x"9D",x"40",x"11",x"89",x"06",x"FF",x"21",x"B7", -- 0x2858
    x"40",x"36",x"0D",x"2C",x"36",x"0A",x"2C",x"36", -- 0x2860
    x"06",x"C9",x"21",x"7C",x"42",x"7E",x"0F",x"D0", -- 0x2868
    x"23",x"3A",x"BB",x"40",x"C6",x"02",x"96",x"FE", -- 0x2870
    x"05",x"D0",x"2C",x"2C",x"7E",x"FE",x"6E",x"D0", -- 0x2878
    x"FE",x"69",x"3F",x"C9",x"AF",x"32",x"BA",x"40", -- 0x2880
    x"32",x"7C",x"42",x"21",x"BB",x"40",x"35",x"7E", -- 0x2888
    x"47",x"2F",x"C6",x"80",x"32",x"38",x"40",x"32", -- 0x2890
    x"3A",x"40",x"78",x"FE",x"08",x"C0",x"CD",x"62", -- 0x2898
    x"2A",x"21",x"B7",x"40",x"34",x"2C",x"36",x"64", -- 0x28A0
    x"C9",x"21",x"B8",x"40",x"35",x"C0",x"3E",x"01", -- 0x28A8
    x"32",x"00",x"41",x"32",x"B7",x"40",x"C9",x"21", -- 0x28B0
    x"B8",x"40",x"35",x"C0",x"E5",x"21",x"E0",x"58", -- 0x28B8
    x"CB",x"C6",x"E1",x"AF",x"32",x"BA",x"40",x"32", -- 0x28C0
    x"7C",x"42",x"36",x"0A",x"CD",x"62",x"2A",x"2D", -- 0x28C8
    x"34",x"C9",x"21",x"B8",x"40",x"35",x"C0",x"36", -- 0x28D0
    x"0A",x"CD",x"75",x"2A",x"2D",x"34",x"C9",x"21", -- 0x28D8
    x"B9",x"40",x"35",x"20",x"17",x"CD",x"62",x"2A", -- 0x28E0
    x"11",x"AB",x"40",x"AF",x"12",x"1C",x"12",x"1C", -- 0x28E8
    x"12",x"E5",x"CD",x"31",x"29",x"E1",x"36",x"64", -- 0x28F0
    x"2D",x"2D",x"34",x"C9",x"2D",x"2D",x"36",x"0D", -- 0x28F8
    x"C9",x"21",x"B9",x"40",x"35",x"C0",x"11",x"8A", -- 0x2900
    x"06",x"FF",x"36",x"0A",x"2D",x"2D",x"34",x"C9", -- 0x2908
    x"21",x"B9",x"40",x"35",x"C0",x"36",x"0A",x"CD", -- 0x2910
    x"9B",x"2A",x"38",x"0C",x"CD",x"31",x"29",x"CD", -- 0x2918
    x"AD",x"2A",x"21",x"E0",x"58",x"CB",x"CE",x"C9", -- 0x2920
    x"21",x"B7",x"40",x"34",x"2C",x"2C",x"36",x"46", -- 0x2928
    x"C9",x"3A",x"BC",x"40",x"47",x"3E",x"0A",x"90", -- 0x2930
    x"07",x"07",x"07",x"07",x"E6",x"F0",x"00",x"00", -- 0x2938
    x"21",x"AB",x"40",x"86",x"27",x"77",x"23",x"3E", -- 0x2940
    x"00",x"8E",x"27",x"77",x"2D",x"7E",x"E6",x"0F", -- 0x2948
    x"32",x"CD",x"51",x"7E",x"0F",x"0F",x"0F",x"0F", -- 0x2950
    x"E6",x"0F",x"32",x"ED",x"51",x"2C",x"7E",x"E6", -- 0x2958
    x"F0",x"28",x"0E",x"0F",x"0F",x"0F",x"0F",x"32", -- 0x2960
    x"2D",x"52",x"7E",x"E6",x"0F",x"32",x"0D",x"52", -- 0x2968
    x"C9",x"7E",x"E6",x"0F",x"C8",x"32",x"0D",x"52", -- 0x2970
    x"C9",x"21",x"B9",x"40",x"35",x"C0",x"11",x"8A", -- 0x2978
    x"06",x"FF",x"11",x"00",x"03",x"FF",x"2D",x"2D", -- 0x2980
    x"3E",x"01",x"77",x"32",x"00",x"41",x"AF",x"32", -- 0x2988
    x"16",x"41",x"C9",x"11",x"65",x"06",x"3A",x"13", -- 0x2990
    x"41",x"0F",x"38",x"11",x"3A",x"14",x"41",x"FE", -- 0x2998
    x"05",x"20",x"05",x"3E",x"04",x"32",x"14",x"41", -- 0x29A0
    x"C6",x"20",x"F6",x"40",x"5F",x"FF",x"21",x"B8", -- 0x29A8
    x"40",x"36",x"00",x"2D",x"34",x"C9",x"21",x"B8", -- 0x29B0
    x"40",x"35",x"C0",x"11",x"A5",x"06",x"FF",x"3E", -- 0x29B8
    x"05",x"32",x"0A",x"40",x"C9",x"21",x"B9",x"40", -- 0x29C0
    x"36",x"08",x"2D",x"36",x"32",x"2D",x"34",x"E5", -- 0x29C8
    x"21",x"A0",x"58",x"CB",x"DE",x"E1",x"11",x"26", -- 0x29D0
    x"06",x"FF",x"AF",x"32",x"3A",x"40",x"C9",x"21", -- 0x29D8
    x"B8",x"40",x"35",x"C0",x"36",x"0F",x"11",x"27", -- 0x29E0
    x"06",x"FF",x"11",x"26",x"06",x"FF",x"2D",x"34", -- 0x29E8
    x"C9",x"21",x"B8",x"40",x"35",x"C0",x"36",x"0F", -- 0x29F0
    x"E5",x"21",x"A0",x"58",x"CB",x"9E",x"E1",x"11", -- 0x29F8
    x"A7",x"06",x"FF",x"11",x"A6",x"06",x"FF",x"2D", -- 0x2A00
    x"34",x"C9",x"21",x"B9",x"40",x"35",x"28",x"05", -- 0x2A08
    x"2D",x"2D",x"36",x"16",x"C9",x"21",x"96",x"10", -- 0x2A10
    x"11",x"04",x"41",x"01",x"0C",x"00",x"ED",x"B0", -- 0x2A18
    x"21",x"B2",x"10",x"11",x"20",x"41",x"01",x"C0", -- 0x2A20
    x"00",x"ED",x"B0",x"11",x"60",x"06",x"FF",x"AF", -- 0x2A28
    x"21",x"13",x"41",x"77",x"2C",x"77",x"2C",x"77", -- 0x2A30
    x"32",x"12",x"41",x"32",x"1C",x"41",x"32",x"16", -- 0x2A38
    x"41",x"3E",x"2E",x"32",x"11",x"41",x"3E",x"60", -- 0x2A40
    x"32",x"1A",x"41",x"21",x"B7",x"40",x"34",x"2C", -- 0x2A48
    x"36",x"00",x"C9",x"21",x"B8",x"40",x"35",x"C0", -- 0x2A50
    x"11",x"A0",x"06",x"FF",x"3E",x"05",x"32",x"0A", -- 0x2A58
    x"40",x"C9",x"E5",x"06",x"06",x"21",x"AC",x"51", -- 0x2A60
    x"11",x"1F",x"00",x"36",x"10",x"23",x"36",x"10", -- 0x2A68
    x"19",x"10",x"F8",x"E1",x"C9",x"E5",x"06",x"06", -- 0x2A70
    x"21",x"AC",x"51",x"11",x"20",x"00",x"DD",x"21", -- 0x2A78
    x"D8",x"02",x"DD",x"7E",x"00",x"77",x"19",x"DD", -- 0x2A80
    x"23",x"10",x"F7",x"06",x"06",x"21",x"AD",x"51", -- 0x2A88
    x"DD",x"7E",x"00",x"77",x"19",x"DD",x"23",x"10", -- 0x2A90
    x"F7",x"E1",x"C9",x"06",x"30",x"21",x"20",x"41", -- 0x2A98
    x"CB",x"4E",x"20",x"05",x"23",x"10",x"F9",x"37", -- 0x2AA0
    x"C9",x"CB",x"8E",x"A7",x"C9",x"21",x"55",x"41", -- 0x2AA8
    x"11",x"06",x"00",x"4B",x"06",x"18",x"CB",x"4E", -- 0x2AB0
    x"20",x"0B",x"19",x"10",x"F9",x"7D",x"D6",x"91", -- 0x2AB8
    x"6F",x"0D",x"20",x"F0",x"C9",x"36",x"01",x"21", -- 0x2AC0
    x"1A",x"41",x"34",x"C9",x"3E",x"03",x"32",x"06", -- 0x2AC8
    x"68",x"0F",x"32",x"07",x"68",x"3A",x"F3",x"58", -- 0x2AD0
    x"32",x"05",x"68",x"0F",x"32",x"03",x"68",x"0F", -- 0x2AD8
    x"32",x"00",x"68",x"32",x"01",x"68",x"32",x"02", -- 0x2AE0
    x"68",x"21",x"A0",x"42",x"11",x"20",x"00",x"06", -- 0x2AE8
    x"08",x"AF",x"B6",x"19",x"10",x"FC",x"0F",x"38", -- 0x2AF0
    x"05",x"21",x"C0",x"58",x"CB",x"96",x"21",x"B1", -- 0x2AF8
    x"2D",x"DD",x"21",x"C0",x"58",x"FD",x"21",x"F3", -- 0x2B00
    x"58",x"CD",x"36",x"2D",x"21",x"E1",x"2D",x"DD", -- 0x2B08
    x"21",x"90",x"58",x"FD",x"21",x"F1",x"58",x"CD", -- 0x2B10
    x"1A",x"2C",x"21",x"F1",x"2D",x"DD",x"21",x"B0", -- 0x2B18
    x"58",x"FD",x"21",x"F0",x"58",x"CD",x"1A",x"2C", -- 0x2B20
    x"21",x"11",x"2E",x"DD",x"21",x"E0",x"58",x"FD", -- 0x2B28
    x"21",x"F5",x"58",x"CD",x"1A",x"2C",x"21",x"B2", -- 0x2B30
    x"2D",x"DD",x"21",x"A0",x"58",x"FD",x"21",x"F2", -- 0x2B38
    x"58",x"CD",x"92",x"2B",x"06",x"00",x"21",x"F5", -- 0x2B40
    x"58",x"CD",x"6D",x"2B",x"21",x"F6",x"58",x"CD", -- 0x2B48
    x"6D",x"2B",x"21",x"F0",x"58",x"CD",x"6D",x"2B", -- 0x2B50
    x"21",x"F2",x"58",x"CD",x"6D",x"2B",x"21",x"F1", -- 0x2B58
    x"58",x"CD",x"6D",x"2B",x"CB",x"40",x"C0",x"3E", -- 0x2B60
    x"FF",x"32",x"00",x"78",x"C9",x"7E",x"A7",x"C8", -- 0x2B68
    x"CB",x"C0",x"32",x"00",x"78",x"C9",x"85",x"6F", -- 0x2B70
    x"3E",x"00",x"8C",x"67",x"7E",x"C9",x"78",x"87", -- 0x2B78
    x"CD",x"76",x"2B",x"5F",x"23",x"56",x"EB",x"C9", -- 0x2B80
    x"E1",x"87",x"CD",x"76",x"2B",x"5F",x"23",x"56", -- 0x2B88
    x"EB",x"E9",x"DD",x"7E",x"00",x"A7",x"CA",x"20", -- 0x2B90
    x"2C",x"4F",x"06",x"08",x"1E",x"80",x"7B",x"A1", -- 0x2B98
    x"20",x"05",x"CB",x"3B",x"10",x"F8",x"C9",x"DD", -- 0x2BA0
    x"7E",x"02",x"A3",x"20",x"09",x"DD",x"73",x"02", -- 0x2BA8
    x"05",x"CD",x"7E",x"2B",x"18",x"0C",x"DD",x"35", -- 0x2BB0
    x"0C",x"C2",x"13",x"2C",x"DD",x"6E",x"06",x"DD", -- 0x2BB8
    x"66",x"07",x"7E",x"23",x"DD",x"75",x"06",x"DD", -- 0x2BC0
    x"74",x"07",x"FE",x"F0",x"38",x"2A",x"21",x"BC", -- 0x2BC8
    x"2B",x"E5",x"E6",x"0F",x"CD",x"88",x"2B",x"14", -- 0x2BD0
    x"2D",x"24",x"2D",x"F7",x"2B",x"F7",x"2B",x"F7", -- 0x2BD8
    x"2B",x"F7",x"2B",x"F7",x"2B",x"F7",x"2B",x"F7", -- 0x2BE0
    x"2B",x"F7",x"2B",x"F7",x"2B",x"F7",x"2B",x"F7", -- 0x2BE8
    x"2B",x"F7",x"2B",x"F7",x"2B",x"A0",x"2D",x"C9", -- 0x2BF0
    x"47",x"07",x"07",x"07",x"E6",x"07",x"21",x"BA", -- 0x2BF8
    x"2D",x"CD",x"76",x"2B",x"DD",x"77",x"0C",x"78", -- 0x2C00
    x"E6",x"1F",x"21",x"C2",x"2D",x"CD",x"76",x"2B", -- 0x2C08
    x"DD",x"77",x"0E",x"DD",x"7E",x"0E",x"FD",x"77", -- 0x2C10
    x"00",x"C9",x"DD",x"7E",x"00",x"A7",x"20",x"23", -- 0x2C18
    x"DD",x"7E",x"02",x"A7",x"3E",x"00",x"FD",x"77", -- 0x2C20
    x"00",x"C8",x"DD",x"36",x"00",x"00",x"DD",x"36", -- 0x2C28
    x"02",x"00",x"DD",x"36",x"0D",x"00",x"DD",x"36", -- 0x2C30
    x"0E",x"00",x"DD",x"36",x"0F",x"00",x"FD",x"36", -- 0x2C38
    x"00",x"00",x"C9",x"4F",x"06",x"08",x"1E",x"80", -- 0x2C40
    x"7B",x"A1",x"20",x"05",x"CB",x"3B",x"10",x"F8", -- 0x2C48
    x"C9",x"DD",x"7E",x"02",x"A3",x"20",x"3F",x"DD", -- 0x2C50
    x"73",x"02",x"05",x"78",x"07",x"07",x"07",x"4F", -- 0x2C58
    x"06",x"00",x"E5",x"09",x"DD",x"E5",x"D1",x"13", -- 0x2C60
    x"13",x"13",x"01",x"08",x"00",x"ED",x"B0",x"E1", -- 0x2C68
    x"DD",x"7E",x"06",x"E6",x"7F",x"DD",x"77",x"0C", -- 0x2C70
    x"DD",x"7E",x"04",x"DD",x"77",x"0E",x"DD",x"7E", -- 0x2C78
    x"09",x"47",x"0F",x"0F",x"0F",x"0F",x"E6",x"0F", -- 0x2C80
    x"DD",x"77",x"0B",x"E6",x"08",x"20",x"07",x"DD", -- 0x2C88
    x"70",x"0F",x"DD",x"36",x"0D",x"00",x"DD",x"35", -- 0x2C90
    x"0C",x"20",x"5A",x"DD",x"7E",x"08",x"A7",x"28", -- 0x2C98
    x"10",x"DD",x"35",x"08",x"20",x"0B",x"7B",x"2F", -- 0x2CA0
    x"DD",x"A6",x"00",x"DD",x"77",x"00",x"C3",x"1A", -- 0x2CA8
    x"2C",x"DD",x"7E",x"06",x"E6",x"7F",x"DD",x"77", -- 0x2CB0
    x"0C",x"DD",x"CB",x"06",x"7E",x"28",x"16",x"DD", -- 0x2CB8
    x"7E",x"05",x"ED",x"44",x"DD",x"77",x"05",x"DD", -- 0x2CC0
    x"CB",x"0D",x"46",x"DD",x"CB",x"0D",x"C6",x"28", -- 0x2CC8
    x"24",x"DD",x"CB",x"0D",x"86",x"DD",x"7E",x"04", -- 0x2CD0
    x"DD",x"86",x"07",x"DD",x"77",x"04",x"DD",x"77", -- 0x2CD8
    x"0E",x"DD",x"7E",x"09",x"DD",x"86",x"0A",x"DD", -- 0x2CE0
    x"77",x"09",x"47",x"DD",x"7E",x"0B",x"E6",x"08", -- 0x2CE8
    x"20",x"03",x"DD",x"70",x"0F",x"DD",x"7E",x"0E", -- 0x2CF0
    x"DD",x"86",x"05",x"DD",x"77",x"0E",x"6F",x"26", -- 0x2CF8
    x"00",x"DD",x"7E",x"03",x"E6",x"70",x"28",x"08", -- 0x2D00
    x"0F",x"0F",x"0F",x"0F",x"47",x"29",x"10",x"FD", -- 0x2D08
    x"FD",x"75",x"00",x"C9",x"DD",x"6E",x"06",x"DD", -- 0x2D10
    x"66",x"07",x"7E",x"DD",x"77",x"06",x"23",x"7E", -- 0x2D18
    x"DD",x"77",x"07",x"C9",x"DD",x"6E",x"06",x"DD", -- 0x2D20
    x"66",x"07",x"7E",x"23",x"DD",x"75",x"06",x"DD", -- 0x2D28
    x"74",x"07",x"32",x"F4",x"58",x"C9",x"CD",x"40", -- 0x2D30
    x"2D",x"CD",x"64",x"2D",x"CD",x"88",x"2D",x"C9", -- 0x2D38
    x"DD",x"7E",x"00",x"CB",x"47",x"28",x"0A",x"DD", -- 0x2D40
    x"CB",x"00",x"86",x"3E",x"08",x"DD",x"77",x"01", -- 0x2D48
    x"C9",x"DD",x"7E",x"01",x"A7",x"28",x"08",x"DD", -- 0x2D50
    x"35",x"01",x"FD",x"CB",x"00",x"C6",x"C9",x"FD", -- 0x2D58
    x"CB",x"00",x"86",x"C9",x"DD",x"7E",x"00",x"CB", -- 0x2D60
    x"4F",x"28",x"0A",x"DD",x"CB",x"00",x"8E",x"3E", -- 0x2D68
    x"1D",x"DD",x"77",x"02",x"C9",x"DD",x"7E",x"02", -- 0x2D70
    x"A7",x"28",x"08",x"DD",x"35",x"02",x"FD",x"CB", -- 0x2D78
    x"00",x"CE",x"C9",x"FD",x"CB",x"00",x"8E",x"C9", -- 0x2D80
    x"DD",x"7E",x"00",x"CB",x"57",x"28",x"0C",x"3A", -- 0x2D88
    x"A0",x"58",x"CB",x"47",x"20",x"05",x"FD",x"CB", -- 0x2D90
    x"00",x"D6",x"C9",x"FD",x"CB",x"00",x"96",x"C9", -- 0x2D98
    x"DD",x"7E",x"02",x"2F",x"DD",x"A6",x"00",x"AF", -- 0x2DA0
    x"FD",x"77",x"00",x"DD",x"77",x"00",x"C3",x"20", -- 0x2DA8
    x"2C",x"00",x"21",x"2E",x"40",x"2E",x"6F",x"2E", -- 0x2DB0
    x"85",x"2E",x"01",x"02",x"04",x"08",x"10",x"20", -- 0x2DB8
    x"40",x"00",x"FF",x"00",x"40",x"55",x"5F",x"68", -- 0x2DC0
    x"70",x"80",x"8E",x"9A",x"A0",x"AA",x"B4",x"B8", -- 0x2DC8
    x"C0",x"C7",x"CD",x"D0",x"D5",x"DA",x"DC",x"E0", -- 0x2DD0
    x"1C",x"35",x"87",x"A5",x"C4",x"D3",x"CA",x"E3", -- 0x2DD8
    x"E6",x"20",x"40",x"10",x"87",x"00",x"0A",x"FF", -- 0x2DE0
    x"FF",x"40",x"20",x"FF",x"90",x"00",x"01",x"FF", -- 0x2DE8
    x"FF",x"40",x"20",x"FB",x"87",x"00",x"01",x"FF", -- 0x2DF0
    x"FF",x"40",x"20",x"FB",x"87",x"00",x"01",x"FF", -- 0x2DF8
    x"FF",x"20",x"70",x"FB",x"87",x"00",x"02",x"FF", -- 0x2E00
    x"FF",x"20",x"70",x"FB",x"87",x"00",x"02",x"FF", -- 0x2E08
    x"FF",x"80",x"20",x"F4",x"87",x"FE",x"10",x"FF", -- 0x2E10
    x"FF",x"80",x"20",x"F4",x"87",x"04",x"01",x"FF", -- 0x2E18
    x"FF",x"68",x"00",x"68",x"6A",x"6C",x"8B",x"88", -- 0x2E20
    x"00",x"68",x"00",x"68",x"67",x"6A",x"88",x"88", -- 0x2E28
    x"00",x"68",x"00",x"68",x"6A",x"6C",x"8B",x"8F", -- 0x2E30
    x"6E",x"00",x"6E",x"6C",x"6A",x"8F",x"8F",x"FF", -- 0x2E38
    x"80",x"6C",x"6B",x"8C",x"6B",x"6A",x"8B",x"6A", -- 0x2E40
    x"69",x"8A",x"69",x"68",x"89",x"65",x"67",x"88", -- 0x2E48
    x"4A",x"00",x"4A",x"00",x"4A",x"88",x"6C",x"6B", -- 0x2E50
    x"8C",x"6B",x"6A",x"8B",x"6A",x"69",x"8A",x"69", -- 0x2E58
    x"68",x"89",x"65",x"67",x"88",x"4A",x"00",x"4A", -- 0x2E60
    x"00",x"4A",x"88",x"A0",x"A0",x"10",x"FF",x"80", -- 0x2E68
    x"60",x"69",x"00",x"69",x"00",x"69",x"87",x"87", -- 0x2E70
    x"87",x"68",x"00",x"68",x"00",x"68",x"86",x"86", -- 0x2E78
    x"86",x"A0",x"A0",x"10",x"FF",x"65",x"67",x"67", -- 0x2E80
    x"65",x"68",x"87",x"00",x"87",x"60",x"65",x"68", -- 0x2E88
    x"00",x"68",x"65",x"69",x"88",x"00",x"88",x"60", -- 0x2E90
    x"A0",x"A0",x"A0",x"A0",x"A0",x"10",x"FF",x"FF", -- 0x2E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3428
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3448
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3468
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3610
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3620
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3638
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3648
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3650
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3658
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3668
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3678
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3688
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3690
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3698
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3708
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3710
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3718
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3728
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3738
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3748
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3750
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3758
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3768
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3778
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3788
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3798
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3828
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3838
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
       DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
