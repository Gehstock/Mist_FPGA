library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_spr_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_spr_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"07",X"03",X"03",X"02",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"F1",X"F8",X"7D",X"1F",X"3F",X"3F",X"37",X"21",X"30",X"30",X"18",X"4F",
		X"80",X"80",X"82",X"8F",X"8F",X"0F",X"0E",X"C0",X"C0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"31",X"39",X"19",X"19",X"1C",X"1C",X"0E",X"0E",X"0E",X"06",X"06",X"04",X"04",X"04",X"06",X"02",
		X"C0",X"E0",X"E0",X"A0",X"A0",X"A0",X"A0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0C",X"0E",X"0F",X"0F",X"07",X"03",X"03",X"02",X"08",
		X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"E0",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"98",X"88",X"80",X"C8",X"48",X"24",X"34",X"3E",X"3F",X"7F",
		X"00",X"00",X"00",X"20",X"70",X"70",X"38",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"0E",X"FC",X"FE",X"DE",X"8F",X"87",X"87",X"43",X"33",X"39",X"1D",X"0C",X"08",X"08",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"27",X"37",X"3F",X"1F",X"0F",X"0C",X"08",X"30",X"60",X"C0",X"C4",
		X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"C2",X"42",X"40",X"40",X"00",X"40",X"40",X"40",X"A0",X"F8",X"F8",X"D8",X"D8",X"CC",
		X"80",X"C0",X"C3",X"62",X"20",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"30",X"38",X"3C",X"9C",X"CC",X"FE",X"FE",X"76",X"77",X"33",X"3B",X"9D",X"CF",X"EF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"00",X"01",X"03",X"03",X"03",X"03",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"F8",X"F8",X"FC",X"FC",X"FC",X"F8",X"78",X"7C",X"F8",X"F0",X"E0",X"80",X"80",X"80",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"B0",X"19",X"4E",X"00",X"00",X"00",X"A0",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"78",X"7C",X"3C",X"3E",X"DE",X"CF",X"E7",X"73",X"79",X"3C",X"1F",X"0F",X"CF",X"C3",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"E0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"07",X"07",X"0F",X"07",X"03",X"03",X"07",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"30",X"70",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"7E",X"7C",X"3C",X"1A",X"06",X"06",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"09",X"19",X"11",X"03",X"11",X"10",X"28",X"78",X"F8",X"7C",X"64",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"7B",X"F7",X"F6",X"FC",X"FC",X"EC",X"CC",X"DC",X"D8",X"D8",X"D8",X"D8",X"D0",X"D0",X"F0",X"F0",
		X"01",X"01",X"03",X"03",X"03",X"01",X"01",X"03",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"FC",X"FC",X"FC",X"E4",X"EC",X"FC",X"F8",X"F0",X"F0",X"E0",X"04",X"02",X"03",X"03",
		X"00",X"00",X"61",X"23",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"C1",X"A1",X"23",X"02",X"00",X"04",X"05",X"C9",X"FD",X"FF",X"FF",X"7E",X"7E",X"72",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",
		X"00",X"11",X"11",X"23",X"23",X"27",X"67",X"4F",X"4E",X"DE",X"9C",X"BC",X"BC",X"38",X"78",X"78",
		X"1F",X"1F",X"3F",X"3F",X"3F",X"1F",X"1E",X"3E",X"1F",X"0F",X"07",X"01",X"01",X"01",X"00",X"04",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"0D",X"98",X"70",X"00",X"00",X"04",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"02",X"06",X"07",X"0E",X"0E",
		X"06",X"1F",X"3F",X"3E",X"7E",X"7C",X"FC",X"F8",X"F1",X"F3",X"2F",X"4E",X"9C",X"1C",X"38",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"06",X"04",X"0C",X"0C",X"1C",X"1C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"F1",X"F8",X"7D",X"1F",X"3F",X"3F",X"37",X"21",X"30",X"30",X"18",X"4F",
		X"80",X"80",X"82",X"8F",X"8F",X"0F",X"0E",X"C0",X"C0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"40",X"40",X"60",X"78",X"3E",X"38",X"30",X"30",X"31",X"39",X"19",X"19",X"1C",X"1C",X"0E",X"0E",
		X"00",X"80",X"90",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"A0",X"A0",X"A0",X"A0",X"E0",
		X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"70",X"70",X"70",X"70",X"30",X"30",X"B0",X"B0",X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"10",X"30",X"30",X"71",X"71",X"71",X"79",X"78",X"78",X"7C",X"34",X"02",X"03",X"03",X"03",X"07",
		X"00",X"00",X"00",X"02",X"07",X"07",X"83",X"83",X"00",X"80",X"80",X"40",X"40",X"E0",X"F8",X"F0",
		X"4E",X"46",X"66",X"66",X"7F",X"00",X"00",X"00",X"04",X"1F",X"0F",X"0F",X"06",X"06",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"F0",X"F8",X"78",X"3C",X"1C",X"1C",X"0C",
		X"06",X"06",X"06",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"20",X"B0",X"B0",X"B0",X"B0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"C4",X"E4",X"66",X"62",X"72",X"72",X"70",X"62",X"3A",X"0A",X"0D",X"07",X"07",X"06",X"06",X"06",
		X"04",X"0E",X"16",X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"60",
		X"EE",X"F8",X"00",X"00",X"00",X"01",X"13",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"10",X"38",X"FE",X"FF",X"AF",X"03",X"01",X"01",X"C0",X"70",X"1E",X"07",X"03",X"03",
		X"63",X"31",X"18",X"0E",X"07",X"07",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"60",X"20",X"30",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"7E",
		X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"A0",X"B0",X"90",X"C4",X"CE",X"E7",X"73",X"3F",X"03",X"03",X"01",X"01",X"01",X"00",
		X"E0",X"F0",X"F8",X"D8",X"D0",X"E0",X"C0",X"01",X"01",X"03",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"3C",X"3F",X"FF",X"CC",X"C0",X"80",X"80",X"E0",X"30",X"0F",X"01",
		X"70",X"38",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"48",X"0C",X"84",X"EE",X"FE",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"E0",X"E0",X"C1",X"C1",X"A0",X"61",X"61",X"42",X"07",X"0F",X"07",X"06",
		X"00",X"00",X"00",X"80",X"98",X"98",X"98",X"1C",X"3E",X"1E",X"0C",X"80",X"80",X"80",X"C0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"1F",X"1E",X"3D",X"3D",X"3F",X"7F",X"7B",X"73",X"77",
		X"64",X"C4",X"CC",X"7C",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"20",X"30",X"68",X"C8",X"80",X"00",X"01",X"01",X"32",X"3F",X"3F",X"3F",X"1F",X"1F",X"1C",X"19",
		X"47",X"47",X"4E",X"CE",X"9E",X"1E",X"1E",X"7E",X"4C",X"40",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"01",X"20",X"20",X"70",X"78",X"F3",X"EE",X"F0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"E4",X"38",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"06",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7E",
		X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"04",X"04",X"0D",X"19",X"13",X"67",X"EA",X"D8",X"B0",X"F0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",
		X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"04",X"0C",X"0E",X"3F",X"7F",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"3F",X"1F",X"1F",X"0B",X"03",X"C3",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"11",X"33",X"27",X"7F",X"7F",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"10",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"1C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"70",X"1C",X"03",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"78",X"08",X"07",
		X"00",X"00",X"00",X"08",X"04",X"04",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"06",X"1C",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"80",X"00",X"80",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"08",X"80",X"00",X"80",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"08",X"80",X"80",X"08",X"80",X"80",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"01",X"23",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"02",X"02",X"02",X"66",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"02",X"02",X"02",X"02",X"E6",X"3F",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"07",X"FC",
		X"00",X"00",X"00",X"00",X"01",X"05",X"01",X"00",X"00",X"02",X"02",X"02",X"02",X"86",X"F4",X"1F",
		X"00",X"00",X"04",X"0C",X"04",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"03",X"06",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"02",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"06",X"06",X"EC",X"3F",
		X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"03",X"00",
		X"00",X"01",X"05",X"01",X"00",X"00",X"00",X"02",X"02",X"02",X"03",X"03",X"07",X"06",X"EC",X"3F",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",
		X"C0",X"80",X"80",X"00",X"00",X"40",X"C0",X"40",X"00",X"00",X"00",X"10",X"30",X"60",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"D0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",X"04",X"04",X"0C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"60",X"E0",X"EC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"04",X"05",X"0D",X"18",X"39",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"E4",X"EC",X"FE",
		X"00",X"00",X"04",X"04",X"0C",X"08",X"18",X"18",X"1A",X"32",X"71",X"E1",X"3B",X"7F",X"1C",X"08",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C4",X"CE",X"FC",X"F6",X"FC",X"2A",
		X"02",X"04",X"04",X"04",X"0C",X"0C",X"19",X"39",X"78",X"F0",X"61",X"3F",X"1F",X"37",X"C2",X"02",
		X"40",X"40",X"40",X"40",X"40",X"40",X"60",X"62",X"E1",X"E1",X"E2",X"FF",X"FF",X"DE",X"0A",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"0C",X"0C",X"0C",X"18",X"38",X"79",X"F9",X"F0",X"F1",X"E0",X"79",X"3F",X"7F",X"DF",X"0E",X"35",
		X"60",X"60",X"60",X"60",X"60",X"61",X"71",X"70",X"F0",X"F1",X"F3",X"FF",X"FF",X"8B",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"80",X"00",X"80",X"C0",X"80",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"01",X"03",X"01",X"00",X"02",X"00",X"01",X"06",X"00",X"01",
		X"38",X"38",X"78",X"F0",X"F1",X"F1",X"F0",X"E1",X"E0",X"C0",X"79",X"DF",X"0F",X"07",X"3F",X"C6",
		X"20",X"20",X"70",X"70",X"70",X"70",X"78",X"78",X"F8",X"F8",X"FF",X"FF",X"FE",X"F1",X"02",X"80",
		X"00",X"00",X"00",X"00",X"60",X"30",X"28",X"30",X"60",X"C0",X"E0",X"F8",X"D0",X"40",X"20",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"07",
		X"00",X"00",X"03",X"1F",X"3F",X"7F",X"FE",X"FC",X"FC",X"FE",X"7F",X"00",X"00",X"00",X"03",X"FF",
		X"00",X"00",X"C0",X"F8",X"FC",X"FE",X"7F",X"7F",X"7F",X"7F",X"FE",X"00",X"00",X"00",X"C0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"03",X"0F",X"1F",X"1F",X"3E",X"2E",X"4E",X"4F",X"80",X"80",X"00",X"03",X"FF",
		X"00",X"00",X"7C",X"FF",X"FF",X"FF",X"3F",X"3F",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"C0",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"40",X"40",X"40",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"1E",X"16",X"26",X"47",X"40",X"80",X"00",X"07",X"FF",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"3F",X"3F",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"80",X"FF",
		X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"40",X"40",X"40",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0C",X"08",X"10",X"21",X"40",X"80",X"00",X"0F",X"FF",
		X"00",X"00",X"07",X"3F",X"FF",X"FF",X"3F",X"3F",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"20",X"40",X"40",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"30",X"43",X"80",X"00",X"00",X"1E",X"FF",
		X"00",X"00",X"03",X"1F",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"FF",
		X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"F0",X"F0",X"E0",X"40",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"08",X"30",X"7F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0C",X"18",X"11",X"21",X"C7",X"00",X"00",X"00",X"78",X"FF",
		X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"02",X"FC",
		X"00",X"00",X"F8",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"10",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"08",X"09",X"31",X"47",X"80",X"00",X"00",X"F0",X"FF",
		X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"06",X"08",X"F0",
		X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0E",X"10",X"E3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"02",X"13",X"EF",X"00",X"00",X"00",X"F0",X"FF",
		X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"06",X"08",X"F0",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"38",X"C7",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"04",X"05",X"7F",X"00",X"00",X"00",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"06",X"18",X"E0",
		X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F8",X"F8",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"0E",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3E",
		X"00",X"00",X"00",X"04",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"04",X"08",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"07",X"4F",X"2F",X"0F",X"07",X"06",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"F2",X"F4",X"F0",X"F0",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"07",X"4F",X"2F",X"0F",X"07",X"06",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"F2",X"F4",X"F0",X"F0",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"4F",X"4F",X"4F",X"0E",X"07",X"57",X"7B",X"2F",
		X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F8",X"F4",X"F4",X"74",X"60",X"C2",X"C2",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"1F",X"0F",X"20",X"30",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"E0",X"00",X"00",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"06",X"07",X"0F",X"07",X"07",X"03",X"07",
		X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"F0",X"E0",X"C0",X"80",X"00",
		X"1F",X"40",X"40",X"60",X"70",X"7F",X"3E",X"3C",X"3D",X"19",X"19",X"1D",X"0D",X"08",X"08",X"0C",
		X"80",X"00",X"00",X"80",X"F0",X"F0",X"E0",X"E0",X"E0",X"A0",X"20",X"20",X"A0",X"A0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"06",X"06",
		X"0F",X"0F",X"0F",X"0E",X"0F",X"07",X"03",X"03",X"02",X"00",X"00",X"E1",X"E2",X"12",X"12",X"14",
		X"F0",X"F0",X"F0",X"70",X"70",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",
		X"7F",X"7F",X"3C",X"38",X"18",X"1C",X"0F",X"07",X"03",X"07",X"06",X"06",X"06",X"06",X"03",X"03",
		X"F8",X"B0",X"F0",X"E0",X"E0",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"70",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"86",X"C6",X"7E",X"7E",X"7E",
		X"03",X"03",X"10",X"22",X"62",X"E4",X"87",X"0C",X"08",X"00",X"11",X"1B",X"3C",X"3E",X"3E",X"7F",
		X"E0",X"E0",X"C0",X"00",X"00",X"80",X"08",X"10",X"30",X"60",X"C0",X"00",X"40",X"00",X"00",X"00",
		X"1F",X"1F",X"1E",X"1E",X"0F",X"0F",X"0F",X"06",X"06",X"0E",X"0C",X"0C",X"0C",X"0C",X"04",X"06",
		X"E4",X"FC",X"FC",X"7C",X"78",X"78",X"78",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"07",X"0F",X"1F",X"1F",X"1F",X"1E",X"1F",X"0F",X"0C",X"04",X"06",X"0F",X"07",X"00",X"04",X"38",
		X"80",X"C0",X"F0",X"E0",X"F0",X"C0",X"A0",X"A0",X"C0",X"00",X"00",X"80",X"00",X"10",X"20",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"F8",X"FF",X"7F",X"3F",X"0F",X"03",X"01",X"07",X"0F",X"1F",X"1F",X"1E",X"3A",X"37",X"6F",
		X"00",X"00",X"80",X"F8",X"DC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"6F",X"6F",X"DF",X"EF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"7F",X"FF",X"FE",X"FE",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"12",X"0E",X"0C",X"19",X"00",X"30",X"60",X"C2",X"C3",X"C0",X"C2",X"C7",X"EC",X"EF",
		X"80",X"00",X"00",X"40",X"80",X"00",X"20",X"30",X"18",X"0C",X"0E",X"07",X"0F",X"9F",X"1E",X"8C",
		X"38",X"3C",X"3C",X"3C",X"18",X"18",X"1E",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"60",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"40",X"40",X"40",X"C0",X"A0",X"A0",X"60",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"03",X"05",X"04",X"06",X"04",X"02",X"01",X"01",X"03",X"00",X"04",X"0C",X"08",X"18",
		X"F8",X"F8",X"78",X"A8",X"10",X"10",X"00",X"40",X"D0",X"A0",X"48",X"0C",X"07",X"03",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"04",X"06",X"02",X"02",X"02",X"02",X"03",X"03",X"03",
		X"3E",X"3C",X"3C",X"3C",X"78",X"78",X"F8",X"70",X"70",X"60",X"60",X"60",X"60",X"30",X"30",X"30",
		X"00",X"00",X"07",X"FF",X"FE",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"13",X"0F",X"18",X"00",X"0F",X"70",X"8F",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",X"1F",X"0C",X"30",X"C0",X"00",X"00",
		X"04",X"06",X"06",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",
		X"04",X"06",X"06",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"C0",X"81",X"80",X"00",
		X"0C",X"0E",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E8",X"F0",X"D0",X"80",
		X"0C",X"0E",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"D8",X"E8",X"E0",X"C0",X"80",
		X"03",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"FE",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"00",X"3F",X"3F",X"1F",X"1F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"00",X"FC",X"FC",X"F8",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"03",X"FF",X"FF",X"7F",X"7F",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"FE",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"FF",X"3F",X"3F",X"1F",X"1F",X"39",X"1D",X"1F",X"1F",X"1F",X"0F",X"06",X"00",X"00",
		X"88",X"92",X"D0",X"D8",X"D0",X"D0",X"E0",X"E0",X"C0",X"08",X"08",X"F0",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"00",X"83",X"67",X"0F",X"0F",X"0F",X"07",X"07",X"0E",X"07",X"07",X"07",X"03",X"00",X"00",
		X"01",X"01",X"E1",X"E1",X"F2",X"F2",X"F2",X"F6",X"F4",X"74",X"63",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",
		X"07",X"1F",X"1F",X"0F",X"0F",X"0F",X"2F",X"1F",X"0F",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"80",X"C0",X"C0",X"C4",X"C8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",
		X"07",X"1F",X"1F",X"0F",X"0F",X"0F",X"2F",X"1F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"C0",X"C0",X"C0",X"C4",X"C8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"10",X"18",X"31",X"38",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"00",
		X"04",X"04",X"84",X"80",X"88",X"F0",X"00",X"F0",X"F0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F0",X"00",
		X"0F",X"0F",X"0F",X"0E",X"4F",X"57",X"07",X"4B",X"47",X"60",X"20",X"30",X"18",X"1C",X"34",X"38",
		X"F0",X"F0",X"F0",X"70",X"6C",X"F8",X"C0",X"80",X"00",X"02",X"04",X"84",X"88",X"98",X"F0",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0C",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"07",X"07",X"3B",X"67",X"00",X"00",X"C0",X"70",X"10",X"00",X"08",X"0D",X"1D",X"3F",X"3F",X"3F",
		X"E0",X"C0",X"9C",X"06",X"00",X"00",X"83",X"8E",X"88",X"80",X"00",X"90",X"B0",X"F0",X"E0",X"E0",
		X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"E0",X"E0",X"60",X"20",X"20",X"20",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"E0",X"E0",X"E0",
		X"00",X"00",X"80",X"80",X"C0",X"70",X"70",X"18",X"08",X"1D",X"3D",X"3F",X"3F",X"3E",X"38",X"3C",
		X"00",X"00",X"00",X"80",X"84",X"8E",X"8E",X"00",X"C0",X"C0",X"F0",X"E0",X"80",X"80",X"C0",X"E0",
		X"0E",X"0E",X"06",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"60",X"60",X"60",X"60",X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0C",X"0C",X"0C",X"0C",X"6C",X"3E",X"1E",X"1F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"30",X"3C",X"3F",X"7F",X"7F",X"EF",X"CF",X"C7",X"47",X"67",X"3F",X"00",X"00",X"80",X"E2",
		X"60",X"E0",X"20",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",X"A0",X"20",X"30",X"10",X"10",X"10",X"10",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"70",X"70",X"70",X"30",X"30",X"B0",X"B0",X"B0",X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"02",X"03",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"7C",X"7C",X"F8",X"F8",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"1F",X"03",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FE",X"FC",X"FC",X"F8",X"F8",X"18",X"00",X"00",X"00",X"50",X"79",X"3F",X"3F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"84",X"C6",X"C6",X"E6",
		X"0E",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3E",X"3E",X"3C",X"18",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"3C",X"70",X"70",X"70",X"30",X"3B",X"3F",X"1F",X"3A",X"36",X"64",X"60",X"01",X"01",X"01",
		X"F1",X"61",X"20",X"40",X"70",X"F8",X"F0",X"C2",X"00",X"00",X"18",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"3F",X"7F",X"FF",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"E7",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"7F",X"3F",X"7F",X"1B",X"2D",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"40",X"80",
		X"5E",X"1E",X"3C",X"2C",X"2C",X"2E",X"07",X"00",X"3C",X"78",X"70",X"70",X"38",X"38",X"18",X"18",
		X"10",X"10",X"48",X"08",X"08",X"38",X"C0",X"08",X"10",X"10",X"30",X"70",X"F0",X"E0",X"60",X"60",
		X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"7C",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",
		X"38",X"38",X"70",X"71",X"7B",X"77",X"77",X"77",X"07",X"03",X"0C",X"0F",X"0E",X"0E",X"0C",X"0C",
		X"80",X"71",X"C1",X"E1",X"DC",X"80",X"10",X"02",X"02",X"C3",X"7F",X"00",X"01",X"07",X"0E",X"1E",
		X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"B0",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FE",X"FE",X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0D",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
