library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity draw_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of draw_bg_bits_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"BF",X"FE",X"BE",X"BE",X"AA",X"FE",X"AB",X"FA",X"AF",X"EA",X"BF",X"AA",X"BE",X"BE",X"BF",X"FE",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7D",X"55",X"7D",X"55",X"55",
		X"55",X"55",X"57",X"55",X"5D",X"D5",X"75",X"75",X"FF",X"FD",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"5D",X"D5",X"55",X"D5",X"55",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"55",X"FF",X"D5",X"D5",X"55",X"D5",X"55",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"FF",X"D5",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"D7",X"FD",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"FF",X"FD",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"55",X"FD",X"55",X"75",X"55",X"75",X"D5",X"75",X"D5",X"75",X"FF",X"F5",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D5",X"75",X"FF",X"D5",X"D5",X"75",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"5D",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"F5",X"7D",X"DD",X"DD",X"D7",X"5D",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"F5",X"5D",X"DD",X"5D",X"D7",X"5D",X"D5",X"DD",X"D5",X"7D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"BF",X"FE",X"BE",X"BE",X"AA",X"FE",X"AB",X"FA",X"AF",X"EA",X"BF",X"AA",X"BE",X"BE",X"BF",X"FE",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"FF",X"FD",X"55",X"5D",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D7",X"5D",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"75",X"75",X"75",X"75",X"5D",X"D5",X"5D",X"D5",X"57",X"55",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D7",X"5D",X"D7",X"5D",X"DD",X"DD",X"DD",X"DD",X"75",X"75",X"55",X"55",
		X"55",X"55",X"F5",X"7D",X"7D",X"F5",X"5F",X"D5",X"7D",X"F5",X"F5",X"7D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"75",X"75",X"5D",X"D5",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",
		X"55",X"D5",X"7F",X"FD",X"75",X"D5",X"7F",X"FD",X"55",X"DD",X"55",X"DD",X"7F",X"FD",X"55",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"53",X"FF",X"4F",X"FF",X"3F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"95",X"FF",X"C5",X"FF",X"F1",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"4F",X"FF",X"53",X"FF",X"54",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FC",X"FF",X"F1",X"FF",X"C5",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"BF",X"FE",X"BE",X"BE",X"AA",X"FE",X"AB",X"FA",X"AF",X"EA",X"BF",X"AA",X"BE",X"BE",X"BF",X"FE",
		X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"51",X"55",X"45",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"51",X"55",X"45",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"15",X"55",X"45",X"55",X"51",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"45",X"55",X"51",X"55",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"40",X"00",X"00",
		X"54",X"00",X"53",X"FF",X"4F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"15",X"FF",X"C5",X"FF",X"F1",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"4F",X"FF",X"53",X"FF",X"54",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F1",X"FF",X"C5",X"00",X"15",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"40",X"00",X"01",
		X"00",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"15",X"55",
		X"55",X"55",X"55",X"75",X"55",X"F5",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"55",X"5D",X"7F",X"FD",X"D5",X"55",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"5D",X"57",X"F5",X"55",X"5D",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"55",X"75",X"D5",X"75",X"D5",X"75",X"FF",X"FD",X"55",X"75",X"55",X"75",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"FF",X"FD",X"55",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"7F",X"FD",X"D5",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"7F",X"F5",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"7F",X"FD",X"55",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"BF",X"FE",X"BE",X"BE",X"AA",X"FE",X"AB",X"FA",X"AF",X"EA",X"BF",X"AA",X"BE",X"BE",X"BF",X"FE",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"FF",X"55",X"D5",X"55",X"D5",X"55",X"55",
		X"55",X"55",X"5D",X"FF",X"5D",X"D5",X"5D",X"FF",X"FD",X"D5",X"5D",X"D5",X"5D",X"FF",X"55",X"55",
		X"55",X"55",X"F5",X"D5",X"55",X"D5",X"D5",X"D5",X"55",X"D5",X"55",X"D5",X"FD",X"FF",X"55",X"55",
		X"55",X"55",X"55",X"FF",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"5D",X"D5",X"FD",X"FF",X"55",X"55",
		X"55",X"55",X"F5",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"01",X"55",
		X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"05",X"55",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"00",X"55",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",
		X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"01",X"55",X"00",X"55",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"00",X"15",X"00",X"15",X"00",X"55",X"01",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"55",X"5D",X"D5",X"75",X"75",X"FF",X"FD",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"5D",X"D5",X"55",X"D5",X"55",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"55",X"FF",X"D5",X"D5",X"55",X"D5",X"55",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"55",X"FF",X"D5",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"D5",X"FD",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"FF",X"FD",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"5F",X"FD",X"55",X"75",X"55",X"75",X"D5",X"75",X"D5",X"75",X"7F",X"D5",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D5",X"75",X"FF",X"D5",X"D5",X"75",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"F5",X"7D",X"DD",X"DD",X"D7",X"5D",X"D5",X"5D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"F5",X"5D",X"DD",X"5D",X"D7",X"5D",X"D5",X"DD",X"D5",X"7D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"FF",X"F5",X"D5",X"75",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"FF",X"FD",X"55",X"5D",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"75",X"75",X"75",X"75",X"5D",X"D5",X"5D",X"D5",X"57",X"55",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"D7",X"5D",X"D7",X"5D",X"D7",X"5D",X"DD",X"DD",X"75",X"75",X"55",X"55",
		X"55",X"55",X"D5",X"5D",X"75",X"75",X"5D",X"D5",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",
		X"55",X"55",X"F5",X"7D",X"7D",X"F5",X"5F",X"D5",X"7D",X"F5",X"F5",X"7D",X"D5",X"5D",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"55",X"75",X"55",X"F5",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"55",X"5D",X"7F",X"FD",X"D5",X"55",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"5D",X"57",X"F5",X"55",X"5D",X"D5",X"5D",X"FF",X"FD",X"55",X"55",
		X"55",X"55",X"55",X"75",X"D5",X"75",X"D5",X"75",X"FF",X"FD",X"55",X"75",X"55",X"75",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"55",X"FF",X"FD",X"55",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"7F",X"FD",X"D5",X"55",X"FF",X"F5",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"FF",X"FD",X"D5",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"7F",X"F5",X"D5",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"7F",X"F5",X"D5",X"5D",X"7F",X"FD",X"55",X"5D",X"D5",X"5D",X"7F",X"F5",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7D",X"55",X"7D",X"55",X"55",
		X"57",X"55",X"7F",X"FD",X"77",X"55",X"7F",X"FD",X"57",X"5D",X"57",X"5D",X"7F",X"FD",X"57",X"55",
		X"AA",X"95",X"AA",X"A5",X"A5",X"A9",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",
		X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"A9",X"AA",X"A5",X"AA",X"95",
		X"AA",X"A9",X"AA",X"A9",X"A5",X"69",X"A5",X"69",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"A5",
		X"AA",X"A5",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"69",X"A5",X"69",X"AA",X"A9",X"AA",X"A9",
		X"5A",X"95",X"6A",X"A5",X"69",X"A5",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"AA",X"A9",
		X"AA",X"A9",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"AA",X"95",X"AA",X"A5",X"A5",X"A9",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A5",X"69",X"AA",X"A5",
		X"A5",X"5A",X"A5",X"5A",X"A5",X"5A",X"A5",X"5A",X"A6",X"9A",X"A6",X"9A",X"A6",X"9A",X"A6",X"9A",
		X"A6",X"9A",X"A6",X"9A",X"AA",X"AA",X"AA",X"AA",X"A9",X"6A",X"A9",X"6A",X"A5",X"5A",X"A5",X"5A",
		X"AA",X"A9",X"AA",X"A9",X"A5",X"69",X"A5",X"69",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"A9",
		X"AA",X"A9",X"55",X"69",X"55",X"69",X"55",X"69",X"A5",X"69",X"A5",X"69",X"AA",X"A9",X"AA",X"A9",
		X"AA",X"AA",X"AA",X"AA",X"96",X"96",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",
		X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",
		X"A5",X"69",X"A5",X"69",X"A5",X"69",X"A9",X"69",X"A9",X"69",X"A9",X"69",X"AA",X"69",X"A6",X"69",
		X"A6",X"69",X"A6",X"A9",X"A5",X"A9",X"A5",X"A9",X"A5",X"A9",X"A5",X"69",X"A5",X"69",X"A5",X"69",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"69",X"A5",X"69",X"AA",X"A9",X"AA",X"A9",
		X"5F",X"D5",X"7F",X"F5",X"FD",X"FD",X"F5",X"7D",X"F5",X"55",X"FD",X"55",X"7F",X"55",X"5F",X"D5",
		X"57",X"F5",X"55",X"FD",X"55",X"7D",X"F5",X"7D",X"F5",X"7D",X"FD",X"FD",X"7F",X"F5",X"5F",X"D5",
		X"FF",X"FF",X"FF",X"FF",X"D7",X"D7",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"FD",X"7D",X"FD",X"7D",X"FD",X"7D",X"FF",X"7D",X"F7",X"7D",
		X"F7",X"7D",X"F7",X"FD",X"F5",X"FD",X"F5",X"FD",X"F5",X"FD",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",
		X"5F",X"D5",X"5F",X"D5",X"7D",X"F5",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"FF",X"FD",
		X"FF",X"FD",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",
		X"FF",X"55",X"FF",X"D5",X"F5",X"F5",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",
		X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"FD",X"FF",X"F5",X"FF",X"D5",
		X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"55",X"00",X"55",
		X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",X"55",X"55",X"55",X"55",
		X"55",X"F5",X"57",X"F5",X"5F",X"F5",X"5F",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",
		X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"5F",X"D5",X"7F",X"F5",X"FD",X"FD",X"F5",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"F5",
		X"57",X"F5",X"5F",X"D5",X"7F",X"55",X"FD",X"55",X"F5",X"55",X"F5",X"7D",X"FF",X"FD",X"FF",X"FD",
		X"5F",X"D5",X"7F",X"F5",X"FD",X"FD",X"F5",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"FD",X"5F",X"F5",
		X"5F",X"F5",X"55",X"FD",X"55",X"7D",X"55",X"7D",X"F5",X"7D",X"FD",X"FD",X"7F",X"F5",X"5F",X"D5",
		X"55",X"F5",X"55",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",
		X"FF",X"FD",X"FF",X"FD",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",
		X"FF",X"FD",X"FF",X"FD",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F7",X"D5",X"FF",X"F5",
		X"FD",X"FD",X"F5",X"7D",X"55",X"7D",X"55",X"7D",X"F5",X"7D",X"FD",X"FD",X"7F",X"F5",X"5F",X"D5",
		X"50",X"15",X"40",X"05",X"01",X"01",X"05",X"41",X"05",X"41",X"05",X"55",X"05",X"55",X"00",X"15",
		X"00",X"05",X"01",X"01",X"05",X"41",X"05",X"41",X"05",X"41",X"01",X"01",X"40",X"05",X"50",X"15",
		X"00",X"01",X"00",X"01",X"05",X"41",X"05",X"41",X"55",X"41",X"55",X"05",X"55",X"05",X"55",X"05",
		X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",
		X"50",X"15",X"40",X"05",X"01",X"01",X"05",X"41",X"05",X"41",X"01",X"01",X"40",X"05",X"50",X"15",
		X"40",X"05",X"01",X"01",X"05",X"41",X"05",X"41",X"05",X"41",X"01",X"01",X"40",X"05",X"50",X"15",
		X"50",X"15",X"40",X"05",X"01",X"01",X"05",X"41",X"05",X"41",X"05",X"41",X"01",X"01",X"40",X"01",
		X"50",X"01",X"55",X"41",X"55",X"41",X"05",X"41",X"05",X"41",X"01",X"01",X"40",X"01",X"50",X"05",
		X"50",X"15",X"40",X"05",X"01",X"01",X"05",X"41",X"05",X"41",X"05",X"41",X"05",X"41",X"05",X"41",
		X"05",X"41",X"05",X"41",X"05",X"41",X"05",X"41",X"05",X"41",X"01",X"01",X"40",X"05",X"50",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"05",X"54",X"05",X"54",X"05",
		X"50",X"15",X"40",X"05",X"00",X"01",X"04",X"41",X"04",X"41",X"04",X"55",X"00",X"05",X"40",X"01",
		X"54",X"41",X"04",X"41",X"00",X"01",X"00",X"01",X"40",X"05",X"50",X"15",X"55",X"55",X"55",X"55",
		X"FD",X"FD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"FD",X"FD",X"5D",X"D5",X"FD",X"FD",X"D5",X"5D",X"D5",X"5D",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"FD",X"FD",X"D5",X"DD",X"FD",X"DD",X"5D",X"DD",X"5D",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"FD",X"FD",X"5D",X"D5",X"5D",X"FD",X"5D",X"5D",X"5D",X"5D",X"5D",X"FD",X"55",X"55",X"FF",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"55",X"55",X"55",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FD",X"FD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",X"55",X"55",
		X"FF",X"D5",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"FD",X"FD",X"7D",X"F5",
		X"5F",X"D5",X"5F",X"D5",X"5F",X"D5",X"5F",X"D5",X"5F",X"D5",X"5F",X"D5",X"5F",X"D5",X"5F",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",
		X"55",X"55",X"55",X"55",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"55",X"55",X"55",X"55",X"95",X"95",X"95",X"A9",X"95",X"55",X"95",X"55",X"95",X"95",X"95",X"95",
		X"55",X"55",X"55",X"56",X"95",X"56",X"99",X"5A",X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"59",
		X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"5A",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"95",X"95",X"95",X"95",X"55",X"95",X"55",X"9A",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"53",X"FF",X"4F",X"FF",X"3F",X"FF",X"3A",X"BF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FC",X"00",X"F3",X"FF",X"CF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FD",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FD",X"FD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"55",X"55",X"FD",X"FD",X"5D",X"D5",X"FD",X"FD",X"D5",X"5D",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"55",X"55",X"FD",X"FD",X"D5",X"DD",X"FD",X"DD",X"5D",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"5F",X"D5",X"7F",X"F5",X"FD",X"FD",X"F5",X"7D",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"7D",X"FD",X"FD",X"7F",X"F5",X"5F",X"D5",
		X"5F",X"D5",X"7F",X"F5",X"FD",X"FD",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",
		X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"FD",X"FD",X"7F",X"F5",X"5F",X"D5",
		X"7F",X"FD",X"7F",X"FD",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"7F",X"FD",X"7F",X"FD",
		X"FF",X"D5",X"FF",X"F5",X"F5",X"FD",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"FD",X"FF",X"F5",
		X"FF",X"F5",X"F5",X"FD",X"F5",X"7D",X"F5",X"7D",X"F5",X"7D",X"F5",X"FD",X"FF",X"F5",X"FF",X"D5",
		X"FF",X"FD",X"FF",X"FD",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"FF",X"F5",
		X"FF",X"F5",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"FF",X"FD",X"FF",X"FD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"F5",X"75",X"5D",X"D7",X"D7",X"DD",X"57",X"DD",X"57",X"D7",X"D7",X"75",X"5D",X"5F",X"F5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"54",X"00",X"54",X"15",X"54",X"15",X"54",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"54",X"15",X"54",X"15",X"54",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"15",X"00",X"15",X"54",X"15",X"54",X"15",X"54",X"15",
		X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"15",
		X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"00",X"54",X"00",X"54",X"15",X"54",X"15",X"54",X"15",
		X"54",X"15",X"54",X"15",X"54",X"15",X"00",X"00",X"00",X"00",X"54",X"15",X"54",X"15",X"54",X"15",
		X"54",X"15",X"54",X"15",X"54",X"15",X"00",X"15",X"00",X"15",X"54",X"15",X"54",X"15",X"54",X"15",
		X"54",X"15",X"54",X"15",X"54",X"15",X"54",X"00",X"54",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"15",X"54",X"15",X"54",X"15",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"15",X"54",X"15",X"54",X"15",X"00",X"15",X"00",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FD",X"FD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"55",X"55",X"FD",X"FD",X"5D",X"D5",X"FD",X"FD",X"D5",X"5D",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"55",X"55",X"FD",X"FD",X"D5",X"DD",X"FD",X"DD",X"5D",X"DD",X"FD",X"FD",X"55",X"55",X"FF",X"FD",
		X"55",X"55",X"FD",X"FD",X"5D",X"D5",X"5D",X"FD",X"5D",X"5D",X"5D",X"FD",X"55",X"55",X"FF",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
