library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"C0",X"4F",X"C3",X"0A",X"01",X"FF",X"77",X"23",X"32",X"C0",X"50",X"10",X"F9",X"0D",
		X"20",X"F6",X"C9",X"3A",X"76",X"4C",X"3D",X"C9",X"D5",X"11",X"20",X"00",X"19",X"D1",X"C9",X"FF",
		X"D5",X"11",X"E0",X"FF",X"19",X"D1",X"C9",X"FF",X"E1",X"87",X"85",X"6F",X"3E",X"00",X"8C",X"67",
		X"7E",X"5F",X"23",X"7E",X"57",X"EB",X"E9",X"FF",X"F5",X"E5",X"D5",X"C5",X"DD",X"E5",X"FD",X"E5",
		X"AF",X"32",X"00",X"50",X"DD",X"21",X"00",X"4C",X"CD",X"6A",X"00",X"DD",X"23",X"CD",X"00",X"02",
		X"DD",X"23",X"CD",X"50",X"02",X"32",X"C0",X"50",X"CD",X"24",X"03",X"FB",X"3E",X"01",X"32",X"00",
		X"50",X"FD",X"E1",X"DD",X"E1",X"C1",X"D1",X"E1",X"F1",X"C9",X"DD",X"7E",X"00",X"CB",X"47",X"28",
		X"2C",X"21",X"0F",X"4C",X"11",X"51",X"50",X"01",X"05",X"00",X"ED",X"B0",X"DD",X"7E",X"1E",X"32",
		X"45",X"50",X"DD",X"7E",X"13",X"A7",X"28",X"06",X"CD",X"D6",X"8A",X"DD",X"77",X"13",X"DD",X"7E",
		X"21",X"3D",X"DD",X"77",X"21",X"C0",X"00",X"00",X"DD",X"CB",X"00",X"86",X"C9",X"CB",X"4F",X"20",
		X"0C",X"2A",X"03",X"4C",X"22",X"05",X"4C",X"3E",X"02",X"DD",X"77",X"00",X"C9",X"2A",X"05",X"4C",
		X"CD",X"BE",X"00",X"A7",X"28",X"F3",X"22",X"05",X"4C",X"DD",X"CB",X"00",X"C6",X"C9",X"7C",X"A7",
		X"20",X"03",X"C3",X"EC",X"02",X"7E",X"FE",X"10",X"20",X"02",X"AF",X"C9",X"DD",X"77",X"1E",X"DD",
		X"E5",X"C1",X"0C",X"11",X"0A",X"4C",X"13",X"13",X"13",X"13",X"13",X"0D",X"20",X"F8",X"23",X"06",
		X"02",X"7E",X"4F",X"CD",X"9E",X"02",X"E6",X"0F",X"12",X"13",X"79",X"12",X"13",X"23",X"10",X"F1",
		X"7E",X"12",X"23",X"7E",X"CD",X"3C",X"32",X"23",X"3E",X"01",X"C9",X"0F",X"0F",X"0F",X"0F",X"C9",
		X"21",X"00",X"40",X"01",X"04",X"00",X"3E",X"40",X"CF",X"C9",X"CD",X"00",X"01",X"00",X"36",X"00",
		X"23",X"32",X"C0",X"50",X"7C",X"FE",X"48",X"20",X"F5",X"21",X"00",X"40",X"01",X"04",X"00",X"3E",
		X"80",X"CF",X"21",X"00",X"44",X"3E",X"12",X"01",X"04",X"00",X"CF",X"21",X"00",X"4C",X"AF",X"01",
		X"02",X"00",X"CF",X"21",X"00",X"50",X"36",X"00",X"23",X"7C",X"FE",X"51",X"20",X"F8",X"CD",X"21",
		X"32",X"00",X"00",X"00",X"00",X"00",X"3E",X"01",X"32",X"01",X"50",X"3E",X"01",X"32",X"00",X"50",
		X"18",X"4E",X"20",X"03",X"3E",X"20",X"B0",X"21",X"2D",X"4C",X"CB",X"CE",X"32",X"2E",X"4C",X"C9",
		X"0B",X"00",X"3A",X"00",X"50",X"E6",X"0F",X"FE",X"0E",X"28",X"27",X"FE",X"0B",X"28",X"26",X"FE",
		X"07",X"28",X"25",X"FE",X"0D",X"28",X"24",X"3E",X"0F",X"32",X"2E",X"4C",X"3A",X"40",X"50",X"CB",
		X"47",X"CA",X"AD",X"06",X"21",X"2D",X"4C",X"CB",X"8E",X"3A",X"47",X"4C",X"C3",X"5A",X"11",X"00",
		X"00",X"11",X"3E",X"00",X"11",X"3E",X"01",X"11",X"3E",X"02",X"11",X"3E",X"03",X"C3",X"A4",X"02",
		X"ED",X"56",X"FB",X"00",X"00",X"00",X"CD",X"13",X"90",X"CD",X"00",X"90",X"CD",X"1E",X"35",X"00",
		X"00",X"CD",X"62",X"80",X"18",X"F0",X"CD",X"BF",X"01",X"CD",X"BF",X"01",X"CD",X"BF",X"01",X"3E",
		X"80",X"32",X"2C",X"4C",X"32",X"C0",X"50",X"3A",X"26",X"4C",X"A7",X"C2",X"0D",X"90",X"3A",X"2C",
		X"4C",X"A7",X"20",X"F3",X"C9",X"1A",X"47",X"13",X"1A",X"FE",X"FF",X"C8",X"CD",X"E2",X"01",X"2B",
		X"18",X"F5",X"D5",X"E5",X"11",X"00",X"04",X"19",X"70",X"E1",X"D1",X"77",X"C9",X"1A",X"47",X"13",
		X"1A",X"FE",X"FF",X"C8",X"CD",X"E2",X"01",X"C5",X"01",X"20",X"00",X"ED",X"42",X"C1",X"18",X"EF",
		X"DD",X"7E",X"00",X"CB",X"47",X"28",X"2C",X"CB",X"C7",X"21",X"14",X"4C",X"11",X"56",X"50",X"01",
		X"05",X"00",X"ED",X"B0",X"3A",X"2F",X"4C",X"32",X"4A",X"50",X"DD",X"7E",X"17",X"A7",X"28",X"06",
		X"CD",X"D6",X"8A",X"DD",X"77",X"17",X"DD",X"7E",X"21",X"3D",X"DD",X"77",X"21",X"C0",X"DD",X"CB",
		X"00",X"86",X"C9",X"CB",X"4F",X"20",X"09",X"2A",X"07",X"4C",X"22",X"09",X"4C",X"C3",X"2C",X"04",
		X"2A",X"09",X"4C",X"CD",X"BE",X"00",X"A7",X"CA",X"A9",X"00",X"22",X"09",X"4C",X"C3",X"B9",X"00",
		X"DD",X"7E",X"00",X"CB",X"47",X"28",X"2A",X"21",X"19",X"4C",X"11",X"5B",X"50",X"01",X"05",X"00",
		X"ED",X"B0",X"DD",X"7E",X"1E",X"32",X"4F",X"50",X"DD",X"7E",X"1B",X"A7",X"28",X"06",X"CD",X"D6",
		X"8A",X"DD",X"77",X"1B",X"DD",X"7E",X"21",X"3D",X"DD",X"77",X"21",X"C0",X"DD",X"CB",X"00",X"86",
		X"C9",X"CB",X"4F",X"20",X"09",X"2A",X"0B",X"4C",X"22",X"0D",X"4C",X"C3",X"A7",X"00",X"2A",X"0D",
		X"4C",X"CD",X"BE",X"00",X"A7",X"CA",X"38",X"04",X"22",X"0D",X"4C",X"C3",X"B9",X"00",X"32",X"C0",
		X"50",X"C3",X"FB",X"00",X"47",X"3A",X"40",X"50",X"CB",X"47",X"C2",X"B4",X"06",X"3A",X"2D",X"4C",
		X"CB",X"4F",X"78",X"C3",X"52",X"01",X"3A",X"40",X"50",X"CB",X"6F",X"20",X"15",X"3A",X"24",X"4C",
		X"CB",X"67",X"C0",X"CB",X"E7",X"CD",X"09",X"03",X"00",X"E6",X"10",X"06",X"0F",X"B0",X"32",X"24",
		X"4C",X"C9",X"3A",X"24",X"4C",X"CB",X"A7",X"A7",X"C8",X"00",X"3D",X"32",X"24",X"4C",X"21",X"1D",
		X"80",X"22",X"0B",X"4C",X"C9",X"21",X"00",X"00",X"22",X"0B",X"4C",X"C9",X"7D",X"A7",X"C2",X"C5",
		X"00",X"DD",X"E5",X"C1",X"0C",X"11",X"50",X"50",X"13",X"13",X"13",X"13",X"13",X"0D",X"20",X"F8",
		X"21",X"27",X"4C",X"01",X"01",X"00",X"ED",X"B0",X"C9",X"F5",X"3A",X"25",X"4C",X"3C",X"32",X"25",
		X"4C",X"47",X"3A",X"80",X"50",X"E6",X"03",X"3C",X"B8",X"20",X"07",X"21",X"26",X"4C",X"34",X"2B",
		X"36",X"00",X"F1",X"C9",X"CD",X"B6",X"02",X"CD",X"F2",X"06",X"CD",X"00",X"80",X"35",X"3A",X"26",
		X"4C",X"FE",X"0A",X"30",X"05",X"21",X"14",X"40",X"77",X"C9",X"3E",X"46",X"18",X"F7",X"01",X"54",
		X"48",X"41",X"4E",X"4B",X"40",X"59",X"4F",X"55",X"40",X"5B",X"FF",X"02",X"01",X"40",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"40",X"50",X"55",X"53",X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",
		X"5B",X"5B",X"FF",X"07",X"54",X"48",X"49",X"53",X"40",X"4D",X"41",X"43",X"48",X"49",X"4E",X"45",
		X"FF",X"07",X"49",X"53",X"FF",X"07",X"4F",X"4E",X"4C",X"59",X"40",X"4F",X"4E",X"45",X"40",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"FF",X"06",X"48",X"41",X"4E",X"53",X"48",X"49",X"4E",X"40",X"47",
		X"4F",X"52",X"41",X"4B",X"55",X"FF",X"0F",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"FF",X"07",
		X"40",X"40",X"42",X"59",X"40",X"26",X"50",X"45",X"4E",X"49",X"26",X"FF",X"3E",X"03",X"84",X"42",
		X"4B",X"03",X"09",X"43",X"63",X"03",X"AD",X"42",X"71",X"03",X"0F",X"42",X"75",X"03",X"D1",X"42",
		X"86",X"03",X"7D",X"43",X"9F",X"03",X"BD",X"41",X"E7",X"03",X"DF",X"40",X"FF",X"FF",X"DB",X"3A",
		X"D5",X"0A",X"5F",X"03",X"0A",X"57",X"03",X"0A",X"6F",X"03",X"0A",X"67",X"C5",X"CD",X"ED",X"01",
		X"C1",X"D1",X"03",X"15",X"20",X"EA",X"C9",X"0F",X"01",X"09",X"08",X"03",X"FF",X"31",X"C0",X"4F",
		X"CD",X"00",X"01",X"01",X"AC",X"03",X"16",X"08",X"CD",X"D0",X"03",X"21",X"1B",X"40",X"11",X"96",
		X"03",X"CD",X"D5",X"01",X"3A",X"2C",X"4C",X"CB",X"5F",X"20",X"1D",X"3E",X"06",X"21",X"7D",X"47",
		X"06",X"0E",X"77",X"11",X"20",X"00",X"ED",X"52",X"10",X"F8",X"3A",X"40",X"50",X"CB",X"77",X"20",
		X"E3",X"21",X"26",X"4C",X"35",X"C3",X"41",X"04",X"3E",X"02",X"18",X"E1",X"F5",X"ED",X"5F",X"E6",
		X"07",X"32",X"2F",X"4C",X"F1",X"C3",X"A7",X"00",X"21",X"00",X"00",X"22",X"0B",X"4C",X"C3",X"A9",
		X"00",X"CD",X"9D",X"06",X"AF",X"77",X"23",X"77",X"23",X"77",X"CD",X"D7",X"04",X"3A",X"80",X"50",
		X"E6",X"0C",X"0F",X"0F",X"3C",X"32",X"3F",X"4C",X"CD",X"93",X"20",X"18",X"77",X"CD",X"DD",X"9A",
		X"00",X"EF",X"72",X"04",X"2E",X"09",X"3A",X"09",X"6F",X"94",X"46",X"09",X"46",X"09",X"46",X"09",
		X"46",X"09",X"CD",X"74",X"20",X"22",X"41",X"4C",X"21",X"DC",X"43",X"11",X"C3",X"04",X"CD",X"D5",
		X"01",X"21",X"D4",X"43",X"11",X"CA",X"04",X"CD",X"D5",X"01",X"21",X"40",X"44",X"3E",X"0E",X"CD",
		X"7C",X"20",X"CF",X"21",X"40",X"40",X"ED",X"5B",X"41",X"4C",X"01",X"02",X"C0",X"C5",X"D5",X"1A",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"F6",X"F0",X"77",X"13",X"23",X"10",X"F2",X"0D",X"20",X"EF",
		X"D1",X"C1",X"1A",X"E6",X"0F",X"F6",X"F0",X"77",X"13",X"23",X"10",X"F6",X"0D",X"20",X"F3",X"CD",
		X"20",X"14",X"C9",X"0F",X"53",X"43",X"4F",X"52",X"45",X"FF",X"0F",X"48",X"49",X"40",X"53",X"43",
		X"4F",X"52",X"45",X"FF",X"C3",X"BD",X"06",X"3E",X"01",X"32",X"40",X"4C",X"C9",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"00",X"00",X"0C",X"0E",X"BE",X"0E",X"0E",X"0B",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"BB",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"A0",X"00",X"00",X"0A",X"00",X"B0",X"00",X"00",X"0D",
		X"0F",X"8F",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"00",X"0D",X"0F",X"0F",X"BB",X"00",X"00",X"0D",
		X"0F",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0C",
		X"0E",X"7E",X"0E",X"0E",X"0B",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0E",X"BB",X"00",X"00",X"0C",
		X"0E",X"0E",X"0E",X"0B",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"F9",X"F0",X"D0",X"F0",X"F0",X"0A",
		X"00",X"00",X"00",X"00",X"0D",X"0F",X"0F",X"0F",X"0F",X"0B",X"00",X"00",X"BB",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"C9",X"E0",X"E0",X"ED",X"EF",X"CF",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0E",X"0B",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"AB",X"00",X"00",X"0E",X"0E",X"AE",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"0B",X"D0",X"F0",X"F0",X"F0",X"BA",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"9D",X"0F",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"D9",
		X"F0",X"F0",X"F0",X"F0",X"FA",X"C0",X"E0",X"E0",X"E0",X"D0",X"F0",X"F0",X"BB",X"00",X"00",X"00",
		X"09",X"00",X"00",X"BC",X"0E",X"0E",X"0E",X"9B",X"00",X"00",X"90",X"00",X"0B",X"00",X"00",X"CB",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"B0",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"BB",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"DA",X"F0",X"F0",X"F0",X"BB",X"00",X"00",X"D0",X"F0",X"FB",X"F0",X"F0",X"BA",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"A0",X"00",X"00",X"BB",X"00",X"00",X"90",
		X"0A",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"BD",X"0F",X"0F",X"CF",X"EF",X"ED",X"EF",X"EF",X"AF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"BF",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"BB",X"00",X"00",X"D0",
		X"F0",X"F0",X"F0",X"B0",X"00",X"00",X"00",X"BC",X"0E",X"0E",X"BE",X"0E",X"0C",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"AE",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"BB",X"00",X"00",X"C0",
		X"E0",X"E0",X"E0",X"A0",X"00",X"00",X"00",X"DA",X"F0",X"F0",X"B0",X"00",X"0B",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"BB",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"B0",X"00",X"0B",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"BB",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B9",X"00",X"00",X"D0",X"F0",X"FB",X"F0",X"F0",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"BB",X"CD",X"00",X"01",
		X"21",X"1B",X"40",X"11",X"96",X"03",X"CD",X"D5",X"01",X"21",X"3C",X"4C",X"C9",X"3A",X"2E",X"4C",
		X"47",X"C3",X"AD",X"02",X"78",X"21",X"2D",X"4C",X"CB",X"8E",X"C3",X"5C",X"01",X"CD",X"12",X"0D",
		X"CD",X"01",X"07",X"CD",X"E0",X"06",X"CD",X"0C",X"0A",X"CD",X"14",X"10",X"CD",X"ED",X"13",X"CD",
		X"B7",X"16",X"C3",X"B9",X"1C",X"CD",X"62",X"01",X"3A",X"2E",X"4C",X"FE",X"0F",X"C0",X"E1",X"C9",
		X"21",X"66",X"18",X"22",X"3A",X"4C",X"21",X"20",X"0E",X"22",X"FC",X"4F",X"21",X"2D",X"4C",X"CB",
		X"C6",X"C9",X"CD",X"5F",X"07",X"21",X"30",X"4C",X"11",X"62",X"50",X"01",X"0C",X"00",X"ED",X"B0",
		X"C9",X"CD",X"C4",X"8F",X"22",X"03",X"4C",X"21",X"92",X"83",X"22",X"07",X"4C",X"C9",X"2A",X"3A",
		X"4C",X"45",X"4C",X"C5",X"79",X"3D",X"2F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"4F",X"78",X"D6",
		X"06",X"CB",X"3F",X"CB",X"3F",X"E6",X"FE",X"0F",X"0F",X"0F",X"0F",X"5F",X"E6",X"0F",X"26",X"40",
		X"B4",X"67",X"7B",X"E6",X"F0",X"B1",X"6F",X"C1",X"C9",X"F5",X"7D",X"E6",X"1F",X"CB",X"27",X"CB",
		X"27",X"CB",X"27",X"ED",X"44",X"4F",X"7C",X"E6",X"03",X"0F",X"0F",X"0F",X"0F",X"57",X"7D",X"E6",
		X"E0",X"0F",X"0F",X"0F",X"0F",X"B2",X"CB",X"27",X"CB",X"27",X"C6",X"06",X"47",X"F1",X"C9",X"3A",
		X"2D",X"4C",X"CB",X"47",X"C8",X"3A",X"43",X"4C",X"A7",X"C2",X"73",X"08",X"CD",X"7F",X"1B",X"CB",
		X"6F",X"C2",X"FF",X"1A",X"F5",X"CD",X"0E",X"07",X"22",X"45",X"4C",X"F1",X"EF",X"85",X"07",X"FD",
		X"07",X"2A",X"08",X"42",X"08",X"2A",X"45",X"4C",X"23",X"7E",X"FE",X"FC",X"28",X"04",X"FE",X"FE",
		X"C0",X"00",X"21",X"44",X"4C",X"CB",X"C6",X"AF",X"32",X"47",X"4C",X"3E",X"08",X"C3",X"C5",X"0F",
		X"28",X"3A",X"2E",X"4C",X"E6",X"0F",X"EF",X"AF",X"07",X"C4",X"07",X"D7",X"07",X"EA",X"07",X"3A",
		X"48",X"4C",X"3C",X"32",X"48",X"4C",X"CB",X"47",X"28",X"06",X"3E",X"2C",X"32",X"FC",X"4F",X"C9",
		X"3E",X"30",X"18",X"F8",X"3A",X"49",X"4C",X"3C",X"32",X"49",X"4C",X"CB",X"47",X"28",X"04",X"3E",
		X"22",X"18",X"E9",X"3E",X"26",X"18",X"E5",X"3A",X"4A",X"4C",X"3C",X"32",X"4A",X"4C",X"CB",X"47",
		X"28",X"04",X"3E",X"2C",X"18",X"D6",X"3E",X"30",X"18",X"D2",X"3A",X"4B",X"4C",X"3C",X"32",X"4B",
		X"4C",X"CB",X"47",X"28",X"04",X"3E",X"20",X"18",X"C3",X"3E",X"24",X"18",X"BF",X"2A",X"45",X"4C",
		X"23",X"23",X"CD",X"64",X"09",X"28",X"1C",X"FE",X"F6",X"CD",X"39",X"26",X"FE",X"CA",X"28",X"05",
		X"FE",X"CF",X"C2",X"91",X"1C",X"7C",X"CD",X"0A",X"09",X"CD",X"92",X"0A",X"CB",X"86",X"3E",X"01",
		X"C3",X"98",X"07",X"CD",X"D3",X"14",X"CB",X"CE",X"18",X"F4",X"CD",X"05",X"09",X"23",X"7E",X"FE",
		X"FC",X"28",X"05",X"FE",X"FE",X"C2",X"FE",X"0B",X"21",X"44",X"4C",X"CB",X"C6",X"3E",X"02",X"C3",
		X"98",X"07",X"2A",X"45",X"4C",X"23",X"23",X"E7",X"CD",X"6E",X"09",X"28",X"1F",X"FE",X"F6",X"D2",
		X"88",X"1C",X"7D",X"FE",X"40",X"D2",X"88",X"1C",X"00",X"00",X"00",X"00",X"7C",X"FE",X"40",X"CA",
		X"19",X"09",X"CD",X"A1",X"0A",X"CB",X"86",X"3E",X"03",X"C3",X"98",X"07",X"CD",X"D3",X"14",X"CB",
		X"CE",X"18",X"F4",X"21",X"44",X"4C",X"CB",X"4E",X"28",X"1F",X"FE",X"01",X"20",X"1B",X"3A",X"89",
		X"4C",X"3D",X"32",X"89",X"4C",X"00",X"2A",X"3A",X"4C",X"25",X"22",X"3A",X"4C",X"CD",X"DB",X"14",
		X"00",X"21",X"44",X"4C",X"CB",X"8E",X"CB",X"E6",X"C9",X"3D",X"32",X"43",X"4C",X"CD",X"2C",X"1B",
		X"EF",X"A9",X"08",X"C9",X"08",X"E4",X"08",X"EA",X"08",X"2A",X"3A",X"4C",X"24",X"3A",X"43",X"4C",
		X"FE",X"06",X"30",X"0D",X"FE",X"03",X"30",X"0D",X"3E",X"2C",X"32",X"FC",X"4F",X"22",X"3A",X"4C",
		X"C9",X"3E",X"30",X"18",X"F5",X"3E",X"34",X"18",X"F1",X"2A",X"3A",X"4C",X"2C",X"3A",X"43",X"4C",
		X"FE",X"06",X"30",X"08",X"FE",X"03",X"30",X"08",X"3E",X"22",X"18",X"DE",X"3E",X"26",X"18",X"DA",
		X"3E",X"2A",X"18",X"D6",X"2A",X"3A",X"4C",X"25",X"18",X"C3",X"2A",X"3A",X"4C",X"2D",X"3A",X"43",
		X"4C",X"FE",X"06",X"30",X"08",X"FE",X"03",X"30",X"08",X"3E",X"20",X"18",X"BD",X"3E",X"24",X"18",
		X"B9",X"3E",X"28",X"18",X"B5",X"2A",X"45",X"4C",X"23",X"C9",X"FE",X"43",X"C0",X"E1",X"3E",X"01",
		X"32",X"47",X"4C",X"3E",X"28",X"32",X"43",X"4C",X"C9",X"3E",X"03",X"32",X"47",X"4C",X"3E",X"28",
		X"32",X"43",X"4C",X"C9",X"21",X"52",X"9C",X"22",X"4C",X"4C",X"21",X"DD",X"04",X"C9",X"21",X"64",
		X"22",X"22",X"4C",X"4C",X"21",X"96",X"20",X"C3",X"1D",X"26",X"21",X"2E",X"8A",X"22",X"4C",X"4C",
		X"21",X"6E",X"88",X"C3",X"89",X"8A",X"21",X"64",X"34",X"22",X"4C",X"4C",X"21",X"A4",X"32",X"C3",
		X"CC",X"34",X"CD",X"5D",X"04",X"2A",X"4C",X"4C",X"46",X"23",X"7E",X"5F",X"23",X"56",X"23",X"7E",
		X"12",X"10",X"F6",X"C9",X"7E",X"FE",X"FE",X"28",X"03",X"FE",X"F0",X"C9",X"E1",X"C9",X"7E",X"FE",
		X"FF",X"28",X"03",X"FE",X"F0",X"C9",X"E1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3A",X"44",X"4C",X"CB",X"6F",X"C0",X"CB",X"57",X"C0",X"3A",X"47",X"4C",X"E6",X"0F",X"FE",
		X"01",X"28",X"26",X"CD",X"0E",X"07",X"23",X"E7",X"E7",X"7E",X"FE",X"0A",X"CD",X"52",X"0A",X"22",
		X"51",X"4C",X"CD",X"E4",X"0A",X"CB",X"D6",X"CB",X"9E",X"3E",X"0C",X"32",X"FC",X"4F",X"21",X"F3",
		X"09",X"CD",X"76",X"26",X"AF",X"32",X"02",X"4C",X"C9",X"CD",X"0E",X"07",X"23",X"DF",X"7E",X"FE",
		X"0A",X"CD",X"72",X"0A",X"00",X"22",X"51",X"4C",X"CD",X"E4",X"0A",X"CB",X"D6",X"CB",X"DE",X"3E",
		X"0E",X"18",X"D8",X"07",X"D2",X"00",X"0F",X"1F",X"10",X"21",X"B1",X"43",X"06",X"0A",X"36",X"14",
		X"E5",X"11",X"00",X"04",X"19",X"36",X"0F",X"E1",X"23",X"10",X"F3",X"C9",X"3A",X"50",X"4C",X"A7",
		X"28",X"05",X"3D",X"32",X"50",X"4C",X"C9",X"3E",X"10",X"32",X"50",X"4C",X"3A",X"44",X"4C",X"CB",
		X"57",X"C2",X"9A",X"0B",X"CB",X"6F",X"C2",X"F5",X"0A",X"3A",X"4E",X"4C",X"A7",X"28",X"05",X"3D",
		X"32",X"4E",X"4C",X"C9",X"3E",X"10",X"32",X"4E",X"4C",X"3A",X"4F",X"4C",X"FE",X"0A",X"20",X"01",
		X"AF",X"3C",X"32",X"4F",X"4C",X"CD",X"F9",X"09",X"21",X"BA",X"47",X"36",X"01",X"2B",X"3D",X"20",
		X"FA",X"C9",X"30",X"1A",X"E5",X"3A",X"3A",X"4C",X"FE",X"27",X"D2",X"A7",X"22",X"E1",X"C1",X"2B",
		X"00",X"22",X"51",X"4C",X"CD",X"B0",X"0A",X"CB",X"EE",X"CB",X"96",X"C3",X"C7",X"09",X"E1",X"C3",
		X"C9",X"09",X"30",X"1A",X"E5",X"3A",X"3A",X"4C",X"FE",X"E6",X"DA",X"B3",X"22",X"00",X"E1",X"C1",
		X"2B",X"22",X"51",X"4C",X"CD",X"B0",X"0A",X"CB",X"EE",X"CB",X"96",X"C3",X"ED",X"09",X"E1",X"C3",
		X"EF",X"09",X"2B",X"DF",X"7E",X"FE",X"0A",X"30",X"04",X"E1",X"C3",X"96",X"0B",X"21",X"44",X"4C",
		X"C9",X"2B",X"E7",X"7E",X"FE",X"0A",X"30",X"04",X"E1",X"C3",X"8E",X"0B",X"21",X"44",X"4C",X"C9",
		X"3E",X"28",X"32",X"53",X"4C",X"23",X"7E",X"36",X"F0",X"2B",X"CD",X"F2",X"0C",X"68",X"61",X"22",
		X"38",X"4C",X"CD",X"D1",X"0A",X"32",X"FA",X"4F",X"3E",X"08",X"32",X"FB",X"4F",X"21",X"44",X"4C",
		X"C9",X"32",X"54",X"4C",X"06",X"38",X"A7",X"28",X"09",X"F5",X"3E",X"04",X"80",X"47",X"F1",X"3D",
		X"20",X"F7",X"78",X"C9",X"3A",X"4F",X"4C",X"06",X"08",X"F5",X"3E",X"08",X"80",X"47",X"F1",X"3D",
		X"20",X"F7",X"78",X"18",X"BD",X"3A",X"44",X"4C",X"CB",X"5F",X"20",X"66",X"3A",X"53",X"4C",X"3D",
		X"32",X"53",X"4C",X"2A",X"38",X"4C",X"FE",X"28",X"30",X"1E",X"FE",X"20",X"30",X"1D",X"FE",X"10",
		X"30",X"1D",X"FE",X"08",X"30",X"1C",X"A7",X"20",X"0A",X"3A",X"44",X"4C",X"00",X"00",X"CB",X"AF",
		X"C3",X"36",X"0B",X"25",X"22",X"38",X"4C",X"C9",X"24",X"18",X"F9",X"24",X"2C",X"18",X"F5",X"2C",
		X"18",X"F2",X"2C",X"25",X"18",X"EE",X"32",X"44",X"4C",X"E5",X"CD",X"89",X"0B",X"23",X"23",X"CD",
		X"E0",X"0C",X"28",X"11",X"2B",X"CD",X"FC",X"0C",X"77",X"E1",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E1",X"25",X"22",X"38",X"4C",X"21",X"44",X"4C",X"CB",X"F6",X"CB",
		X"D6",X"C9",X"3A",X"53",X"4C",X"3D",X"32",X"53",X"4C",X"2A",X"38",X"4C",X"FE",X"28",X"30",X"B8",
		X"FE",X"20",X"30",X"0A",X"FE",X"10",X"30",X"0A",X"FE",X"08",X"30",X"09",X"18",X"98",X"24",X"2D",
		X"18",X"A2",X"2D",X"18",X"9F",X"2D",X"25",X"18",X"9B",X"45",X"4C",X"C3",X"13",X"07",X"3E",X"03",
		X"32",X"47",X"4C",X"C3",X"67",X"0C",X"3E",X"01",X"18",X"F6",X"CB",X"77",X"CA",X"DB",X"0B",X"CD",
		X"73",X"11",X"3A",X"55",X"4C",X"A7",X"28",X"09",X"25",X"3D",X"32",X"55",X"4C",X"22",X"38",X"4C",
		X"C9",X"CD",X"89",X"0B",X"23",X"23",X"7E",X"CD",X"81",X"0C",X"00",X"3E",X"08",X"32",X"55",X"4C",
		X"C9",X"2B",X"CD",X"54",X"1A",X"77",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3A",X"44",X"4C",X"E6",X"9B",X"32",X"44",X"4C",X"C9",X"CB",X"5F",X"28",X"52",X"3A",
		X"53",X"4C",X"3D",X"32",X"53",X"4C",X"FE",X"08",X"D2",X"26",X"0C",X"2A",X"38",X"4C",X"CD",X"89",
		X"0B",X"23",X"23",X"7E",X"FE",X"F6",X"30",X"7A",X"DF",X"7E",X"FE",X"F6",X"18",X"0B",X"FE",X"0A",
		X"D2",X"A1",X"07",X"C3",X"38",X"08",X"FF",X"FF",X"FF",X"AF",X"32",X"53",X"4C",X"32",X"55",X"4C",
		X"21",X"44",X"4C",X"CB",X"F6",X"C9",X"2B",X"3A",X"54",X"4C",X"77",X"21",X"00",X"00",X"22",X"FA",
		X"4F",X"22",X"38",X"4C",X"18",X"AC",X"CD",X"73",X"11",X"2A",X"38",X"4C",X"2C",X"C3",X"B0",X"0C",
		X"FE",X"3A",X"53",X"4C",X"3D",X"32",X"53",X"4C",X"FE",X"08",X"30",X"20",X"2A",X"38",X"4C",X"CD",
		X"89",X"0B",X"23",X"23",X"7E",X"FE",X"F6",X"30",X"29",X"E7",X"7E",X"FE",X"F6",X"30",X"BA",X"CD",
		X"78",X"0C",X"CB",X"97",X"00",X"00",X"CB",X"EF",X"32",X"44",X"4C",X"C9",X"CD",X"73",X"11",X"2A",
		X"38",X"4C",X"2D",X"C3",X"8B",X"0C",X"C9",X"3A",X"44",X"4C",X"CB",X"87",X"32",X"44",X"4C",X"C3",
		X"A1",X"07",X"FE",X"FE",X"38",X"A0",X"18",X"80",X"3E",X"10",X"32",X"53",X"4C",X"3A",X"44",X"4C",
		X"C9",X"FE",X"15",X"D8",X"FE",X"FE",X"D0",X"00",X"C3",X"8F",X"0D",X"7D",X"FE",X"17",X"D8",X"22",
		X"38",X"4C",X"CD",X"D5",X"0C",X"FE",X"08",X"28",X"03",X"00",X"A7",X"C0",X"CD",X"89",X"0B",X"23",
		X"E7",X"7E",X"FE",X"0A",X"D0",X"DF",X"23",X"7E",X"FE",X"F6",X"DA",X"09",X"0C",X"C3",X"16",X"0C",
		X"7D",X"FE",X"EF",X"D0",X"22",X"38",X"4C",X"CD",X"D5",X"0C",X"FE",X"08",X"28",X"03",X"00",X"A7",
		X"C0",X"CD",X"89",X"0B",X"23",X"DF",X"7E",X"FE",X"0A",X"D0",X"E7",X"23",X"7E",X"FE",X"F6",X"DA",
		X"09",X"0C",X"C3",X"16",X"0C",X"3A",X"53",X"4C",X"E6",X"0F",X"C9",X"32",X"44",X"4C",X"3E",X"09",
		X"7E",X"FE",X"15",X"38",X"0B",X"FE",X"F0",X"28",X"07",X"FE",X"FE",X"30",X"03",X"AF",X"3D",X"C9",
		X"AF",X"C9",X"F5",X"E5",X"7E",X"23",X"77",X"E1",X"F1",X"C3",X"39",X"07",X"E5",X"3A",X"38",X"4C",
		X"FE",X"16",X"38",X"09",X"FE",X"EE",X"30",X"05",X"CD",X"54",X"1A",X"E1",X"C9",X"E1",X"C1",X"C3",
		X"49",X"0B",X"CD",X"53",X"0D",X"21",X"58",X"0D",X"3D",X"23",X"20",X"FC",X"7E",X"32",X"56",X"4C",
		X"32",X"57",X"4C",X"21",X"5F",X"0D",X"CD",X"53",X"0D",X"3D",X"23",X"20",X"FC",X"5E",X"23",X"16",
		X"0D",X"EB",X"11",X"30",X"4C",X"01",X"0A",X"00",X"ED",X"B0",X"CD",X"9F",X"0D",X"11",X"F2",X"4F",
		X"01",X"0A",X"00",X"ED",X"B0",X"CD",X"53",X"0D",X"21",X"96",X"0D",X"3D",X"23",X"20",X"FC",X"7E",
		X"C3",X"27",X"10",X"CD",X"87",X"0D",X"E6",X"07",X"C9",X"80",X"60",X"55",X"50",X"40",X"35",X"30",
		X"67",X"6F",X"77",X"77",X"7F",X"7F",X"7F",X"36",X"98",X"26",X"C0",X"C6",X"98",X"D6",X"C0",X"26",
		X"98",X"26",X"C0",X"86",X"C0",X"C6",X"D8",X"2E",X"80",X"86",X"A8",X"66",X"F8",X"C6",X"C0",X"4E",
		X"F0",X"4E",X"98",X"8E",X"B8",X"96",X"98",X"3A",X"40",X"4C",X"E6",X"07",X"C0",X"3C",X"C9",X"FE",
		X"F0",X"C8",X"C1",X"C3",X"C1",X"0B",X"FF",X"09",X"08",X"08",X"07",X"06",X"06",X"06",X"FF",X"3A",
		X"40",X"4C",X"CB",X"47",X"28",X"04",X"21",X"AE",X"0D",X"C9",X"21",X"B6",X"0D",X"C9",X"12",X"08",
		X"16",X"0A",X"14",X"0D",X"10",X"05",X"18",X"08",X"1C",X"0A",X"18",X"0D",X"1C",X"05",X"3A",X"57",
		X"4C",X"3D",X"32",X"57",X"4C",X"C0",X"3A",X"56",X"4C",X"32",X"57",X"4C",X"DD",X"21",X"30",X"4C",
		X"CD",X"52",X"0E",X"DD",X"23",X"DD",X"23",X"DD",X"E5",X"E1",X"7D",X"FE",X"38",X"20",X"F1",X"C9",
		X"CD",X"0E",X"07",X"EB",X"D5",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"CD",X"13",X"07",X"D1",X"E5",
		X"D5",X"7D",X"E6",X"1F",X"6F",X"7B",X"E6",X"1F",X"BD",X"28",X"4D",X"38",X"41",X"DD",X"CB",X"31",
		X"86",X"DD",X"CB",X"31",X"CE",X"D1",X"E1",X"7C",X"BA",X"28",X"17",X"ED",X"52",X"FA",X"19",X"0E",
		X"DD",X"CB",X"31",X"D6",X"DD",X"CB",X"31",X"9E",X"C9",X"DD",X"CB",X"31",X"DE",X"DD",X"CB",X"31",
		X"96",X"C9",X"7D",X"93",X"F2",X"29",X"0E",X"3D",X"2F",X"FE",X"20",X"38",X"08",X"18",X"DC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"7E",X"31",X"E6",X"F3",X"DD",X"77",X"31",X"C9",X"DD",X"CB",
		X"31",X"C6",X"DD",X"CB",X"31",X"8E",X"18",X"BD",X"DD",X"7E",X"31",X"E6",X"FC",X"DD",X"77",X"31",
		X"18",X"B3",X"CD",X"63",X"23",X"CB",X"4F",X"C2",X"CC",X"11",X"CB",X"7F",X"C0",X"CB",X"47",X"C2",
		X"40",X"12",X"CB",X"57",X"C2",X"FA",X"11",X"CD",X"E9",X"36",X"CD",X"3C",X"15",X"FE",X"06",X"28",
		X"04",X"FE",X"0E",X"20",X"0A",X"7C",X"E6",X"0F",X"FE",X"08",X"28",X"49",X"A7",X"28",X"46",X"DD",
		X"7E",X"2A",X"CB",X"7F",X"20",X"12",X"E6",X"03",X"EF",X"91",X"0E",X"B3",X"0E",X"B9",X"0E",X"BF",
		X"0E",X"DD",X"7E",X"01",X"3C",X"DD",X"77",X"01",X"DD",X"7E",X"3E",X"3C",X"DD",X"77",X"3E",X"FE",
		X"04",X"C0",X"DD",X"7E",X"32",X"CB",X"57",X"20",X"06",X"CB",X"D7",X"CD",X"00",X"10",X"C9",X"CB",
		X"97",X"18",X"F8",X"DD",X"7E",X"00",X"C3",X"E1",X"0F",X"DD",X"7E",X"01",X"3D",X"18",X"D6",X"DD",
		X"7E",X"00",X"C3",X"E8",X"0F",X"CD",X"E0",X"0D",X"DD",X"7E",X"31",X"E6",X"0F",X"CC",X"DE",X"36",
		X"F6",X"FF",X"DD",X"77",X"3E",X"CD",X"2C",X"11",X"18",X"A5",X"DD",X"46",X"00",X"DD",X"4E",X"01",
		X"CD",X"13",X"07",X"22",X"6C",X"4C",X"DD",X"7E",X"2A",X"E6",X"01",X"20",X"04",X"CD",X"C6",X"10",
		X"C0",X"CD",X"DB",X"10",X"CB",X"6F",X"C2",X"32",X"10",X"CB",X"67",X"C2",X"32",X"10",X"E6",X"03",
		X"CA",X"A0",X"0F",X"2A",X"6C",X"4C",X"CD",X"D6",X"0F",X"28",X"43",X"2A",X"6C",X"4C",X"CD",X"FE",
		X"10",X"CA",X"F2",X"0F",X"CD",X"EB",X"0F",X"EF",X"20",X"0F",X"33",X"0F",X"3C",X"0F",X"45",X"0F",
		X"DD",X"7E",X"31",X"CB",X"FF",X"CB",X"B7",X"DD",X"77",X"31",X"78",X"3C",X"3C",X"E6",X"03",X"DD",
		X"77",X"2A",X"C9",X"DD",X"7E",X"31",X"CB",X"E7",X"CB",X"AF",X"18",X"EB",X"DD",X"7E",X"31",X"CB",
		X"F7",X"CB",X"BF",X"18",X"E2",X"DD",X"7E",X"31",X"CB",X"EF",X"CB",X"A7",X"18",X"D9",X"DD",X"7E",
		X"31",X"CB",X"47",X"28",X"05",X"AF",X"DD",X"77",X"2A",X"C9",X"3E",X"02",X"DD",X"77",X"2A",X"C9",
		X"DD",X"7E",X"31",X"E6",X"0C",X"28",X"35",X"CB",X"57",X"23",X"23",X"20",X"0B",X"DF",X"7E",X"FE",
		X"FE",X"38",X"56",X"AF",X"3D",X"C9",X"AF",X"C9",X"E7",X"E7",X"18",X"F2",X"CB",X"47",X"23",X"28",
		X"0E",X"7E",X"FE",X"FC",X"28",X"07",X"FE",X"FE",X"28",X"03",X"AF",X"3D",X"C9",X"AF",X"C9",X"23",
		X"7E",X"FE",X"FC",X"28",X"F8",X"FE",X"FE",X"28",X"F4",X"AF",X"3D",X"C9",X"C3",X"EF",X"10",X"28",
		X"2A",X"6C",X"4C",X"CD",X"60",X"0F",X"28",X"0C",X"CD",X"14",X"0F",X"DD",X"7E",X"29",X"CB",X"DF",
		X"DD",X"77",X"29",X"C9",X"DD",X"7E",X"31",X"CB",X"57",X"20",X"06",X"3E",X"01",X"DD",X"77",X"2A",
		X"C9",X"3E",X"03",X"18",X"F8",X"32",X"43",X"4C",X"C9",X"FE",X"F6",X"38",X"A6",X"AF",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"7E",X"29",X"CB",X"67",X"C0",X"DD",X"7E",X"31",X"18",
		X"9B",X"3C",X"DD",X"77",X"00",X"C3",X"98",X"0E",X"3D",X"18",X"F7",X"DD",X"7E",X"2A",X"47",X"E6",
		X"03",X"C9",X"DD",X"7E",X"29",X"CB",X"A7",X"DD",X"77",X"29",X"C3",X"8A",X"10",X"FF",X"FF",X"FF",
		X"DD",X"77",X"32",X"21",X"62",X"4C",X"11",X"F2",X"4F",X"01",X"04",X"00",X"ED",X"A0",X"23",X"13",
		X"EA",X"0C",X"10",X"C9",X"3A",X"6A",X"4C",X"A7",X"28",X"05",X"3D",X"CD",X"D6",X"12",X"C9",X"3E",
		X"01",X"32",X"6A",X"4C",X"C3",X"BE",X"0D",X"32",X"58",X"4C",X"21",X"F2",X"4F",X"11",X"62",X"4C",
		X"18",X"D7",X"DD",X"7E",X"29",X"CB",X"5F",X"2A",X"6C",X"4C",X"C2",X"50",X"10",X"DD",X"7E",X"31",
		X"CD",X"DC",X"0F",X"20",X"3C",X"DD",X"7E",X"31",X"E6",X"CF",X"DD",X"77",X"31",X"C3",X"4E",X"0F",
		X"ED",X"5F",X"CB",X"57",X"2A",X"6C",X"4C",X"23",X"20",X"1E",X"CD",X"8F",X"0F",X"C2",X"81",X"10",
		X"3E",X"02",X"DD",X"77",X"2A",X"DD",X"7E",X"29",X"00",X"00",X"CB",X"E7",X"DD",X"77",X"29",X"DD",
		X"7E",X"31",X"E6",X"CF",X"DD",X"77",X"31",X"C9",X"CD",X"81",X"0F",X"C2",X"81",X"10",X"AF",X"18",
		X"E1",X"2A",X"6C",X"4C",X"CD",X"A3",X"10",X"C2",X"BB",X"10",X"DD",X"7E",X"2A",X"CB",X"47",X"C0",
		X"00",X"DD",X"7E",X"31",X"CB",X"57",X"20",X"06",X"3E",X"01",X"DD",X"77",X"2A",X"C9",X"3E",X"03",
		X"18",X"F8",X"C9",X"DD",X"7E",X"2A",X"23",X"23",X"FE",X"01",X"20",X"0B",X"DF",X"7E",X"FE",X"F6",
		X"30",X"03",X"AF",X"3D",X"C9",X"AF",X"C9",X"E7",X"E7",X"18",X"F2",X"DD",X"7E",X"29",X"CB",X"DF",
		X"DD",X"77",X"29",X"C3",X"14",X"0F",X"DD",X"7E",X"31",X"E6",X"03",X"28",X"03",X"C3",X"60",X"0F",
		X"DD",X"7E",X"29",X"CB",X"EF",X"DD",X"77",X"29",X"C3",X"60",X"0F",X"DD",X"7E",X"29",X"CB",X"6F",
		X"20",X"04",X"DD",X"7E",X"31",X"C9",X"CB",X"AF",X"CB",X"E7",X"DD",X"77",X"29",X"18",X"F3",X"CD",
		X"26",X"11",X"7E",X"FE",X"FE",X"30",X"04",X"FE",X"F6",X"30",X"10",X"AF",X"3D",X"C9",X"DD",X"7E",
		X"31",X"E6",X"0C",X"28",X"1D",X"CD",X"91",X"10",X"C3",X"1C",X"11",X"ED",X"5F",X"CB",X"47",X"20",
		X"07",X"3E",X"01",X"DD",X"77",X"2A",X"AF",X"C9",X"3E",X"03",X"18",X"F7",X"2A",X"6C",X"4C",X"C3",
		X"A3",X"10",X"C1",X"C3",X"14",X"0F",X"2A",X"6C",X"4C",X"23",X"23",X"C9",X"CD",X"DA",X"0E",X"DD",
		X"7E",X"2A",X"CB",X"47",X"00",X"00",X"FE",X"01",X"28",X"11",X"3A",X"40",X"4C",X"CB",X"47",X"28",
		X"06",X"3E",X"10",X"C3",X"00",X"10",X"00",X"3E",X"18",X"18",X"F8",X"3A",X"40",X"4C",X"CB",X"47",
		X"28",X"04",X"3E",X"12",X"18",X"ED",X"3E",X"1A",X"18",X"E9",X"E6",X"0F",X"EF",X"65",X"11",X"6B",
		X"11",X"65",X"11",X"6F",X"11",X"3E",X"2C",X"32",X"FC",X"4F",X"C9",X"3E",X"22",X"18",X"F8",X"3E",
		X"20",X"18",X"F4",X"2A",X"38",X"4C",X"E5",X"DD",X"21",X"30",X"4C",X"DD",X"56",X"00",X"DD",X"5E",
		X"01",X"CD",X"92",X"11",X"DD",X"23",X"DD",X"23",X"DD",X"E5",X"D1",X"7B",X"FE",X"38",X"20",X"EB",
		X"E1",X"C9",X"DD",X"7E",X"29",X"CB",X"4F",X"C0",X"7C",X"93",X"F2",X"9F",X"11",X"ED",X"44",X"FE",
		X"09",X"D0",X"7D",X"92",X"28",X"0C",X"38",X"18",X"7D",X"92",X"F2",X"B1",X"11",X"ED",X"44",X"FE",
		X"09",X"D0",X"DD",X"7E",X"29",X"CB",X"57",X"C0",X"CD",X"9A",X"1E",X"CB",X"CF",X"C3",X"83",X"13",
		X"7D",X"92",X"F2",X"C7",X"11",X"ED",X"44",X"FE",X"11",X"D0",X"18",X"E6",X"DD",X"7E",X"3E",X"3C",
		X"DD",X"77",X"3E",X"CB",X"47",X"C0",X"DD",X"7E",X"3F",X"3D",X"DD",X"77",X"3F",X"06",X"E0",X"28",
		X"0D",X"F5",X"3E",X"04",X"80",X"47",X"F1",X"3D",X"20",X"F7",X"78",X"C3",X"00",X"10",X"DD",X"7E",
		X"29",X"CB",X"8F",X"CB",X"D7",X"DD",X"77",X"29",X"18",X"F0",X"DD",X"7E",X"01",X"FE",X"19",X"DA",
		X"15",X"12",X"3D",X"DD",X"77",X"01",X"CD",X"2F",X"11",X"DD",X"7E",X"32",X"3C",X"3C",X"3C",X"DD",
		X"77",X"32",X"C3",X"00",X"10",X"DD",X"7E",X"29",X"CB",X"C7",X"CB",X"97",X"DD",X"77",X"29",X"CD",
		X"70",X"12",X"CD",X"50",X"13",X"2E",X"FF",X"DD",X"75",X"46",X"CD",X"70",X"12",X"DD",X"70",X"32",
		X"C3",X"03",X"10",X"DD",X"7E",X"29",X"CB",X"FF",X"DD",X"77",X"29",X"21",X"4D",X"81",X"C9",X"4F",
		X"14",X"00",X"DD",X"7E",X"46",X"3D",X"DD",X"77",X"46",X"28",X"51",X"FE",X"55",X"30",X"07",X"ED",
		X"5F",X"E6",X"07",X"CD",X"91",X"12",X"DD",X"7E",X"00",X"FE",X"1E",X"28",X"0F",X"3D",X"DD",X"77",
		X"00",X"CB",X"4F",X"DD",X"7E",X"01",X"20",X"05",X"3C",X"DD",X"77",X"01",X"C9",X"3D",X"18",X"F9",
		X"3A",X"40",X"4C",X"21",X"87",X"12",X"3D",X"23",X"23",X"20",X"FB",X"00",X"00",X"7D",X"FE",X"91",
		X"38",X"03",X"21",X"8F",X"12",X"7E",X"23",X"46",X"C9",X"30",X"60",X"40",X"64",X"50",X"68",X"60",
		X"6C",X"3C",X"DD",X"E5",X"E1",X"11",X"C3",X"03",X"19",X"77",X"C9",X"A9",X"3A",X"58",X"4C",X"3D",
		X"CD",X"7C",X"13",X"FE",X"04",X"DD",X"7E",X"29",X"30",X"05",X"CB",X"F7",X"C3",X"E2",X"13",X"E6",
		X"FE",X"DD",X"77",X"29",X"3E",X"01",X"DD",X"77",X"2A",X"CD",X"2F",X"11",X"21",X"1E",X"18",X"DD",
		X"75",X"00",X"DD",X"74",X"01",X"C9",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"C9",X"CB",X"D6",X"CD",
		X"60",X"32",X"32",X"9E",X"4C",X"C9",X"32",X"6A",X"4C",X"3A",X"BE",X"4C",X"CB",X"57",X"C8",X"3A",
		X"9E",X"4C",X"C3",X"73",X"32",X"32",X"58",X"4C",X"C9",X"C3",X"63",X"94",X"11",X"7E",X"4C",X"1A",
		X"86",X"27",X"77",X"23",X"13",X"1A",X"8E",X"27",X"77",X"23",X"13",X"1A",X"8E",X"27",X"77",X"11",
		X"F7",X"43",X"AF",X"12",X"1E",X"FD",X"21",X"3E",X"4C",X"7E",X"4F",X"E6",X"F0",X"28",X"05",X"0F",
		X"0F",X"0F",X"0F",X"12",X"1B",X"79",X"E6",X"0F",X"28",X"01",X"12",X"06",X"02",X"4E",X"2B",X"1B",
		X"79",X"A7",X"7E",X"20",X"05",X"E6",X"F0",X"28",X"08",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"12",X"1B",X"79",X"A7",X"20",X"0A",X"7E",X"E6",X"F0",X"20",X"05",X"7E",X"E6",X"0F",X"28",X"04",
		X"7E",X"E6",X"0F",X"12",X"10",X"D7",X"21",X"7E",X"4C",X"AF",X"77",X"23",X"77",X"23",X"18",X"06",
		X"32",X"7E",X"4C",X"C3",X"E9",X"12",X"77",X"3A",X"81",X"4C",X"CB",X"47",X"C0",X"3A",X"3D",X"4C",
		X"FE",X"10",X"D8",X"3E",X"FA",X"CD",X"F2",X"9A",X"00",X"CD",X"CD",X"12",X"3A",X"3F",X"4C",X"3C",
		X"32",X"3F",X"4C",X"CD",X"48",X"1E",X"21",X"81",X"4C",X"CB",X"C6",X"C9",X"FE",X"02",X"C8",X"C3",
		X"E5",X"12",X"12",X"DD",X"77",X"29",X"3E",X"08",X"DD",X"77",X"3F",X"CD",X"1C",X"90",X"22",X"0B",
		X"4C",X"AF",X"32",X"02",X"4C",X"C9",X"05",X"A7",X"00",X"0F",X"04",X"05",X"98",X"00",X"0F",X"04",
		X"05",X"89",X"00",X"0F",X"04",X"05",X"77",X"00",X"0F",X"04",X"05",X"68",X"00",X"0F",X"04",X"05",
		X"59",X"00",X"0F",X"04",X"05",X"27",X"00",X"0F",X"04",X"05",X"38",X"00",X"0F",X"04",X"05",X"49",
		X"00",X"0F",X"04",X"05",X"57",X"00",X"0F",X"04",X"05",X"68",X"00",X"0F",X"04",X"05",X"79",X"00",
		X"0F",X"04",X"05",X"87",X"00",X"0F",X"04",X"05",X"98",X"00",X"0F",X"04",X"05",X"A9",X"00",X"0F",
		X"04",X"10",X"E6",X"FE",X"DD",X"77",X"29",X"21",X"16",X"18",X"C3",X"43",X"15",X"CD",X"CC",X"14",
		X"3D",X"32",X"84",X"4C",X"C0",X"3E",X"05",X"32",X"84",X"4C",X"3A",X"82",X"4C",X"3D",X"32",X"82",
		X"4C",X"C0",X"3E",X"F0",X"32",X"82",X"4C",X"3A",X"83",X"4C",X"3C",X"32",X"83",X"4C",X"CB",X"47",
		X"3E",X"18",X"28",X"02",X"3E",X"0D",X"21",X"9E",X"46",X"06",X"0A",X"77",X"DF",X"10",X"FC",X"C9",
		X"CD",X"F9",X"09",X"3A",X"58",X"4C",X"21",X"9F",X"46",X"06",X"0A",X"36",X"0F",X"DF",X"10",X"FB",
		X"2A",X"85",X"4C",X"22",X"87",X"4C",X"CD",X"48",X"1E",X"CD",X"0F",X"26",X"21",X"60",X"41",X"11",
		X"5C",X"14",X"C3",X"5C",X"94",X"29",X"21",X"00",X"11",X"22",X"85",X"4C",X"C3",X"24",X"09",X"FF",
		X"FF",X"FF",X"FF",X"04",X"BE",X"40",X"69",X"40",X"09",X"42",X"C1",X"41",X"0F",X"54",X"49",X"4D",
		X"45",X"FF",X"11",X"87",X"4C",X"21",X"73",X"14",X"1A",X"96",X"27",X"12",X"23",X"13",X"1A",X"9E",
		X"27",X"12",X"C9",X"01",X"00",X"3A",X"81",X"4C",X"CB",X"4F",X"C0",X"3A",X"AF",X"4C",X"3D",X"32",
		X"AF",X"4C",X"C0",X"3D",X"32",X"AF",X"4C",X"3A",X"B0",X"4C",X"3D",X"32",X"B0",X"4C",X"C0",X"3E",
		X"04",X"32",X"B0",X"4C",X"CD",X"62",X"14",X"11",X"87",X"4C",X"21",X"60",X"40",X"CD",X"B2",X"14",
		X"CD",X"4D",X"32",X"AF",X"21",X"87",X"4C",X"BE",X"C0",X"23",X"BE",X"C0",X"21",X"81",X"4C",X"C3",
		X"69",X"32",X"06",X"02",X"1A",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"77",X"D5",X"E7",X"D1",X"1A",
		X"E6",X"0F",X"77",X"13",X"D5",X"DF",X"DF",X"DF",X"D1",X"10",X"E9",X"C9",X"CD",X"75",X"14",X"3A",
		X"84",X"4C",X"C9",X"AF",X"32",X"89",X"4C",X"CD",X"07",X"15",X"C9",X"CD",X"16",X"15",X"23",X"23",
		X"7E",X"FE",X"F1",X"30",X"02",X"E1",X"C9",X"3A",X"89",X"4C",X"FE",X"C0",X"38",X"0D",X"21",X"EC",
		X"9A",X"CD",X"8E",X"13",X"21",X"44",X"4C",X"CB",X"8E",X"E1",X"C9",X"21",X"00",X"00",X"C3",X"D6",
		X"24",X"01",X"FF",X"00",X"0F",X"01",X"10",X"21",X"01",X"15",X"11",X"8A",X"4C",X"01",X"06",X"00",
		X"ED",X"B0",X"21",X"44",X"4C",X"C9",X"3A",X"90",X"4C",X"3D",X"32",X"90",X"4C",X"CB",X"57",X"C2",
		X"11",X"07",X"3A",X"8B",X"4C",X"0F",X"0F",X"0F",X"0F",X"3D",X"0F",X"0F",X"0F",X"0F",X"32",X"8B",
		X"4C",X"E5",X"21",X"8A",X"4C",X"CD",X"8E",X"13",X"E1",X"C3",X"11",X"07",X"CD",X"C6",X"12",X"7D",
		X"E6",X"0F",X"C9",X"CD",X"BF",X"12",X"3A",X"81",X"4C",X"CB",X"57",X"C0",X"CB",X"D7",X"E6",X"C7",
		X"CB",X"DF",X"32",X"81",X"4C",X"CD",X"33",X"12",X"22",X"07",X"4C",X"AF",X"32",X"01",X"4C",X"DD",
		X"22",X"91",X"4C",X"3C",X"32",X"95",X"4C",X"2A",X"91",X"4C",X"11",X"FE",X"F0",X"73",X"C3",X"04",
		X"18",X"3A",X"81",X"4C",X"CB",X"5F",X"C8",X"3A",X"95",X"4C",X"A7",X"28",X"07",X"3D",X"32",X"95",
		X"4C",X"C2",X"C7",X"16",X"CD",X"6F",X"1C",X"CB",X"77",X"C2",X"A7",X"19",X"CB",X"67",X"C2",X"01",
		X"19",X"CB",X"6F",X"C2",X"27",X"18",X"CD",X"4A",X"19",X"CA",X"70",X"19",X"00",X"3A",X"3B",X"4C",
		X"47",X"0E",X"F8",X"FE",X"C0",X"30",X"03",X"C6",X"30",X"4F",X"CD",X"DE",X"15",X"7C",X"B8",X"38",
		X"06",X"B9",X"30",X"6F",X"C3",X"34",X"16",X"CD",X"D9",X"15",X"28",X"62",X"3E",X"03",X"06",X"00",
		X"CD",X"E6",X"15",X"28",X"04",X"78",X"32",X"94",X"4C",X"CD",X"D9",X"15",X"E6",X"01",X"32",X"93",
		X"4C",X"3E",X"0D",X"32",X"95",X"4C",X"00",X"00",X"C9",X"ED",X"5F",X"CB",X"67",X"C9",X"2A",X"91",
		X"4C",X"5E",X"23",X"56",X"EB",X"C9",X"32",X"94",X"4C",X"A7",X"20",X"03",X"11",X"08",X"08",X"3D",
		X"20",X"03",X"11",X"08",X"F8",X"3D",X"20",X"03",X"11",X"F8",X"F8",X"3D",X"20",X"03",X"11",X"F8",
		X"08",X"7D",X"83",X"6F",X"7C",X"82",X"67",X"7D",X"FE",X"0E",X"38",X"0F",X"FE",X"F7",X"30",X"0B",
		X"7C",X"FE",X"18",X"38",X"06",X"FE",X"F9",X"30",X"02",X"AF",X"C9",X"AF",X"3D",X"C9",X"06",X"03",
		X"AF",X"18",X"9D",X"CD",X"D9",X"15",X"28",X"06",X"3E",X"01",X"06",X"02",X"18",X"92",X"3E",X"02",
		X"06",X"01",X"18",X"8C",X"2A",X"3A",X"4C",X"7D",X"FE",X"5E",X"38",X"3E",X"FE",X"AE",X"30",X"3E",
		X"F5",X"D6",X"40",X"47",X"F1",X"C6",X"40",X"4F",X"7C",X"FE",X"C0",X"30",X"38",X"F5",X"C6",X"40",
		X"57",X"F1",X"C6",X"20",X"5F",X"D5",X"CD",X"DE",X"15",X"D1",X"7D",X"B8",X"38",X"2C",X"B9",X"30",
		X"29",X"7C",X"BB",X"38",X"25",X"BA",X"30",X"22",X"3A",X"81",X"4C",X"CB",X"EF",X"32",X"81",X"4C",
		X"CD",X"D9",X"15",X"E6",X"07",X"3C",X"32",X"96",X"4C",X"C9",X"06",X"16",X"18",X"C7",X"0E",X"EE",
		X"D6",X"40",X"47",X"18",X"C3",X"16",X"F8",X"7C",X"18",X"C8",X"ED",X"5B",X"3A",X"4C",X"7D",X"93",
		X"38",X"13",X"CD",X"D9",X"15",X"28",X"07",X"3E",X"03",X"06",X"02",X"C3",X"C0",X"15",X"3E",X"02",
		X"06",X"03",X"C3",X"C0",X"15",X"CD",X"D9",X"15",X"20",X"07",X"3E",X"01",X"06",X"00",X"C3",X"C0",
		X"15",X"AF",X"06",X"01",X"C3",X"C0",X"15",X"CD",X"6E",X"23",X"3D",X"32",X"98",X"4C",X"C0",X"3E",
		X"A0",X"32",X"98",X"4C",X"C3",X"71",X"15",X"00",X"CD",X"08",X"1C",X"3A",X"81",X"4C",X"CB",X"67",
		X"C2",X"26",X"19",X"3A",X"94",X"4C",X"EF",X"DF",X"16",X"CE",X"17",X"E0",X"17",X"F2",X"17",X"3A",
		X"93",X"4C",X"A7",X"28",X"3C",X"21",X"07",X"17",X"CD",X"FF",X"16",X"D5",X"CD",X"DE",X"15",X"D1",
		X"7D",X"83",X"6F",X"7C",X"82",X"67",X"EB",X"2A",X"91",X"4C",X"73",X"23",X"C3",X"0C",X"18",X"3A",
		X"95",X"4C",X"87",X"85",X"6F",X"5E",X"23",X"56",X"C9",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"21",X"24",X"17",X"18",X"C2",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"FF",
		X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",
		X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"3A",X"93",
		X"4C",X"A7",X"28",X"06",X"21",X"54",X"17",X"C3",X"E8",X"16",X"21",X"3C",X"17",X"C3",X"E8",X"16",
		X"3A",X"93",X"4C",X"A7",X"28",X"06",X"21",X"84",X"17",X"C3",X"E8",X"16",X"21",X"6C",X"17",X"C3",
		X"E8",X"16",X"3A",X"93",X"4C",X"A7",X"28",X"06",X"21",X"B4",X"17",X"C3",X"E8",X"16",X"21",X"9C",
		X"17",X"C3",X"E8",X"16",X"23",X"72",X"3E",X"70",X"32",X"97",X"4C",X"C9",X"72",X"3A",X"95",X"4C",
		X"FE",X"07",X"3E",X"70",X"30",X"02",X"3E",X"74",X"DD",X"2A",X"91",X"4C",X"DD",X"77",X"32",X"3A",
		X"81",X"4C",X"CB",X"77",X"C3",X"EE",X"19",X"3A",X"96",X"4C",X"3D",X"32",X"96",X"4C",X"20",X"30",
		X"CD",X"DE",X"15",X"ED",X"5B",X"3A",X"4C",X"7D",X"BB",X"38",X"1B",X"CD",X"D9",X"15",X"3E",X"03",
		X"28",X"02",X"3E",X"02",X"32",X"94",X"4C",X"3E",X"0D",X"32",X"95",X"4C",X"CD",X"D9",X"15",X"CD",
		X"F5",X"18",X"32",X"96",X"4C",X"C9",X"CD",X"D9",X"15",X"3E",X"01",X"28",X"E7",X"AF",X"18",X"E4",
		X"CD",X"DE",X"15",X"7D",X"FE",X"0E",X"38",X"67",X"FE",X"FE",X"30",X"63",X"2A",X"3A",X"4C",X"7D",
		X"FE",X"3E",X"38",X"65",X"FE",X"C6",X"30",X"65",X"F5",X"D6",X"28",X"47",X"F1",X"C6",X"28",X"4F",
		X"7C",X"FE",X"C0",X"30",X"5F",X"F5",X"C6",X"40",X"57",X"F1",X"5F",X"D5",X"CD",X"DE",X"15",X"D1",
		X"7D",X"B8",X"38",X"54",X"B9",X"30",X"51",X"7C",X"BB",X"38",X"4D",X"BA",X"30",X"4A",X"3A",X"81",
		X"4C",X"CB",X"AF",X"CB",X"E7",X"32",X"81",X"4C",X"ED",X"5B",X"3A",X"4C",X"7D",X"BB",X"28",X"3E",
		X"38",X"40",X"3E",X"02",X"32",X"94",X"4C",X"3E",X"09",X"32",X"95",X"4C",X"CD",X"D9",X"15",X"E6",
		X"07",X"3C",X"32",X"96",X"4C",X"3A",X"98",X"4C",X"D6",X"65",X"00",X"32",X"98",X"4C",X"C9",X"3A",
		X"94",X"4C",X"3C",X"3C",X"E6",X"03",X"C3",X"44",X"18",X"06",X"16",X"18",X"A0",X"0E",X"EE",X"D6",
		X"28",X"47",X"18",X"9C",X"16",X"F8",X"18",X"A2",X"3E",X"0D",X"32",X"95",X"4C",X"C9",X"3E",X"01",
		X"18",X"C2",X"AF",X"18",X"BF",X"F5",X"0F",X"E6",X"01",X"32",X"93",X"4C",X"F1",X"E6",X"07",X"3C",
		X"C9",X"3A",X"96",X"4C",X"3D",X"32",X"96",X"4C",X"28",X"13",X"CD",X"4A",X"19",X"CA",X"70",X"19",
		X"3E",X"09",X"32",X"95",X"4C",X"CD",X"DE",X"15",X"7C",X"FE",X"21",X"30",X"A8",X"3A",X"81",X"4C",
		X"CB",X"A7",X"32",X"81",X"4C",X"C9",X"3A",X"94",X"4C",X"EF",X"30",X"19",X"38",X"19",X"3F",X"19",
		X"CD",X"DE",X"15",X"25",X"2C",X"C3",X"44",X"19",X"CD",X"DE",X"15",X"25",X"C3",X"44",X"19",X"CD",
		X"DE",X"15",X"25",X"2D",X"CD",X"C5",X"18",X"C3",X"F6",X"16",X"CD",X"23",X"1D",X"ED",X"5B",X"3A",
		X"4C",X"7C",X"92",X"38",X"17",X"FE",X"09",X"30",X"13",X"7B",X"F5",X"C6",X"08",X"47",X"F1",X"D6",
		X"08",X"4F",X"7D",X"B9",X"38",X"05",X"B8",X"30",X"02",X"AF",X"C9",X"AF",X"3D",X"C9",X"00",X"00",
		X"CD",X"D9",X"15",X"3E",X"03",X"28",X"01",X"AF",X"32",X"94",X"4C",X"CD",X"D9",X"15",X"0F",X"E6",
		X"01",X"32",X"93",X"4C",X"3A",X"81",X"4C",X"CB",X"F7",X"E6",X"CF",X"CD",X"36",X"1A",X"21",X"2D",
		X"4C",X"CB",X"86",X"21",X"69",X"85",X"22",X"03",X"4C",X"21",X"0A",X"86",X"22",X"07",X"4C",X"AF",
		X"32",X"00",X"4C",X"32",X"01",X"4C",X"C9",X"3A",X"96",X"4C",X"3D",X"32",X"96",X"4C",X"3E",X"0D",
		X"32",X"95",X"4C",X"28",X"1B",X"CD",X"19",X"1A",X"28",X"0F",X"21",X"2D",X"4C",X"CD",X"3C",X"1A",
		X"3A",X"81",X"4C",X"CB",X"B7",X"CD",X"E4",X"9A",X"C9",X"CD",X"FC",X"19",X"18",X"EC",X"00",X"00",
		X"CD",X"D9",X"15",X"3E",X"03",X"20",X"01",X"AF",X"32",X"94",X"4C",X"CD",X"D9",X"15",X"E6",X"07",
		X"3C",X"32",X"96",X"4C",X"CD",X"D9",X"15",X"0F",X"E6",X"01",X"C3",X"2A",X"1A",X"B9",X"C8",X"CD",
		X"DE",X"15",X"7C",X"D6",X"10",X"57",X"5D",X"ED",X"53",X"3A",X"4C",X"C9",X"3A",X"3B",X"4C",X"FE",
		X"E8",X"D0",X"3A",X"3A",X"4C",X"FE",X"1E",X"D8",X"FE",X"E6",X"D0",X"C1",X"C9",X"21",X"4D",X"81",
		X"22",X"03",X"4C",X"21",X"92",X"83",X"C3",X"9C",X"19",X"CD",X"D9",X"15",X"47",X"3A",X"2C",X"4C",
		X"80",X"FE",X"10",X"30",X"03",X"AF",X"3D",X"C9",X"AF",X"C9",X"32",X"93",X"4C",X"CD",X"FC",X"19",
		X"C3",X"BA",X"19",X"00",X"00",X"00",X"32",X"81",X"4C",X"C3",X"EF",X"19",X"CB",X"C6",X"3E",X"08",
		X"32",X"43",X"4C",X"CD",X"0D",X"1A",X"CD",X"0E",X"07",X"CD",X"39",X"07",X"68",X"61",X"CD",X"EA",
		X"1A",X"C3",X"E4",X"1A",X"3A",X"54",X"4C",X"47",X"7E",X"FE",X"0A",X"78",X"30",X"68",X"3A",X"44",
		X"4C",X"CB",X"5F",X"06",X"00",X"20",X"4B",X"E7",X"7E",X"04",X"FE",X"0A",X"38",X"F9",X"CD",X"CC",
		X"1A",X"E5",X"DF",X"7E",X"E1",X"77",X"DF",X"10",X"F8",X"3A",X"9B",X"4C",X"C9",X"3A",X"54",X"4C",
		X"32",X"9B",X"4C",X"E5",X"23",X"7E",X"E1",X"FE",X"F0",X"20",X"13",X"7E",X"36",X"F0",X"00",X"E5",
		X"CD",X"DE",X"1A",X"CB",X"F6",X"CB",X"D6",X"E1",X"3E",X"08",X"32",X"55",X"4C",X"C9",X"E5",X"21",
		X"00",X"00",X"22",X"FA",X"4F",X"22",X"38",X"4C",X"3A",X"44",X"4C",X"E6",X"9B",X"32",X"44",X"4C",
		X"E1",X"C9",X"DF",X"7E",X"04",X"FE",X"0A",X"38",X"F9",X"CD",X"D2",X"1A",X"E5",X"E7",X"7E",X"E1",
		X"77",X"E7",X"10",X"F8",X"18",X"B3",X"F5",X"CD",X"9E",X"1A",X"F1",X"C9",X"DF",X"CD",X"D8",X"1A",
		X"E7",X"C9",X"E7",X"CD",X"D8",X"1A",X"DF",X"C9",X"C5",X"CD",X"7D",X"1A",X"C1",X"C9",X"CD",X"39",
		X"07",X"C3",X"BD",X"0A",X"21",X"44",X"4C",X"CB",X"CE",X"C9",X"7D",X"FE",X"17",X"38",X"08",X"FE",
		X"EE",X"30",X"08",X"22",X"3A",X"4C",X"C9",X"2E",X"1E",X"18",X"F8",X"2E",X"E6",X"18",X"F4",X"CD",
		X"79",X"1B",X"FE",X"0F",X"CA",X"A1",X"09",X"CB",X"47",X"CA",X"A1",X"09",X"CB",X"4F",X"3A",X"44",
		X"4C",X"CB",X"FF",X"CB",X"9F",X"20",X"02",X"CB",X"DF",X"32",X"44",X"4C",X"3E",X"20",X"32",X"43",
		X"4C",X"21",X"A6",X"1B",X"22",X"0B",X"4C",X"AF",X"32",X"02",X"4C",X"C9",X"3A",X"44",X"4C",X"CB",
		X"7F",X"20",X"04",X"3A",X"47",X"4C",X"C9",X"E1",X"47",X"3A",X"43",X"4C",X"A7",X"78",X"20",X"05",
		X"CB",X"BF",X"32",X"44",X"4C",X"CB",X"5F",X"2A",X"3A",X"4C",X"7D",X"28",X"15",X"FE",X"EE",X"3A",
		X"44",X"4C",X"30",X"09",X"32",X"44",X"4C",X"CD",X"D8",X"1B",X"C3",X"BA",X"08",X"CB",X"9F",X"C3",
		X"FD",X"1B",X"FE",X"17",X"3A",X"44",X"4C",X"38",X"08",X"CD",X"F1",X"1B",X"3E",X"0C",X"C3",X"BA",
		X"08",X"CB",X"DF",X"32",X"44",X"4C",X"C3",X"F7",X"1B",X"3A",X"2E",X"4C",X"E6",X"0F",X"C9",X"CD",
		X"0E",X"07",X"7C",X"FE",X"43",X"20",X"10",X"7D",X"FE",X"C8",X"CA",X"D5",X"06",X"FE",X"CD",X"CA",
		X"D5",X"06",X"FE",X"BD",X"CA",X"85",X"1C",X"23",X"23",X"7E",X"FE",X"F0",X"C2",X"D5",X"06",X"E7",
		X"7E",X"FE",X"F0",X"C3",X"A2",X"1C",X"04",X"69",X"10",X"0F",X"02",X"04",X"0F",X"00",X"0F",X"02",
		X"02",X"CC",X"00",X"0F",X"0A",X"07",X"6B",X"00",X"0F",X"02",X"04",X"A7",X"00",X"0F",X"02",X"07",
		X"D2",X"00",X"0F",X"02",X"10",X"3A",X"43",X"4C",X"FE",X"1B",X"30",X"09",X"FE",X"05",X"30",X"03",
		X"2C",X"25",X"C9",X"2C",X"C9",X"2C",X"24",X"C9",X"CD",X"C5",X"1B",X"3E",X"0E",X"C9",X"3A",X"43",
		X"4C",X"FE",X"1B",X"30",X"09",X"FE",X"05",X"30",X"03",X"2D",X"25",X"C9",X"2D",X"C9",X"2D",X"24",
		X"C9",X"32",X"44",X"4C",X"C3",X"DE",X"1B",X"CD",X"C5",X"1B",X"C3",X"6C",X"1B",X"32",X"44",X"4C",
		X"CD",X"DE",X"1B",X"3E",X"0E",X"C3",X"BA",X"08",X"CD",X"6A",X"1C",X"DD",X"7E",X"29",X"CB",X"57",
		X"C8",X"E1",X"3A",X"81",X"4C",X"CB",X"7F",X"20",X"19",X"DD",X"7E",X"01",X"FE",X"19",X"38",X"08",
		X"3D",X"DD",X"77",X"01",X"C3",X"AB",X"1C",X"B1",X"3E",X"00",X"32",X"9D",X"4C",X"CD",X"D4",X"1E",
		X"CB",X"FE",X"3A",X"9D",X"4C",X"3D",X"32",X"9D",X"4C",X"28",X"10",X"CB",X"57",X"3E",X"7C",X"20",
		X"02",X"3E",X"78",X"CD",X"1A",X"1D",X"AF",X"32",X"98",X"4C",X"C9",X"AF",X"32",X"95",X"4C",X"3E",
		X"06",X"CD",X"91",X"12",X"DD",X"7E",X"29",X"CB",X"97",X"DD",X"77",X"29",X"3A",X"81",X"4C",X"E6",
		X"0F",X"32",X"81",X"4C",X"21",X"EE",X"E8",X"C3",X"9A",X"1C",X"DD",X"2A",X"91",X"4C",X"C9",X"CD",
		X"6A",X"1C",X"DD",X"7E",X"29",X"CB",X"4F",X"3A",X"81",X"4C",X"C8",X"E1",X"C9",X"CB",X"4F",X"3E",
		X"03",X"C0",X"3E",X"01",X"C9",X"3E",X"23",X"C9",X"CD",X"28",X"26",X"CC",X"BF",X"22",X"C3",X"62",
		X"08",X"CD",X"28",X"26",X"CC",X"BF",X"22",X"C3",X"19",X"08",X"CD",X"BF",X"12",X"3E",X"06",X"C3",
		X"00",X"10",X"C2",X"D5",X"06",X"3A",X"47",X"4C",X"C3",X"7D",X"1C",X"32",X"95",X"4C",X"CB",X"57",
		X"3E",X"73",X"20",X"02",X"3E",X"77",X"C3",X"00",X"10",X"CD",X"79",X"23",X"3A",X"81",X"4C",X"CB",
		X"4F",X"C2",X"59",X"1D",X"3A",X"44",X"4C",X"CB",X"67",X"C2",X"F1",X"1D",X"CD",X"20",X"23",X"C3",
		X"C6",X"06",X"AF",X"CD",X"60",X"32",X"CD",X"D6",X"24",X"C3",X"05",X"1F",X"FF",X"FF",X"E1",X"21",
		X"2D",X"4C",X"CB",X"86",X"21",X"4A",X"87",X"22",X"03",X"4C",X"21",X"D7",X"87",X"CD",X"E8",X"34",
		X"06",X"08",X"3E",X"08",X"CD",X"01",X"1D",X"3E",X"0E",X"CD",X"01",X"1D",X"10",X"F4",X"C3",X"35",
		X"1F",X"C5",X"21",X"40",X"44",X"01",X"04",X"80",X"CF",X"CD",X"0E",X"1D",X"C1",X"C9",X"3E",X"1A",
		X"32",X"2C",X"4C",X"3A",X"2C",X"4C",X"A7",X"20",X"FA",X"C9",X"CD",X"00",X"10",X"3E",X"90",X"32",
		X"95",X"4C",X"C9",X"DD",X"2A",X"91",X"4C",X"DD",X"7E",X"29",X"CB",X"4F",X"20",X"05",X"CB",X"57",
		X"CA",X"DE",X"15",X"E1",X"AF",X"3D",X"C9",X"FB",X"CD",X"84",X"26",X"3A",X"81",X"4C",X"32",X"A4",
		X"4C",X"21",X"43",X"4C",X"01",X"01",X"60",X"AF",X"CF",X"3A",X"A4",X"4C",X"E6",X"01",X"32",X"81",
		X"4C",X"3E",X"80",X"CD",X"10",X"1D",X"C3",X"58",X"04",X"CD",X"EB",X"1D",X"21",X"AD",X"42",X"11",
		X"F7",X"1D",X"CD",X"08",X"1E",X"21",X"30",X"4C",X"01",X"01",X"08",X"AF",X"CF",X"3E",X"20",X"CD",
		X"10",X"1D",X"06",X"10",X"CD",X"C3",X"80",X"32",X"7E",X"4C",X"3E",X"0E",X"32",X"FD",X"4F",X"3E",
		X"80",X"32",X"FC",X"4F",X"3E",X"05",X"CD",X"10",X"1D",X"3E",X"84",X"32",X"FC",X"4F",X"3E",X"05",
		X"CD",X"10",X"1D",X"10",X"EA",X"3A",X"3F",X"4C",X"3D",X"32",X"3F",X"4C",X"CA",X"C2",X"26",X"CD",
		X"48",X"1E",X"21",X"5F",X"0D",X"CD",X"53",X"0D",X"3D",X"23",X"20",X"FC",X"5E",X"CD",X"03",X"1E",
		X"11",X"30",X"4C",X"01",X"0A",X"00",X"ED",X"B0",X"21",X"45",X"4C",X"01",X"01",X"07",X"AF",X"CF",
		X"32",X"43",X"4C",X"3A",X"44",X"4C",X"E6",X"44",X"32",X"44",X"4C",X"CD",X"E0",X"06",X"3A",X"7E",
		X"4C",X"3A",X"81",X"4C",X"E6",X"BD",X"32",X"81",X"4C",X"2A",X"85",X"4C",X"22",X"87",X"4C",X"21",
		X"60",X"40",X"11",X"87",X"4C",X"CD",X"B2",X"14",X"C3",X"FD",X"1E",X"21",X"2D",X"4C",X"CB",X"86",
		X"C9",X"CD",X"EB",X"1D",X"C3",X"65",X"1D",X"07",X"F0",X"54",X"49",X"4D",X"45",X"F0",X"4F",X"55",
		X"54",X"F0",X"FF",X"23",X"16",X"0D",X"EB",X"C9",X"E5",X"D5",X"CD",X"2B",X"1E",X"D1",X"E1",X"CD",
		X"ED",X"01",X"3E",X"B0",X"CD",X"10",X"1D",X"11",X"A4",X"4C",X"21",X"AD",X"42",X"C3",X"86",X"1E",
		X"E5",X"C1",X"3E",X"04",X"80",X"47",X"0A",X"32",X"B3",X"4C",X"C9",X"CD",X"20",X"1E",X"06",X"0B",
		X"11",X"A4",X"4C",X"7E",X"12",X"13",X"E7",X"10",X"FA",X"C9",X"06",X"0B",X"1A",X"77",X"13",X"E7",
		X"10",X"FA",X"C9",X"E5",X"C1",X"3E",X"04",X"C9",X"21",X"04",X"40",X"3E",X"40",X"CD",X"75",X"1E",
		X"2E",X"24",X"CD",X"75",X"1E",X"2E",X"03",X"3A",X"3F",X"4C",X"3D",X"C8",X"47",X"23",X"23",X"3D",
		X"20",X"FB",X"3E",X"16",X"E5",X"77",X"2B",X"3C",X"77",X"3C",X"DF",X"77",X"3C",X"23",X"77",X"E1",
		X"2B",X"2B",X"10",X"EE",X"C9",X"C5",X"06",X"08",X"77",X"23",X"10",X"FC",X"C1",X"C9",X"CD",X"43",
		X"1E",X"80",X"47",X"C5",X"E1",X"C9",X"E5",X"CD",X"7E",X"1E",X"CD",X"90",X"1E",X"E1",X"18",X"AA",
		X"06",X"0B",X"3A",X"B3",X"4C",X"77",X"E7",X"10",X"FC",X"C9",X"CB",X"7F",X"C8",X"F5",X"CD",X"C6",
		X"12",X"CD",X"11",X"07",X"E5",X"CD",X"20",X"1E",X"06",X"02",X"CD",X"30",X"1E",X"E1",X"E5",X"23",
		X"06",X"02",X"CD",X"33",X"1E",X"E1",X"11",X"D0",X"1E",X"E5",X"CD",X"ED",X"01",X"E1",X"22",X"B1",
		X"4C",X"3E",X"01",X"32",X"7F",X"4C",X"3E",X"50",X"32",X"7E",X"4C",X"CD",X"E9",X"12",X"F1",X"C9",
		X"02",X"1A",X"1B",X"FF",X"2A",X"B1",X"4C",X"E5",X"CD",X"7E",X"1E",X"06",X"02",X"E5",X"CD",X"92",
		X"1E",X"E1",X"23",X"06",X"02",X"CD",X"92",X"1E",X"E1",X"E5",X"06",X"02",X"11",X"A4",X"4C",X"CD",
		X"3C",X"1E",X"E1",X"23",X"06",X"02",X"CD",X"3C",X"1E",X"21",X"81",X"4C",X"C9",X"3E",X"80",X"CD",
		X"10",X"1D",X"C3",X"06",X"87",X"21",X"BE",X"43",X"06",X"06",X"C5",X"3E",X"09",X"CD",X"10",X"1D",
		X"00",X"06",X"0A",X"E5",X"CD",X"30",X"1E",X"E1",X"E5",X"06",X"0A",X"36",X"F0",X"E7",X"10",X"FB",
		X"3E",X"01",X"CD",X"10",X"1D",X"E1",X"2B",X"E5",X"11",X"A4",X"4C",X"06",X"0A",X"CD",X"3C",X"1E",
		X"E1",X"C1",X"10",X"D6",X"C9",X"21",X"BE",X"43",X"CD",X"97",X"1F",X"21",X"40",X"40",X"01",X"04",
		X"80",X"3E",X"F0",X"CF",X"21",X"BE",X"43",X"11",X"A4",X"4C",X"06",X"0A",X"CD",X"3C",X"1E",X"21",
		X"30",X"4C",X"01",X"01",X"0C",X"AF",X"CF",X"CD",X"D2",X"1C",X"CD",X"6B",X"1F",X"CD",X"5E",X"20",
		X"3E",X"20",X"CD",X"10",X"1D",X"CD",X"FC",X"23",X"C3",X"38",X"1D",X"06",X"03",X"C5",X"E5",X"3E",
		X"09",X"CD",X"10",X"1D",X"06",X"0A",X"CD",X"30",X"1E",X"E1",X"E5",X"06",X"0A",X"36",X"F0",X"E7",
		X"10",X"FB",X"3E",X"01",X"CD",X"10",X"1D",X"E1",X"E7",X"E5",X"11",X"A4",X"4C",X"06",X"0A",X"CD",
		X"3C",X"1E",X"E1",X"C1",X"10",X"D7",X"C9",X"06",X"0A",X"C3",X"30",X"1E",X"06",X"09",X"21",X"94",
		X"43",X"3E",X"2A",X"CD",X"2D",X"20",X"06",X"09",X"21",X"F4",X"41",X"3E",X"2B",X"CD",X"2D",X"20",
		X"3E",X"0A",X"21",X"44",X"43",X"CD",X"33",X"20",X"3E",X"0A",X"21",X"46",X"43",X"CD",X"46",X"20",
		X"3E",X"07",X"21",X"48",X"43",X"CD",X"33",X"20",X"3E",X"07",X"21",X"4A",X"43",X"CD",X"46",X"20",
		X"3E",X"05",X"21",X"4C",X"43",X"CD",X"33",X"20",X"3E",X"05",X"21",X"4E",X"43",X"CD",X"46",X"20",
		X"3E",X"03",X"21",X"50",X"43",X"CD",X"33",X"20",X"3E",X"03",X"21",X"52",X"43",X"CD",X"46",X"20",
		X"3E",X"01",X"21",X"54",X"43",X"CD",X"33",X"20",X"21",X"34",X"41",X"06",X"03",X"C5",X"E5",X"06",
		X"09",X"AF",X"CD",X"2D",X"20",X"E1",X"C1",X"DF",X"10",X"F3",X"21",X"AA",X"41",X"06",X"04",X"3E",
		X"01",X"CD",X"2D",X"20",X"C3",X"CA",X"96",X"21",X"94",X"41",X"06",X"09",X"1A",X"77",X"2B",X"2B",
		X"13",X"10",X"F9",X"C9",X"01",X"05",X"05",X"08",X"08",X"00",X"00",X"05",X"05",X"77",X"2B",X"2B",
		X"10",X"FB",X"C9",X"06",X"0A",X"A7",X"28",X"0A",X"F5",X"78",X"3D",X"77",X"F1",X"3D",X"E7",X"10",
		X"F4",X"C9",X"36",X"3B",X"18",X"F8",X"06",X"00",X"A7",X"28",X"0C",X"70",X"3D",X"04",X"E7",X"F5",
		X"78",X"FE",X"0A",X"20",X"06",X"F1",X"C9",X"36",X"3B",X"18",X"F2",X"F1",X"18",X"EA",X"3E",X"06",
		X"06",X"14",X"21",X"34",X"45",X"E5",X"C5",X"06",X"09",X"CD",X"2D",X"20",X"C1",X"E1",X"DF",X"10",
		X"F4",X"C3",X"5A",X"22",X"3E",X"0E",X"32",X"2E",X"4C",X"C3",X"46",X"14",X"01",X"04",X"80",X"3A",
		X"2E",X"4C",X"C9",X"3E",X"0F",X"32",X"2E",X"4C",X"C3",X"75",X"04",X"3E",X"0D",X"18",X"F6",X"3E",
		X"08",X"18",X"F2",X"C3",X"52",X"09",X"00",X"00",X"0D",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"00",
		X"BC",X"0E",X"0E",X"0C",X"0E",X"AE",X"0D",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"BB",X"00",X"00",X"0C",X"0E",X"0E",X"0D",X"0F",X"0F",X"0F",X"0F",
		X"DB",X"F0",X"F0",X"FA",X"F0",X"F0",X"9C",X"0E",X"0E",X"0E",X"0E",X"0E",X"8E",X"0E",X"0E",X"0E",
		X"0E",X"0C",X"0E",X"0E",X"0E",X"BB",X"00",X"00",X"0A",X"00",X"00",X"0C",X"DE",X"FE",X"FE",X"FE",
		X"EB",X"E0",X"E0",X"E0",X"E0",X"E0",X"AB",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"0A",X"C0",X"E0",X"E0",X"E0",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"80",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"6D",X"0F",X"0F",X"7F",X"00",X"0D",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"0D",X"0F",X"9F",X"00",X"00",X"0D",X"0F",X"0F",
		X"D9",X"F0",X"F0",X"F0",X"F0",X"F0",X"7C",X"0E",X"0E",X"0E",X"00",X"0C",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0A",X"00",X"00",X"00",X"BB",X"00",X"00",X"0C",X"0E",X"DE",X"F0",X"F0",X"FC",X"0E",X"0E",
		X"CB",X"E0",X"E0",X"E0",X"E0",X"E0",X"0A",X"00",X"00",X"00",X"00",X"0A",X"90",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"00",X"C0",X"E0",X"E0",X"EA",X"00",X"00",
		X"AB",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"F0",
		X"F0",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"0A",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"B0",X"00",X"00",X"00",X"D0",X"F0",X"F9",X"F0",X"F0",X"C0",X"E0",X"E0",X"E0",
		X"E0",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"C0",X"E0",X"EA",X"E0",X"E0",X"B0",X"00",X"00",X"00",
		X"00",X"D0",X"F0",X"F0",X"F0",X"BB",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"A0",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"BB",X"00",X"00",X"90",X"00",X"07",X"B0",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"90",X"00",X"0B",X"90",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"BB",X"00",X"00",X"B0",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",
		X"DB",X"F0",X"F0",X"D0",X"F0",X"FB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"3A",X"40",X"4C",X"3C",X"32",X"40",
		X"4C",X"C3",X"32",X"80",X"16",X"01",X"43",X"09",X"94",X"42",X"09",X"CF",X"40",X"09",X"01",X"42",
		X"08",X"3A",X"41",X"08",X"C9",X"41",X"07",X"09",X"41",X"07",X"5A",X"42",X"06",X"6F",X"42",X"06",
		X"29",X"43",X"05",X"B5",X"41",X"05",X"BA",X"41",X"04",X"69",X"42",X"04",X"D5",X"41",X"03",X"70",
		X"41",X"03",X"2C",X"42",X"02",X"35",X"41",X"02",X"32",X"43",X"01",X"55",X"41",X"01",X"F4",X"42",
		X"00",X"9A",X"42",X"00",X"C6",X"42",X"00",X"E1",X"E5",X"E7",X"7E",X"FE",X"0A",X"DA",X"5D",X"0A",
		X"E1",X"2B",X"C9",X"E1",X"E5",X"DF",X"7E",X"FE",X"0A",X"DA",X"7E",X"0A",X"E1",X"2B",X"C9",X"E5",
		X"CD",X"6C",X"26",X"21",X"69",X"85",X"22",X"03",X"4C",X"21",X"0A",X"86",X"CD",X"9C",X"19",X"CD",
		X"EF",X"22",X"3A",X"9A",X"4C",X"CB",X"47",X"20",X"05",X"00",X"00",X"CD",X"5B",X"26",X"3E",X"13",
		X"E1",X"32",X"B4",X"4C",X"11",X"F3",X"4F",X"06",X"04",X"12",X"13",X"13",X"10",X"FB",X"C9",X"CD",
		X"DD",X"9A",X"EF",X"03",X"23",X"06",X"23",X"09",X"23",X"0C",X"23",X"0F",X"23",X"12",X"23",X"15",
		X"23",X"15",X"23",X"3E",X"60",X"11",X"3E",X"50",X"11",X"3E",X"48",X"11",X"3E",X"46",X"11",X"3E",
		X"44",X"11",X"3E",X"3F",X"11",X"3E",X"32",X"32",X"B6",X"4C",X"3E",X"FF",X"32",X"B5",X"4C",X"C9",
		X"3A",X"9A",X"4C",X"CB",X"47",X"C8",X"3A",X"2C",X"4C",X"CB",X"47",X"C8",X"3A",X"B5",X"4C",X"3D",
		X"32",X"B5",X"4C",X"F5",X"3A",X"B6",X"4C",X"FE",X"10",X"30",X"0B",X"CB",X"47",X"3A",X"B4",X"4C",
		X"20",X"01",X"AF",X"CD",X"E4",X"22",X"F1",X"C0",X"3D",X"32",X"B5",X"4C",X"3A",X"B6",X"4C",X"3D",
		X"32",X"B6",X"4C",X"C0",X"21",X"9A",X"4C",X"CB",X"86",X"CD",X"01",X"07",X"11",X"F3",X"4F",X"C3",
		X"4E",X"26",X"00",X"3A",X"9A",X"4C",X"CB",X"47",X"DD",X"7E",X"29",X"C8",X"E1",X"C9",X"3A",X"9A",
		X"4C",X"CB",X"47",X"3A",X"98",X"4C",X"C8",X"E1",X"C9",X"3A",X"00",X"50",X"CB",X"67",X"CA",X"A8",
		X"96",X"3A",X"B7",X"4C",X"A7",X"28",X"05",X"3D",X"32",X"B7",X"4C",X"C9",X"0E",X"00",X"3D",X"32",
		X"B7",X"4C",X"21",X"40",X"40",X"23",X"06",X"1B",X"7E",X"FE",X"0A",X"30",X"02",X"0C",X"00",X"23",
		X"10",X"F6",X"23",X"23",X"23",X"23",X"7D",X"FE",X"C0",X"20",X"EA",X"7C",X"FE",X"43",X"20",X"E5",
		X"3A",X"44",X"4C",X"CB",X"57",X"C0",X"C3",X"D7",X"34",X"06",X"2A",X"F0",X"3D",X"3D",X"3B",X"3B",
		X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"F0",X"2B",X"F0",X"F0",X"F0",X"3D",X"3D",X"30",X"FF",X"07",
		X"59",X"4F",X"55",X"52",X"F0",X"42",X"4F",X"4E",X"55",X"53",X"F0",X"F0",X"2B",X"FF",X"21",X"96",
		X"43",X"11",X"B9",X"23",X"CD",X"ED",X"01",X"21",X"7A",X"43",X"11",X"CF",X"23",X"CD",X"ED",X"01",
		X"C3",X"9C",X"1F",X"0A",X"0A",X"07",X"07",X"05",X"05",X"03",X"03",X"01",X"CD",X"D6",X"24",X"11",
		X"F3",X"23",X"1A",X"47",X"CD",X"90",X"24",X"CA",X"15",X"25",X"13",X"23",X"23",X"7B",X"FE",X"FC",
		X"20",X"F0",X"3E",X"01",X"21",X"58",X"47",X"E5",X"F5",X"21",X"80",X"25",X"22",X"03",X"4C",X"C3",
		X"A0",X"25",X"E1",X"06",X"02",X"77",X"E7",X"3C",X"F5",X"3E",X"03",X"CD",X"10",X"1D",X"F1",X"10",
		X"F4",X"FE",X"19",X"20",X"DF",X"21",X"58",X"43",X"18",X"06",X"3A",X"87",X"4C",X"E6",X"F0",X"C9",
		X"CD",X"6E",X"24",X"B0",X"0F",X"0F",X"0F",X"0F",X"4F",X"E7",X"CD",X"6E",X"24",X"B0",X"B1",X"32",
		X"7E",X"4C",X"21",X"7A",X"41",X"11",X"7E",X"4C",X"CD",X"66",X"24",X"3E",X"20",X"CD",X"10",X"1D",
		X"CD",X"69",X"94",X"C3",X"AA",X"25",X"CD",X"B2",X"14",X"AF",X"32",X"3A",X"41",X"C9",X"7E",X"06",
		X"00",X"FE",X"0A",X"D8",X"78",X"C9",X"11",X"58",X"43",X"1A",X"CD",X"98",X"24",X"4F",X"7E",X"B9",
		X"20",X"0B",X"CD",X"CE",X"24",X"E7",X"EB",X"E7",X"EB",X"10",X"EE",X"AF",X"C9",X"AF",X"3D",X"C9",
		X"E5",X"D5",X"CD",X"76",X"24",X"D1",X"E1",X"C9",X"C5",X"F5",X"E5",X"D5",X"3E",X"04",X"84",X"67",
		X"3E",X"04",X"82",X"57",X"D5",X"DD",X"E1",X"DD",X"46",X"00",X"7E",X"4F",X"16",X"07",X"3E",X"00",
		X"DD",X"77",X"00",X"77",X"F5",X"3E",X"04",X"CD",X"10",X"1D",X"F1",X"71",X"CD",X"E3",X"24",X"F5",
		X"3E",X"02",X"CD",X"10",X"1D",X"F1",X"15",X"20",X"E5",X"D1",X"E1",X"F1",X"C1",X"C9",X"F5",X"3E",
		X"09",X"CD",X"00",X"25",X"F1",X"C9",X"21",X"00",X"00",X"22",X"03",X"4C",X"CD",X"9C",X"19",X"21",
		X"44",X"43",X"C9",X"E5",X"F5",X"21",X"F5",X"24",X"22",X"0B",X"4C",X"AF",X"32",X"02",X"4C",X"F1",
		X"E1",X"DD",X"70",X"00",X"C9",X"06",X"6B",X"00",X"0F",X"02",X"07",X"6B",X"00",X"05",X"02",X"10",
		X"CD",X"10",X"1D",X"E5",X"21",X"00",X"00",X"22",X"0B",X"4C",X"AF",X"32",X"02",X"4C",X"3E",X"01",
		X"CD",X"10",X"1D",X"E1",X"C9",X"11",X"60",X"FE",X"19",X"E5",X"D1",X"CD",X"D9",X"96",X"CD",X"6E",
		X"24",X"B0",X"0F",X"0F",X"0F",X"0F",X"4F",X"E7",X"CD",X"6E",X"24",X"B0",X"B1",X"C3",X"07",X"26",
		X"E5",X"21",X"5A",X"25",X"22",X"03",X"4C",X"21",X"6A",X"25",X"CD",X"9C",X"19",X"EB",X"3E",X"04",
		X"84",X"67",X"3E",X"01",X"E5",X"06",X"05",X"77",X"E7",X"F5",X"3E",X"03",X"CD",X"10",X"1D",X"F1",
		X"3C",X"10",X"F4",X"FE",X"2E",X"E1",X"20",X"EC",X"18",X"20",X"07",X"27",X"00",X"0F",X"07",X"07",
		X"88",X"00",X"0F",X"07",X"07",X"6B",X"00",X"0F",X"07",X"10",X"06",X"6B",X"00",X"0F",X"07",X"06",
		X"2E",X"00",X"0F",X"07",X"06",X"E0",X"10",X"0F",X"07",X"10",X"E1",X"3E",X"20",X"C3",X"10",X"1D",
		X"07",X"56",X"00",X"0F",X"02",X"07",X"A7",X"00",X"0F",X"02",X"07",X"79",X"00",X"0F",X"02",X"10",
		X"06",X"CC",X"00",X"0F",X"05",X"06",X"0F",X"00",X"0F",X"05",X"06",X"F2",X"10",X"0F",X"05",X"10",
		X"21",X"90",X"25",X"CD",X"9C",X"19",X"F1",X"C3",X"22",X"24",X"CD",X"D6",X"24",X"21",X"BE",X"25",
		X"22",X"03",X"4C",X"21",X"C9",X"25",X"CD",X"D4",X"25",X"3E",X"10",X"C3",X"10",X"1D",X"02",X"88",
		X"00",X"0F",X"0F",X"02",X"6B",X"00",X"0F",X"0F",X"10",X"06",X"CC",X"00",X"0F",X"0F",X"06",X"2E",
		X"00",X"0F",X"0F",X"10",X"CD",X"9C",X"19",X"3E",X"5A",X"CD",X"10",X"1D",X"21",X"00",X"00",X"22",
		X"03",X"4C",X"22",X"07",X"4C",X"C9",X"CD",X"DD",X"9A",X"00",X"EF",X"FB",X"25",X"FB",X"25",X"FF",
		X"25",X"FF",X"25",X"03",X"26",X"03",X"26",X"03",X"26",X"03",X"26",X"21",X"53",X"14",X"C9",X"21",
		X"94",X"8A",X"C9",X"21",X"BF",X"34",X"C9",X"32",X"7F",X"4C",X"E7",X"C3",X"40",X"24",X"09",X"CD",
		X"F3",X"34",X"3E",X"10",X"46",X"23",X"5E",X"23",X"56",X"12",X"10",X"F9",X"C9",X"E5",X"21",X"00",
		X"15",X"22",X"85",X"4C",X"E1",X"C3",X"83",X"20",X"E5",X"2A",X"45",X"4C",X"23",X"7E",X"FE",X"10",
		X"28",X"34",X"E1",X"AF",X"3D",X"C9",X"AF",X"3D",X"C9",X"30",X"02",X"7D",X"C9",X"C1",X"C3",X"91",
		X"1C",X"06",X"04",X"21",X"B8",X"4C",X"1A",X"13",X"13",X"77",X"23",X"10",X"F9",X"C9",X"06",X"04",
		X"21",X"B8",X"4C",X"7E",X"12",X"13",X"13",X"23",X"10",X"F9",X"C9",X"CB",X"C7",X"32",X"9A",X"4C",
		X"11",X"F3",X"4F",X"C3",X"41",X"26",X"22",X"BC",X"4C",X"E1",X"AF",X"C9",X"2A",X"BC",X"4C",X"36",
		X"F0",X"3E",X"95",X"C3",X"50",X"13",X"22",X"0B",X"4C",X"3A",X"44",X"4C",X"CB",X"6F",X"C8",X"3E",
		X"01",X"C3",X"50",X"13",X"21",X"7C",X"43",X"11",X"5D",X"14",X"06",X"04",X"CD",X"B6",X"26",X"11",
		X"D4",X"23",X"06",X"09",X"CD",X"B6",X"26",X"CD",X"7B",X"25",X"21",X"7C",X"41",X"CD",X"39",X"80",
		X"CD",X"B2",X"14",X"2A",X"87",X"4C",X"CD",X"43",X"80",X"3E",X"40",X"CD",X"10",X"1D",X"CD",X"69",
		X"94",X"3E",X"50",X"C3",X"10",X"1D",X"1A",X"77",X"E7",X"3E",X"03",X"CD",X"10",X"1D",X"13",X"10",
		X"F5",X"C9",X"3E",X"40",X"CD",X"10",X"1D",X"21",X"AE",X"42",X"11",X"E5",X"26",X"06",X"0B",X"CD",
		X"B6",X"26",X"21",X"6D",X"80",X"22",X"03",X"4C",X"21",X"AB",X"86",X"CD",X"9C",X"19",X"3E",X"80",
		X"CD",X"10",X"1D",X"18",X"15",X"40",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"40",
		X"21",X"40",X"40",X"01",X"04",X"80",X"3E",X"40",X"CF",X"C9",X"CD",X"F0",X"26",X"CD",X"62",X"80",
		X"3A",X"3E",X"4C",X"21",X"0F",X"4E",X"06",X"05",X"4E",X"B9",X"38",X"0E",X"C3",X"99",X"97",X"2B",
		X"5E",X"2A",X"3C",X"4C",X"ED",X"52",X"F2",X"23",X"27",X"E1",X"11",X"10",X"00",X"19",X"10",X"E8",
		X"C3",X"A1",X"8A",X"E1",X"CD",X"A6",X"97",X"E5",X"7D",X"D6",X"0F",X"6F",X"FE",X"40",X"28",X"20",
		X"22",X"E3",X"4C",X"21",X"30",X"4E",X"11",X"40",X"4E",X"01",X"10",X"00",X"E5",X"C5",X"ED",X"B0",
		X"C1",X"E1",X"7D",X"ED",X"5B",X"E3",X"4C",X"BB",X"28",X"06",X"5F",X"D6",X"10",X"6F",X"18",X"E9",
		X"E1",X"11",X"3E",X"4C",X"06",X"03",X"1A",X"77",X"2B",X"1B",X"10",X"FA",X"3A",X"40",X"4C",X"77",
		X"2B",X"06",X"0C",X"3E",X"40",X"77",X"2B",X"10",X"FA",X"00",X"00",X"00",X"21",X"E5",X"42",X"3E",
		X"3B",X"06",X"04",X"E5",X"C5",X"06",X"08",X"77",X"E7",X"E7",X"3C",X"10",X"FA",X"C1",X"E1",X"23",
		X"23",X"23",X"10",X"EF",X"21",X"F1",X"42",X"11",X"A1",X"27",X"CD",X"ED",X"01",X"11",X"A6",X"27",
		X"21",X"71",X"42",X"CD",X"ED",X"01",X"11",X"AB",X"27",X"21",X"75",X"43",X"CD",X"ED",X"01",X"18",
		X"23",X"10",X"52",X"55",X"42",X"FF",X"07",X"45",X"4E",X"44",X"FF",X"06",X"59",X"4F",X"55",X"52",
		X"40",X"4E",X"41",X"4D",X"45",X"40",X"40",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",
		X"3B",X"3B",X"3B",X"FF",X"21",X"29",X"42",X"22",X"04",X"4D",X"21",X"15",X"42",X"22",X"06",X"4D",
		X"2A",X"00",X"4D",X"7D",X"D6",X"0F",X"6F",X"22",X"08",X"4D",X"21",X"FF",X"00",X"22",X"0A",X"4D",
		X"21",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"AF",X"32",X"0C",X"4D",
		X"2A",X"0A",X"4D",X"01",X"01",X"00",X"ED",X"42",X"22",X"0A",X"4D",X"C3",X"00",X"30",X"AB",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"30",X"10",X"21",X"FF",X"00",X"22",X"0A",X"4D",X"3A",X"0C",X"4D",X"3D",X"32",X"0C",X"4D",X"CA",
		X"F1",X"30",X"CD",X"2D",X"32",X"FE",X"0F",X"28",X"1F",X"21",X"0D",X"4D",X"CB",X"46",X"20",X"1D",
		X"2A",X"04",X"4D",X"36",X"40",X"FE",X"00",X"28",X"35",X"FE",X"01",X"28",X"46",X"FE",X"02",X"28",
		X"50",X"FE",X"03",X"28",X"59",X"C3",X"9C",X"30",X"21",X"0D",X"4D",X"CB",X"86",X"3A",X"2C",X"4C",
		X"CB",X"67",X"28",X"0D",X"2A",X"04",X"4D",X"36",X"81",X"2A",X"06",X"4D",X"36",X"80",X"C3",X"F0",
		X"27",X"2A",X"04",X"4D",X"36",X"40",X"2A",X"06",X"4D",X"36",X"40",X"C3",X"F0",X"27",X"7D",X"E6",
		X"1F",X"FE",X"06",X"28",X"07",X"7D",X"D6",X"03",X"6F",X"22",X"04",X"4D",X"21",X"0D",X"4D",X"CB",
		X"C6",X"18",X"CA",X"7C",X"FE",X"42",X"20",X"05",X"7D",X"FE",X"E0",X"30",X"EF",X"DF",X"DF",X"18",
		X"E8",X"7D",X"E6",X"1F",X"FE",X"12",X"28",X"E4",X"7D",X"C6",X"03",X"6F",X"18",X"DB",X"7C",X"FE",
		X"41",X"20",X"05",X"7D",X"FE",X"60",X"38",X"D4",X"E7",X"E7",X"18",X"CD",X"2A",X"04",X"4D",X"7C",
		X"FE",X"42",X"20",X"11",X"7D",X"FE",X"F2",X"28",X"2F",X"FE",X"B2",X"28",X"2B",X"FE",X"72",X"28",
		X"40",X"FE",X"32",X"28",X"3C",X"EB",X"2A",X"06",X"4D",X"7C",X"FE",X"40",X"20",X"05",X"7D",X"FE",
		X"B5",X"28",X"A9",X"EB",X"2B",X"7E",X"2A",X"08",X"4D",X"77",X"23",X"22",X"08",X"4D",X"2A",X"06",
		X"4D",X"77",X"E7",X"22",X"06",X"4D",X"18",X"94",X"2A",X"06",X"4D",X"7C",X"FE",X"42",X"28",X"8C",
		X"36",X"3B",X"DF",X"22",X"06",X"4D",X"2A",X"08",X"4D",X"36",X"40",X"2B",X"22",X"08",X"4D",X"18",
		X"E5",X"CD",X"F0",X"26",X"CD",X"02",X"31",X"3E",X"FF",X"CD",X"10",X"1D",X"CD",X"D6",X"24",X"C3",
		X"AF",X"01",X"CD",X"6B",X"31",X"DD",X"21",X"00",X"4E",X"0E",X"01",X"3E",X"07",X"06",X"05",X"FD",
		X"21",X"A7",X"43",X"FD",X"E5",X"E1",X"11",X"00",X"04",X"19",X"CD",X"9D",X"31",X"FD",X"71",X"00",
		X"F5",X"DD",X"7E",X"0C",X"CD",X"A8",X"31",X"F1",X"FD",X"E5",X"E1",X"11",X"20",X"FF",X"19",X"DD",
		X"E5",X"D1",X"E5",X"EB",X"11",X"0F",X"00",X"19",X"EB",X"E1",X"C5",X"F5",X"06",X"03",X"CD",X"CB",
		X"31",X"F1",X"C1",X"DD",X"E5",X"D1",X"FD",X"E5",X"E1",X"D5",X"11",X"00",X"FE",X"19",X"D1",X"C5",
		X"F5",X"06",X"0C",X"1A",X"77",X"E7",X"13",X"10",X"FA",X"F1",X"C1",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"11",X"10",X"00",X"DD",X"19",X"0C",X"3D",X"10",X"A9",X"C9",X"CD",X"00",X"01",X"11",X"89",
		X"31",X"21",X"45",X"41",X"CD",X"ED",X"01",X"11",X"8F",X"31",X"21",X"65",X"43",X"CD",X"ED",X"01",
		X"11",X"96",X"31",X"21",X"A5",X"42",X"C3",X"ED",X"01",X"12",X"4E",X"41",X"4D",X"45",X"FF",X"12",
		X"52",X"4F",X"55",X"4E",X"44",X"FF",X"12",X"53",X"43",X"4F",X"52",X"45",X"FF",X"F5",X"C5",X"06",
		X"1C",X"77",X"E7",X"10",X"FC",X"C1",X"F1",X"C9",X"F5",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"FD",
		X"77",X"A0",X"F1",X"E6",X"0F",X"FD",X"77",X"80",X"C9",X"1A",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"77",X"E7",X"1A",X"E6",X"0F",X"77",X"E7",X"1B",X"10",X"EF",X"C9",X"CD",X"B9",X"31",X"36",X"00",
		X"C9",X"4E",X"4F",X"4E",X"50",X"45",X"40",X"3D",X"40",X"40",X"40",X"40",X"40",X"03",X"70",X"32",
		X"00",X"54",X"41",X"4B",X"41",X"53",X"48",X"49",X"40",X"48",X"41",X"52",X"41",X"03",X"57",X"10",
		X"00",X"46",X"55",X"4D",X"49",X"4B",X"4F",X"40",X"59",X"41",X"4D",X"41",X"3D",X"01",X"60",X"09",
		X"00",X"52",X"45",X"49",X"4B",X"4F",X"40",X"49",X"5A",X"55",X"4D",X"49",X"40",X"01",X"54",X"05",
		X"00",X"41",X"54",X"53",X"55",X"4B",X"4F",X"40",X"4B",X"49",X"42",X"41",X"40",X"01",X"32",X"04",
		X"00",X"21",X"D1",X"31",X"11",X"00",X"4E",X"01",X"50",X"00",X"ED",X"B0",X"C9",X"06",X"A0",X"10",
		X"FE",X"CD",X"62",X"01",X"3A",X"2E",X"4C",X"06",X"F0",X"10",X"FE",X"C9",X"E5",X"F5",X"DD",X"E5",
		X"E1",X"7D",X"C6",X"FD",X"6F",X"46",X"F1",X"E1",X"80",X"DD",X"77",X"21",X"C9",X"3A",X"9A",X"4C",
		X"CB",X"4F",X"C0",X"3A",X"88",X"4C",X"C3",X"99",X"32",X"3E",X"FD",X"21",X"9A",X"4C",X"18",X"20",
		X"32",X"FD",X"4C",X"32",X"FE",X"4C",X"C3",X"9F",X"19",X"CB",X"CE",X"21",X"9A",X"4C",X"CB",X"8E",
		X"AF",X"18",X"1D",X"3D",X"32",X"9E",X"4C",X"C0",X"21",X"BE",X"4C",X"CB",X"96",X"AF",X"18",X"10",
		X"CB",X"CE",X"CD",X"60",X"32",X"00",X"00",X"21",X"00",X"00",X"22",X"07",X"4C",X"C3",X"9F",X"19",
		X"CD",X"60",X"32",X"CD",X"01",X"07",X"C3",X"9F",X"19",X"FE",X"01",X"28",X"BC",X"FE",X"00",X"3E",
		X"FC",X"28",X"B8",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"0D",
		X"0F",X"0F",X"0F",X"BC",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0B",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"0C",
		X"0E",X"0E",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0F",X"0F",X"BB",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"09",X"00",X"60",X"00",X"00",X"09",X"00",X"00",X"00",
		X"0C",X"0E",X"0E",X"BB",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"07",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0F",X"6F",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"0C",X"0E",X"7E",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B8",X"00",X"00",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"FB",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"B6",X"00",X"00",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E6",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"C8",X"E0",X"E0",X"E0",X"EA",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"B6",X"00",X"00",X"00",X"00",X"B0",X"00",X"08",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"A0",X"00",X"06",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"60",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"70",X"00",X"00",X"0B",X"90",
		X"00",X"00",X"00",X"D6",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"90",X"00",X"00",X"B7",X"1E",X"C3",X"40",X"09",X"63",X"42",X"09",X"C8",X"42",X"09",X"4A",X"42",
		X"08",X"96",X"41",X"08",X"17",X"43",X"08",X"CE",X"42",X"07",X"2E",X"41",X"07",X"52",X"43",X"07",
		X"B2",X"42",X"06",X"77",X"42",X"06",X"43",X"41",X"06",X"C3",X"41",X"05",X"8C",X"41",X"05",X"89",
		X"43",X"05",X"CE",X"40",X"04",X"52",X"42",X"04",X"7B",X"42",X"04",X"49",X"40",X"03",X"25",X"43",
		X"03",X"CE",X"41",X"03",X"4E",X"40",X"02",X"43",X"42",X"02",X"4E",X"42",X"02",X"EA",X"41",X"01",
		X"D6",X"41",X"01",X"AE",X"43",X"01",X"4E",X"41",X"40",X"23",X"41",X"00",X"E8",X"42",X"00",X"06",
		X"94",X"40",X"7E",X"41",X"72",X"43",X"AC",X"41",X"C6",X"41",X"E5",X"42",X"E5",X"21",X"00",X"25",
		X"22",X"85",X"4C",X"E1",X"C3",X"8F",X"20",X"CB",X"6F",X"C0",X"CB",X"77",X"C0",X"79",X"FE",X"01",
		X"CA",X"DC",X"25",X"A7",X"C0",X"C3",X"DE",X"1C",X"CD",X"9C",X"19",X"3E",X"10",X"CD",X"10",X"1D",
		X"C3",X"DC",X"25",X"21",X"C9",X"43",X"11",X"8F",X"31",X"CD",X"D5",X"01",X"3A",X"40",X"4C",X"2E",
		X"E6",X"47",X"E6",X"0F",X"77",X"23",X"78",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"77",X"11",X"EF",
		X"43",X"21",X"0F",X"4E",X"AF",X"12",X"1E",X"F5",X"CD",X"09",X"13",X"C3",X"E6",X"25",X"AF",X"32",
		X"2D",X"4C",X"3C",X"32",X"40",X"4C",X"CD",X"CF",X"9B",X"CD",X"00",X"01",X"CD",X"52",X"09",X"CD",
		X"12",X"0D",X"CD",X"5B",X"35",X"CD",X"77",X"35",X"CD",X"9F",X"36",X"CD",X"D6",X"9B",X"06",X"0E",
		X"CD",X"45",X"35",X"18",X"F0",X"3A",X"26",X"4C",X"A7",X"20",X"03",X"10",X"F8",X"C9",X"21",X"30",
		X"4C",X"06",X"0C",X"36",X"00",X"23",X"10",X"FB",X"C3",X"0D",X"90",X"CD",X"E0",X"06",X"CB",X"86",
		X"3E",X"30",X"CD",X"C1",X"01",X"AF",X"32",X"44",X"4C",X"3C",X"32",X"81",X"4C",X"32",X"42",X"4C",
		X"21",X"08",X"37",X"CD",X"99",X"37",X"C9",X"3A",X"41",X"4C",X"A7",X"28",X"05",X"3D",X"32",X"41",
		X"4C",X"C9",X"3E",X"40",X"32",X"41",X"4C",X"3A",X"43",X"4C",X"A7",X"C2",X"14",X"36",X"2A",X"45",
		X"4C",X"3A",X"42",X"4C",X"3D",X"28",X"03",X"23",X"18",X"FA",X"3A",X"42",X"4C",X"3C",X"32",X"42",
		X"4C",X"7E",X"47",X"E6",X"0F",X"32",X"47",X"4C",X"78",X"E6",X"F0",X"C2",X"F8",X"35",X"CD",X"0E",
		X"36",X"3E",X"08",X"32",X"43",X"4C",X"C9",X"AF",X"CD",X"0E",X"36",X"3A",X"47",X"4C",X"FE",X"01",
		X"28",X"0B",X"CD",X"26",X"36",X"3E",X"01",X"32",X"01",X"50",X"C9",X"AE",X"35",X"AF",X"CD",X"D6",
		X"24",X"CD",X"42",X"36",X"18",X"EF",X"AF",X"CD",X"D6",X"24",X"3A",X"47",X"4C",X"FE",X"01",X"3A",
		X"44",X"4C",X"CB",X"9F",X"20",X"02",X"CB",X"DF",X"CB",X"FF",X"CB",X"8F",X"32",X"44",X"4C",X"3E",
		X"20",X"32",X"43",X"4C",X"00",X"00",X"00",X"C9",X"CB",X"77",X"20",X"0B",X"CB",X"6F",X"20",X"B7",
		X"CB",X"67",X"20",X"D2",X"C3",X"6E",X"37",X"21",X"44",X"4C",X"CB",X"CE",X"18",X"A3",X"21",X"44",
		X"4C",X"CB",X"8E",X"C9",X"F5",X"3A",X"44",X"4C",X"CB",X"4F",X"20",X"04",X"00",X"C3",X"79",X"37",
		X"F1",X"3D",X"32",X"43",X"4C",X"C9",X"CD",X"0E",X"07",X"23",X"E7",X"E7",X"7E",X"FE",X"0A",X"CD",
		X"5B",X"36",X"22",X"51",X"4C",X"CD",X"E4",X"0A",X"CB",X"D6",X"CB",X"9E",X"3E",X"0C",X"32",X"FC",
		X"4F",X"C9",X"CD",X"0E",X"07",X"23",X"DF",X"7E",X"FE",X"0A",X"CD",X"7A",X"36",X"22",X"51",X"4C",
		X"CD",X"E4",X"0A",X"CB",X"D6",X"CB",X"DE",X"3E",X"0E",X"18",X"E3",X"30",X"19",X"E5",X"E7",X"7E",
		X"FE",X"0A",X"E1",X"38",X"02",X"2B",X"C9",X"C1",X"2B",X"22",X"51",X"4C",X"CD",X"B0",X"0A",X"CB",
		X"EE",X"CB",X"96",X"C3",X"3A",X"36",X"E1",X"C3",X"3C",X"36",X"30",X"19",X"E5",X"DF",X"7E",X"FE",
		X"0A",X"E1",X"38",X"02",X"2B",X"C9",X"C1",X"2B",X"22",X"51",X"4C",X"CD",X"B0",X"0A",X"CB",X"EE",
		X"CB",X"96",X"C3",X"55",X"36",X"E1",X"C3",X"57",X"36",X"CD",X"0C",X"0A",X"C3",X"14",X"10",X"3A",
		X"44",X"4C",X"CB",X"67",X"C8",X"21",X"30",X"4C",X"06",X"08",X"36",X"00",X"23",X"10",X"FB",X"3E",
		X"20",X"CD",X"C1",X"01",X"3A",X"FD",X"4F",X"32",X"7E",X"4F",X"3E",X"11",X"32",X"FD",X"4F",X"06",
		X"10",X"3E",X"80",X"32",X"FC",X"4F",X"3E",X"05",X"CD",X"C1",X"01",X"3E",X"84",X"32",X"FC",X"4F",
		X"3E",X"05",X"CD",X"C1",X"01",X"10",X"EA",X"3E",X"80",X"CD",X"C1",X"01",X"C1",X"C9",X"F5",X"3A",
		X"44",X"4C",X"CB",X"E7",X"32",X"44",X"4C",X"F1",X"C9",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"2A",
		X"3A",X"4C",X"7C",X"92",X"F2",X"F9",X"36",X"ED",X"44",X"FE",X"09",X"D0",X"7D",X"93",X"F2",X"03",
		X"37",X"ED",X"44",X"FE",X"09",X"38",X"D7",X"C9",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"21",
		X"40",X"01",X"21",X"40",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"21",X"40",X"40",X"01",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"40",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"11",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"13",X"01",X"00",X"00",X"00",X"00",
		X"23",X"40",X"03",X"03",X"23",X"40",X"03",X"03",X"03",X"13",X"03",X"03",X"23",X"03",X"02",X"02",
		X"02",X"02",X"03",X"13",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"80",X"21",X"44",
		X"4C",X"CB",X"C6",X"3E",X"F0",X"32",X"43",X"4C",X"C9",X"CB",X"47",X"20",X"04",X"F1",X"C3",X"99",
		X"08",X"F1",X"3D",X"32",X"43",X"4C",X"3A",X"3B",X"4C",X"3D",X"32",X"3B",X"4C",X"CD",X"0E",X"07",
		X"23",X"23",X"7E",X"FE",X"F6",X"D8",X"C3",X"DE",X"36",X"ED",X"5F",X"CB",X"4F",X"28",X"03",X"21",
		X"A6",X"37",X"22",X"45",X"4C",X"C9",X"03",X"03",X"03",X"00",X"00",X"00",X"03",X"21",X"01",X"01",
		X"11",X"01",X"01",X"23",X"03",X"03",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"23",X"03",
		X"03",X"03",X"03",X"23",X"01",X"11",X"03",X"23",X"40",X"03",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"03",X"23",X"03",X"03",X"23",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"11",X"01",X"01",X"01",X"11",X"01",X"01",X"11",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
