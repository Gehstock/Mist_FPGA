library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj_7n is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj_7n is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"00",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"D0",X"BC",X"BC",X"FC",X"F0",X"E0",X"C0",X"E0",X"F0",X"80",X"DC",
		X"00",X"00",X"00",X"E0",X"E0",X"E0",X"F0",X"60",X"FC",X"FF",X"FF",X"C3",X"E0",X"F0",X"80",X"DC",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"F0",X"FC",X"FE",X"FE",X"84",X"E0",X"F0",X"80",X"DC",
		X"00",X"00",X"3C",X"FC",X"FC",X"FA",X"FF",X"6F",X"FE",X"FC",X"F0",X"E0",X"E0",X"F0",X"80",X"DC",
		X"00",X"F8",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"DE",X"FF",X"FB",X"F3",X"E0",X"F0",X"F8",X"40",X"EE",X"BC",
		X"00",X"00",X"38",X"F8",X"F8",X"F8",X"FC",X"F8",X"F8",X"F0",X"E0",X"F0",X"F8",X"40",X"EE",X"BC",
		X"00",X"00",X"00",X"FE",X"FE",X"FF",X"77",X"FF",X"FE",X"F0",X"80",X"DE",X"FC",X"F8",X"C0",X"00",
		X"FC",X"1C",X"DC",X"38",X"78",X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F8",X"F8",X"78",X"E0",X"F0",X"F0",X"F0",X"B8",X"F8",X"1C",X"7C",
		X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"71",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FE",X"FE",X"FC",X"F0",X"F0",
		X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"F0",X"F8",X"F8",X"F0",X"F8",X"BC",X"FE",X"FE",X"EE",X"DE",X"8C",X"C0",X"00",X"70",
		X"00",X"20",X"F0",X"F8",X"F8",X"F0",X"F8",X"BC",X"FE",X"F8",X"EE",X"DE",X"8C",X"C0",X"00",X"70",
		X"00",X"20",X"F0",X"F8",X"F8",X"F0",X"F8",X"BC",X"FE",X"FE",X"EE",X"DE",X"8C",X"C0",X"00",X"70",
		X"00",X"3C",X"FC",X"FC",X"F8",X"FB",X"EF",X"FF",X"FE",X"F0",X"80",X"DC",X"38",X"20",X"F8",X"C0",
		X"00",X"FC",X"FC",X"FB",X"EF",X"FF",X"FE",X"70",X"80",X"DE",X"3C",X"F8",X"C0",X"00",X"00",X"00",
		X"B0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F8",X"F8",X"DC",X"FC",X"FC",X"F8",X"F8",X"FC",X"1C",X"CE",X"CF",X"DB",X"92",X"90",
		X"C0",X"E0",X"F8",X"F8",X"DC",X"FD",X"FF",X"F7",X"FE",X"FE",X"1C",X"C8",X"C8",X"D8",X"90",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"68",X"FA",X"FF",X"FF",X"FF",X"F0",X"88",X"80",
		X"EE",X"9C",X"10",X"00",X"90",X"E8",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"F8",X"FC",X"FC",X"F8",X"F0",X"FE",X"BE",X"FE",X"F8",X"F0",X"E0",X"F0",X"80",X"DC",
		X"00",X"08",X"78",X"FC",X"FC",X"FC",X"FC",X"DF",X"FF",X"FC",X"F8",X"F0",X"F8",X"40",X"EE",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"70",X"B8",X"FC",X"4C",X"06",X"06",X"06",X"06",X"06",X"06",X"0C",X"1C",X"38",X"F0",X"C0",
		X"38",X"DD",X"EA",X"C0",X"40",X"60",X"A4",X"A0",X"F0",X"F0",X"72",X"B0",X"B8",X"D8",X"D8",X"F0",
		X"B0",X"F0",X"F8",X"FC",X"8C",X"06",X"06",X"06",X"06",X"06",X"06",X"0C",X"1C",X"38",X"F0",X"C0",
		X"6B",X"77",X"D6",X"60",X"69",X"E0",X"F0",X"70",X"B0",X"B8",X"D8",X"D8",X"F8",X"F0",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"52",X"52",X"F7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"10",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"7E",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"F0",X"F0",
		X"00",X"00",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"F1",X"52",X"54",X"65",X"42",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"42",X"4C",X"50",X"52",X"8C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"5E",X"4A",X"4A",X"4C",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"50",X"50",X"5C",X"44",X"9C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"52",X"52",X"4C",X"52",X"8C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"54",X"54",X"54",X"54",X"26",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"54",X"54",X"74",X"14",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"14",X"64",X"83",X"94",X"67",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"E8",X"FC",X"FC",X"FF",X"7C",X"BC",X"60",X"E0",X"E0",X"20",X"80",X"97",X"77",X"E4",X"E0",
		X"C8",X"E8",X"FC",X"FC",X"FF",X"7D",X"BF",X"63",X"E0",X"E0",X"20",X"80",X"90",X"70",X"E0",X"E0",
		X"0E",X"7C",X"D0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"9A",X"8B",X"0B",X"13",X"F0",X"88",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"86",X"86",X"86",X"86",X"86",X"06",X"06",X"06",X"0E",X"0C",X"1C",X"38",X"F8",X"E0",X"80",X"00",
		X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",
		X"00",X"80",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"DE",X"BE",X"1A",X"50",X"78",X"78",X"70",X"30",
		X"00",X"80",X"80",X"C0",X"EC",X"FE",X"FF",X"FF",X"CD",X"A8",X"3C",X"BC",X"D8",X"D8",X"C0",X"00",
		X"F0",X"E0",X"C0",X"F0",X"FC",X"F0",X"F0",X"B3",X"3F",X"7F",X"67",X"4E",X"4E",X"04",X"00",X"00",
		X"E0",X"E0",X"C0",X"80",X"F0",X"F8",X"FC",X"FB",X"B7",X"7F",X"67",X"4E",X"4E",X"04",X"00",X"00",
		X"C0",X"C0",X"80",X"F0",X"F8",X"FC",X"FB",X"B7",X"7F",X"67",X"4E",X"4E",X"04",X"00",X"00",X"00",
		X"00",X"78",X"F0",X"C0",X"F0",X"F8",X"FC",X"FB",X"B7",X"7F",X"67",X"4E",X"4E",X"04",X"00",X"00",
		X"78",X"F0",X"C0",X"F0",X"F8",X"FC",X"FB",X"B7",X"7F",X"67",X"4E",X"4E",X"04",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"C0",X"00",X"E0",X"E0",X"30",X"00",X"CC",X"9C",X"FC",X"FC",X"1C",X"18",X"80",
		X"C0",X"80",X"00",X"00",X"00",X"E0",X"E0",X"30",X"00",X"CC",X"9C",X"FC",X"FC",X"1C",X"18",X"80",
		X"F0",X"E0",X"00",X"00",X"F0",X"F0",X"18",X"80",X"E6",X"CE",X"FE",X"FE",X"8E",X"8C",X"40",X"00",
		X"78",X"70",X"E0",X"00",X"00",X"0E",X"7C",X"78",X"80",X"CC",X"9C",X"FC",X"AC",X"AC",X"88",X"C0",
		X"C0",X"80",X"00",X"08",X"0E",X"0E",X"06",X"82",X"00",X"00",X"D8",X"F8",X"F8",X"38",X"30",X"00",
		X"EE",X"FE",X"EC",X"F8",X"F8",X"F8",X"FB",X"FF",X"FE",X"FC",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"E0",X"F0",X"E8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"C0",X"F0",X"E8",X"E8",X"E8",X"F8",X"F0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"C0",X"E0",X"F8",X"F0",X"F4",X"D4",X"9A",X"3E",X"9E",X"0C",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",
		X"00",X"00",X"00",X"20",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",X"00",
		X"00",X"20",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"C0",X"00",X"40",X"40",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"08",X"10",X"20",X"C0",X"00",X"40",X"40",X"40",X"A0",X"50",X"20",X"00",X"00",X"00",
		X"00",X"0A",X"12",X"26",X"46",X"8C",X"04",X"40",X"40",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"40",X"70",X"00",X"40",X"10",X"10",X"10",X"08",X"00",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"08",X"5C",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"04",X"1C",X"88",X"02",X"00",X"00",X"60",X"22",X"04",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"18",X"F0",X"11",X"31",X"73",X"F2",X"F4",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"33",X"C3",X"07",X"0F",X"0F",X"1F",X"3C",X"30",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"08",X"F0",X"01",X"07",X"1F",X"FF",X"FE",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"06",X"03",X"01",X"FF",X"FF",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"18",X"E0",X"01",X"07",X"1F",X"FF",X"FE",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"EE",X"EE",X"EE",X"EE",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"EE",X"EE",X"EE",X"EE",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"66",X"77",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"22",X"66",X"76",X"7F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"22",X"66",X"76",X"7F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"02",X"04",X"48",X"F8",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"01",X"02",X"8E",X"FC",X"14",X"4E",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"8F",X"F9",X"F2",X"E6",X"CF",X"11",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"3C",X"3C",X"3C",X"7E",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"19",X"E3",X"03",X"03",X"C3",X"C6",X"C4",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"03",X"0C",X"30",X"C0",X"0C",X"3C",X"3E",X"3F",X"3C",X"70",X"C0",X"00",
		X"00",X"E0",X"F0",X"C8",X"80",X"80",X"80",X"C4",X"60",X"70",X"30",X"32",X"60",X"C0",X"80",X"00",
		X"00",X"60",X"F0",X"98",X"0C",X"6C",X"6C",X"6C",X"4C",X"9C",X"38",X"F8",X"F0",X"E0",X"00",X"00",
		X"00",X"E0",X"F0",X"38",X"98",X"CC",X"EC",X"2C",X"8C",X"EC",X"FC",X"78",X"70",X"60",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"98",X"58",X"58",X"38",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"30",X"B0",X"30",X"B0",X"E0",X"60",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"B0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"E0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"08",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"48",X"08",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"10",X"E8",X"68",X"A8",X"A8",X"A8",X"A8",X"E8",X"10",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"0A",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"2A",X"12",X"C4",X"F8",X"E0",X"DC",X"C6",X"8E",X"D4",X"C8",X"D0",X"C0",X"00",X"00",X"00",
		X"20",X"29",X"12",X"C2",X"F8",X"E0",X"D8",X"C4",X"8E",X"CE",X"CA",X"C0",X"C0",X"00",X"00",X"00",
		X"94",X"54",X"54",X"14",X"C0",X"F8",X"E0",X"DC",X"CE",X"8B",X"C9",X"C5",X"C0",X"C0",X"00",X"00",
		X"29",X"29",X"72",X"66",X"78",X"60",X"F8",X"CC",X"C6",X"8F",X"DF",X"7B",X"E3",X"C6",X"5C",X"38",
		X"52",X"52",X"64",X"70",X"60",X"6E",X"F7",X"CF",X"CB",X"8A",X"C2",X"46",X"C4",X"C0",X"40",X"20",
		X"48",X"24",X"64",X"60",X"78",X"60",X"FC",X"C6",X"CF",X"9F",X"DB",X"56",X"C6",X"CC",X"40",X"20",
		X"E0",X"04",X"EA",X"EA",X"CF",X"E7",X"FB",X"EE",X"E0",X"D8",X"24",X"12",X"09",X"00",X"00",X"00",
		X"E0",X"04",X"EA",X"EA",X"CF",X"E7",X"FB",X"EE",X"E0",X"D0",X"20",X"28",X"48",X"08",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"C0",X"9C",X"BE",X"E0",X"E0",X"E0",X"F0",X"F1",X"FF",X"1F",X"3F",X"3E",X"5E",X"1C",X"18",
		X"0E",X"1C",X"08",X"04",X"6C",X"FC",X"FC",X"FC",X"F8",X"F8",X"78",X"30",X"30",X"20",X"40",X"00",
		X"1E",X"38",X"1E",X"1C",X"1C",X"9C",X"F8",X"F0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"3B",X"36",X"3E",X"7E",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",X"E0",X"60",X"00",X"00",X"00",X"00",
		X"FF",X"EF",X"EF",X"EF",X"E0",X"0F",X"E0",X"20",X"20",X"20",X"20",X"E1",X"EF",X"2F",X"21",X"F0",
		X"5F",X"5F",X"5F",X"2F",X"17",X"08",X"07",X"00",X"00",X"80",X"E0",X"FF",X"3F",X"00",X"00",X"00",
		X"2F",X"2F",X"2F",X"E0",X"DE",X"0E",X"46",X"52",X"5A",X"1A",X"82",X"1A",X"5A",X"52",X"46",X"0E",
		X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"7C",X"BC",X"5E",X"5E",X"5E",X"5E",X"5E",X"DE",X"00",
		X"5E",X"5F",X"5F",X"2F",X"17",X"0B",X"04",X"03",X"00",X"80",X"E0",X"FF",X"3F",X"00",X"00",X"00",
		X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"DE",X"00",X"2F",X"2F",X"2F",X"E0",
		X"00",X"2F",X"2F",X"2F",X"E0",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",
		X"00",X"60",X"80",X"7F",X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"1E",X"1F",X"FF",
		X"FF",X"EF",X"EF",X"EF",X"E0",X"0F",X"E0",X"20",X"20",X"20",X"20",X"E1",X"EF",X"2F",X"21",X"F0",
		X"FF",X"EF",X"EF",X"EF",X"60",X"8F",X"60",X"20",X"20",X"20",X"20",X"61",X"EF",X"AF",X"21",X"70",
		X"EF",X"EF",X"EF",X"E0",X"0F",X"E0",X"A0",X"20",X"20",X"20",X"20",X"E1",X"EF",X"EF",X"2F",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"24",X"68",X"70",X"64",X"6C",X"ED",X"D9",X"FB",X"BB",X"FE",X"DE",X"DE",X"CC",X"48",X"20",
		X"40",X"20",X"A0",X"A0",X"80",X"80",X"80",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"80",
		X"50",X"48",X"08",X"F0",X"F0",X"E0",X"EC",X"C6",X"83",X"47",X"6D",X"6A",X"4A",X"44",X"0C",X"00",
		X"40",X"20",X"A0",X"A0",X"80",X"80",X"80",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"80",
		X"00",X"80",X"40",X"40",X"E0",X"B0",X"B0",X"E0",X"80",X"00",X"40",X"30",X"D8",X"E0",X"F8",X"70",
		X"00",X"80",X"40",X"40",X"E0",X"B0",X"B0",X"E0",X"90",X"1C",X"5E",X"1E",X"8E",X"04",X"00",X"00",
		X"00",X"80",X"40",X"40",X"E0",X"B8",X"B2",X"E6",X"9E",X"1C",X"40",X"00",X"80",X"00",X"00",X"00",
		X"C0",X"20",X"E2",X"D6",X"3C",X"68",X"80",X"10",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"03",X"4F",X"1E",X"90",X"E0",X"B0",X"B0",X"E0",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"03",X"4F",X"1E",X"90",X"E0",X"B0",X"B0",X"E0",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"A0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"18",X"18",X"18",X"F0",X"F0",X"A0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"FE",X"AE",X"5C",X"FC",X"18",X"18",X"18",X"F0",X"F0",X"A0",X"80",X"80",X"00",
		X"FC",X"06",X"FA",X"AE",X"5E",X"FC",X"FC",X"18",X"18",X"18",X"F0",X"F0",X"A0",X"80",X"80",X"00",
		X"FC",X"06",X"FA",X"FE",X"AE",X"5C",X"FC",X"18",X"18",X"18",X"F0",X"F0",X"A0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"06",X"03",X"FF",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FE",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"10",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"10",X"00",
		X"00",X"30",X"30",X"30",X"30",X"32",X"32",X"32",X"32",X"32",X"32",X"30",X"30",X"30",X"30",X"00",
		X"40",X"60",X"60",X"64",X"64",X"66",X"66",X"66",X"66",X"66",X"66",X"64",X"64",X"60",X"60",X"40",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"48",X"08",X"10",X"00",X"80",X"80",X"80",
		X"00",X"00",X"E0",X"10",X"E8",X"68",X"A8",X"A8",X"A8",X"A8",X"E8",X"10",X"E0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"E0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"F8",X"C0",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"80",X"80",X"80",X"E0",X"F0",X"B8",X"D8",X"FF",X"D8",X"B8",X"F0",X"E0",X"80",X"80",X"80",X"80",
		X"80",X"80",X"F0",X"F8",X"9C",X"CC",X"EC",X"FF",X"EC",X"CC",X"9C",X"F8",X"F0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"10",X"00",X"C0",X"E0",X"E4",X"E0",X"C0",X"00",X"00",X"10",X"80",X"00",X"00",
		X"80",X"00",X"04",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",X"00",
		X"00",X"00",X"00",X"40",X"60",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"C0",X"E0",X"00",
		X"80",X"80",X"80",X"80",X"90",X"B0",X"B8",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B8",X"B8",X"B0",
		X"80",X"80",X"90",X"90",X"90",X"90",X"FC",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B8",X"B8",X"B0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"A0",X"A0",X"B0",X"B0",X"B0",X"B8",X"B8",X"B0",
		X"00",X"80",X"80",X"C0",X"EC",X"FE",X"FF",X"FF",X"CD",X"A8",X"3C",X"BC",X"D8",X"D8",X"C0",X"00",
		X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"F0",X"F0",X"78",X"F8",X"80",X"60",X"00",
		X"20",X"70",X"70",X"39",X"3E",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"78",X"00",X"00",
		X"00",X"00",X"84",X"8E",X"CE",X"CC",X"FC",X"FE",X"FF",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",
		X"C0",X"E0",X"E0",X"E0",X"C0",X"10",X"F8",X"F8",X"E4",X"FE",X"FE",X"FC",X"FC",X"FC",X"F0",X"EC",
		X"00",X"20",X"66",X"F7",X"F3",X"FF",X"CF",X"DE",X"8C",X"C0",X"E0",X"F0",X"60",X"00",X"00",X"00",
		X"70",X"54",X"72",X"7E",X"C7",X"E3",X"EA",X"E6",X"F0",X"EC",X"12",X"09",X"04",X"00",X"00",X"00",
		X"60",X"F0",X"B0",X"EC",X"6E",X"96",X"DC",X"EC",X"E2",X"F3",X"E0",X"E4",X"56",X"5C",X"0E",X"00",
		X"04",X"0E",X"5F",X"57",X"14",X"C4",X"E2",X"E0",X"E8",X"FC",X"F6",X"DE",X"EC",X"B0",X"F0",X"60",
		X"00",X"00",X"00",X"10",X"92",X"A4",X"10",X"C0",X"CE",X"F3",X"E7",X"CF",X"EA",X"EA",X"A4",X"E8",
		X"80",X"00",X"00",X"C0",X"00",X"10",X"94",X"C0",X"D8",X"C0",X"F8",X"CC",X"1C",X"28",X"18",X"60",
		X"08",X"1C",X"66",X"1E",X"04",X"98",X"C0",X"D8",X"E0",X"D4",X"90",X"00",X"C0",X"00",X"00",X"80",
		X"00",X"40",X"00",X"90",X"E6",X"BF",X"BF",X"E6",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"D0",X"E4",X"B8",X"70",X"D4",X"B8",X"E8",X"5C",X"3C",X"D4",X"34",X"2C",X"18",X"00",
		X"00",X"0C",X"1E",X"18",X"D2",X"3C",X"5C",X"E8",X"B8",X"D4",X"70",X"B8",X"E4",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"10",X"F1",X"5D",X"5B",X"7E",X"CC",X"80",X"A0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"20",X"A0",X"C0",X"C0",X"F0",X"B8",X"98",X"50",
		X"30",X"F8",X"98",X"E8",X"C0",X"C0",X"A0",X"20",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"98",X"90",X"30",X"60",X"60",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"28",X"60",X"50",X"E0",X"A0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"CC",X"98",X"90",X"A0",X"20",X"40",X"40",X"C0",X"40",X"40",X"00",X"A4",X"F8",X"FC",X"78",X"30",
		X"CC",X"98",X"30",X"60",X"E0",X"40",X"C0",X"80",X"00",X"04",X"00",X"81",X"07",X"1E",X"0C",X"00",
		X"70",X"C0",X"82",X"00",X"00",X"00",X"18",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"8C",X"52",X"22",X"32",X"2C",X"20",X"10",X"08",X"05",X"03",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"6D",X"AF",X"AB",X"A9",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"B0",X"80",X"80",X"F0",X"30",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D8",X"D8",X"58",X"58",X"58",X"58",X"D8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"26",X"26",X"E6",X"26",X"26",X"26",X"26",X"FE",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"42",X"42",X"72",X"66",X"5E",X"52",X"42",X"FE",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1B",X"9B",X"9B",X"9F",X"8F",X"87",X"8F",X"9B",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"01",X"01",X"00",X"83",X"C3",X"CF",X"D3",X"D3",X"D3",X"D3",X"8F",X"00",X"01",X"01",X"FE",
		X"00",X"00",X"00",X"FE",X"01",X"01",X"00",X"83",X"CF",X"D3",X"D3",X"8F",X"00",X"01",X"01",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"01",X"01",X"CF",X"D3",X"DF",X"01",X"01",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
