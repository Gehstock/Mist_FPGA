library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mw05 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mw05 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"40",X"40",X"6D",X"40",X"B0",X"40",X"EB",X"40",X"1C",X"41",X"A4",X"41",X"DF",X"41",X"12",X"42",
		X"45",X"42",X"78",X"42",X"21",X"46",X"A4",X"42",X"85",X"43",X"62",X"44",X"CA",X"44",X"F6",X"44",
		X"22",X"45",X"A3",X"45",X"E4",X"45",X"2D",X"46",X"34",X"49",X"99",X"49",X"FD",X"49",X"27",X"4B",
		X"4F",X"4C",X"49",X"4D",X"41",X"4E",X"69",X"4E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D0",X"70",X"DB",X"17",X"02",X"0F",X"20",X"01",X"FE",X"00",X"28",X"CD",X"53",X"40",X"01",X"FD",
		X"01",X"30",X"76",X"D0",X"70",X"1B",X"18",X"02",X"0F",X"02",X"01",X"FE",X"00",X"20",X"01",X"FE",
		X"01",X"00",X"F8",X"00",X"01",X"FE",X"01",X"18",X"01",X"FF",X"FF",X"20",X"76",X"D0",X"30",X"DB",
		X"17",X"02",X"0F",X"20",X"01",X"FE",X"00",X"10",X"CD",X"90",X"40",X"01",X"FE",X"01",X"08",X"01",
		X"FE",X"FF",X"08",X"01",X"FD",X"01",X"10",X"AF",X"FE",X"FF",X"06",X"01",X"FE",X"01",X"10",X"76",
		X"D0",X"30",X"1B",X"18",X"02",X"0F",X"02",X"01",X"FE",X"01",X"18",X"01",X"FE",X"FF",X"10",X"01",
		X"FE",X"00",X"10",X"AF",X"FE",X"FF",X"08",X"01",X"FE",X"FF",X"08",X"01",X"FE",X"01",X"10",X"76",
		X"D0",X"A0",X"DB",X"17",X"02",X"0F",X"20",X"01",X"FE",X"00",X"18",X"CD",X"C7",X"40",X"01",X"FD",
		X"00",X"08",X"01",X"FD",X"FF",X"18",X"76",X"D0",X"A0",X"1B",X"18",X"02",X"0F",X"02",X"01",X"FE",
		X"00",X"18",X"01",X"FE",X"01",X"08",X"01",X"FE",X"FF",X"08",X"01",X"FE",X"00",X"10",X"AF",X"FE",
		X"FF",X"08",X"01",X"FE",X"01",X"10",X"01",X"FE",X"FF",X"10",X"76",X"D0",X"D0",X"DB",X"17",X"02",
		X"0F",X"20",X"01",X"FE",X"00",X"10",X"CD",X"0E",X"41",X"01",X"FE",X"00",X"10",X"AF",X"FF",X"FF",
		X"10",X"01",X"FE",X"FF",X"08",X"01",X"FE",X"01",X"10",X"01",X"FD",X"00",X"18",X"76",X"D0",X"D0",
		X"1B",X"18",X"02",X"0F",X"02",X"01",X"FE",X"00",X"20",X"C3",X"5E",X"40",X"D0",X"88",X"5B",X"18",
		X"02",X"0F",X"10",X"CD",X"3C",X"41",X"CD",X"51",X"41",X"01",X"FE",X"FF",X"0A",X"AF",X"FE",X"FF",
		X"02",X"01",X"FE",X"01",X"0A",X"AF",X"FE",X"01",X"02",X"C3",X"29",X"41",X"D0",X"76",X"5B",X"18",
		X"02",X"0F",X"10",X"AF",X"00",X"00",X"12",X"CD",X"66",X"41",X"01",X"FF",X"FF",X"10",X"C3",X"29",
		X"41",X"D0",X"9A",X"5B",X"18",X"02",X"0F",X"10",X"AF",X"00",X"00",X"12",X"CD",X"77",X"41",X"01",
		X"FF",X"01",X"10",X"C3",X"29",X"41",X"D0",X"5C",X"5B",X"18",X"02",X"0F",X"10",X"AF",X"00",X"00",
		X"12",X"CD",X"88",X"41",X"C3",X"4A",X"41",X"D0",X"B4",X"5B",X"18",X"02",X"0F",X"10",X"AF",X"00",
		X"00",X"12",X"CD",X"96",X"41",X"C3",X"5F",X"41",X"D0",X"40",X"5B",X"18",X"02",X"0F",X"10",X"AF",
		X"00",X"00",X"12",X"C3",X"4A",X"41",X"D0",X"CE",X"5B",X"18",X"02",X"0F",X"10",X"AF",X"00",X"00",
		X"12",X"C3",X"5F",X"41",X"D0",X"30",X"5B",X"19",X"01",X"0B",X"50",X"CD",X"B9",X"41",X"01",X"FE",
		X"01",X"14",X"01",X"FE",X"FF",X"14",X"C3",X"AE",X"41",X"D0",X"40",X"75",X"19",X"01",X"0B",X"50",
		X"AF",X"00",X"00",X"10",X"CD",X"CA",X"41",X"C3",X"AE",X"41",X"D0",X"40",X"68",X"19",X"01",X"0B",
		X"50",X"AF",X"00",X"00",X"10",X"01",X"FE",X"00",X"28",X"CD",X"40",X"40",X"C3",X"AE",X"41",X"D0",
		X"50",X"82",X"19",X"01",X"0B",X"50",X"CD",X"EC",X"41",X"C3",X"AE",X"41",X"D0",X"60",X"75",X"19",
		X"01",X"0B",X"50",X"AF",X"00",X"00",X"18",X"CD",X"FD",X"41",X"C3",X"AE",X"41",X"D0",X"50",X"68",
		X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",X"10",X"01",X"FE",X"00",X"28",X"CD",X"6D",X"40",X"C3",
		X"AE",X"41",X"D0",X"70",X"5B",X"19",X"01",X"0B",X"50",X"CD",X"1F",X"42",X"C3",X"AE",X"41",X"D0",
		X"80",X"68",X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",X"10",X"CD",X"30",X"42",X"C3",X"AE",X"41",
		X"D0",X"70",X"75",X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",X"10",X"01",X"FE",X"00",X"28",X"CD",
		X"B0",X"40",X"C3",X"AE",X"41",X"D0",X"90",X"82",X"19",X"01",X"0B",X"50",X"CD",X"52",X"42",X"C3",
		X"AE",X"41",X"D0",X"A0",X"68",X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",X"10",X"CD",X"63",X"42",
		X"C3",X"AE",X"41",X"D0",X"90",X"75",X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",X"10",X"01",X"FE",
		X"00",X"20",X"CD",X"EB",X"40",X"C3",X"AE",X"41",X"D0",X"B0",X"5B",X"19",X"01",X"0B",X"50",X"CD",
		X"85",X"42",X"C3",X"AE",X"41",X"D0",X"C0",X"5B",X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",X"10",
		X"CD",X"96",X"42",X"C3",X"AE",X"41",X"D0",X"B0",X"5B",X"19",X"01",X"0B",X"50",X"AF",X"00",X"00",
		X"18",X"C3",X"AE",X"41",X"D0",X"80",X"9B",X"18",X"02",X"0F",X"30",X"CD",X"E9",X"42",X"01",X"FF",
		X"FF",X"10",X"01",X"FF",X"01",X"10",X"CD",X"1F",X"43",X"01",X"FF",X"00",X"10",X"CD",X"2B",X"43",
		X"01",X"FF",X"00",X"10",X"AF",X"FF",X"FF",X"10",X"01",X"FF",X"FF",X"10",X"CD",X"35",X"43",X"01",
		X"FF",X"FF",X"10",X"CD",X"3F",X"43",X"01",X"FF",X"FF",X"10",X"CD",X"49",X"43",X"01",X"FF",X"00",
		X"10",X"CD",X"53",X"43",X"01",X"FF",X"00",X"30",X"76",X"D0",X"60",X"9B",X"18",X"02",X"0F",X"30",
		X"AF",X"00",X"00",X"60",X"01",X"FF",X"FF",X"10",X"01",X"FF",X"01",X"10",X"CD",X"5D",X"43",X"01",
		X"FF",X"00",X"10",X"CD",X"67",X"43",X"01",X"FF",X"00",X"20",X"AF",X"FF",X"01",X"10",X"01",X"FF",
		X"01",X"10",X"CD",X"71",X"43",X"01",X"FF",X"00",X"10",X"CD",X"7B",X"43",X"C3",X"E4",X"42",X"A0",
		X"80",X"01",X"1C",X"02",X"05",X"66",X"01",X"FD",X"00",X"30",X"76",X"90",X"8A",X"01",X"1C",X"02",
		X"05",X"66",X"C3",X"26",X"43",X"60",X"60",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"50",
		X"58",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"40",X"40",X"01",X"1C",X"02",X"05",X"66",
		X"C3",X"26",X"43",X"30",X"4A",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"A0",X"60",X"01",
		X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"90",X"6A",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",
		X"43",X"50",X"80",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"38",X"70",X"01",X"1C",X"02",
		X"05",X"66",X"C3",X"26",X"43",X"D0",X"A0",X"9B",X"18",X"02",X"0F",X"30",X"CD",X"C8",X"43",X"01",
		X"FF",X"00",X"10",X"CD",X"FE",X"43",X"01",X"FF",X"00",X"10",X"CD",X"08",X"44",X"01",X"FF",X"00",
		X"10",X"AF",X"FF",X"00",X"10",X"01",X"FF",X"01",X"10",X"CD",X"12",X"44",X"01",X"FF",X"01",X"10",
		X"CD",X"1C",X"44",X"01",X"FF",X"01",X"08",X"AF",X"FF",X"01",X"10",X"01",X"FF",X"01",X"08",X"CD",
		X"26",X"44",X"CD",X"30",X"44",X"C3",X"E4",X"42",X"D0",X"C0",X"9B",X"18",X"02",X"0F",X"30",X"AF",
		X"00",X"00",X"50",X"01",X"FF",X"00",X"10",X"CD",X"3A",X"44",X"01",X"FF",X"00",X"10",X"CD",X"44",
		X"44",X"01",X"FF",X"FF",X"10",X"AF",X"FF",X"00",X"10",X"01",X"FF",X"01",X"10",X"01",X"FF",X"FF",
		X"10",X"CD",X"4E",X"44",X"01",X"FF",X"FF",X"10",X"CD",X"58",X"44",X"C3",X"E4",X"42",X"A0",X"A0",
		X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"A0",X"AA",X"01",X"1C",X"02",X"05",X"66",X"C3",
		X"26",X"43",X"60",X"C0",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"60",X"CA",X"01",X"1C",
		X"02",X"05",X"66",X"C3",X"26",X"43",X"40",X"E0",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",
		X"40",X"EA",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"A0",X"C0",X"01",X"1C",X"02",X"05",
		X"66",X"C3",X"26",X"43",X"A0",X"CA",X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"50",X"A0",
		X"01",X"1C",X"02",X"05",X"66",X"C3",X"26",X"43",X"50",X"AA",X"01",X"1C",X"02",X"05",X"66",X"C3",
		X"26",X"43",X"D0",X"40",X"1B",X"18",X"02",X"0F",X"02",X"CD",X"AB",X"44",X"01",X"FE",X"00",X"12",
		X"01",X"FE",X"01",X"04",X"EB",X"6A",X"1F",X"02",X"0B",X"10",X"01",X"FE",X"01",X"04",X"01",X"FE",
		X"01",X"04",X"EB",X"7E",X"4E",X"02",X"07",X"20",X"01",X"FE",X"01",X"04",X"AF",X"00",X"04",X"01",
		X"EB",X"8E",X"4E",X"02",X"07",X"30",X"01",X"FE",X"02",X"03",X"01",X"FE",X"01",X"03",X"01",X"FE",
		X"00",X"08",X"01",X"FE",X"FF",X"08",X"01",X"FE",X"FE",X"30",X"76",X"D0",X"44",X"1B",X"18",X"02",
		X"0F",X"02",X"AF",X"00",X"00",X"20",X"CD",X"BC",X"44",X"C3",X"6C",X"44",X"D0",X"38",X"1B",X"18",
		X"02",X"0F",X"02",X"AF",X"00",X"00",X"20",X"C3",X"6C",X"44",X"D0",X"80",X"1B",X"18",X"02",X"0F",
		X"02",X"CD",X"D7",X"44",X"C3",X"6C",X"44",X"D0",X"84",X"1B",X"18",X"02",X"0F",X"02",X"AF",X"00",
		X"00",X"20",X"CD",X"E8",X"44",X"C3",X"6C",X"44",X"D0",X"78",X"1B",X"18",X"02",X"0F",X"02",X"AF",
		X"00",X"00",X"20",X"C3",X"6C",X"44",X"D0",X"C0",X"1B",X"18",X"02",X"0F",X"02",X"CD",X"03",X"45",
		X"C3",X"6C",X"44",X"D0",X"C4",X"1B",X"18",X"02",X"0F",X"02",X"AF",X"00",X"00",X"20",X"CD",X"14",
		X"45",X"C3",X"6C",X"44",X"D0",X"B8",X"1B",X"18",X"02",X"0F",X"02",X"AF",X"00",X"00",X"20",X"C3",
		X"6C",X"44",X"D0",X"30",X"9E",X"4E",X"02",X"05",X"20",X"CD",X"79",X"45",X"CD",X"87",X"45",X"CD",
		X"95",X"45",X"01",X"FF",X"01",X"10",X"EB",X"AA",X"4E",X"02",X"07",X"20",X"01",X"FF",X"01",X"08",
		X"EB",X"BA",X"4E",X"02",X"09",X"20",X"01",X"FE",X"01",X"08",X"EB",X"CE",X"4E",X"02",X"0B",X"20",
		X"01",X"FE",X"01",X"04",X"EB",X"E6",X"4E",X"02",X"0D",X"20",X"01",X"FE",X"01",X"02",X"EB",X"DB",
		X"17",X"02",X"0F",X"20",X"01",X"FE",X"00",X"08",X"AF",X"FE",X"FF",X"08",X"01",X"FD",X"FF",X"08",
		X"01",X"FE",X"01",X"10",X"01",X"FD",X"01",X"16",X"76",X"D0",X"50",X"9E",X"4E",X"02",X"05",X"20",
		X"01",X"00",X"00",X"08",X"C3",X"32",X"45",X"D0",X"70",X"9E",X"4E",X"02",X"05",X"20",X"01",X"00",
		X"00",X"10",X"C3",X"32",X"45",X"D0",X"90",X"9E",X"4E",X"02",X"05",X"20",X"01",X"00",X"00",X"18",
		X"C3",X"32",X"45",X"D0",X"30",X"9E",X"4E",X"02",X"05",X"20",X"CD",X"BA",X"45",X"CD",X"C8",X"45",
		X"CD",X"D6",X"45",X"AF",X"00",X"00",X"20",X"C3",X"32",X"45",X"D0",X"50",X"9E",X"4E",X"02",X"05",
		X"20",X"AF",X"00",X"00",X"28",X"C3",X"32",X"45",X"D0",X"70",X"9E",X"4E",X"02",X"05",X"20",X"AF",
		X"00",X"00",X"30",X"C3",X"32",X"45",X"D0",X"90",X"9E",X"4E",X"02",X"05",X"20",X"AF",X"00",X"00",
		X"38",X"C3",X"32",X"45",X"C0",X"BD",X"23",X"1B",X"02",X"28",X"40",X"01",X"FF",X"FF",X"41",X"CD",
		X"F7",X"45",X"01",X"00",X"00",X"FF",X"76",X"77",X"8C",X"75",X"1B",X"01",X"0B",X"40",X"CD",X"06",
		X"46",X"01",X"00",X"00",X"FF",X"76",X"23",X"90",X"82",X"1B",X"0B",X"01",X"40",X"CD",X"15",X"46",
		X"01",X"00",X"00",X"FF",X"76",X"23",X"92",X"82",X"1B",X"0B",X"01",X"40",X"01",X"00",X"00",X"FF",
		X"76",X"C0",X"F0",X"8F",X"19",X"05",X"28",X"70",X"01",X"FD",X"FD",X"40",X"76",X"80",X"B0",X"82",
		X"1F",X"02",X"11",X"38",X"01",X"00",X"00",X"01",X"CD",X"82",X"47",X"CD",X"8E",X"47",X"CD",X"98",
		X"47",X"CD",X"A4",X"47",X"CD",X"AE",X"47",X"AF",X"00",X"FE",X"04",X"CD",X"B8",X"47",X"01",X"00",
		X"FE",X"04",X"CD",X"C2",X"47",X"01",X"00",X"FE",X"04",X"CD",X"CC",X"47",X"AF",X"00",X"FE",X"04",
		X"CD",X"D6",X"47",X"01",X"00",X"FE",X"04",X"CD",X"E0",X"47",X"01",X"00",X"FE",X"04",X"CD",X"EA",
		X"47",X"AF",X"00",X"FF",X"08",X"CD",X"F4",X"47",X"01",X"00",X"FE",X"04",X"CD",X"FE",X"47",X"01",
		X"00",X"FE",X"04",X"CD",X"08",X"48",X"01",X"00",X"FF",X"08",X"CD",X"12",X"48",X"CD",X"1C",X"48",
		X"AF",X"00",X"FE",X"04",X"CD",X"26",X"48",X"01",X"00",X"FE",X"04",X"CD",X"30",X"48",X"01",X"00",
		X"FE",X"04",X"CD",X"3A",X"48",X"01",X"00",X"FE",X"04",X"CD",X"44",X"48",X"01",X"00",X"FE",X"04",
		X"CD",X"4E",X"48",X"01",X"00",X"FE",X"04",X"CD",X"58",X"48",X"01",X"00",X"FE",X"04",X"CD",X"62",
		X"48",X"01",X"00",X"02",X"04",X"CD",X"6C",X"48",X"AF",X"00",X"02",X"04",X"CD",X"76",X"48",X"01",
		X"00",X"02",X"04",X"CD",X"80",X"48",X"AF",X"00",X"02",X"04",X"CD",X"30",X"48",X"01",X"00",X"02",
		X"04",X"CD",X"8A",X"48",X"01",X"00",X"01",X"08",X"CD",X"94",X"48",X"AF",X"00",X"01",X"08",X"CD",
		X"1C",X"48",X"01",X"00",X"02",X"04",X"CD",X"9E",X"48",X"01",X"00",X"02",X"04",X"CD",X"F4",X"47",
		X"AF",X"00",X"02",X"04",X"CD",X"A8",X"48",X"01",X"00",X"02",X"04",X"CD",X"B2",X"48",X"01",X"00",
		X"02",X"04",X"CD",X"D6",X"47",X"01",X"00",X"02",X"04",X"CD",X"BC",X"48",X"01",X"00",X"02",X"04",
		X"CD",X"C6",X"48",X"AF",X"00",X"02",X"04",X"CD",X"D0",X"48",X"01",X"00",X"02",X"04",X"CD",X"8E",
		X"47",X"01",X"00",X"02",X"04",X"CD",X"DA",X"48",X"01",X"00",X"02",X"04",X"CD",X"AE",X"47",X"AF",
		X"00",X"02",X"04",X"CD",X"E4",X"48",X"01",X"00",X"02",X"04",X"CD",X"EE",X"48",X"01",X"00",X"02",
		X"04",X"CD",X"F8",X"48",X"01",X"00",X"01",X"08",X"CD",X"02",X"49",X"01",X"00",X"02",X"08",X"CD",
		X"0C",X"49",X"01",X"00",X"FE",X"08",X"CD",X"16",X"49",X"01",X"00",X"FE",X"04",X"CD",X"20",X"49",
		X"01",X"00",X"FE",X"04",X"CD",X"2A",X"49",X"AF",X"00",X"FE",X"0C",X"01",X"00",X"FE",X"04",X"C3",
		X"34",X"46",X"70",X"AC",X"66",X"1F",X"02",X"01",X"64",X"01",X"FC",X"00",X"18",X"76",X"70",X"B2",
		X"66",X"1F",X"02",X"01",X"64",X"C3",X"89",X"47",X"70",X"B6",X"01",X"1C",X"02",X"05",X"66",X"01",
		X"FD",X"00",X"20",X"76",X"70",X"BE",X"66",X"1F",X"02",X"01",X"64",X"C3",X"89",X"47",X"70",X"C4",
		X"66",X"1F",X"02",X"01",X"64",X"C3",X"89",X"47",X"70",X"AA",X"01",X"1C",X"02",X"05",X"66",X"C3",
		X"9F",X"47",X"70",X"A2",X"01",X"1C",X"02",X"05",X"66",X"C3",X"9F",X"47",X"70",X"9A",X"01",X"1C",
		X"02",X"05",X"66",X"C3",X"9F",X"47",X"70",X"94",X"66",X"1F",X"02",X"01",X"64",X"C3",X"89",X"47",
		X"70",X"8A",X"01",X"1C",X"02",X"05",X"66",X"C3",X"9F",X"47",X"70",X"82",X"01",X"1C",X"02",X"05",
		X"66",X"C3",X"9F",X"47",X"70",X"7C",X"66",X"1F",X"02",X"01",X"64",X"C3",X"89",X"47",X"70",X"72");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
