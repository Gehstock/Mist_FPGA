-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity PISCES_ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of PISCES_ROM_PGM_0 is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"AF",x"32",x"01",x"70",x"31",x"FF",x"43",x"C3", -- 0x0000
    x"72",x"02",x"F5",x"DD",x"E5",x"FD",x"E5",x"C5", -- 0x0008
    x"D5",x"E5",x"AF",x"32",x"01",x"70",x"3A",x"00", -- 0x0010
    x"78",x"21",x"6A",x"41",x"11",x"00",x"58",x"01", -- 0x0018
    x"80",x"00",x"ED",x"B0",x"2A",x"14",x"41",x"2B", -- 0x0020
    x"22",x"14",x"41",x"2A",x"32",x"41",x"2B",x"C2", -- 0x0028
    x"9B",x"00",x"3A",x"31",x"41",x"2F",x"21",x"FF", -- 0x0030
    x"FF",x"0F",x"CB",x"1C",x"0F",x"CB",x"1C",x"22", -- 0x0038
    x"32",x"41",x"CD",x"03",x"01",x"CD",x"58",x"01", -- 0x0040
    x"CD",x"C1",x"01",x"3A",x"00",x"40",x"FE",x"06", -- 0x0048
    x"D2",x"DB",x"00",x"3A",x"08",x"40",x"A7",x"CA", -- 0x0050
    x"DB",x"00",x"CD",x"00",x"00",x"CD",x"00",x"00", -- 0x0058
    x"AF",x"32",x"06",x"70",x"32",x"07",x"F5",x"DD", -- 0x0060
    x"E5",x"FD",x"E5",x"C5",x"D5",x"E5",x"AF",x"32", -- 0x0068
    x"01",x"70",x"3A",x"00",x"78",x"21",x"6A",x"41", -- 0x0070
    x"11",x"00",x"58",x"01",x"80",x"00",x"ED",x"B0", -- 0x0078
    x"2A",x"14",x"41",x"2B",x"22",x"14",x"41",x"2A", -- 0x0080
    x"32",x"41",x"2B",x"C2",x"9B",x"00",x"3A",x"31", -- 0x0088
    x"41",x"2F",x"21",x"FF",x"FF",x"0F",x"CB",x"1C", -- 0x0090
    x"0F",x"CB",x"1C",x"22",x"32",x"41",x"CD",x"03", -- 0x0098
    x"01",x"CD",x"58",x"01",x"CD",x"C1",x"01",x"3A", -- 0x00A0
    x"00",x"40",x"FE",x"06",x"D2",x"DB",x"00",x"3A", -- 0x00A8
    x"08",x"40",x"A7",x"CA",x"DB",x"00",x"CD",x"FC", -- 0x00B0
    x"26",x"CD",x"B1",x"26",x"AF",x"32",x"06",x"70", -- 0x00B8
    x"32",x"07",x"70",x"21",x"EF",x"52",x"11",x"5F", -- 0x00C0
    x"02",x"CD",x"E7",x"26",x"3E",x"04",x"32",x"A9", -- 0x00C8
    x"41",x"3E",x"01",x"32",x"8E",x"40",x"3E",x"06", -- 0x00D0
    x"32",x"00",x"40",x"21",x"F5",x"00",x"E5",x"21", -- 0x00D8
    x"85",x"28",x"ED",x"4B",x"06",x"41",x"09",x"5E", -- 0x00E0
    x"23",x"56",x"EB",x"ED",x"4B",x"00",x"40",x"09", -- 0x00E8
    x"5E",x"23",x"56",x"EB",x"E9",x"E1",x"D1",x"C1", -- 0x00F0
    x"FD",x"E1",x"DD",x"E1",x"3E",x"01",x"32",x"01", -- 0x00F8
    x"70",x"F1",x"C9",x"3A",x"00",x"68",x"4F",x"32", -- 0x0100
    x"04",x"40",x"3A",x"00",x"60",x"47",x"32",x"06", -- 0x0108
    x"40",x"3A",x"00",x"40",x"FE",x"04",x"C2",x"43", -- 0x0110
    x"01",x"3A",x"05",x"40",x"47",x"21",x"9B",x"40", -- 0x0118
    x"35",x"C2",x"39",x"01",x"CD",x"09",x"28",x"E6", -- 0x0120
    x"1F",x"3C",x"32",x"9B",x"40",x"CD",x"09",x"28", -- 0x0128
    x"E6",x"01",x"06",x"04",x"CA",x"39",x"01",x"06", -- 0x0130
    x"08",x"CD",x"09",x"28",x"E6",x"10",x"B0",x"32", -- 0x0138
    x"05",x"40",x"C9",x"3A",x"00",x"68",x"CB",x"7F", -- 0x0140
    x"CA",x"53",x"01",x"3A",x"00",x"40",x"FE",x"18", -- 0x0148
    x"79",x"28",x"01",x"78",x"32",x"05",x"40",x"C9", -- 0x0150
    x"21",x"07",x"40",x"D9",x"11",x"09",x"40",x"21", -- 0x0158
    x"06",x"40",x"CB",x"4E",x"EB",x"CA",x"6C",x"01", -- 0x0160
    x"34",x"C3",x"7D",x"01",x"7E",x"36",x"00",x"FE", -- 0x0168
    x"02",x"DA",x"7D",x"01",x"D9",x"3E",x"01",x"86", -- 0x0170
    x"77",x"D9",x"CD",x"B6",x"01",x"23",x"EB",x"CB", -- 0x0178
    x"46",x"EB",x"CA",x"89",x"01",x"34",x"C3",x"99", -- 0x0180
    x"01",x"7E",x"36",x"00",x"FE",x"02",x"DA",x"99", -- 0x0188
    x"01",x"D9",x"3E",x"06",x"86",x"77",x"CD",x"B6", -- 0x0190
    x"01",x"11",x"08",x"40",x"1A",x"FE",x"99",x"C8", -- 0x0198
    x"21",x"07",x"40",x"3A",x"0B",x"40",x"BE",x"D0", -- 0x01A0
    x"2F",x"86",x"77",x"EB",x"3E",x"01",x"86",x"27", -- 0x01A8
    x"D8",x"77",x"EB",x"C3",x"A3",x"01",x"D5",x"E5", -- 0x01B0
    x"11",x"03",x"2A",x"CD",x"1F",x"27",x"E1",x"D1", -- 0x01B8
    x"C9",x"21",x"02",x"40",x"35",x"C0",x"2A",x"0C", -- 0x01C0
    x"40",x"7C",x"B5",x"C8",x"3A",x"00",x"40",x"FE", -- 0x01C8
    x"04",x"CA",x"07",x"02",x"7E",x"E6",x"3F",x"3C", -- 0x01D0
    x"32",x"02",x"40",x"7E",x"07",x"32",x"06",x"68", -- 0x01D8
    x"07",x"32",x"07",x"68",x"23",x"7E",x"FE",x"FE", -- 0x01E0
    x"CA",x"07",x"02",x"FE",x"FD",x"CA",x"17",x"02", -- 0x01E8
    x"FE",x"FC",x"CA",x"26",x"02",x"FE",x"FB",x"CA", -- 0x01F0
    x"3B",x"02",x"FE",x"FA",x"CA",x"4A",x"02",x"32", -- 0x01F8
    x"00",x"78",x"23",x"22",x"0C",x"40",x"C9",x"CD", -- 0x0200
    x"12",x"27",x"2A",x"0E",x"40",x"22",x"0C",x"40", -- 0x0208
    x"21",x"00",x"00",x"22",x"0E",x"40",x"C9",x"23", -- 0x0210
    x"7E",x"32",x"1B",x"40",x"23",x"7E",x"32",x"1C", -- 0x0218
    x"40",x"23",x"22",x"0C",x"40",x"C9",x"23",x"3A", -- 0x0220
    x"1B",x"40",x"86",x"32",x"00",x"78",x"32",x"1B", -- 0x0228
    x"40",x"23",x"BE",x"C2",x"50",x"02",x"23",x"22", -- 0x0230
    x"0C",x"40",x"C9",x"23",x"7E",x"32",x"1C",x"40", -- 0x0238
    x"23",x"7E",x"32",x"1B",x"40",x"23",x"22",x"0C", -- 0x0240
    x"40",x"C9",x"3A",x"1B",x"40",x"32",x"00",x"78", -- 0x0248
    x"3A",x"1B",x"40",x"47",x"3A",x"1C",x"40",x"32", -- 0x0250
    x"1B",x"40",x"78",x"32",x"1C",x"40",x"C9",x"50", -- 0x0258
    x"55",x"53",x"48",x"20",x"53",x"54",x"41",x"52", -- 0x0260
    x"54",x"20",x"42",x"55",x"54",x"54",x"4F",x"4E", -- 0x0268
    x"FF",x"25",x"21",x"00",x"40",x"55",x"72",x"23", -- 0x0270
    x"7C",x"FE",x"44",x"20",x"F9",x"21",x"00",x"50", -- 0x0278
    x"06",x"04",x"0E",x"10",x"71",x"2C",x"20",x"FC", -- 0x0280
    x"24",x"3A",x"00",x"78",x"10",x"F6",x"CD",x"B1", -- 0x0288
    x"26",x"21",x"00",x"60",x"06",x"04",x"AF",x"77", -- 0x0290
    x"23",x"10",x"FC",x"3C",x"06",x"04",x"77",x"23", -- 0x0298
    x"10",x"FC",x"3E",x"03",x"32",x"6D",x"41",x"3D", -- 0x02A0
    x"32",x"A9",x"41",x"32",x"79",x"41",x"32",x"9D", -- 0x02A8
    x"41",x"07",x"32",x"9B",x"41",x"3E",x"07",x"32", -- 0x02B0
    x"A3",x"41",x"32",x"A5",x"41",x"32",x"6B",x"41", -- 0x02B8
    x"3E",x"04",x"32",x"A7",x"41",x"32",x"A9",x"41", -- 0x02C0
    x"AF",x"06",x"08",x"21",x"00",x"68",x"77",x"23", -- 0x02C8
    x"10",x"FC",x"32",x"06",x"70",x"32",x"07",x"70", -- 0x02D0
    x"3D",x"32",x"00",x"78",x"3A",x"00",x"68",x"CB", -- 0x02D8
    x"77",x"3E",x"03",x"CA",x"E8",x"02",x"3E",x"04", -- 0x02E0
    x"32",x"69",x"40",x"3A",x"00",x"68",x"CB",x"7F", -- 0x02E8
    x"3E",x"01",x"C2",x"F6",x"02",x"AF",x"32",x"8F", -- 0x02F0
    x"40",x"3A",x"00",x"70",x"CB",x"47",x"3E",x"10", -- 0x02F8
    x"CA",x"05",x"03",x"3E",x"20",x"32",x"68",x"40", -- 0x0300
    x"3A",x"00",x"70",x"CB",x"4F",x"3E",x"00",x"CA", -- 0x0308
    x"14",x"03",x"3E",x"01",x"32",x"0B",x"40",x"3A", -- 0x0310
    x"00",x"78",x"11",x"EB",x"03",x"21",x"40",x"53", -- 0x0318
    x"CD",x"E7",x"26",x"11",x"F5",x"03",x"21",x"80", -- 0x0320
    x"52",x"CD",x"E7",x"26",x"11",x"F0",x"03",x"21", -- 0x0328
    x"00",x"51",x"CD",x"E7",x"26",x"AF",x"32",x"01", -- 0x0330
    x"53",x"32",x"41",x"50",x"32",x"61",x"50",x"32", -- 0x0338
    x"A1",x"51",x"32",x"C1",x"51",x"3E",x"01",x"32", -- 0x0340
    x"04",x"70",x"32",x"01",x"70",x"DD",x"21",x"A1", -- 0x0348
    x"53",x"21",x"02",x"41",x"01",x"E0",x"FF",x"CD", -- 0x0350
    x"BA",x"03",x"DD",x"21",x"E1",x"50",x"21",x"05", -- 0x0358
    x"41",x"CD",x"BA",x"03",x"DD",x"21",x"41",x"52", -- 0x0360
    x"21",x"23",x"40",x"CD",x"BA",x"03",x"21",x"5F", -- 0x0368
    x"51",x"3A",x"8E",x"40",x"A7",x"C2",x"8B",x"03", -- 0x0370
    x"11",x"E0",x"FF",x"06",x"09",x"7E",x"FE",x"2C", -- 0x0378
    x"D2",x"85",x"03",x"36",x"10",x"19",x"10",x"F5", -- 0x0380
    x"C3",x"AB",x"03",x"11",x"00",x"04",x"CD",x"E7", -- 0x0388
    x"26",x"21",x"08",x"40",x"7E",x"0F",x"0F",x"0F", -- 0x0390
    x"0F",x"E6",x"0F",x"C2",x"A0",x"03",x"3E",x"10", -- 0x0398
    x"11",x"7F",x"50",x"12",x"7E",x"E6",x"0F",x"11", -- 0x03A0
    x"5F",x"50",x"12",x"21",x"67",x"40",x"ED",x"5F", -- 0x03A8
    x"E6",x"0F",x"86",x"77",x"CD",x"09",x"28",x"C3", -- 0x03B0
    x"4D",x"03",x"11",x"10",x"00",x"7E",x"CD",x"DE", -- 0x03B8
    x"03",x"2B",x"7E",x"0F",x"0F",x"0F",x"0F",x"CD", -- 0x03C0
    x"DE",x"03",x"7E",x"CD",x"DE",x"03",x"2B",x"7E", -- 0x03C8
    x"0F",x"0F",x"0F",x"0F",x"CD",x"DE",x"03",x"7E", -- 0x03D0
    x"E6",x"0F",x"DD",x"77",x"00",x"C9",x"E6",x"0F", -- 0x03D8
    x"CA",x"E4",x"03",x"5A",x"B3",x"DD",x"77",x"00", -- 0x03E0
    x"DD",x"09",x"C9",x"31",x"20",x"55",x"50",x"FF", -- 0x03E8
    x"32",x"20",x"55",x"50",x"FF",x"48",x"49",x"47", -- 0x03F0
    x"48",x"40",x"53",x"43",x"4F",x"52",x"45",x"FF", -- 0x03F8
    x"43",x"52",x"45",x"44",x"49",x"54",x"40",x"FF", -- 0x0400
    x"3A",x"08",x"41",x"FE",x"08",x"CA",x"1F",x"05", -- 0x0408
    x"FE",x"0C",x"CA",x"A8",x"04",x"FE",x"0A",x"CA", -- 0x0410
    x"CC",x"04",x"FE",x"10",x"CA",x"0F",x"05",x"FE", -- 0x0418
    x"06",x"CA",x"25",x"04",x"C9",x"3A",x"05",x"40", -- 0x0420
    x"E6",x"0C",x"CA",x"50",x"04",x"FE",x"0C",x"CA", -- 0x0428
    x"50",x"04",x"CB",x"57",x"21",x"A2",x"41",x"7E", -- 0x0430
    x"C2",x"47",x"04",x"FE",x"68",x"CA",x"50",x"04", -- 0x0438
    x"34",x"23",x"23",x"34",x"C3",x"50",x"04",x"FE", -- 0x0440
    x"96",x"CA",x"50",x"04",x"35",x"23",x"23",x"35", -- 0x0448
    x"3A",x"65",x"40",x"3C",x"E6",x"03",x"32",x"65", -- 0x0450
    x"40",x"CA",x"25",x"04",x"DD",x"21",x"EA",x"41", -- 0x0458
    x"FD",x"21",x"AA",x"41",x"3A",x"29",x"41",x"47", -- 0x0460
    x"DD",x"7E",x"00",x"FE",x"0E",x"D2",x"7D",x"04", -- 0x0468
    x"11",x"24",x"00",x"DD",x"19",x"11",x"04",x"00", -- 0x0470
    x"FD",x"19",x"10",x"EC",x"C9",x"FD",x"7E",x"03", -- 0x0478
    x"D6",x"D9",x"FE",x"13",x"D2",x"70",x"04",x"3A", -- 0x0480
    x"A2",x"41",x"4F",x"FD",x"7E",x"00",x"DD",x"86", -- 0x0488
    x"1A",x"C6",x"7F",x"91",x"D2",x"99",x"04",x"ED", -- 0x0490
    x"44",x"DD",x"BE",x"1D",x"D2",x"70",x"04",x"CD", -- 0x0498
    x"40",x"07",x"3E",x"0C",x"32",x"08",x"41",x"C9", -- 0x04A0
    x"3E",x"07",x"32",x"A7",x"41",x"32",x"A9",x"41", -- 0x04A8
    x"3A",x"00",x"40",x"FE",x"04",x"CA",x"BD",x"04", -- 0x04B0
    x"3E",x"01",x"32",x"03",x"68",x"21",x"3C",x"52", -- 0x04B8
    x"36",x"B8",x"3E",x"0A",x"32",x"08",x"41",x"21", -- 0x04C0
    x"03",x"40",x"36",x"01",x"21",x"03",x"40",x"35", -- 0x04C8
    x"C0",x"36",x"0A",x"21",x"3C",x"52",x"7E",x"C6", -- 0x04D0
    x"08",x"FE",x"E0",x"CA",x"EC",x"04",x"FE",x"D0", -- 0x04D8
    x"C2",x"E8",x"04",x"21",x"03",x"68",x"36",x"00", -- 0x04E0
    x"CD",x"FD",x"06",x"C9",x"3E",x"04",x"32",x"A7", -- 0x04E8
    x"41",x"32",x"A9",x"41",x"21",x"3C",x"52",x"11", -- 0x04F0
    x"DF",x"FF",x"3E",x"10",x"06",x"04",x"77",x"23", -- 0x04F8
    x"77",x"19",x"10",x"FA",x"3E",x"80",x"32",x"0A", -- 0x0500
    x"41",x"3E",x"10",x"32",x"08",x"41",x"C9",x"21", -- 0x0508
    x"0A",x"41",x"35",x"C0",x"3E",x"80",x"32",x"0A", -- 0x0510
    x"41",x"3E",x"0E",x"32",x"08",x"41",x"C9",x"21", -- 0x0518
    x"0A",x"41",x"35",x"C0",x"36",x"80",x"3E",x"FF", -- 0x0520
    x"32",x"A2",x"41",x"32",x"A4",x"41",x"3E",x"07", -- 0x0528
    x"32",x"A3",x"41",x"32",x"A5",x"41",x"3E",x"60", -- 0x0530
    x"32",x"FC",x"51",x"3C",x"32",x"FD",x"51",x"3C", -- 0x0538
    x"32",x"1C",x"52",x"3C",x"32",x"1D",x"52",x"3E", -- 0x0540
    x"06",x"32",x"08",x"41",x"C9",x"3A",x"0D",x"41", -- 0x0548
    x"21",x"13",x"41",x"BE",x"D2",x"DC",x"05",x"3A", -- 0x0550
    x"08",x"41",x"FE",x"06",x"C2",x"DC",x"05",x"3A", -- 0x0558
    x"05",x"40",x"CB",x"67",x"C2",x"6E",x"05",x"AF", -- 0x0560
    x"32",x"7B",x"40",x"C3",x"DC",x"05",x"3A",x"7B", -- 0x0568
    x"40",x"A7",x"C2",x"DC",x"05",x"3A",x"00",x"40", -- 0x0570
    x"FE",x"04",x"3E",x"01",x"CA",x"82",x"05",x"32", -- 0x0578
    x"05",x"68",x"32",x"7B",x"40",x"21",x"0D",x"41", -- 0x0580
    x"34",x"21",x"C7",x"41",x"11",x"04",x"00",x"3A", -- 0x0588
    x"A2",x"41",x"C6",x"7F",x"06",x"07",x"0E",x"07", -- 0x0590
    x"19",x"BE",x"C2",x"9F",x"05",x"CB",x"89",x"3C", -- 0x0598
    x"BE",x"C2",x"A6",x"05",x"CB",x"81",x"3C",x"BE", -- 0x05A0
    x"C2",x"AD",x"05",x"CB",x"91",x"D6",x"02",x"10", -- 0x05A8
    x"E7",x"3C",x"CB",x"41",x"C2",x"C5",x"05",x"3D", -- 0x05B0
    x"CB",x"49",x"C2",x"C5",x"05",x"C6",x"02",x"CB", -- 0x05B8
    x"51",x"C2",x"C5",x"05",x"3D",x"47",x"21",x"EA", -- 0x05C0
    x"41",x"11",x"FC",x"FF",x"AF",x"19",x"BE",x"C2", -- 0x05C8
    x"CD",x"05",x"36",x"FF",x"23",x"70",x"23",x"23", -- 0x05D0
    x"3A",x"20",x"41",x"77",x"DD",x"21",x"E6",x"41", -- 0x05D8
    x"3E",x"03",x"08",x"DD",x"22",x"6C",x"40",x"DD", -- 0x05E0
    x"CB",x"00",x"7E",x"CA",x"EE",x"06",x"DD",x"7E", -- 0x05E8
    x"03",x"21",x"1B",x"41",x"AE",x"C6",x"06",x"AE", -- 0x05F0
    x"DD",x"77",x"03",x"AE",x"FE",x"08",x"DA",x"C3", -- 0x05F8
    x"06",x"DD",x"35",x"00",x"DD",x"7E",x"00",x"FE", -- 0x0600
    x"FC",x"C2",x"11",x"06",x"21",x"05",x"68",x"36", -- 0x0608
    x"00",x"FE",x"DD",x"CA",x"C3",x"06",x"DD",x"56", -- 0x0610
    x"01",x"3A",x"1B",x"41",x"DD",x"AE",x"03",x"5F", -- 0x0618
    x"DD",x"21",x"EA",x"41",x"FD",x"21",x"AA",x"41", -- 0x0620
    x"3A",x"29",x"41",x"47",x"DD",x"7E",x"00",x"FE", -- 0x0628
    x"0E",x"DA",x"DE",x"06",x"7B",x"FD",x"86",x"03", -- 0x0630
    x"C6",x"14",x"FE",x"0F",x"D2",x"DE",x"06",x"FD", -- 0x0638
    x"7E",x"00",x"DD",x"86",x"1A",x"92",x"D2",x"4B", -- 0x0640
    x"06",x"ED",x"44",x"DD",x"BE",x"1B",x"D2",x"DE", -- 0x0648
    x"06",x"DD",x"BE",x"1C",x"DA",x"C0",x"06",x"3E", -- 0x0650
    x"02",x"CD",x"2B",x"28",x"4A",x"11",x"0D",x"2A", -- 0x0658
    x"CD",x"1F",x"27",x"CD",x"4A",x"28",x"DD",x"7E", -- 0x0660
    x"00",x"FE",x"18",x"CA",x"C3",x"06",x"CD",x"09", -- 0x0668
    x"28",x"E6",x"0F",x"C6",x"08",x"DD",x"77",x"21", -- 0x0670
    x"FD",x"7E",x"00",x"DD",x"86",x"1A",x"91",x"DA", -- 0x0678
    x"A0",x"06",x"DD",x"36",x"1F",x"80",x"FD",x"36", -- 0x0680
    x"01",x"94",x"DD",x"6E",x"18",x"DD",x"66",x"19", -- 0x0688
    x"23",x"3E",x"14",x"BE",x"CA",x"C3",x"06",x"36", -- 0x0690
    x"93",x"DD",x"36",x"00",x"1C",x"C3",x"C3",x"06", -- 0x0698
    x"DD",x"36",x"20",x"80",x"3E",x"94",x"FD",x"BE", -- 0x06A0
    x"01",x"CA",x"B0",x"06",x"FD",x"36",x"01",x"13", -- 0x06A8
    x"DD",x"6E",x"18",x"DD",x"66",x"19",x"23",x"36", -- 0x06B0
    x"14",x"DD",x"36",x"00",x"1C",x"C3",x"C3",x"06", -- 0x06B8
    x"CD",x"0E",x"07",x"AF",x"32",x"05",x"68",x"DD", -- 0x06C0
    x"2A",x"6C",x"40",x"DD",x"36",x"00",x"00",x"DD", -- 0x06C8
    x"36",x"01",x"00",x"DD",x"36",x"03",x"00",x"21", -- 0x06D0
    x"0D",x"41",x"35",x"C3",x"EE",x"06",x"D5",x"11", -- 0x06D8
    x"24",x"00",x"DD",x"19",x"11",x"04",x"00",x"FD", -- 0x06E0
    x"19",x"D1",x"05",x"C2",x"2C",x"06",x"DD",x"2A", -- 0x06E8
    x"6C",x"40",x"11",x"FC",x"FF",x"DD",x"19",x"08", -- 0x06F0
    x"3D",x"C2",x"E2",x"05",x"C9",x"11",x"DF",x"FF", -- 0x06F8
    x"21",x"3C",x"52",x"06",x"04",x"77",x"23",x"3C", -- 0x0700
    x"77",x"3C",x"19",x"10",x"F8",x"C9",x"DD",x"7E", -- 0x0708
    x"00",x"FE",x"14",x"C2",x"40",x"07",x"DD",x"36", -- 0x0710
    x"00",x"20",x"FD",x"36",x"02",x"05",x"DD",x"7E", -- 0x0718
    x"0D",x"CD",x"2B",x"28",x"3A",x"0B",x"41",x"FE", -- 0x0720
    x"03",x"3E",x"80",x"DA",x"3A",x"07",x"3A",x"67", -- 0x0728
    x"40",x"E6",x"30",x"C2",x"38",x"07",x"3E",x"10", -- 0x0730
    x"F6",x"80",x"DD",x"77",x"0D",x"C3",x"68",x"07", -- 0x0738
    x"FD",x"36",x"01",x"1C",x"DD",x"36",x"0A",x"07", -- 0x0740
    x"FD",x"36",x"02",x"07",x"DD",x"7E",x"00",x"DD", -- 0x0748
    x"36",x"00",x"0C",x"FE",x"12",x"DA",x"6B",x"07", -- 0x0750
    x"FE",x"16",x"DA",x"68",x"07",x"CA",x"6B",x"07", -- 0x0758
    x"FE",x"1E",x"DC",x"C2",x"0B",x"C3",x"6B",x"07", -- 0x0760
    x"CD",x"24",x"0D",x"11",x"EF",x"29",x"CD",x"1F", -- 0x0768
    x"27",x"CD",x"4A",x"28",x"C9",x"B1",x"07",x"B1", -- 0x0770
    x"07",x"B1",x"07",x"B9",x"07",x"44",x"09",x"C6", -- 0x0778
    x"07",x"FA",x"08",x"B1",x"07",x"B1",x"07",x"B4", -- 0x0780
    x"09",x"B4",x"09",x"9C",x"09",x"9C",x"09",x"9C", -- 0x0788
    x"09",x"43",x"08",x"DC",x"08",x"8C",x"09",x"DD", -- 0x0790
    x"21",x"EA",x"41",x"FD",x"21",x"AA",x"41",x"3A", -- 0x0798
    x"29",x"41",x"47",x"21",x"75",x"07",x"DD",x"5E", -- 0x07A0
    x"00",x"16",x"00",x"19",x"5E",x"23",x"56",x"EB", -- 0x07A8
    x"E9",x"DD",x"22",x"72",x"40",x"FD",x"22",x"74", -- 0x07B0
    x"40",x"11",x"24",x"00",x"DD",x"19",x"11",x"04", -- 0x07B8
    x"00",x"FD",x"19",x"10",x"DE",x"C9",x"DD",x"35", -- 0x07C0
    x"11",x"C2",x"B9",x"07",x"FD",x"7E",x"02",x"FE", -- 0x07C8
    x"07",x"3E",x"12",x"CA",x"D8",x"07",x"3E",x"14", -- 0x07D0
    x"DD",x"77",x"00",x"FD",x"36",x"01",x"12",x"FD", -- 0x07D8
    x"36",x"00",x"00",x"DD",x"6E",x"0F",x"DD",x"66", -- 0x07E0
    x"10",x"11",x"06",x"00",x"19",x"7E",x"FD",x"77", -- 0x07E8
    x"03",x"23",x"7E",x"DD",x"77",x"0C",x"DD",x"36", -- 0x07F0
    x"12",x"01",x"21",x"99",x"29",x"22",x"0C",x"40", -- 0x07F8
    x"21",x"00",x"00",x"22",x"0E",x"40",x"3E",x"01", -- 0x0800
    x"32",x"02",x"40",x"DD",x"7E",x"0E",x"E6",x"03", -- 0x0808
    x"C2",x"EB",x"0B",x"C5",x"DD",x"7E",x"0F",x"21", -- 0x0810
    x"D5",x"41",x"11",x"A9",x"41",x"01",x"24",x"00", -- 0x0818
    x"09",x"EB",x"01",x"04",x"00",x"09",x"EB",x"BE", -- 0x0820
    x"C2",x"1D",x"08",x"1A",x"FD",x"77",x"03",x"01", -- 0x0828
    x"F2",x"FF",x"09",x"DD",x"E5",x"D1",x"13",x"06", -- 0x0830
    x"0B",x"7E",x"12",x"23",x"13",x"10",x"FA",x"C1", -- 0x0838
    x"C3",x"B9",x"07",x"DD",x"7E",x"1F",x"A7",x"CA", -- 0x0840
    x"70",x"08",x"DD",x"35",x"1F",x"C2",x"69",x"08", -- 0x0848
    x"DD",x"36",x"21",x"00",x"21",x"30",x"41",x"3A", -- 0x0850
    x"0B",x"41",x"BE",x"DA",x"B6",x"08",x"FD",x"36", -- 0x0858
    x"01",x"13",x"DD",x"7E",x"20",x"A7",x"CA",x"94", -- 0x0860
    x"08",x"DD",x"7E",x"20",x"A7",x"CA",x"9F",x"08", -- 0x0868
    x"DD",x"35",x"20",x"C2",x"9F",x"08",x"DD",x"36", -- 0x0870
    x"21",x"00",x"21",x"30",x"41",x"3A",x"0B",x"41", -- 0x0878
    x"BE",x"DA",x"B6",x"08",x"DD",x"6E",x"18",x"DD", -- 0x0880
    x"66",x"19",x"23",x"36",x"93",x"DD",x"7E",x"1F", -- 0x0888
    x"A7",x"C2",x"9F",x"08",x"DD",x"36",x"00",x"1A", -- 0x0890
    x"DD",x"36",x"21",x"00",x"C3",x"B9",x"07",x"3A", -- 0x0898
    x"0B",x"41",x"21",x"30",x"41",x"BE",x"D2",x"D0", -- 0x08A0
    x"08",x"DD",x"7E",x"21",x"A7",x"CA",x"B6",x"08", -- 0x08A8
    x"DD",x"35",x"21",x"C2",x"D0",x"08",x"FD",x"7E", -- 0x08B0
    x"03",x"C6",x"06",x"FE",x"08",x"DA",x"91",x"0B", -- 0x08B8
    x"FD",x"77",x"03",x"DD",x"6E",x"18",x"DD",x"66", -- 0x08C0
    x"19",x"23",x"23",x"23",x"77",x"C3",x"B9",x"07", -- 0x08C8
    x"ED",x"5F",x"E6",x"02",x"3D",x"DD",x"36",x"12", -- 0x08D0
    x"01",x"C3",x"12",x"0A",x"DD",x"35",x"0A",x"C2", -- 0x08D8
    x"B9",x"07",x"DD",x"36",x"0A",x"06",x"FD",x"7E", -- 0x08E0
    x"02",x"EE",x"01",x"FD",x"77",x"02",x"DD",x"35", -- 0x08E8
    x"0C",x"C2",x"B9",x"07",x"CD",x"40",x"07",x"C3", -- 0x08F0
    x"B9",x"07",x"DD",x"35",x"0A",x"C2",x"B9",x"07", -- 0x08F8
    x"DD",x"36",x"0A",x"07",x"FD",x"34",x"01",x"FD", -- 0x0900
    x"7E",x"01",x"FE",x"20",x"C2",x"B9",x"07",x"DD", -- 0x0908
    x"7E",x"0D",x"E6",x"7F",x"C2",x"19",x"09",x"F6", -- 0x0910
    x"80",x"CD",x"2B",x"28",x"CD",x"4A",x"28",x"DD", -- 0x0918
    x"CB",x"0D",x"7E",x"CA",x"4A",x"09",x"DD",x"7E", -- 0x0920
    x"0D",x"0F",x"0F",x"0F",x"0F",x"E6",x"03",x"0E", -- 0x0928
    x"20",x"81",x"FD",x"77",x"01",x"FD",x"36",x"02", -- 0x0930
    x"05",x"DD",x"36",x"0A",x"20",x"DD",x"36",x"00", -- 0x0938
    x"08",x"C3",x"B9",x"07",x"DD",x"35",x"0A",x"C2", -- 0x0940
    x"B9",x"07",x"FD",x"36",x"01",x"00",x"FD",x"36", -- 0x0948
    x"00",x"00",x"FD",x"36",x"03",x"00",x"DD",x"36", -- 0x0950
    x"00",x"00",x"21",x"0C",x"41",x"35",x"2B",x"35", -- 0x0958
    x"20",x"0D",x"3A",x"00",x"40",x"FE",x"04",x"C2", -- 0x0960
    x"B9",x"07",x"36",x"08",x"C3",x"B9",x"07",x"7E", -- 0x0968
    x"21",x"30",x"41",x"BE",x"D2",x"B9",x"07",x"3A", -- 0x0970
    x"06",x"41",x"FE",x"04",x"C2",x"B9",x"07",x"CD", -- 0x0978
    x"09",x"28",x"E6",x"0F",x"C6",x"08",x"DD",x"77", -- 0x0980
    x"21",x"C3",x"B9",x"07",x"FD",x"7E",x"03",x"C6", -- 0x0988
    x"06",x"FD",x"77",x"03",x"FE",x"08",x"DA",x"80", -- 0x0990
    x"0B",x"C3",x"B9",x"07",x"FD",x"7E",x"00",x"CB", -- 0x0998
    x"7F",x"CA",x"A5",x"09",x"2F",x"07",x"07",x"07", -- 0x09A0
    x"E6",x"03",x"C2",x"AE",x"09",x"3C",x"DD",x"77", -- 0x09A8
    x"12",x"C3",x"C6",x"09",x"DD",x"35",x"23",x"C2", -- 0x09B0
    x"C6",x"09",x"DD",x"36",x"23",x"07",x"FD",x"7E", -- 0x09B8
    x"01",x"EE",x"06",x"FD",x"77",x"01",x"AF",x"57", -- 0x09C0
    x"5F",x"DD",x"BE",x"05",x"CA",x"D3",x"09",x"DD", -- 0x09C8
    x"35",x"05",x"1D",x"DD",x"BE",x"06",x"CA",x"DD", -- 0x09D0
    x"09",x"DD",x"35",x"06",x"15",x"B2",x"B3",x"C2", -- 0x09D8
    x"F1",x"09",x"DD",x"7E",x"03",x"DD",x"77",x"05", -- 0x09E0
    x"DD",x"7E",x"04",x"DD",x"77",x"06",x"C3",x"C6", -- 0x09E8
    x"09",x"DD",x"7E",x"09",x"07",x"E6",x"02",x"3D", -- 0x09F0
    x"A3",x"FD",x"86",x"00",x"DD",x"BE",x"14",x"CA", -- 0x09F8
    x"62",x"0B",x"DD",x"BE",x"15",x"CA",x"62",x"0B", -- 0x0A00
    x"FD",x"77",x"00",x"DD",x"7E",x"09",x"E6",x"02", -- 0x0A08
    x"3D",x"A2",x"FD",x"86",x"03",x"CA",x"91",x"0B", -- 0x0A10
    x"FE",x"10",x"D2",x"30",x"0A",x"DD",x"7E",x"0C", -- 0x0A18
    x"EE",x"AA",x"DD",x"77",x"0C",x"DD",x"7E",x"09", -- 0x0A20
    x"EE",x"AA",x"DD",x"77",x"09",x"C3",x"6B",x"0A", -- 0x0A28
    x"FD",x"77",x"03",x"FE",x"E0",x"C2",x"6B",x"0A", -- 0x0A30
    x"DD",x"7E",x"00",x"FE",x"14",x"C2",x"6B",x"0A", -- 0x0A38
    x"FD",x"7E",x"00",x"FE",x"40",x"DA",x"6B",x"0A", -- 0x0A40
    x"FE",x"C0",x"D2",x"6B",x"0A",x"21",x"66",x"40", -- 0x0A48
    x"BE",x"CA",x"6B",x"0A",x"77",x"ED",x"5F",x"E6", -- 0x0A50
    x"FE",x"3C",x"DD",x"77",x"0C",x"DD",x"36",x"0A", -- 0x0A58
    x"06",x"DD",x"36",x"00",x"1E",x"CD",x"24",x"0D", -- 0x0A60
    x"C3",x"B9",x"07",x"DD",x"7E",x"00",x"FE",x"18", -- 0x0A68
    x"DA",x"86",x"0A",x"DD",x"6E",x"18",x"DD",x"66", -- 0x0A70
    x"19",x"FD",x"7E",x"00",x"C6",x"0F",x"77",x"23", -- 0x0A78
    x"23",x"23",x"FD",x"7E",x"03",x"77",x"DD",x"35", -- 0x0A80
    x"12",x"C2",x"C6",x"09",x"21",x"30",x"41",x"3A", -- 0x0A88
    x"0B",x"41",x"BE",x"3E",x"01",x"D2",x"99",x"0A", -- 0x0A90
    x"3C",x"DD",x"77",x"12",x"DD",x"35",x"0B",x"C2", -- 0x0A98
    x"8C",x"0C",x"DD",x"7E",x"00",x"FE",x"16",x"DA", -- 0x0AA0
    x"B3",x"0A",x"ED",x"5F",x"E6",x"1F",x"C6",x"08", -- 0x0AA8
    x"C3",x"BB",x"0A",x"DD",x"6E",x"0F",x"DD",x"66", -- 0x0AB0
    x"10",x"23",x"7E",x"DD",x"77",x"0B",x"DD",x"6E", -- 0x0AB8
    x"01",x"DD",x"66",x"02",x"23",x"DD",x"75",x"01", -- 0x0AC0
    x"DD",x"74",x"02",x"7E",x"A7",x"CA",x"DA",x"0B", -- 0x0AC8
    x"0F",x"0F",x"0F",x"0F",x"E6",x"0F",x"DD",x"77", -- 0x0AD0
    x"03",x"DD",x"77",x"05",x"7E",x"E6",x"0F",x"DD", -- 0x0AD8
    x"77",x"04",x"DD",x"77",x"06",x"DD",x"CB",x"09", -- 0x0AE0
    x"0E",x"DD",x"CB",x"09",x"0E",x"DD",x"35",x"0A", -- 0x0AE8
    x"C2",x"0B",x"0B",x"DD",x"36",x"0A",x"04",x"DD", -- 0x0AF0
    x"6E",x"07",x"DD",x"66",x"08",x"23",x"DD",x"75", -- 0x0AF8
    x"07",x"DD",x"74",x"08",x"7E",x"DD",x"AE",x"0C", -- 0x0B00
    x"DD",x"77",x"09",x"CD",x"11",x"0B",x"C3",x"B9", -- 0x0B08
    x"07",x"DD",x"7E",x"00",x"FE",x"1A",x"C0",x"DD", -- 0x0B10
    x"7E",x"03",x"A7",x"CA",x"54",x"0B",x"DD",x"96", -- 0x0B18
    x"04",x"D2",x"26",x"0B",x"ED",x"44",x"DD",x"BE", -- 0x0B20
    x"03",x"CA",x"54",x"0B",x"FE",x"03",x"DA",x"54", -- 0x0B28
    x"0B",x"DD",x"CB",x"09",x"46",x"C2",x"46",x"0B", -- 0x0B30
    x"FD",x"36",x"01",x"96",x"DD",x"6E",x"18",x"DD", -- 0x0B38
    x"66",x"19",x"23",x"36",x"95",x"C9",x"FD",x"36", -- 0x0B40
    x"01",x"15",x"DD",x"6E",x"18",x"DD",x"66",x"19", -- 0x0B48
    x"23",x"36",x"16",x"C9",x"FD",x"36",x"01",x"13", -- 0x0B50
    x"DD",x"6E",x"18",x"DD",x"66",x"19",x"23",x"36", -- 0x0B58
    x"93",x"C9",x"DD",x"7E",x"00",x"FE",x"16",x"DA", -- 0x0B60
    x"91",x"0B",x"3E",x"55",x"DD",x"AE",x"0C",x"DD", -- 0x0B68
    x"77",x"0C",x"3E",x"55",x"DD",x"AE",x"09",x"DD", -- 0x0B70
    x"77",x"09",x"CD",x"11",x"0B",x"C3",x"6B",x"0A", -- 0x0B78
    x"21",x"0B",x"41",x"35",x"C2",x"91",x"0B",x"3A", -- 0x0B80
    x"00",x"40",x"FE",x"04",x"C2",x"91",x"0B",x"36", -- 0x0B88
    x"10",x"FD",x"36",x"01",x"00",x"FD",x"36",x"00", -- 0x0B90
    x"00",x"FD",x"36",x"03",x"00",x"FD",x"36",x"02", -- 0x0B98
    x"00",x"DD",x"7E",x"00",x"FE",x"16",x"DA",x"B4", -- 0x0BA0
    x"0B",x"CA",x"B7",x"0B",x"FE",x"1E",x"DC",x"C2", -- 0x0BA8
    x"0B",x"C3",x"B7",x"0B",x"CD",x"24",x"0D",x"DD", -- 0x0BB0
    x"36",x"00",x"00",x"21",x"0C",x"41",x"35",x"C3", -- 0x0BB8
    x"B9",x"07",x"DD",x"6E",x"16",x"DD",x"66",x"17", -- 0x0BC0
    x"36",x"00",x"DD",x"6E",x"18",x"DD",x"66",x"19", -- 0x0BC8
    x"0E",x"04",x"36",x"00",x"23",x"0D",x"C2",x"D2", -- 0x0BD0
    x"0B",x"C9",x"DD",x"7E",x"00",x"FE",x"16",x"DA", -- 0x0BD8
    x"EB",x"0B",x"CD",x"7D",x"27",x"CD",x"11",x"0B", -- 0x0BE0
    x"C3",x"B9",x"07",x"DD",x"5E",x"0F",x"DD",x"56", -- 0x0BE8
    x"10",x"13",x"DD",x"CB",x"0E",x"46",x"C2",x"32", -- 0x0BF0
    x"0C",x"EB",x"7E",x"DD",x"77",x"0B",x"23",x"5E", -- 0x0BF8
    x"DD",x"73",x"07",x"23",x"56",x"DD",x"72",x"08", -- 0x0C00
    x"1A",x"DD",x"AE",x"0C",x"DD",x"77",x"09",x"23", -- 0x0C08
    x"5E",x"DD",x"73",x"01",x"23",x"56",x"DD",x"72", -- 0x0C10
    x"02",x"1A",x"0F",x"0F",x"0F",x"0F",x"E6",x"0F", -- 0x0C18
    x"DD",x"77",x"03",x"DD",x"77",x"05",x"1A",x"E6", -- 0x0C20
    x"0F",x"DD",x"77",x"04",x"DD",x"77",x"06",x"C3", -- 0x0C28
    x"B9",x"07",x"C5",x"ED",x"5F",x"E6",x"0F",x"C6", -- 0x0C30
    x"08",x"DD",x"77",x"0B",x"12",x"13",x"ED",x"5F", -- 0x0C38
    x"E6",x"0C",x"4F",x"06",x"00",x"21",x"68",x"2B", -- 0x0C40
    x"09",x"7E",x"23",x"12",x"13",x"4F",x"DD",x"77", -- 0x0C48
    x"07",x"7E",x"23",x"47",x"12",x"13",x"DD",x"77", -- 0x0C50
    x"08",x"0A",x"DD",x"AE",x"0C",x"DD",x"77",x"09", -- 0x0C58
    x"DD",x"36",x"0A",x"04",x"7E",x"23",x"4F",x"12", -- 0x0C60
    x"13",x"DD",x"77",x"01",x"7E",x"47",x"12",x"DD", -- 0x0C68
    x"77",x"02",x"0A",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x0C70
    x"0F",x"DD",x"77",x"03",x"DD",x"77",x"05",x"0A", -- 0x0C78
    x"E6",x"0F",x"DD",x"77",x"04",x"DD",x"77",x"06", -- 0x0C80
    x"C1",x"C3",x"B9",x"07",x"DD",x"35",x"13",x"C2", -- 0x0C88
    x"B9",x"07",x"DD",x"36",x"13",x"50",x"DD",x"7E", -- 0x0C90
    x"00",x"FE",x"18",x"CA",x"02",x"0D",x"FE",x"16", -- 0x0C98
    x"C2",x"B9",x"07",x"2A",x"72",x"40",x"7C",x"B5", -- 0x0CA0
    x"CA",x"B9",x"07",x"11",x"00",x"00",x"ED",x"53", -- 0x0CA8
    x"72",x"40",x"ED",x"5B",x"74",x"40",x"36",x"06", -- 0x0CB0
    x"DD",x"75",x"16",x"DD",x"74",x"17",x"DD",x"73", -- 0x0CB8
    x"18",x"DD",x"72",x"19",x"DD",x"36",x"14",x"08", -- 0x0CC0
    x"DD",x"36",x"15",x"F0",x"FD",x"7E",x"00",x"D6", -- 0x0CC8
    x"08",x"FD",x"77",x"00",x"C6",x"0F",x"12",x"13", -- 0x0CD0
    x"FD",x"34",x"01",x"FD",x"7E",x"01",x"F6",x"80", -- 0x0CD8
    x"12",x"13",x"FD",x"7E",x"02",x"12",x"13",x"FD", -- 0x0CE0
    x"7E",x"03",x"12",x"DD",x"36",x"1A",x"0F",x"DD", -- 0x0CE8
    x"36",x"1B",x"0B",x"DD",x"36",x"1C",x"05",x"DD", -- 0x0CF0
    x"36",x"1D",x"11",x"DD",x"36",x"00",x"18",x"C3", -- 0x0CF8
    x"B9",x"07",x"FD",x"34",x"01",x"DD",x"6E",x"18", -- 0x0D00
    x"DD",x"66",x"19",x"23",x"34",x"DD",x"36",x"1A", -- 0x0D08
    x"0F",x"DD",x"36",x"1B",x"10",x"DD",x"36",x"1C", -- 0x0D10
    x"05",x"DD",x"36",x"1D",x"16",x"DD",x"36",x"00", -- 0x0D18
    x"1A",x"C3",x"B9",x"07",x"DD",x"6E",x"0F",x"DD", -- 0x0D20
    x"66",x"10",x"DD",x"36",x"0F",x"00",x"35",x"C8", -- 0x0D28
    x"DD",x"CB",x"0E",x"46",x"C8",x"7D",x"11",x"24", -- 0x0D30
    x"00",x"21",x"D5",x"41",x"19",x"BE",x"C2",x"3C", -- 0x0D38
    x"0D",x"2B",x"CB",x"C6",x"C9",x"DD",x"21",x"AA", -- 0x0D40
    x"41",x"3A",x"05",x"40",x"E6",x"0C",x"CA",x"7C", -- 0x0D48
    x"0D",x"FE",x"0C",x"CA",x"7C",x"0D",x"CB",x"57", -- 0x0D50
    x"21",x"A2",x"41",x"DD",x"7E",x"00",x"C2",x"70", -- 0x0D58
    x"0D",x"FE",x"E1",x"CA",x"7C",x"0D",x"DD",x"34", -- 0x0D60
    x"00",x"34",x"DD",x"34",x"04",x"C3",x"7C",x"0D", -- 0x0D68
    x"FE",x"0F",x"CA",x"7C",x"0D",x"DD",x"35",x"00", -- 0x0D70
    x"35",x"DD",x"35",x"04",x"3A",x"65",x"40",x"3C", -- 0x0D78
    x"E6",x"03",x"32",x"65",x"40",x"CA",x"49",x"0D", -- 0x0D80
    x"21",x"76",x"40",x"35",x"C2",x"A5",x"0D",x"3A", -- 0x0D88
    x"78",x"40",x"77",x"DD",x"35",x"03",x"DD",x"35", -- 0x0D90
    x"07",x"EB",x"21",x"20",x"41",x"3A",x"1B",x"41", -- 0x0D98
    x"37",x"17",x"86",x"77",x"EB",x"23",x"35",x"C2", -- 0x0DA0
    x"B5",x"0D",x"36",x"0F",x"23",x"35",x"7E",x"FE", -- 0x0DA8
    x"02",x"D2",x"B5",x"0D",x"34",x"21",x"6E",x"40", -- 0x0DB0
    x"35",x"C2",x"C6",x"0D",x"36",x"03",x"DD",x"7E", -- 0x0DB8
    x"05",x"EE",x"34",x"DD",x"77",x"05",x"3A",x"10", -- 0x0DC0
    x"40",x"DD",x"46",x"03",x"FE",x"00",x"CA",x"E0", -- 0x0DC8
    x"0D",x"FE",x"01",x"CA",x"E6",x"0D",x"FE",x"02", -- 0x0DD0
    x"C0",x"78",x"FE",x"E0",x"C0",x"C3",x"E6",x"0D", -- 0x0DD8
    x"78",x"A7",x"CA",x"E6",x"0D",x"C9",x"21",x"10", -- 0x0DE0
    x"40",x"34",x"C9",x"21",x"1D",x"40",x"35",x"C0", -- 0x0DE8
    x"36",x"08",x"3A",x"08",x"41",x"FE",x"06",x"C0", -- 0x0DF0
    x"3A",x"1E",x"40",x"21",x"27",x"41",x"BE",x"C8", -- 0x0DF8
    x"3A",x"0C",x"41",x"A7",x"C8",x"47",x"DD",x"21", -- 0x0E00
    x"C6",x"41",x"FD",x"21",x"A6",x"41",x"11",x"24", -- 0x0E08
    x"00",x"DD",x"19",x"11",x"04",x"00",x"FD",x"19", -- 0x0E10
    x"DD",x"7E",x"00",x"1E",x"00",x"FE",x"12",x"CA", -- 0x0E18
    x"2D",x"0E",x"1D",x"FE",x"1A",x"CA",x"2D",x"0E", -- 0x0E20
    x"FE",x"1C",x"C2",x"93",x"0E",x"FD",x"7E",x"00", -- 0x0E28
    x"FE",x"0A",x"DA",x"93",x"0E",x"FE",x"E7",x"D2", -- 0x0E30
    x"93",x"0E",x"FD",x"7E",x"03",x"FE",x"A0",x"D2", -- 0x0E38
    x"93",x"0E",x"3A",x"A2",x"41",x"FD",x"96",x"00", -- 0x0E40
    x"C6",x"89",x"FE",x"21",x"D2",x"93",x"0E",x"FD", -- 0x0E48
    x"7E",x"00",x"DD",x"86",x"1E",x"4F",x"ED",x"5F", -- 0x0E50
    x"E6",x"07",x"D6",x"04",x"A3",x"81",x"21",x"C7", -- 0x0E58
    x"41",x"11",x"04",x"00",x"0E",x"07",x"19",x"BE", -- 0x0E60
    x"CA",x"93",x"0E",x"0D",x"C2",x"66",x"0E",x"DD", -- 0x0E68
    x"21",x"C6",x"41",x"47",x"DD",x"19",x"DD",x"7E", -- 0x0E70
    x"01",x"DD",x"B6",x"03",x"C2",x"74",x"0E",x"DD", -- 0x0E78
    x"70",x"01",x"3E",x"F5",x"FD",x"96",x"03",x"21", -- 0x0E80
    x"1B",x"41",x"AE",x"DD",x"77",x"03",x"21",x"1E", -- 0x0E88
    x"40",x"34",x"C9",x"DD",x"7E",x"00",x"FE",x"08", -- 0x0E90
    x"DA",x"0E",x"0E",x"05",x"C2",x"0E",x"0E",x"C9", -- 0x0E98
    x"3A",x"1E",x"40",x"A7",x"C8",x"47",x"DD",x"21", -- 0x0EA0
    x"C6",x"41",x"11",x"04",x"00",x"DD",x"19",x"DD", -- 0x0EA8
    x"7E",x"03",x"A7",x"CA",x"AD",x"0E",x"21",x"1B", -- 0x0EB0
    x"41",x"AE",x"D6",x"03",x"AE",x"DD",x"77",x"03", -- 0x0EB8
    x"AE",x"FE",x"1B",x"D2",x"05",x"0F",x"3A",x"08", -- 0x0EC0
    x"41",x"FE",x"06",x"C2",x"ED",x"0E",x"3A",x"A2", -- 0x0EC8
    x"41",x"C6",x"87",x"DD",x"96",x"01",x"FE",x"0D", -- 0x0ED0
    x"D2",x"ED",x"0E",x"DD",x"36",x"01",x"00",x"DD", -- 0x0ED8
    x"36",x"03",x"00",x"21",x"1E",x"40",x"35",x"3E", -- 0x0EE0
    x"0C",x"32",x"08",x"41",x"C9",x"DD",x"7E",x"03", -- 0x0EE8
    x"21",x"1B",x"41",x"AE",x"FE",x"0F",x"D2",x"05", -- 0x0EF0
    x"0F",x"DD",x"36",x"03",x"00",x"DD",x"36",x"01", -- 0x0EF8
    x"00",x"21",x"1E",x"40",x"35",x"10",x"A6",x"C9", -- 0x0F00
    x"3A",x"08",x"41",x"FE",x"06",x"C0",x"3A",x"0C", -- 0x0F08
    x"41",x"21",x"29",x"41",x"BE",x"C8",x"47",x"3A", -- 0x0F10
    x"0B",x"41",x"90",x"C8",x"4F",x"CD",x"09",x"28", -- 0x0F18
    x"47",x"3A",x"0B",x"41",x"21",x"34",x"41",x"BE", -- 0x0F20
    x"78",x"D2",x"32",x"0F",x"E6",x"01",x"3C",x"C3", -- 0x0F28
    x"35",x"0F",x"E6",x"03",x"86",x"47",x"79",x"90", -- 0x0F30
    x"D8",x"3A",x"0C",x"41",x"80",x"21",x"29",x"41", -- 0x0F38
    x"3D",x"BE",x"D0",x"3C",x"32",x"0C",x"41",x"21", -- 0x0F40
    x"1C",x"40",x"11",x"08",x"00",x"AF",x"19",x"BE", -- 0x0F48
    x"C2",x"4E",x"0F",x"70",x"CD",x"09",x"28",x"4F", -- 0x0F50
    x"CB",x"3F",x"A1",x"2F",x"F6",x"01",x"E6",x"03", -- 0x0F58
    x"4F",x"DD",x"21",x"C6",x"41",x"FD",x"21",x"A6", -- 0x0F60
    x"41",x"11",x"24",x"00",x"DD",x"19",x"11",x"04", -- 0x0F68
    x"00",x"FD",x"19",x"DD",x"7E",x"00",x"FE",x"00", -- 0x0F70
    x"C2",x"69",x"0F",x"ED",x"5F",x"E6",x"03",x"80", -- 0x0F78
    x"DD",x"36",x"0D",x"08",x"16",x"07",x"FE",x"03", -- 0x0F80
    x"D2",x"91",x"0F",x"16",x"04",x"DD",x"36",x"0D", -- 0x0F88
    x"05",x"FD",x"72",x"02",x"DD",x"71",x"0E",x"DD", -- 0x0F90
    x"71",x"11",x"DD",x"75",x"0F",x"DD",x"74",x"10", -- 0x0F98
    x"DD",x"36",x"0A",x"04",x"DD",x"36",x"00",x"0A", -- 0x0FA0
    x"DD",x"36",x"14",x"00",x"DD",x"36",x"15",x"00", -- 0x0FA8
    x"DD",x"36",x"1A",x"07",x"DD",x"36",x"1B",x"08", -- 0x0FB0
    x"DD",x"36",x"1C",x"08",x"DD",x"36",x"1D",x"0E", -- 0x0FB8
    x"DD",x"36",x"1E",x"08",x"DD",x"36",x"22",x"FF", -- 0x0FC0
    x"DD",x"36",x"23",x"07",x"3E",x"28",x"81",x"E6", -- 0x0FC8
    x"FE",x"4F",x"10",x"95",x"11",x"06",x"00",x"19", -- 0x0FD0
    x"ED",x"5F",x"E6",x"7F",x"4F",x"ED",x"5F",x"E6", -- 0x0FD8
    x"3F",x"81",x"C6",x"1C",x"77",x"FE",x"60",x"DA", -- 0x0FE0
    x"EC",x"0F",x"CB",x"C8",x"ED",x"5F",x"E6",x"01", -- 0x0FE8
    x"B0",x"47",x"07",x"07",x"B0",x"47",x"07",x"07", -- 0x0FF0
    x"07",x"07",x"B0",x"23",x"77",x"C9",x"3A",x"08", -- 0x0FF8
    x"41",x"FE",x"06",x"C0",x"21",x"0C",x"41",x"3A", -- 0x1000
    x"29",x"41",x"BE",x"C8",x"3A",x"0B",x"41",x"BE", -- 0x1008
    x"C8",x"34",x"21",x"00",x"00",x"22",x"72",x"40", -- 0x1010
    x"DD",x"21",x"C6",x"41",x"FD",x"21",x"A6",x"41", -- 0x1018
    x"01",x"24",x"00",x"11",x"04",x"00",x"DD",x"09", -- 0x1020
    x"FD",x"19",x"DD",x"7E",x"00",x"FE",x"00",x"C2", -- 0x1028
    x"26",x"10",x"FD",x"36",x"01",x"11",x"ED",x"5F", -- 0x1030
    x"E6",x"3F",x"C6",x"10",x"FD",x"77",x"03",x"ED", -- 0x1038
    x"5F",x"E6",x"7F",x"C6",x"40",x"FD",x"77",x"00", -- 0x1040
    x"DD",x"36",x"0D",x"10",x"21",x"30",x"41",x"3A", -- 0x1048
    x"0B",x"41",x"BE",x"3E",x"07",x"D2",x"69",x"10", -- 0x1050
    x"DD",x"36",x"0D",x"15",x"FE",x"01",x"3E",x"04", -- 0x1058
    x"C2",x"69",x"10",x"3E",x"02",x"DD",x"36",x"0D", -- 0x1060
    x"20",x"FD",x"77",x"02",x"DD",x"CB",x"0E",x"C6", -- 0x1068
    x"DD",x"36",x"1E",x"10",x"DD",x"36",x"13",x"50", -- 0x1070
    x"DD",x"36",x"14",x"12",x"DD",x"36",x"15",x"E8", -- 0x1078
    x"DD",x"36",x"1A",x"07",x"DD",x"36",x"1B",x"08", -- 0x1080
    x"DD",x"36",x"1C",x"08",x"DD",x"36",x"1D",x"0E", -- 0x1088
    x"CD",x"09",x"28",x"E6",x"01",x"5F",x"3A",x"31", -- 0x1090
    x"41",x"3C",x"07",x"2F",x"E6",x"07",x"C2",x"A2", -- 0x1098
    x"10",x"3C",x"83",x"DD",x"77",x"11",x"DD",x"36", -- 0x10A0
    x"22",x"FF",x"CD",x"7D",x"27",x"DD",x"36",x"00", -- 0x10A8
    x"16",x"C9",x"CD",x"FC",x"26",x"CD",x"B1",x"26", -- 0x10B0
    x"AF",x"32",x"06",x"70",x"32",x"07",x"70",x"3E", -- 0x10B8
    x"01",x"32",x"02",x"60",x"21",x"47",x"52",x"11", -- 0x10C0
    x"C2",x"18",x"CD",x"E7",x"26",x"21",x"39",x"53", -- 0x10C8
    x"11",x"FB",x"18",x"CD",x"E7",x"26",x"21",x"38", -- 0x10D0
    x"53",x"11",x"11",x"19",x"CD",x"E7",x"26",x"21", -- 0x10D8
    x"37",x"53",x"11",x"27",x"19",x"CD",x"E7",x"26", -- 0x10E0
    x"21",x"36",x"53",x"11",x"3C",x"19",x"CD",x"E7", -- 0x10E8
    x"26",x"3E",x"02",x"32",x"00",x"40",x"C9",x"21", -- 0x10F0
    x"1F",x"40",x"35",x"C0",x"3E",x"04",x"32",x"00", -- 0x10F8
    x"40",x"CD",x"FC",x"26",x"3E",x"00",x"32",x"02", -- 0x1100
    x"60",x"CD",x"41",x"27",x"CD",x"BF",x"12",x"CD", -- 0x1108
    x"09",x"28",x"E6",x"1F",x"3C",x"32",x"9B",x"40", -- 0x1110
    x"3A",x"9C",x"40",x"EE",x"04",x"32",x"9C",x"40", -- 0x1118
    x"EE",x"04",x"32",x"06",x"41",x"A7",x"CA",x"2D", -- 0x1120
    x"11",x"CD",x"6F",x"15",x"C9",x"CD",x"2D",x"18", -- 0x1128
    x"C9",x"3A",x"04",x"40",x"CB",x"4F",x"C2",x"4D", -- 0x1130
    x"11",x"CB",x"47",x"C8",x"3A",x"08",x"40",x"C6", -- 0x1138
    x"99",x"27",x"32",x"08",x"40",x"CD",x"FC",x"26", -- 0x1140
    x"3E",x"08",x"C3",x"65",x"11",x"3A",x"08",x"40", -- 0x1148
    x"C6",x"98",x"27",x"D0",x"32",x"08",x"40",x"CD", -- 0x1150
    x"FC",x"26",x"21",x"8F",x"52",x"11",x"C9",x"18", -- 0x1158
    x"CD",x"E7",x"26",x"3E",x"0A",x"32",x"00",x"40", -- 0x1160
    x"AF",x"32",x"8E",x"40",x"3E",x"80",x"32",x"11", -- 0x1168
    x"41",x"C9",x"CD",x"08",x"04",x"CD",x"84",x"28", -- 0x1170
    x"3A",x"08",x"41",x"FE",x"0E",x"CA",x"AD",x"11", -- 0x1178
    x"CD",x"4D",x"05",x"CD",x"08",x"0F",x"CD",x"97", -- 0x1180
    x"07",x"CD",x"EB",x"0D",x"CD",x"A0",x"0E",x"3A", -- 0x1188
    x"0B",x"41",x"A7",x"C0",x"3A",x"1E",x"40",x"A7", -- 0x1190
    x"C0",x"3A",x"08",x"41",x"FE",x"06",x"C0",x"3A", -- 0x1198
    x"00",x"40",x"C6",x"FA",x"32",x"00",x"40",x"21", -- 0x11A0
    x"06",x"41",x"34",x"34",x"C9",x"3A",x"00",x"40", -- 0x11A8
    x"FE",x"04",x"CA",x"9A",x"14",x"21",x"97",x"29", -- 0x11B0
    x"22",x"0C",x"40",x"21",x"00",x"00",x"22",x"0E", -- 0x11B8
    x"40",x"21",x"60",x"50",x"FE",x"18",x"CA",x"CC", -- 0x11C0
    x"11",x"21",x"A0",x"53",x"35",x"CD",x"B1",x"26", -- 0x11C8
    x"21",x"10",x"41",x"35",x"C2",x"04",x"12",x"CD", -- 0x11D0
    x"FC",x"26",x"21",x"8D",x"52",x"11",x"DF",x"18", -- 0x11D8
    x"CD",x"E7",x"26",x"3A",x"00",x"40",x"FE",x"14", -- 0x11E0
    x"CA",x"FF",x"11",x"21",x"8F",x"52",x"11",x"C9", -- 0x11E8
    x"18",x"FE",x"16",x"CA",x"F9",x"11",x"11",x"D4", -- 0x11F0
    x"18",x"CD",x"E7",x"26",x"3A",x"00",x"40",x"C6", -- 0x11F8
    x"12",x"C3",x"42",x"12",x"3A",x"00",x"40",x"FE", -- 0x1200
    x"14",x"CA",x"3D",x"12",x"CD",x"FC",x"26",x"21", -- 0x1208
    x"8F",x"52",x"11",x"D4",x"18",x"3A",x"00",x"40", -- 0x1210
    x"FE",x"16",x"3A",x"8F",x"40",x"CA",x"24",x"12", -- 0x1218
    x"AF",x"11",x"C9",x"18",x"32",x"06",x"70",x"32", -- 0x1220
    x"07",x"70",x"CD",x"E7",x"26",x"3A",x"20",x"40", -- 0x1228
    x"A7",x"C2",x"3D",x"12",x"21",x"8D",x"52",x"11", -- 0x1230
    x"DF",x"18",x"CD",x"E7",x"26",x"3A",x"00",x"40", -- 0x1238
    x"C6",x"06",x"32",x"00",x"40",x"3E",x"80",x"32", -- 0x1240
    x"11",x"41",x"C9",x"21",x"11",x"41",x"35",x"C0", -- 0x1248
    x"3A",x"00",x"40",x"FE",x"08",x"CA",x"63",x"12", -- 0x1250
    x"3A",x"69",x"40",x"32",x"60",x"50",x"3E",x"64", -- 0x1258
    x"32",x"40",x"50",x"3A",x"69",x"40",x"32",x"A0", -- 0x1260
    x"53",x"3E",x"64",x"32",x"80",x"53",x"11",x"6B", -- 0x1268
    x"29",x"CD",x"1F",x"27",x"CD",x"FC",x"26",x"3E", -- 0x1270
    x"00",x"32",x"02",x"60",x"CD",x"2D",x"18",x"3A", -- 0x1278
    x"00",x"40",x"C6",x"0C",x"32",x"00",x"40",x"CD", -- 0x1280
    x"41",x"27",x"3A",x"8F",x"40",x"3D",x"2F",x"32", -- 0x1288
    x"1B",x"41",x"21",x"03",x"41",x"22",x"0E",x"41", -- 0x1290
    x"3E",x"18",x"32",x"12",x"41",x"3A",x"69",x"40", -- 0x1298
    x"32",x"10",x"41",x"CD",x"BF",x"12",x"CD",x"5F", -- 0x12A0
    x"27",x"AF",x"32",x"1B",x"41",x"21",x"00",x"41", -- 0x12A8
    x"22",x"0E",x"41",x"3A",x"00",x"40",x"32",x"12", -- 0x12B0
    x"41",x"3A",x"69",x"40",x"32",x"10",x"41",x"3E", -- 0x12B8
    x"10",x"32",x"0B",x"41",x"3E",x"03",x"32",x"30", -- 0x12C0
    x"41",x"3E",x"03",x"32",x"34",x"41",x"3E",x"05", -- 0x12C8
    x"32",x"29",x"41",x"3E",x"18",x"21",x"1B",x"41", -- 0x12D0
    x"AE",x"32",x"20",x"41",x"3E",x"03",x"32",x"13", -- 0x12D8
    x"41",x"3E",x"02",x"32",x"27",x"41",x"3E",x"22", -- 0x12E0
    x"32",x"18",x"41",x"3E",x"04",x"32",x"19",x"41", -- 0x12E8
    x"3E",x"03",x"32",x"1A",x"41",x"3E",x"08",x"32", -- 0x12F0
    x"1E",x"41",x"3E",x"0F",x"32",x"1F",x"41",x"3E", -- 0x12F8
    x"05",x"32",x"35",x"41",x"3E",x"25",x"32",x"36", -- 0x1300
    x"41",x"3E",x"05",x"32",x"37",x"41",x"3E",x"08", -- 0x1308
    x"32",x"24",x"41",x"3E",x"20",x"32",x"28",x"41", -- 0x1310
    x"3E",x"50",x"32",x"2B",x"41",x"3E",x"C0",x"32", -- 0x1318
    x"2F",x"41",x"3E",x"1F",x"32",x"2A",x"41",x"3E", -- 0x1320
    x"40",x"32",x"2D",x"41",x"3E",x"02",x"32",x"2E", -- 0x1328
    x"41",x"3E",x"08",x"32",x"08",x"41",x"3E",x"80", -- 0x1330
    x"32",x"0A",x"41",x"3E",x"01",x"32",x"21",x"41", -- 0x1338
    x"3A",x"00",x"70",x"CB",x"57",x"3E",x"01",x"C2", -- 0x1340
    x"4B",x"13",x"AF",x"32",x"31",x"41",x"C9",x"21", -- 0x1348
    x"31",x"41",x"34",x"3E",x"10",x"32",x"0B",x"41", -- 0x1350
    x"3E",x"08",x"32",x"29",x"41",x"3E",x"00",x"32", -- 0x1358
    x"02",x"60",x"3E",x"03",x"32",x"13",x"41",x"CD", -- 0x1360
    x"93",x"18",x"21",x"31",x"41",x"3E",x"03",x"96", -- 0x1368
    x"FE",x"01",x"D2",x"77",x"13",x"3E",x"01",x"32", -- 0x1370
    x"34",x"41",x"3A",x"00",x"40",x"C6",x"06",x"32", -- 0x1378
    x"00",x"40",x"C9",x"21",x"11",x"41",x"35",x"C0", -- 0x1380
    x"3A",x"00",x"40",x"FE",x"1A",x"3E",x"20",x"CA", -- 0x1388
    x"AB",x"13",x"CD",x"FC",x"26",x"3A",x"20",x"40", -- 0x1390
    x"A7",x"CA",x"AF",x"13",x"CD",x"5F",x"27",x"3A", -- 0x1398
    x"00",x"40",x"FE",x"1C",x"3E",x"24",x"CA",x"AB", -- 0x13A0
    x"13",x"3E",x"22",x"32",x"00",x"40",x"C9",x"CD", -- 0x13A8
    x"5F",x"27",x"21",x"8F",x"52",x"11",x"C9",x"18", -- 0x13B0
    x"3A",x"00",x"40",x"FE",x"1C",x"3E",x"1E",x"CA", -- 0x13B8
    x"C7",x"13",x"3E",x"1C",x"11",x"D4",x"18",x"32", -- 0x13C0
    x"00",x"40",x"3A",x"4D",x"41",x"E6",x"01",x"C3", -- 0x13C8
    x"33",x"14",x"C9",x"CD",x"2D",x"18",x"3E",x"00", -- 0x13D0
    x"32",x"02",x"60",x"C3",x"F4",x"13",x"3E",x"01", -- 0x13D8
    x"32",x"00",x"68",x"32",x"01",x"68",x"32",x"02", -- 0x13E0
    x"68",x"3E",x"01",x"32",x"02",x"60",x"21",x"00", -- 0x13E8
    x"00",x"22",x"14",x"41",x"3E",x"08",x"32",x"08", -- 0x13F0
    x"41",x"3A",x"00",x"40",x"C6",x"F4",x"32",x"00", -- 0x13F8
    x"40",x"C9",x"21",x"11",x"41",x"35",x"C0",x"CD", -- 0x1400
    x"FC",x"26",x"3A",x"00",x"40",x"FE",x"26",x"CA", -- 0x1408
    x"42",x"14",x"3A",x"20",x"40",x"A7",x"CA",x"42", -- 0x1410
    x"14",x"3A",x"00",x"40",x"C6",x"F4",x"32",x"00", -- 0x1418
    x"40",x"21",x"8F",x"52",x"11",x"D4",x"18",x"FE", -- 0x1420
    x"1C",x"3A",x"8F",x"40",x"CA",x"33",x"14",x"AF", -- 0x1428
    x"11",x"C9",x"18",x"32",x"06",x"70",x"32",x"07", -- 0x1430
    x"70",x"CD",x"E7",x"26",x"3E",x"80",x"32",x"11", -- 0x1438
    x"41",x"C9",x"A7",x"2A",x"22",x"40",x"ED",x"5B", -- 0x1440
    x"01",x"41",x"ED",x"52",x"DA",x"5D",x"14",x"C2", -- 0x1448
    x"68",x"14",x"3A",x"00",x"41",x"47",x"3A",x"21", -- 0x1450
    x"40",x"90",x"D2",x"68",x"14",x"ED",x"53",x"22", -- 0x1458
    x"40",x"3A",x"00",x"41",x"32",x"21",x"40",x"3F", -- 0x1460
    x"2A",x"22",x"40",x"ED",x"5B",x"04",x"41",x"ED", -- 0x1468
    x"52",x"DA",x"82",x"14",x"C2",x"8C",x"14",x"3A", -- 0x1470
    x"03",x"41",x"47",x"3A",x"21",x"40",x"90",x"D2", -- 0x1478
    x"8C",x"14",x"ED",x"53",x"22",x"40",x"3A",x"03", -- 0x1480
    x"41",x"32",x"21",x"40",x"3E",x"10",x"32",x"A0", -- 0x1488
    x"53",x"32",x"80",x"53",x"32",x"60",x"50",x"32", -- 0x1490
    x"40",x"50",x"AF",x"32",x"A6",x"41",x"32",x"A8", -- 0x1498
    x"41",x"32",x"74",x"41",x"32",x"76",x"41",x"32", -- 0x14A0
    x"78",x"41",x"32",x"7A",x"41",x"3E",x"00",x"32", -- 0x14A8
    x"00",x"40",x"C9",x"DD",x"21",x"AA",x"41",x"3A", -- 0x14B0
    x"1B",x"41",x"E6",x"FE",x"C6",x"79",x"47",x"3A", -- 0x14B8
    x"A2",x"41",x"80",x"47",x"DD",x"77",x"00",x"DD", -- 0x14C0
    x"36",x"03",x"E0",x"DD",x"36",x"01",x"18",x"DD", -- 0x14C8
    x"36",x"02",x"07",x"3E",x"10",x"32",x"FC",x"51", -- 0x14D0
    x"32",x"FD",x"51",x"32",x"1C",x"52",x"32",x"1D", -- 0x14D8
    x"52",x"DD",x"70",x"04",x"DD",x"36",x"07",x"EE", -- 0x14E0
    x"DD",x"36",x"05",x"1B",x"DD",x"36",x"06",x"07", -- 0x14E8
    x"3E",x"0A",x"32",x"78",x"40",x"C6",x"60",x"32", -- 0x14F0
    x"76",x"40",x"3E",x"10",x"32",x"77",x"40",x"3E", -- 0x14F8
    x"03",x"32",x"6E",x"40",x"3E",x"01",x"32",x"03", -- 0x1500
    x"68",x"21",x"37",x"2A",x"22",x"0C",x"40",x"21", -- 0x1508
    x"00",x"00",x"22",x"0E",x"40",x"3E",x"01",x"32", -- 0x1510
    x"02",x"40",x"3E",x"00",x"32",x"10",x"40",x"3A", -- 0x1518
    x"00",x"40",x"C6",x"06",x"32",x"00",x"40",x"CD", -- 0x1520
    x"45",x"0D",x"CD",x"4D",x"05",x"3A",x"10",x"40", -- 0x1528
    x"FE",x"01",x"C2",x"39",x"15",x"CD",x"FC",x"26", -- 0x1530
    x"C9",x"FE",x"03",x"C0",x"AF",x"32",x"03",x"68", -- 0x1538
    x"06",x"08",x"21",x"AA",x"41",x"36",x"00",x"23", -- 0x1540
    x"10",x"FB",x"3A",x"A2",x"41",x"32",x"A4",x"41", -- 0x1548
    x"3E",x"60",x"32",x"FC",x"51",x"3C",x"32",x"FD", -- 0x1550
    x"51",x"3C",x"32",x"1C",x"52",x"3C",x"32",x"1D", -- 0x1558
    x"52",x"21",x"06",x"41",x"34",x"34",x"3A",x"00", -- 0x1560
    x"40",x"C6",x"FA",x"32",x"00",x"40",x"C9",x"3E", -- 0x1568
    x"08",x"32",x"0B",x"41",x"32",x"29",x"41",x"21", -- 0x1570
    x"00",x"00",x"22",x"72",x"40",x"3E",x"01",x"32", -- 0x1578
    x"02",x"60",x"3E",x"01",x"32",x"13",x"41",x"CD", -- 0x1580
    x"93",x"18",x"3A",x"00",x"40",x"FE",x"04",x"C8", -- 0x1588
    x"3E",x"01",x"32",x"00",x"68",x"32",x"01",x"68", -- 0x1590
    x"32",x"02",x"68",x"3A",x"00",x"40",x"C6",x"06", -- 0x1598
    x"32",x"00",x"40",x"C9",x"3E",x"10",x"32",x"0B", -- 0x15A0
    x"41",x"3A",x"31",x"41",x"CB",x"27",x"C6",x"03", -- 0x15A8
    x"FE",x"07",x"DA",x"B7",x"15",x"3E",x"06",x"32", -- 0x15B0
    x"29",x"41",x"3E",x"20",x"32",x"28",x"41",x"3E", -- 0x15B8
    x"01",x"32",x"92",x"40",x"3E",x"60",x"32",x"93", -- 0x15C0
    x"40",x"CD",x"93",x"18",x"3A",x"31",x"41",x"3C", -- 0x15C8
    x"3C",x"FE",x"06",x"DA",x"D8",x"15",x"3E",x"05", -- 0x15D0
    x"32",x"27",x"41",x"3A",x"31",x"41",x"A7",x"CA", -- 0x15D8
    x"E6",x"15",x"AF",x"32",x"2F",x"41",x"3E",x"00", -- 0x15E0
    x"32",x"9D",x"40",x"3E",x"01",x"32",x"00",x"68", -- 0x15E8
    x"32",x"01",x"68",x"32",x"02",x"68",x"3A",x"00", -- 0x15F0
    x"40",x"C6",x"06",x"32",x"00",x"40",x"C9",x"3E", -- 0x15F8
    x"08",x"32",x"08",x"41",x"3E",x"01",x"32",x"92", -- 0x1600
    x"40",x"3E",x"60",x"32",x"93",x"40",x"CD",x"2D", -- 0x1608
    x"18",x"3E",x"00",x"32",x"9D",x"40",x"3E",x"01", -- 0x1610
    x"32",x"00",x"68",x"32",x"01",x"68",x"32",x"02", -- 0x1618
    x"68",x"3E",x"00",x"32",x"02",x"60",x"3A",x"00", -- 0x1620
    x"40",x"C6",x"F4",x"32",x"00",x"40",x"C9",x"CD", -- 0x1628
    x"08",x"04",x"CD",x"84",x"28",x"CD",x"4D",x"05", -- 0x1630
    x"CD",x"91",x"20",x"CD",x"28",x"22",x"CD",x"A0", -- 0x1638
    x"0E",x"CD",x"99",x"22",x"CD",x"48",x"23",x"CD", -- 0x1640
    x"FA",x"24",x"3A",x"08",x"41",x"FE",x"0E",x"CA", -- 0x1648
    x"AD",x"11",x"3A",x"0B",x"41",x"A7",x"C0",x"3A", -- 0x1650
    x"1E",x"40",x"A7",x"C0",x"3A",x"9D",x"40",x"FE", -- 0x1658
    x"04",x"C0",x"CD",x"B1",x"26",x"3A",x"00",x"40", -- 0x1660
    x"C6",x"FA",x"32",x"00",x"40",x"3E",x"00",x"32", -- 0x1668
    x"06",x"41",x"C9",x"3A",x"00",x"40",x"C6",x"FA", -- 0x1670
    x"32",x"00",x"40",x"3E",x"00",x"32",x"06",x"41", -- 0x1678
    x"C9",x"DD",x"21",x"AA",x"41",x"3A",x"1B",x"41", -- 0x1680
    x"E6",x"FE",x"C6",x"79",x"47",x"3A",x"A2",x"41", -- 0x1688
    x"80",x"DD",x"77",x"00",x"DD",x"36",x"03",x"E0", -- 0x1690
    x"DD",x"36",x"02",x"07",x"DD",x"36",x"01",x"18", -- 0x1698
    x"3E",x"10",x"32",x"FC",x"51",x"32",x"FD",x"51", -- 0x16A0
    x"32",x"1C",x"52",x"32",x"1D",x"52",x"3E",x"11", -- 0x16A8
    x"32",x"78",x"40",x"32",x"76",x"40",x"3E",x"10", -- 0x16B0
    x"32",x"77",x"40",x"AF",x"32",x"7E",x"40",x"32", -- 0x16B8
    x"7B",x"40",x"32",x"80",x"40",x"3E",x"0A",x"32", -- 0x16C0
    x"7C",x"40",x"32",x"7D",x"40",x"3E",x"10",x"32", -- 0x16C8
    x"7F",x"40",x"3E",x"00",x"32",x"02",x"60",x"3E", -- 0x16D0
    x"02",x"32",x"08",x"41",x"3E",x"00",x"32",x"91", -- 0x16D8
    x"40",x"3E",x"00",x"32",x"17",x"41",x"AF",x"32", -- 0x16E0
    x"A6",x"41",x"32",x"A8",x"41",x"3E",x"00",x"32", -- 0x16E8
    x"1C",x"41",x"CD",x"79",x"18",x"21",x"31",x"41", -- 0x16F0
    x"3E",x"22",x"96",x"FE",x"1E",x"D2",x"02",x"17", -- 0x16F8
    x"3E",x"1E",x"32",x"18",x"41",x"21",x"19",x"41", -- 0x1700
    x"3A",x"31",x"41",x"C6",x"02",x"E6",x"03",x"CA", -- 0x1708
    x"13",x"17",x"34",x"21",x"1A",x"41",x"3A",x"31", -- 0x1710
    x"41",x"C6",x"02",x"E6",x"04",x"CA",x"2C",x"17", -- 0x1718
    x"7E",x"3D",x"FE",x"01",x"DA",x"2C",x"17",x"35", -- 0x1720
    x"21",x"19",x"41",x"35",x"3A",x"31",x"41",x"CB", -- 0x1728
    x"27",x"47",x"3E",x"08",x"90",x"DA",x"42",x"17", -- 0x1730
    x"FE",x"04",x"D2",x"3F",x"17",x"3E",x"04",x"32", -- 0x1738
    x"1E",x"41",x"3A",x"00",x"40",x"C6",x"06",x"32", -- 0x1740
    x"00",x"40",x"C9",x"3E",x"08",x"32",x"08",x"41", -- 0x1748
    x"CD",x"2D",x"18",x"3E",x"01",x"32",x"91",x"40", -- 0x1750
    x"3E",x"20",x"32",x"90",x"40",x"3E",x"02",x"32", -- 0x1758
    x"17",x"41",x"3E",x"00",x"32",x"02",x"60",x"CD", -- 0x1760
    x"79",x"18",x"3A",x"00",x"40",x"C6",x"F4",x"32", -- 0x1768
    x"00",x"40",x"C9",x"CD",x"08",x"04",x"CD",x"84", -- 0x1770
    x"28",x"CD",x"4D",x"05",x"3A",x"08",x"41",x"FE", -- 0x1778
    x"0E",x"CA",x"AD",x"11",x"CD",x"FE",x"0F",x"CD", -- 0x1780
    x"97",x"07",x"CD",x"EB",x"0D",x"CD",x"A0",x"0E", -- 0x1788
    x"3A",x"08",x"41",x"FE",x"06",x"C0",x"3A",x"0B", -- 0x1790
    x"41",x"A7",x"C0",x"3A",x"1E",x"40",x"A7",x"C0", -- 0x1798
    x"3E",x"01",x"32",x"7B",x"40",x"3A",x"0D",x"41", -- 0x17A0
    x"A7",x"C0",x"AF",x"32",x"00",x"68",x"32",x"01", -- 0x17A8
    x"68",x"32",x"02",x"68",x"3E",x"06",x"32",x"06", -- 0x17B0
    x"41",x"3A",x"00",x"40",x"C6",x"FA",x"32",x"00", -- 0x17B8
    x"40",x"C9",x"CD",x"26",x"1C",x"CD",x"49",x"19", -- 0x17C0
    x"CD",x"99",x"1F",x"CD",x"8C",x"1D",x"CD",x"62", -- 0x17C8
    x"1E",x"CD",x"AF",x"1D",x"3A",x"08",x"41",x"FE", -- 0x17D0
    x"0E",x"C2",x"E8",x"17",x"CD",x"FC",x"26",x"CD", -- 0x17D8
    x"2D",x"18",x"CD",x"54",x"18",x"C3",x"AD",x"11", -- 0x17E0
    x"FE",x"12",x"C0",x"CD",x"FC",x"26",x"CD",x"2D", -- 0x17E8
    x"18",x"3A",x"1B",x"41",x"E6",x"FE",x"C6",x"79", -- 0x17F0
    x"47",x"3A",x"AA",x"41",x"90",x"32",x"A2",x"41", -- 0x17F8
    x"32",x"A4",x"41",x"CD",x"B1",x"26",x"3E",x"60", -- 0x1800
    x"32",x"FC",x"51",x"3C",x"32",x"FD",x"51",x"3C", -- 0x1808
    x"32",x"1C",x"52",x"3C",x"32",x"1D",x"52",x"3E", -- 0x1810
    x"06",x"32",x"08",x"41",x"CD",x"54",x"18",x"3A", -- 0x1818
    x"00",x"40",x"C6",x"FA",x"32",x"00",x"40",x"3E", -- 0x1820
    x"08",x"32",x"06",x"41",x"C9",x"3E",x"04",x"32", -- 0x1828
    x"A7",x"41",x"32",x"A9",x"41",x"3E",x"02",x"32", -- 0x1830
    x"79",x"41",x"21",x"FE",x"53",x"11",x"DF",x"FF", -- 0x1838
    x"06",x"20",x"3E",x"90",x"77",x"23",x"3C",x"77", -- 0x1840
    x"3C",x"FE",x"9A",x"C2",x"50",x"18",x"3E",x"90", -- 0x1848
    x"19",x"10",x"F1",x"C9",x"AF",x"21",x"6E",x"41", -- 0x1850
    x"06",x"34",x"77",x"23",x"10",x"FC",x"3E",x"02", -- 0x1858
    x"32",x"79",x"41",x"32",x"9D",x"41",x"07",x"32", -- 0x1860
    x"9B",x"41",x"3E",x"05",x"32",x"A1",x"41",x"21", -- 0x1868
    x"80",x"52",x"11",x"F5",x"03",x"CD",x"E7",x"26", -- 0x1870
    x"C9",x"21",x"80",x"52",x"11",x"F0",x"18",x"CD", -- 0x1878
    x"E7",x"26",x"21",x"60",x"51",x"22",x"97",x"40", -- 0x1880
    x"3E",x"05",x"32",x"95",x"40",x"3E",x"35",x"32", -- 0x1888
    x"96",x"40",x"C9",x"3A",x"31",x"41",x"C6",x"03", -- 0x1890
    x"FE",x"06",x"DA",x"9F",x"18",x"3E",x"05",x"32", -- 0x1898
    x"27",x"41",x"3A",x"31",x"41",x"3C",x"CB",x"27", -- 0x18A0
    x"32",x"30",x"41",x"3A",x"31",x"41",x"2F",x"21", -- 0x18A8
    x"FF",x"FF",x"0F",x"CB",x"1C",x"0F",x"CB",x"1C", -- 0x18B0
    x"22",x"32",x"41",x"C9",x"C9",x"C9",x"C9",x"C9", -- 0x18B8
    x"C9",x"C9",x"50",x"49",x"53",x"43",x"45",x"53", -- 0x18C0
    x"FF",x"50",x"4C",x"41",x"59",x"45",x"52",x"20", -- 0x18C8
    x"4F",x"4E",x"45",x"FF",x"50",x"4C",x"41",x"59", -- 0x18D0
    x"45",x"52",x"20",x"54",x"57",x"4F",x"FF",x"47", -- 0x18D8
    x"41",x"4D",x"45",x"20",x"20",x"4F",x"56",x"45", -- 0x18E0
    x"52",x"FF",x"20",x"20",x"20",x"20",x"30",x"FF", -- 0x18E8
    x"46",x"55",x"45",x"4C",x"40",x"99",x"99",x"99", -- 0x18F0
    x"99",x"99",x"FF",x"3A",x"3B",x"3C",x"3D",x"3E", -- 0x18F8
    x"3F",x"5C",x"5D",x"5E",x"5F",x"60",x"61",x"62", -- 0x1900
    x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A", -- 0x1908
    x"FF",x"6B",x"6C",x"6D",x"6E",x"6F",x"70",x"71", -- 0x1910
    x"72",x"73",x"BF",x"C0",x"C1",x"C2",x"C3",x"C4", -- 0x1918
    x"C5",x"C6",x"C7",x"C8",x"C9",x"CA",x"FF",x"CB", -- 0x1920
    x"CC",x"CD",x"CE",x"20",x"CF",x"D0",x"D1",x"D2", -- 0x1928
    x"D3",x"D4",x"D5",x"D6",x"20",x"D7",x"D8",x"D9", -- 0x1930
    x"DA",x"DB",x"DC",x"FF",x"DD",x"DE",x"DF",x"E0", -- 0x1938
    x"20",x"20",x"E1",x"20",x"20",x"20",x"E2",x"E3", -- 0x1940
    x"FF",x"DD",x"21",x"AA",x"41",x"3A",x"08",x"41", -- 0x1948
    x"FE",x"00",x"CA",x"47",x"1A",x"FE",x"02",x"CA", -- 0x1950
    x"1B",x"1A",x"FE",x"04",x"CA",x"1B",x"1B",x"FE", -- 0x1958
    x"08",x"CA",x"74",x"19",x"FE",x"0C",x"CA",x"9C", -- 0x1960
    x"19",x"FE",x"0A",x"CA",x"D8",x"19",x"FE",x"10", -- 0x1968
    x"CA",x"0E",x"1A",x"C9",x"21",x"0A",x"41",x"35", -- 0x1970
    x"C0",x"DD",x"36",x"00",x"80",x"DD",x"36",x"03", -- 0x1978
    x"10",x"DD",x"36",x"01",x"18",x"DD",x"36",x"02", -- 0x1980
    x"07",x"3E",x"11",x"32",x"76",x"40",x"32",x"78", -- 0x1988
    x"40",x"3E",x"10",x"32",x"77",x"40",x"3E",x"00", -- 0x1990
    x"32",x"08",x"41",x"C9",x"AF",x"32",x"03",x"68", -- 0x1998
    x"11",x"1D",x"2A",x"CD",x"1F",x"27",x"CD",x"86", -- 0x19A0
    x"20",x"DD",x"7E",x"00",x"DD",x"77",x"04",x"DD", -- 0x19A8
    x"7E",x"03",x"C6",x"08",x"DD",x"77",x"07",x"D6", -- 0x19B0
    x"10",x"DD",x"77",x"03",x"3E",x"38",x"DD",x"77", -- 0x19B8
    x"01",x"3C",x"DD",x"77",x"05",x"DD",x"36",x"02", -- 0x19C0
    x"07",x"DD",x"36",x"06",x"07",x"3E",x"0A",x"32", -- 0x19C8
    x"79",x"40",x"3E",x"0A",x"32",x"08",x"41",x"C9", -- 0x19D0
    x"21",x"79",x"40",x"35",x"C0",x"36",x"0A",x"DD", -- 0x19D8
    x"7E",x"01",x"C6",x"02",x"FE",x"40",x"CA",x"F1", -- 0x19E0
    x"19",x"DD",x"77",x"01",x"3C",x"DD",x"77",x"05", -- 0x19E8
    x"C9",x"21",x"AA",x"41",x"06",x"08",x"AF",x"77", -- 0x19F0
    x"23",x"10",x"FC",x"3E",x"04",x"32",x"A7",x"41", -- 0x19F8
    x"32",x"A9",x"41",x"3E",x"80",x"32",x"0A",x"41", -- 0x1A00
    x"3E",x"10",x"32",x"08",x"41",x"C9",x"21",x"0A", -- 0x1A08
    x"41",x"35",x"C0",x"36",x"80",x"3E",x"0E",x"32", -- 0x1A10
    x"08",x"41",x"C9",x"DD",x"7E",x"03",x"A7",x"C2", -- 0x1A18
    x"29",x"1B",x"CD",x"2D",x"18",x"3E",x"01",x"32", -- 0x1A20
    x"91",x"40",x"3E",x"20",x"32",x"90",x"40",x"3E", -- 0x1A28
    x"02",x"32",x"1C",x"41",x"3A",x"1E",x"41",x"32", -- 0x1A30
    x"1D",x"41",x"3E",x"02",x"32",x"17",x"41",x"3E", -- 0x1A38
    x"00",x"32",x"08",x"41",x"C3",x"29",x"1B",x"DD", -- 0x1A40
    x"7E",x"03",x"FE",x"E0",x"C2",x"29",x"1B",x"DD", -- 0x1A48
    x"46",x"10",x"DD",x"7E",x"11",x"FE",x"27",x"CA", -- 0x1A50
    x"6D",x"1A",x"FE",x"29",x"CA",x"7B",x"1A",x"DD", -- 0x1A58
    x"7E",x"00",x"90",x"D6",x"05",x"FE",x"0C",x"DA", -- 0x1A60
    x"94",x"1A",x"C3",x"86",x"1A",x"DD",x"7E",x"00", -- 0x1A68
    x"90",x"D6",x"02",x"FE",x"0F",x"DA",x"94",x"1A", -- 0x1A70
    x"C3",x"86",x"1A",x"DD",x"7E",x"00",x"90",x"D6", -- 0x1A78
    x"04",x"FE",x"0D",x"DA",x"94",x"1A",x"3E",x"0C", -- 0x1A80
    x"32",x"08",x"41",x"3E",x"07",x"32",x"A7",x"41", -- 0x1A88
    x"32",x"A9",x"41",x"C9",x"3E",x"00",x"32",x"81", -- 0x1A90
    x"40",x"3E",x"04",x"32",x"08",x"41",x"3E",x"00", -- 0x1A98
    x"32",x"1C",x"41",x"21",x"9A",x"40",x"0E",x"00", -- 0x1AA0
    x"71",x"2B",x"71",x"ED",x"5B",x"97",x"40",x"1A", -- 0x1AA8
    x"D6",x"64",x"DA",x"C7",x"1A",x"E6",x"07",x"5F", -- 0x1AB0
    x"3A",x"95",x"40",x"CB",x"27",x"CB",x"27",x"83", -- 0x1AB8
    x"3C",x"11",x"35",x"41",x"CD",x"F2",x"1A",x"DD", -- 0x1AC0
    x"7E",x"15",x"D6",x"26",x"11",x"36",x"41",x"CD", -- 0x1AC8
    x"F2",x"1A",x"3A",x"1E",x"41",x"2F",x"0F",x"0F", -- 0x1AD0
    x"E6",x"07",x"C6",x"04",x"11",x"37",x"41",x"CD", -- 0x1AD8
    x"F2",x"1A",x"CD",x"4A",x"28",x"3E",x"03",x"32", -- 0x1AE0
    x"91",x"40",x"3E",x"04",x"32",x"90",x"40",x"C3", -- 0x1AE8
    x"E9",x"1F",x"01",x"00",x"00",x"08",x"08",x"3D", -- 0x1AF0
    x"CA",x"08",x"1B",x"08",x"1A",x"81",x"27",x"4F", -- 0x1AF8
    x"78",x"CE",x"00",x"27",x"47",x"C3",x"F6",x"1A", -- 0x1B00
    x"79",x"CD",x"2B",x"28",x"78",x"CD",x"18",x"28", -- 0x1B08
    x"79",x"86",x"27",x"77",x"23",x"78",x"8E",x"27", -- 0x1B10
    x"77",x"2B",x"C9",x"21",x"81",x"40",x"35",x"C0", -- 0x1B18
    x"CD",x"86",x"20",x"3E",x"12",x"32",x"08",x"41", -- 0x1B20
    x"C9",x"3A",x"05",x"40",x"E6",x"0C",x"CA",x"85", -- 0x1B28
    x"1B",x"FE",x"0C",x"CA",x"85",x"1B",x"CB",x"57", -- 0x1B30
    x"21",x"7B",x"40",x"C2",x"53",x"1B",x"34",x"7E", -- 0x1B38
    x"FE",x"08",x"DA",x"89",x"1B",x"36",x"00",x"23", -- 0x1B40
    x"3A",x"7E",x"40",x"FE",x"01",x"CA",x"67",x"1B", -- 0x1B48
    x"C3",x"7A",x"1B",x"35",x"7E",x"ED",x"44",x"FE", -- 0x1B50
    x"08",x"DA",x"89",x"1B",x"36",x"00",x"23",x"3A", -- 0x1B58
    x"7E",x"40",x"FE",x"01",x"CA",x"7A",x"1B",x"34", -- 0x1B60
    x"7E",x"FE",x"0B",x"DA",x"89",x"1B",x"35",x"3A", -- 0x1B68
    x"7E",x"40",x"EE",x"01",x"32",x"7E",x"40",x"C3", -- 0x1B70
    x"89",x"1B",x"35",x"7E",x"FE",x"01",x"D2",x"89", -- 0x1B78
    x"1B",x"34",x"C3",x"89",x"1B",x"AF",x"32",x"7B", -- 0x1B80
    x"40",x"21",x"7D",x"40",x"35",x"C2",x"C4",x"1B", -- 0x1B88
    x"3A",x"7E",x"40",x"FE",x"01",x"DD",x"7E",x"00", -- 0x1B90
    x"CA",x"A6",x"1B",x"FE",x"E1",x"CA",x"AB",x"1B", -- 0x1B98
    x"DD",x"34",x"00",x"C3",x"BE",x"1B",x"FE",x"0F", -- 0x1BA0
    x"C2",x"BB",x"1B",x"3E",x"0A",x"32",x"7C",x"40", -- 0x1BA8
    x"3A",x"7E",x"40",x"EE",x"01",x"32",x"7E",x"40", -- 0x1BB0
    x"C3",x"BE",x"1B",x"DD",x"35",x"00",x"3A",x"7C", -- 0x1BB8
    x"40",x"32",x"7D",x"40",x"21",x"7F",x"40",x"35", -- 0x1BC0
    x"C2",x"D9",x"1B",x"36",x"10",x"3A",x"7C",x"40", -- 0x1BC8
    x"FE",x"0A",x"CA",x"D9",x"1B",x"3C",x"32",x"7C", -- 0x1BD0
    x"40",x"21",x"76",x"40",x"35",x"C2",x"FD",x"1B", -- 0x1BD8
    x"3A",x"78",x"40",x"77",x"3A",x"80",x"40",x"FE", -- 0x1BE0
    x"01",x"CA",x"FA",x"1B",x"DD",x"7E",x"03",x"FE", -- 0x1BE8
    x"10",x"CA",x"FD",x"1B",x"DD",x"35",x"03",x"C3", -- 0x1BF0
    x"FD",x"1B",x"DD",x"34",x"03",x"23",x"35",x"C0", -- 0x1BF8
    x"36",x"0F",x"3A",x"80",x"40",x"FE",x"01",x"CA", -- 0x1C00
    x"1C",x"1C",x"23",x"34",x"34",x"7E",x"FE",x"12", -- 0x1C08
    x"D8",x"35",x"35",x"3A",x"80",x"40",x"EE",x"01", -- 0x1C10
    x"32",x"80",x"40",x"C9",x"23",x"35",x"35",x"7E", -- 0x1C18
    x"FE",x"02",x"D0",x"34",x"34",x"C9",x"3A",x"08", -- 0x1C20
    x"41",x"FE",x"03",x"D0",x"DD",x"21",x"AA",x"41", -- 0x1C28
    x"DD",x"7E",x"03",x"CB",x"3F",x"CB",x"3F",x"E6", -- 0x1C30
    x"3E",x"5F",x"CB",x"3F",x"16",x"00",x"FD",x"21", -- 0x1C38
    x"6A",x"41",x"FD",x"19",x"5F",x"16",x"50",x"ED", -- 0x1C40
    x"53",x"85",x"40",x"DD",x"7E",x"03",x"E6",x"07", -- 0x1C48
    x"3C",x"32",x"82",x"40",x"3E",x"03",x"32",x"87", -- 0x1C50
    x"40",x"DD",x"7E",x"00",x"C6",x"02",x"FD",x"96", -- 0x1C58
    x"00",x"06",x"00",x"CB",x"27",x"CB",x"10",x"CB", -- 0x1C60
    x"27",x"CB",x"10",x"E6",x"E0",x"4F",x"21",x"E0", -- 0x1C68
    x"03",x"ED",x"42",x"7C",x"FE",x"04",x"DA",x"7E", -- 0x1C70
    x"1C",x"01",x"0E",x"03",x"ED",x"42",x"ED",x"5B", -- 0x1C78
    x"85",x"40",x"19",x"22",x"89",x"40",x"DD",x"7E", -- 0x1C80
    x"00",x"FD",x"96",x"00",x"ED",x"44",x"C6",x"05", -- 0x1C88
    x"E6",x"07",x"CB",x"27",x"4F",x"06",x"00",x"21", -- 0x1C90
    x"DA",x"2B",x"09",x"22",x"83",x"40",x"3E",x"03", -- 0x1C98
    x"32",x"88",x"40",x"2A",x"89",x"40",x"7E",x"D6", -- 0x1CA0
    x"0A",x"FE",x"06",x"D2",x"42",x"1D",x"CB",x"27", -- 0x1CA8
    x"4F",x"06",x"00",x"21",x"18",x"2C",x"09",x"5E", -- 0x1CB0
    x"23",x"56",x"2A",x"83",x"40",x"3E",x"08",x"47", -- 0x1CB8
    x"32",x"8B",x"40",x"3A",x"87",x"40",x"FE",x"03", -- 0x1CC0
    x"CA",x"FC",x"1C",x"FE",x"02",x"CA",x"1B",x"1D", -- 0x1CC8
    x"23",x"3A",x"82",x"40",x"4F",x"7E",x"06",x"00", -- 0x1CD0
    x"0D",x"CA",x"E3",x"1C",x"CB",x"3F",x"CB",x"18", -- 0x1CD8
    x"C3",x"D8",x"1C",x"EB",x"78",x"AE",x"A0",x"B8", -- 0x1CE0
    x"C2",x"81",x"1D",x"EB",x"23",x"23",x"13",x"3A", -- 0x1CE8
    x"8B",x"40",x"3D",x"32",x"8B",x"40",x"C2",x"D1", -- 0x1CF0
    x"1C",x"C3",x"42",x"1D",x"3A",x"82",x"40",x"4F", -- 0x1CF8
    x"7E",x"0D",x"CA",x"0A",x"1D",x"CB",x"3F",x"C3", -- 0x1D00
    x"01",x"1D",x"EB",x"4F",x"AE",x"A1",x"B9",x"C2", -- 0x1D08
    x"81",x"1D",x"EB",x"23",x"23",x"13",x"10",x"E4", -- 0x1D10
    x"C3",x"42",x"1D",x"3A",x"82",x"40",x"4F",x"7E", -- 0x1D18
    x"23",x"46",x"0D",x"CA",x"2D",x"1D",x"CB",x"3F", -- 0x1D20
    x"CB",x"18",x"C3",x"22",x"1D",x"EB",x"78",x"AE", -- 0x1D28
    x"A0",x"B8",x"C2",x"81",x"1D",x"EB",x"23",x"13", -- 0x1D30
    x"3A",x"8B",x"40",x"3D",x"32",x"8B",x"40",x"C2", -- 0x1D38
    x"1B",x"1D",x"21",x"88",x"40",x"35",x"CA",x"71", -- 0x1D40
    x"1D",x"2A",x"83",x"40",x"01",x"10",x"00",x"09", -- 0x1D48
    x"22",x"83",x"40",x"2A",x"89",x"40",x"7D",x"E6", -- 0x1D50
    x"E0",x"6F",x"7C",x"E6",x"0F",x"B5",x"2A",x"89", -- 0x1D58
    x"40",x"01",x"E0",x"FF",x"C2",x"6A",x"1D",x"01", -- 0x1D60
    x"E0",x"03",x"09",x"22",x"89",x"40",x"C3",x"A6", -- 0x1D68
    x"1C",x"21",x"87",x"40",x"35",x"C8",x"21",x"85", -- 0x1D70
    x"40",x"34",x"FD",x"23",x"FD",x"23",x"C3",x"59", -- 0x1D78
    x"1C",x"2A",x"89",x"40",x"36",x"10",x"3E",x"0C", -- 0x1D80
    x"32",x"08",x"41",x"C9",x"3A",x"1C",x"41",x"FE", -- 0x1D88
    x"02",x"C0",x"21",x"1D",x"41",x"35",x"C0",x"3A", -- 0x1D90
    x"1E",x"41",x"77",x"21",x"A6",x"41",x"34",x"23", -- 0x1D98
    x"23",x"34",x"3A",x"91",x"40",x"FE",x"02",x"C0", -- 0x1DA0
    x"DD",x"34",x"10",x"DD",x"34",x"14",x"C9",x"DD", -- 0x1DA8
    x"21",x"AA",x"41",x"3A",x"91",x"40",x"FE",x"01", -- 0x1DB0
    x"CA",x"21",x"1E",x"FE",x"02",x"CA",x"15",x"1E", -- 0x1DB8
    x"FE",x"03",x"CA",x"FA",x"1D",x"FE",x"04",x"C0", -- 0x1DC0
    x"21",x"90",x"40",x"35",x"C0",x"36",x"04",x"21", -- 0x1DC8
    x"20",x"52",x"11",x"9A",x"40",x"01",x"E0",x"FF", -- 0x1DD0
    x"1A",x"E6",x"0F",x"CA",x"DF",x"1D",x"77",x"09", -- 0x1DD8
    x"1B",x"1A",x"0F",x"0F",x"0F",x"0F",x"E6",x"0F", -- 0x1DE0
    x"00",x"00",x"00",x"77",x"09",x"1A",x"E6",x"0F", -- 0x1DE8
    x"77",x"09",x"36",x"00",x"3E",x"03",x"32",x"91", -- 0x1DF0
    x"40",x"C9",x"21",x"90",x"40",x"35",x"C0",x"36", -- 0x1DF8
    x"04",x"21",x"80",x"52",x"11",x"E0",x"FF",x"06", -- 0x1E00
    x"0A",x"3E",x"10",x"77",x"19",x"10",x"FC",x"3E", -- 0x1E08
    x"04",x"32",x"91",x"40",x"C9",x"DD",x"7E",x"10", -- 0x1E10
    x"FE",x"FF",x"C0",x"3E",x"01",x"32",x"91",x"40", -- 0x1E18
    x"C9",x"21",x"90",x"40",x"35",x"C0",x"CD",x"09", -- 0x1E20
    x"28",x"47",x"3A",x"1F",x"41",x"A0",x"3C",x"77", -- 0x1E28
    x"AF",x"DD",x"77",x"10",x"3E",x"10",x"DD",x"77", -- 0x1E30
    x"14",x"DD",x"36",x"12",x"06",x"DD",x"36",x"16", -- 0x1E38
    x"06",x"DD",x"36",x"13",x"F0",x"DD",x"36",x"17", -- 0x1E40
    x"F0",x"CD",x"09",x"28",x"E6",x"06",x"C2",x"53", -- 0x1E48
    x"1E",x"3C",x"3C",x"C6",x"25",x"DD",x"77",x"11", -- 0x1E50
    x"3C",x"DD",x"77",x"15",x"3E",x"02",x"32",x"91", -- 0x1E58
    x"40",x"C9",x"3A",x"17",x"41",x"FE",x"02",x"CA", -- 0x1E60
    x"70",x"1E",x"FE",x"04",x"CA",x"0E",x"1F",x"C9", -- 0x1E68
    x"DD",x"21",x"EA",x"41",x"FD",x"21",x"A0",x"41", -- 0x1E70
    x"D9",x"11",x"1B",x"50",x"D9",x"06",x"1A",x"3A", -- 0x1E78
    x"1A",x"41",x"4F",x"CD",x"09",x"28",x"E6",x"01", -- 0x1E80
    x"DD",x"77",x"00",x"3A",x"18",x"41",x"90",x"CB", -- 0x1E88
    x"3F",x"DD",x"77",x"02",x"DD",x"77",x"03",x"CD", -- 0x1E90
    x"09",x"28",x"E6",x"07",x"3C",x"3C",x"DD",x"77", -- 0x1E98
    x"05",x"DD",x"36",x"01",x"00",x"DD",x"36",x"04", -- 0x1EA0
    x"00",x"0D",x"C2",x"EE",x"1E",x"CD",x"09",x"28", -- 0x1EA8
    x"E6",x"01",x"4F",x"3A",x"19",x"41",x"81",x"DD", -- 0x1EB0
    x"77",x"04",x"3A",x"1A",x"41",x"4F",x"78",x"FE", -- 0x1EB8
    x"05",x"DA",x"EE",x"1E",x"D9",x"DD",x"46",x"04", -- 0x1EC0
    x"DD",x"70",x"01",x"26",x"00",x"CD",x"09",x"28", -- 0x1EC8
    x"CB",x"27",x"CB",x"14",x"CB",x"27",x"CB",x"14", -- 0x1ED0
    x"E6",x"E0",x"6F",x"19",x"CD",x"09",x"28",x"E6", -- 0x1ED8
    x"07",x"C6",x"0A",x"FE",x"10",x"DA",x"EA",x"1E", -- 0x1EE0
    x"D6",x"02",x"77",x"10",x"DE",x"D9",x"CD",x"09", -- 0x1EE8
    x"28",x"FD",x"77",x"00",x"FD",x"36",x"01",x"06", -- 0x1EF0
    x"FD",x"2B",x"FD",x"2B",x"11",x"06",x"00",x"DD", -- 0x1EF8
    x"19",x"D9",x"1B",x"D9",x"05",x"C2",x"83",x"1E", -- 0x1F00
    x"3E",x"04",x"32",x"17",x"41",x"C9",x"DD",x"21", -- 0x1F08
    x"EA",x"41",x"FD",x"21",x"A0",x"41",x"11",x"1B", -- 0x1F10
    x"50",x"62",x"6B",x"DD",x"35",x"03",x"C2",x"88", -- 0x1F18
    x"1F",x"DD",x"7E",x"02",x"DD",x"77",x"03",x"FD", -- 0x1F20
    x"34",x"00",x"DD",x"CB",x"00",x"46",x"CA",x"37", -- 0x1F28
    x"1F",x"FD",x"35",x"00",x"FD",x"35",x"00",x"FD", -- 0x1F30
    x"7E",x"00",x"E6",x"07",x"C2",x"88",x"1F",x"06", -- 0x1F38
    x"00",x"FD",x"7E",x"00",x"CB",x"27",x"CB",x"10", -- 0x1F40
    x"CB",x"27",x"CB",x"10",x"E6",x"E0",x"4F",x"09", -- 0x1F48
    x"7E",x"36",x"10",x"FE",x"10",x"CA",x"5B",x"1F", -- 0x1F50
    x"DD",x"35",x"01",x"DD",x"7E",x"01",x"DD",x"BE", -- 0x1F58
    x"04",x"D2",x"88",x"1F",x"DD",x"35",x"05",x"C2", -- 0x1F60
    x"88",x"1F",x"CD",x"09",x"28",x"E6",x"07",x"3C", -- 0x1F68
    x"DD",x"77",x"05",x"CD",x"09",x"28",x"0F",x"0F", -- 0x1F70
    x"0F",x"E6",x"07",x"C6",x"0A",x"FE",x"10",x"DA", -- 0x1F78
    x"84",x"1F",x"D6",x"02",x"77",x"DD",x"34",x"01", -- 0x1F80
    x"FD",x"2B",x"FD",x"2B",x"01",x"06",x"00",x"DD", -- 0x1F88
    x"09",x"1B",x"7B",x"FE",x"01",x"C2",x"19",x"1F", -- 0x1F90
    x"C9",x"3A",x"08",x"41",x"FE",x"00",x"C0",x"DD", -- 0x1F98
    x"21",x"AA",x"41",x"DD",x"7E",x"03",x"FE",x"10", -- 0x1FA0
    x"D8",x"DD",x"7E",x"05",x"A7",x"C2",x"E1",x"1F", -- 0x1FA8
    x"3A",x"95",x"40",x"A7",x"C8",x"3A",x"05",x"40", -- 0x1FB0
    x"CB",x"67",x"C8",x"3E",x"05",x"32",x"7A",x"40", -- 0x1FB8
    x"DD",x"36",x"05",x"1B",x"DD",x"36",x"06",x"07", -- 0x1FC0
    x"3E",x"03",x"32",x"6E",x"40",x"DD",x"7E",x"00", -- 0x1FC8
    x"DD",x"77",x"04",x"DD",x"7E",x"03",x"C6",x"0E", -- 0x1FD0
    x"DD",x"77",x"07",x"3E",x"01",x"32",x"03",x"68", -- 0x1FD8
    x"C9",x"3A",x"05",x"40",x"CB",x"67",x"C2",x"F7", -- 0x1FE0
    x"1F",x"21",x"AE",x"41",x"06",x"04",x"AF",x"77", -- 0x1FE8
    x"23",x"10",x"FC",x"32",x"03",x"68",x"C9",x"21", -- 0x1FF0
    x"96",x"40",x"35",x"C2",x"36",x"20",x"36",x"35", -- 0x1FF8
    x"2A",x"97",x"40",x"7E",x"3D",x"FE",x"64",x"C2", -- 0x2000
    x"35",x"20",x"21",x"95",x"40",x"35",x"C2",x"1D", -- 0x2008
    x"20",x"21",x"97",x"29",x"22",x"0C",x"40",x"22", -- 0x2010
    x"0E",x"40",x"C3",x"E9",x"1F",x"7E",x"FE",x"02", -- 0x2018
    x"C2",x"29",x"20",x"11",x"31",x"2A",x"CD",x"1F", -- 0x2020
    x"27",x"2A",x"97",x"40",x"01",x"20",x"00",x"09", -- 0x2028
    x"22",x"97",x"40",x"3E",x"68",x"77",x"DD",x"7E", -- 0x2030
    x"00",x"DD",x"77",x"04",x"DD",x"7E",x"03",x"C6", -- 0x2038
    x"0E",x"DD",x"77",x"07",x"21",x"6E",x"40",x"35", -- 0x2040
    x"C2",x"55",x"20",x"36",x"03",x"DD",x"7E",x"05", -- 0x2048
    x"EE",x"34",x"DD",x"77",x"05",x"21",x"7A",x"40", -- 0x2050
    x"35",x"C0",x"36",x"05",x"3A",x"80",x"40",x"FE", -- 0x2058
    x"01",x"CA",x"6F",x"20",x"3A",x"78",x"40",x"3D", -- 0x2060
    x"3D",x"FE",x"02",x"D8",x"C3",x"82",x"20",x"3A", -- 0x2068
    x"78",x"40",x"3C",x"3C",x"FE",x"12",x"DA",x"82", -- 0x2070
    x"20",x"3A",x"80",x"40",x"EE",x"01",x"32",x"80", -- 0x2078
    x"40",x"C9",x"32",x"78",x"40",x"C9",x"21",x"BA", -- 0x2080
    x"41",x"AF",x"06",x"08",x"77",x"23",x"10",x"FC", -- 0x2088
    x"C9",x"3A",x"92",x"40",x"FE",x"01",x"CA",x"B2", -- 0x2090
    x"21",x"FE",x"03",x"CA",x"B2",x"20",x"FE",x"02", -- 0x2098
    x"C0",x"3A",x"08",x"41",x"FE",x"10",x"C2",x"B2", -- 0x20A0
    x"20",x"AF",x"32",x"94",x"40",x"3E",x"03",x"32", -- 0x20A8
    x"92",x"40",x"DD",x"21",x"C2",x"42",x"FD",x"21", -- 0x20B0
    x"94",x"40",x"21",x"65",x"52",x"06",x"20",x"DD", -- 0x20B8
    x"7E",x"00",x"A7",x"CA",x"EA",x"20",x"DD",x"35", -- 0x20C0
    x"00",x"C2",x"EA",x"20",x"CD",x"09",x"28",x"E6", -- 0x20C8
    x"0E",x"3C",x"DD",x"77",x"00",x"CD",x"09",x"28", -- 0x20D0
    x"DD",x"A6",x"01",x"DD",x"86",x"02",x"FD",x"A6", -- 0x20D8
    x"00",x"C2",x"E9",x"20",x"DD",x"77",x"00",x"3E", -- 0x20E0
    x"10",x"77",x"23",x"78",x"E6",x"03",x"FE",x"01", -- 0x20E8
    x"C2",x"F7",x"20",x"11",x"DC",x"FF",x"19",x"11", -- 0x20F0
    x"03",x"00",x"DD",x"19",x"10",x"C1",x"DD",x"21", -- 0x20F8
    x"AA",x"41",x"21",x"22",x"41",x"35",x"C2",x"22", -- 0x2100
    x"21",x"CD",x"09",x"28",x"E6",x"0F",x"3C",x"77", -- 0x2108
    x"CD",x"09",x"28",x"E6",x"03",x"3C",x"32",x"75", -- 0x2110
    x"41",x"32",x"77",x"41",x"32",x"79",x"41",x"32", -- 0x2118
    x"7B",x"41",x"21",x"23",x"41",x"35",x"C2",x"5C", -- 0x2120
    x"21",x"3A",x"24",x"41",x"77",x"3A",x"9D",x"40", -- 0x2128
    x"FE",x"00",x"C2",x"5C",x"21",x"3A",x"25",x"41", -- 0x2130
    x"A7",x"3A",x"74",x"41",x"CA",x"49",x"21",x"3C", -- 0x2138
    x"DD",x"34",x"18",x"DD",x"34",x"1C",x"C3",x"50", -- 0x2140
    x"21",x"3D",x"DD",x"35",x"18",x"DD",x"35",x"1C", -- 0x2148
    x"32",x"74",x"41",x"32",x"76",x"41",x"32",x"78", -- 0x2150
    x"41",x"32",x"7A",x"41",x"21",x"26",x"41",x"35", -- 0x2158
    x"C2",x"7C",x"21",x"3E",x"30",x"32",x"26",x"41", -- 0x2160
    x"3A",x"A2",x"41",x"D6",x"84",x"47",x"DD",x"7E", -- 0x2168
    x"18",x"90",x"06",x"00",x"D2",x"78",x"21",x"04", -- 0x2170
    x"78",x"32",x"25",x"41",x"3A",x"A2",x"41",x"D6", -- 0x2178
    x"84",x"47",x"DD",x"7E",x"18",x"90",x"06",x"03", -- 0x2180
    x"D2",x"8F",x"21",x"06",x"01",x"ED",x"44",x"FE", -- 0x2188
    x"23",x"D2",x"96",x"21",x"06",x"00",x"3E",x"16", -- 0x2190
    x"A8",x"DD",x"77",x"19",x"3A",x"9D",x"40",x"FE", -- 0x2198
    x"00",x"C0",x"3A",x"08",x"41",x"FE",x"06",x"3E", -- 0x21A0
    x"10",x"CA",x"AE",x"21",x"3E",x"0F",x"DD",x"77", -- 0x21A8
    x"1D",x"C9",x"21",x"93",x"40",x"35",x"C0",x"3E", -- 0x21B0
    x"02",x"32",x"75",x"41",x"32",x"77",x"41",x"32", -- 0x21B8
    x"79",x"41",x"32",x"7B",x"41",x"AF",x"32",x"74", -- 0x21C0
    x"41",x"32",x"76",x"41",x"32",x"78",x"41",x"32", -- 0x21C8
    x"7A",x"41",x"21",x"C2",x"42",x"11",x"54",x"2C", -- 0x21D0
    x"06",x"60",x"1A",x"77",x"23",x"13",x"10",x"FA", -- 0x21D8
    x"DD",x"21",x"AA",x"41",x"DD",x"36",x"18",x"7A", -- 0x21E0
    x"DD",x"36",x"19",x"16",x"DD",x"36",x"1A",x"07", -- 0x21E8
    x"DD",x"36",x"1B",x"30",x"DD",x"36",x"1C",x"7A", -- 0x21F0
    x"DD",x"36",x"1D",x"10",x"DD",x"36",x"1E",x"07", -- 0x21F8
    x"DD",x"36",x"1F",x"34",x"3E",x"10",x"32",x"22", -- 0x2200
    x"41",x"3A",x"24",x"41",x"32",x"23",x"41",x"CD", -- 0x2208
    x"09",x"28",x"E6",x"01",x"32",x"25",x"41",x"3A", -- 0x2210
    x"30",x"00",x"32",x"26",x"41",x"3E",x"FF",x"32", -- 0x2218
    x"94",x"40",x"3E",x"02",x"32",x"92",x"40",x"C9", -- 0x2220
    x"3A",x"08",x"41",x"FE",x"06",x"C0",x"3A",x"92", -- 0x2228
    x"40",x"FE",x"02",x"C0",x"21",x"1D",x"40",x"35", -- 0x2230
    x"C0",x"3A",x"74",x"41",x"47",x"3A",x"A2",x"41", -- 0x2238
    x"90",x"D2",x"46",x"22",x"ED",x"44",x"CB",x"3F", -- 0x2240
    x"CB",x"3F",x"CB",x"3F",x"47",x"CD",x"09",x"28", -- 0x2248
    x"E6",x"0F",x"80",x"3C",x"77",x"3A",x"1E",x"40", -- 0x2250
    x"21",x"27",x"41",x"BE",x"C8",x"3A",x"74",x"41", -- 0x2258
    x"C6",x"6B",x"47",x"CD",x"09",x"28",x"E6",x"2F", -- 0x2260
    x"80",x"21",x"C7",x"41",x"11",x"04",x"00",x"06", -- 0x2268
    x"06",x"19",x"BE",x"CA",x"5D",x"22",x"10",x"F9", -- 0x2270
    x"DD",x"21",x"C6",x"41",x"47",x"DD",x"19",x"DD", -- 0x2278
    x"7E",x"01",x"DD",x"B6",x"03",x"C2",x"7D",x"22", -- 0x2280
    x"DD",x"70",x"01",x"3E",x"B9",x"21",x"1B",x"41", -- 0x2288
    x"AE",x"DD",x"77",x"03",x"21",x"1E",x"40",x"34", -- 0x2290
    x"C9",x"21",x"2C",x"41",x"35",x"C0",x"3A",x"2D", -- 0x2298
    x"41",x"77",x"3A",x"08",x"41",x"FE",x"06",x"C0", -- 0x22A0
    x"3A",x"92",x"40",x"FE",x"02",x"C0",x"21",x"0B", -- 0x22A8
    x"41",x"3A",x"0C",x"41",x"BE",x"D0",x"21",x"29", -- 0x22B0
    x"41",x"BE",x"C8",x"DD",x"21",x"C6",x"41",x"FD", -- 0x22B8
    x"21",x"A6",x"41",x"01",x"24",x"00",x"11",x"04", -- 0x22C0
    x"00",x"DD",x"09",x"FD",x"19",x"DD",x"7E",x"00", -- 0x22C8
    x"FE",x"00",x"C2",x"C9",x"22",x"DD",x"36",x"00", -- 0x22D0
    x"02",x"CD",x"09",x"28",x"E6",x"01",x"DD",x"77", -- 0x22D8
    x"05",x"3A",x"28",x"41",x"DD",x"77",x"06",x"3A", -- 0x22E0
    x"2B",x"41",x"DD",x"77",x"04",x"3A",x"2F",x"41", -- 0x22E8
    x"DD",x"77",x"08",x"CD",x"09",x"28",x"21",x"2A", -- 0x22F0
    x"41",x"A6",x"3C",x"DD",x"77",x"03",x"DD",x"36", -- 0x22F8
    x"01",x"02",x"DD",x"36",x"02",x"01",x"3A",x"2E", -- 0x2300
    x"41",x"DD",x"77",x"07",x"DD",x"36",x"1A",x"07", -- 0x2308
    x"DD",x"36",x"1B",x"08",x"DD",x"36",x"1C",x"08", -- 0x2310
    x"DD",x"36",x"1D",x"0E",x"3A",x"74",x"41",x"C6", -- 0x2318
    x"7A",x"FD",x"77",x"00",x"FD",x"36",x"03",x"38", -- 0x2320
    x"FD",x"36",x"01",x"0B",x"3A",x"75",x"41",x"FD", -- 0x2328
    x"77",x"02",x"21",x"0C",x"41",x"34",x"21",x"CF", -- 0x2330
    x"29",x"22",x"0C",x"40",x"3E",x"01",x"32",x"02", -- 0x2338
    x"40",x"21",x"00",x"00",x"22",x"0E",x"40",x"C9", -- 0x2340
    x"3A",x"0C",x"41",x"A7",x"C8",x"47",x"DD",x"21", -- 0x2348
    x"C6",x"41",x"FD",x"21",x"A6",x"41",x"11",x"24", -- 0x2350
    x"00",x"DD",x"19",x"11",x"04",x"00",x"FD",x"19", -- 0x2358
    x"DD",x"7E",x"00",x"FE",x"00",x"CA",x"56",x"23", -- 0x2360
    x"FE",x"0C",x"C2",x"B5",x"23",x"DD",x"35",x"0A", -- 0x2368
    x"C2",x"F5",x"24",x"DD",x"36",x"0A",x"07",x"FD", -- 0x2370
    x"34",x"01",x"FD",x"7E",x"01",x"FE",x"20",x"C2", -- 0x2378
    x"F5",x"24",x"DD",x"36",x"00",x"00",x"FD",x"36", -- 0x2380
    x"01",x"00",x"FD",x"36",x"00",x"00",x"FD",x"36", -- 0x2388
    x"03",x"00",x"DD",x"7E",x"0D",x"0F",x"0F",x"0F", -- 0x2390
    x"0F",x"E6",x"70",x"CD",x"2B",x"28",x"CD",x"4A", -- 0x2398
    x"28",x"21",x"0C",x"41",x"35",x"2B",x"35",x"7E", -- 0x23A0
    x"FE",x"01",x"C2",x"F5",x"24",x"3E",x"08",x"32", -- 0x23A8
    x"28",x"41",x"C3",x"F5",x"24",x"DD",x"35",x"07", -- 0x23B0
    x"CA",x"C8",x"23",x"21",x"30",x"41",x"3A",x"0B", -- 0x23B8
    x"41",x"BE",x"DA",x"9D",x"24",x"C3",x"F5",x"24", -- 0x23C0
    x"3A",x"2E",x"41",x"DD",x"77",x"07",x"DD",x"7E", -- 0x23C8
    x"00",x"FE",x"05",x"D2",x"FE",x"23",x"DD",x"35", -- 0x23D0
    x"01",x"C2",x"FE",x"23",x"DD",x"36",x"01",x"02", -- 0x23D8
    x"FD",x"7E",x"01",x"DD",x"86",x"02",x"FE",x"0F", -- 0x23E0
    x"D2",x"F0",x"23",x"FE",x"0B",x"D2",x"FB",x"23", -- 0x23E8
    x"DD",x"7E",x"02",x"ED",x"44",x"DD",x"77",x"02", -- 0x23F0
    x"C3",x"E0",x"23",x"FD",x"77",x"01",x"DD",x"35", -- 0x23F8
    x"03",x"C2",x"1F",x"24",x"CD",x"09",x"28",x"21", -- 0x2400
    x"2A",x"41",x"A6",x"3C",x"DD",x"77",x"03",x"FD", -- 0x2408
    x"7E",x"02",x"3C",x"E6",x"03",x"C2",x"19",x"24", -- 0x2410
    x"3C",x"FD",x"77",x"02",x"DD",x"77",x"0D",x"DD", -- 0x2418
    x"7E",x"00",x"FE",x"02",x"C2",x"39",x"24",x"FD", -- 0x2420
    x"35",x"03",x"FD",x"7E",x"03",x"FE",x"10",x"C2", -- 0x2428
    x"9D",x"24",x"DD",x"36",x"00",x"04",x"C3",x"9D", -- 0x2430
    x"24",x"FD",x"34",x"03",x"FD",x"7E",x"03",x"DD", -- 0x2438
    x"BE",x"08",x"DA",x"49",x"24",x"FD",x"34",x"03", -- 0x2440
    x"3C",x"3D",x"FE",x"FE",x"DA",x"5E",x"24",x"3A", -- 0x2448
    x"74",x"41",x"C6",x"7A",x"FD",x"77",x"00",x"DD", -- 0x2450
    x"36",x"00",x"0E",x"C3",x"F5",x"24",x"DD",x"7E", -- 0x2458
    x"00",x"FE",x"04",x"C2",x"7A",x"24",x"FD",x"7E", -- 0x2460
    x"03",x"DD",x"BE",x"04",x"C2",x"7A",x"24",x"FD", -- 0x2468
    x"36",x"01",x"13",x"DD",x"36",x"00",x"10",x"C3", -- 0x2470
    x"9D",x"24",x"DD",x"7E",x"00",x"FE",x"0E",x"C2", -- 0x2478
    x"9D",x"24",x"FD",x"7E",x"03",x"FE",x"38",x"C2", -- 0x2480
    x"F5",x"24",x"DD",x"36",x"00",x"00",x"FD",x"36", -- 0x2488
    x"00",x"00",x"FD",x"36",x"03",x"00",x"21",x"0C", -- 0x2490
    x"41",x"35",x"C3",x"F5",x"24",x"DD",x"7E",x"00", -- 0x2498
    x"FE",x"0E",x"CA",x"F5",x"24",x"3A",x"A2",x"41", -- 0x24A0
    x"C6",x"89",x"4F",x"FD",x"7E",x"00",x"91",x"D2", -- 0x24A8
    x"B4",x"24",x"ED",x"44",x"0F",x"0F",x"0F",x"0F", -- 0x24B0
    x"2F",x"E6",x"03",x"3C",x"DD",x"CB",x"05",x"46", -- 0x24B8
    x"C2",x"C5",x"24",x"ED",x"44",x"FD",x"86",x"00", -- 0x24C0
    x"5F",x"C6",x"1C",x"FE",x"20",x"CB",x"17",x"57", -- 0x24C8
    x"DD",x"AE",x"05",x"DD",x"77",x"05",x"CB",x"42", -- 0x24D0
    x"C2",x"AB",x"24",x"FD",x"73",x"00",x"DD",x"35", -- 0x24D8
    x"06",x"C2",x"F5",x"24",x"3A",x"28",x"41",x"DD", -- 0x24E0
    x"77",x"06",x"FD",x"7E",x"00",x"91",x"CB",x"17", -- 0x24E8
    x"E6",x"01",x"DD",x"77",x"05",x"05",x"C2",x"56", -- 0x24F0
    x"23",x"C9",x"DD",x"21",x"AA",x"41",x"FD",x"21", -- 0x24F8
    x"E6",x"41",x"3A",x"9D",x"40",x"FE",x"01",x"CA", -- 0x2500
    x"16",x"26",x"FE",x"03",x"CA",x"5F",x"26",x"FE", -- 0x2508
    x"02",x"CA",x"36",x"25",x"FE",x"00",x"C0",x"3A", -- 0x2510
    x"0B",x"41",x"A7",x"C0",x"3A",x"08",x"41",x"FE", -- 0x2518
    x"06",x"C0",x"3E",x"20",x"32",x"9E",x"40",x"3E", -- 0x2520
    x"01",x"32",x"9D",x"40",x"AF",x"32",x"94",x"40", -- 0x2528
    x"3E",x"03",x"32",x"92",x"40",x"C9",x"DD",x"7E", -- 0x2530
    x"03",x"FE",x"D8",x"DA",x"53",x"25",x"3A",x"A2", -- 0x2538
    x"41",x"C6",x"83",x"DD",x"96",x"00",x"FE",x"23", -- 0x2540
    x"D2",x"53",x"25",x"3E",x"0C",x"32",x"08",x"41", -- 0x2548
    x"C3",x"7B",x"25",x"DD",x"7E",x"00",x"C6",x"19", -- 0x2550
    x"FD",x"96",x"01",x"FE",x"17",x"D2",x"86",x"25", -- 0x2558
    x"21",x"1B",x"41",x"FD",x"7E",x"03",x"AE",x"DD", -- 0x2560
    x"86",x"03",x"C6",x"10",x"FE",x"08",x"D2",x"86", -- 0x2568
    x"25",x"AF",x"32",x"0D",x"41",x"FD",x"77",x"01", -- 0x2570
    x"FD",x"77",x"03",x"3E",x"20",x"CD",x"2B",x"28", -- 0x2578
    x"CD",x"4A",x"28",x"C3",x"8E",x"25",x"DD",x"7E", -- 0x2580
    x"03",x"FE",x"E0",x"C2",x"B2",x"25",x"3E",x"01", -- 0x2588
    x"32",x"87",x"40",x"32",x"88",x"40",x"3E",x"80", -- 0x2590
    x"32",x"9F",x"40",x"21",x"EF",x"29",x"22",x"0C", -- 0x2598
    x"40",x"21",x"00",x"00",x"22",x"0E",x"40",x"3E", -- 0x25A0
    x"01",x"32",x"02",x"40",x"3E",x"03",x"32",x"9D", -- 0x25A8
    x"40",x"C9",x"DD",x"34",x"03",x"DD",x"34",x"07", -- 0x25B0
    x"DD",x"34",x"1B",x"3A",x"A2",x"41",x"C6",x"70", -- 0x25B8
    x"4F",x"DD",x"7E",x"00",x"91",x"D2",x"CA",x"25", -- 0x25C0
    x"ED",x"44",x"0F",x"0F",x"0F",x"0F",x"E6",x"03", -- 0x25C8
    x"3C",x"3C",x"21",x"72",x"40",x"CB",x"46",x"C2", -- 0x25D0
    x"DC",x"25",x"ED",x"44",x"DD",x"86",x"00",x"5F", -- 0x25D8
    x"C6",x"40",x"FE",x"40",x"CB",x"17",x"47",x"AE", -- 0x25E0
    x"77",x"CB",x"40",x"C2",x"C1",x"25",x"DD",x"73", -- 0x25E8
    x"00",x"3E",x"0F",x"83",x"DD",x"77",x"04",x"3E", -- 0x25F0
    x"07",x"83",x"DD",x"77",x"18",x"21",x"73",x"40", -- 0x25F8
    x"35",x"C0",x"CD",x"09",x"28",x"E6",x"1F",x"C6", -- 0x2600
    x"20",x"77",x"DD",x"7E",x"00",x"91",x"CB",x"17", -- 0x2608
    x"E6",x"01",x"32",x"72",x"40",x"C9",x"21",x"9E", -- 0x2610
    x"40",x"35",x"C0",x"DD",x"7E",x"18",x"D6",x"0F", -- 0x2618
    x"DD",x"77",x"00",x"C6",x"07",x"DD",x"77",x"04", -- 0x2620
    x"DD",x"36",x"03",x"30",x"DD",x"36",x"07",x"30", -- 0x2628
    x"DD",x"36",x"01",x"2D",x"DD",x"36",x"05",x"2E", -- 0x2630
    x"DD",x"36",x"02",x"07",x"DD",x"36",x"06",x"07", -- 0x2638
    x"DD",x"36",x"1C",x"00",x"DD",x"36",x"1F",x"00", -- 0x2640
    x"21",x"A9",x"2A",x"22",x"0C",x"40",x"21",x"00", -- 0x2648
    x"00",x"22",x"0E",x"40",x"3E",x"01",x"32",x"02", -- 0x2650
    x"40",x"3E",x"02",x"32",x"9D",x"40",x"C9",x"21", -- 0x2658
    x"9F",x"40",x"35",x"CA",x"93",x"26",x"21",x"87", -- 0x2660
    x"40",x"35",x"C2",x"7E",x"26",x"CD",x"09",x"28", -- 0x2668
    x"E6",x"0F",x"3C",x"77",x"CD",x"09",x"28",x"E6", -- 0x2670
    x"03",x"C6",x"0B",x"DD",x"77",x"01",x"23",x"35", -- 0x2678
    x"C0",x"CD",x"09",x"28",x"E6",x"0F",x"3C",x"77", -- 0x2680
    x"CD",x"09",x"28",x"E6",x"03",x"C6",x"0B",x"DD", -- 0x2688
    x"77",x"05",x"C9",x"DD",x"36",x"00",x"00",x"DD", -- 0x2690
    x"36",x"04",x"00",x"DD",x"36",x"03",x"00",x"DD", -- 0x2698
    x"36",x"07",x"00",x"DD",x"36",x"18",x"00",x"DD", -- 0x26A0
    x"36",x"1B",x"00",x"3E",x"04",x"32",x"9D",x"40", -- 0x26A8
    x"C9",x"21",x"AA",x"41",x"AF",x"06",x"40",x"77", -- 0x26B0
    x"23",x"10",x"FC",x"32",x"0C",x"41",x"32",x"0D", -- 0x26B8
    x"41",x"32",x"1E",x"40",x"32",x"00",x"68",x"32", -- 0x26C0
    x"01",x"68",x"32",x"02",x"68",x"21",x"EA",x"41", -- 0x26C8
    x"01",x"20",x"01",x"36",x"00",x"23",x"0B",x"78", -- 0x26D0
    x"B1",x"C2",x"D3",x"26",x"21",x"24",x"40",x"06", -- 0x26D8
    x"40",x"36",x"00",x"23",x"10",x"FB",x"C9",x"01", -- 0x26E0
    x"20",x"00",x"1A",x"FE",x"FF",x"C8",x"FE",x"20", -- 0x26E8
    x"CA",x"F6",x"26",x"D6",x"30",x"77",x"ED",x"42", -- 0x26F0
    x"13",x"C3",x"EA",x"26",x"21",x"02",x"50",x"06", -- 0x26F8
    x"20",x"36",x"10",x"23",x"7D",x"E6",x"1F",x"C2", -- 0x2700
    x"01",x"27",x"23",x"23",x"3A",x"00",x"78",x"10", -- 0x2708
    x"F0",x"C9",x"3E",x"FF",x"32",x"00",x"78",x"AF", -- 0x2710
    x"32",x"06",x"68",x"32",x"07",x"68",x"C9",x"C5", -- 0x2718
    x"2A",x"0C",x"40",x"01",x"EF",x"29",x"ED",x"42", -- 0x2720
    x"C1",x"DA",x"31",x"27",x"ED",x"53",x"0C",x"40", -- 0x2728
    x"C9",x"2A",x"0C",x"40",x"22",x"0E",x"40",x"ED", -- 0x2730
    x"53",x"0C",x"40",x"3E",x"01",x"32",x"02",x"40", -- 0x2738
    x"C9",x"21",x"00",x"41",x"01",x"6A",x"00",x"3A", -- 0x2740
    x"00",x"40",x"FE",x"04",x"C2",x"55",x"27",x"21", -- 0x2748
    x"06",x"41",x"01",x"64",x"00",x"36",x"00",x"23", -- 0x2750
    x"0B",x"78",x"B1",x"C2",x"55",x"27",x"C9",x"3A", -- 0x2758
    x"10",x"41",x"32",x"20",x"40",x"21",x"06",x"41", -- 0x2760
    x"11",x"38",x"41",x"01",x"32",x"00",x"7E",x"08", -- 0x2768
    x"1A",x"77",x"08",x"12",x"23",x"13",x"0B",x"78", -- 0x2770
    x"B1",x"C2",x"6E",x"27",x"C9",x"FD",x"7E",x"00", -- 0x2778
    x"FE",x"80",x"1E",x"55",x"D2",x"89",x"27",x"1E", -- 0x2780
    x"00",x"ED",x"5F",x"E6",x"01",x"7B",x"CA",x"93", -- 0x2788
    x"27",x"F6",x"AA",x"DD",x"A6",x"22",x"DD",x"77", -- 0x2790
    x"0C",x"21",x"BA",x"2B",x"DD",x"7E",x"22",x"FE", -- 0x2798
    x"FF",x"C2",x"AA",x"27",x"DD",x"35",x"11",x"C2", -- 0x27A0
    x"C3",x"27",x"21",x"CA",x"2B",x"DD",x"7E",x"0C", -- 0x27A8
    x"E6",x"55",x"DD",x"77",x"0C",x"DD",x"36",x"22", -- 0x27B0
    x"55",x"DD",x"7E",x"11",x"0F",x"DA",x"C3",x"27", -- 0x27B8
    x"DD",x"77",x"11",x"ED",x"5F",x"E6",x"0C",x"5F", -- 0x27C0
    x"16",x"00",x"19",x"5E",x"23",x"56",x"23",x"1A", -- 0x27C8
    x"DD",x"AE",x"0C",x"DD",x"73",x"07",x"DD",x"72", -- 0x27D0
    x"08",x"DD",x"77",x"09",x"5E",x"23",x"56",x"DD", -- 0x27D8
    x"73",x"01",x"DD",x"72",x"02",x"1A",x"0F",x"0F", -- 0x27E0
    x"0F",x"0F",x"E6",x"0F",x"DD",x"77",x"03",x"DD", -- 0x27E8
    x"77",x"05",x"1A",x"E6",x"0F",x"DD",x"77",x"04", -- 0x27F0
    x"DD",x"77",x"06",x"DD",x"36",x"0A",x"04",x"ED", -- 0x27F8
    x"5F",x"E6",x"1F",x"C6",x"08",x"DD",x"77",x"0B", -- 0x2800
    x"C9",x"E5",x"2A",x"8C",x"40",x"23",x"7C",x"E6", -- 0x2808
    x"1F",x"67",x"22",x"8C",x"40",x"7E",x"E1",x"C9", -- 0x2810
    x"D9",x"4F",x"3A",x"00",x"40",x"FE",x"04",x"CA", -- 0x2818
    x"48",x"28",x"79",x"2A",x"0E",x"41",x"23",x"86", -- 0x2820
    x"C3",x"40",x"28",x"D9",x"4F",x"3A",x"00",x"40", -- 0x2828
    x"FE",x"04",x"79",x"CA",x"48",x"28",x"2A",x"0E", -- 0x2830
    x"41",x"86",x"27",x"77",x"23",x"7E",x"CE",x"00", -- 0x2838
    x"27",x"77",x"23",x"7E",x"CE",x"00",x"27",x"77", -- 0x2840
    x"D9",x"C9",x"3A",x"21",x"41",x"A7",x"C8",x"3A", -- 0x2848
    x"00",x"40",x"FE",x"04",x"C8",x"2A",x"0E",x"41", -- 0x2850
    x"23",x"23",x"7E",x"A7",x"C2",x"66",x"28",x"2B", -- 0x2858
    x"7E",x"21",x"68",x"40",x"BE",x"D8",x"3A",x"00", -- 0x2860
    x"40",x"FE",x"18",x"21",x"60",x"50",x"CA",x"74", -- 0x2868
    x"28",x"21",x"A0",x"53",x"34",x"21",x"10",x"41", -- 0x2870
    x"34",x"AF",x"32",x"21",x"41",x"11",x"CB",x"2A", -- 0x2878
    x"CD",x"1F",x"27",x"C9",x"C9",x"8F",x"28",x"BB", -- 0x2880
    x"28",x"E7",x"28",x"13",x"29",x"3F",x"29",x"B2", -- 0x2888
    x"10",x"F7",x"10",x"72",x"11",x"31",x"11",x"4B", -- 0x2890
    x"12",x"4B",x"12",x"4B",x"12",x"4F",x"13",x"4F", -- 0x2898
    x"13",x"4F",x"13",x"72",x"11",x"72",x"11",x"72", -- 0x28A0
    x"11",x"83",x"13",x"83",x"13",x"83",x"13",x"D3", -- 0x28A8
    x"13",x"D3",x"13",x"D3",x"13",x"02",x"14",x"02", -- 0x28B0
    x"14",x"02",x"14",x"00",x"00",x"00",x"00",x"00", -- 0x28B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C0
    x"00",x"B3",x"14",x"B3",x"14",x"B3",x"14",x"27", -- 0x28C8
    x"15",x"27",x"15",x"27",x"15",x"83",x"13",x"83", -- 0x28D0
    x"13",x"83",x"13",x"00",x"00",x"00",x"00",x"00", -- 0x28D8
    x"00",x"02",x"14",x"02",x"14",x"02",x"14",x"B2", -- 0x28E0
    x"10",x"F7",x"10",x"73",x"17",x"31",x"11",x"4B", -- 0x28E8
    x"12",x"4B",x"12",x"4B",x"12",x"6F",x"15",x"6F", -- 0x28F0
    x"15",x"6F",x"15",x"73",x"17",x"73",x"17",x"73", -- 0x28F8
    x"17",x"83",x"13",x"83",x"13",x"83",x"13",x"DE", -- 0x2900
    x"13",x"DE",x"13",x"DE",x"13",x"02",x"14",x"02", -- 0x2908
    x"14",x"02",x"14",x"B2",x"10",x"F7",x"10",x"72", -- 0x2910
    x"11",x"31",x"11",x"4B",x"12",x"4B",x"12",x"4B", -- 0x2918
    x"12",x"81",x"16",x"81",x"16",x"81",x"16",x"C2", -- 0x2920
    x"17",x"C2",x"17",x"C2",x"17",x"83",x"13",x"83", -- 0x2928
    x"13",x"83",x"13",x"4B",x"17",x"4B",x"17",x"4B", -- 0x2930
    x"17",x"02",x"14",x"02",x"14",x"02",x"14",x"B2", -- 0x2938
    x"10",x"F7",x"10",x"72",x"11",x"31",x"11",x"4B", -- 0x2940
    x"12",x"4B",x"12",x"4B",x"12",x"A4",x"15",x"A4", -- 0x2948
    x"15",x"A4",x"15",x"2F",x"16",x"2F",x"16",x"2F", -- 0x2950
    x"16",x"83",x"13",x"83",x"13",x"83",x"13",x"FF", -- 0x2958
    x"15",x"FF",x"15",x"FF",x"15",x"02",x"14",x"02", -- 0x2960
    x"14",x"02",x"14",x"5E",x"4D",x"7C",x"88",x"5E", -- 0x2968
    x"88",x"4A",x"7A",x"4A",x"72",x"4A",x"60",x"7C", -- 0x2970
    x"A6",x"5E",x"88",x"4A",x"7A",x"4A",x"72",x"4A", -- 0x2978
    x"60",x"7C",x"A6",x"5E",x"88",x"4A",x"7A",x"4A", -- 0x2980
    x"72",x"4A",x"7A",x"7C",x"60",x"4F",x"11",x"47", -- 0x2988
    x"FF",x"47",x"11",x"7C",x"4D",x"7C",x"4D",x"00", -- 0x2990
    x"FE",x"41",x"8F",x"41",x"A1",x"41",x"8F",x"41", -- 0x2998
    x"A1",x"41",x"8F",x"41",x"A1",x"05",x"FF",x"41", -- 0x29A0
    x"8F",x"41",x"A1",x"41",x"8F",x"41",x"A1",x"41", -- 0x29A8
    x"8F",x"41",x"A1",x"05",x"FF",x"41",x"8F",x"41", -- 0x29B0
    x"A1",x"41",x"8F",x"41",x"A1",x"41",x"8F",x"41", -- 0x29B8
    x"A1",x"41",x"FD",x"8F",x"A1",x"41",x"FC",x"01", -- 0x29C0
    x"A6",x"41",x"FC",x"FF",x"00",x"00",x"FE",x"C4", -- 0x29C8
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C2",x"FF",x"C4", -- 0x29D0
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C2",x"FF",x"C4", -- 0x29D8
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C1",x"FD",x"E5", -- 0x29E0
    x"D8",x"C1",x"FC",x"FF",x"30",x"00",x"FE",x"C2", -- 0x29E8
    x"1E",x"C2",x"57",x"C2",x"81",x"C2",x"2B",x"C2", -- 0x29F0
    x"60",x"C2",x"88",x"C2",x"37",x"C2",x"69",x"C2", -- 0x29F8
    x"8F",x"00",x"FE",x"C4",x"DC",x"C3",x"D6",x"C2", -- 0x2A00
    x"E5",x"C1",x"E1",x"00",x"FE",x"C2",x"A6",x"C4", -- 0x2A08
    x"B9",x"C2",x"A6",x"C4",x"1E",x"C2",x"A6",x"C4", -- 0x2A10
    x"B9",x"C2",x"A6",x"00",x"FE",x"43",x"11",x"42", -- 0x2A18
    x"1E",x"42",x"11",x"C3",x"4D",x"41",x"37",x"42", -- 0x2A20
    x"81",x"42",x"11",x"C2",x"60",x"43",x"1E",x"00", -- 0x2A28
    x"FE",x"44",x"FB",x"1E",x"11",x"44",x"FA",x"42", -- 0x2A30
    x"4D",x"42",x"7A",x"6C",x"95",x"56",x"95",x"42", -- 0x2A38
    x"69",x"42",x"7A",x"56",x"95",x"42",x"60",x"42", -- 0x2A40
    x"7A",x"56",x"9B",x"42",x"60",x"42",x"7A",x"6C", -- 0x2A48
    x"9B",x"42",x"4D",x"42",x"7A",x"56",x"95",x"42", -- 0x2A50
    x"60",x"42",x"7A",x"61",x"9B",x"42",x"7A",x"4B", -- 0x2A58
    x"95",x"42",x"72",x"56",x"88",x"42",x"60",x"56", -- 0x2A60
    x"7A",x"42",x"4D",x"6C",x"72",x"56",x"72",x"42", -- 0x2A68
    x"72",x"56",x"88",x"42",x"7A",x"42",x"95",x"6C", -- 0x2A70
    x"A6",x"42",x"4D",x"42",x"72",x"6C",x"9B",x"42", -- 0x2A78
    x"7A",x"4B",x"95",x"4B",x"7A",x"42",x"72",x"4B", -- 0x2A80
    x"9B",x"4B",x"88",x"42",x"7A",x"42",x"95",x"56", -- 0x2A88
    x"A6",x"42",x"60",x"42",x"7A",x"56",x"9B",x"42", -- 0x2A90
    x"4D",x"42",x"7A",x"6C",x"95",x"42",x"4D",x"42", -- 0x2A98
    x"72",x"6C",x"88",x"6C",x"7A",x"6C",x"7A",x"00", -- 0x2AA0
    x"FE",x"41",x"FD",x"69",x"72",x"41",x"FC",x"FF", -- 0x2AA8
    x"57",x"41",x"FD",x"42",x"57",x"41",x"FC",x"01", -- 0x2AB0
    x"88",x"41",x"FD",x"95",x"88",x"41",x"FC",x"FF", -- 0x2AB8
    x"1E",x"41",x"FD",x"1E",x"11",x"41",x"FC",x"01", -- 0x2AC0
    x"E5",x"00",x"FE",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x2AC8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x2AD0
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x2AD8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x2AE0
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x2AE8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"00",x"FE",x"F0", -- 0x2AF0
    x"41",x"41",x"53",x"53",x"FF",x"53",x"31",x"F0", -- 0x2AF8
    x"43",x"35",x"0F",x"12",x"12",x"12",x"54",x"52", -- 0x2B00
    x"51",x"F0",x"41",x"35",x"0F",x"15",x"35",x"FF", -- 0x2B08
    x"53",x"53",x"52",x"F0",x"52",x"53",x"41",x"00", -- 0x2B10
    x"FF",x"FF",x"57",x"00",x"80",x"FA",x"FF",x"57", -- 0x2B18
    x"32",x"32",x"32",x"32",x"32",x"32",x"F0",x"21", -- 0x2B20
    x"FF",x"12",x"0F",x"12",x"FF",x"21",x"F0",x"21", -- 0x2B28
    x"FF",x"12",x"0F",x"12",x"FF",x"21",x"F0",x"32", -- 0x2B30
    x"32",x"32",x"32",x"32",x"32",x"00",x"FF",x"7F", -- 0x2B38
    x"15",x"80",x"EA",x"7F",x"55",x"01",x"FF",x"FF", -- 0x2B40
    x"FF",x"21",x"21",x"F0",x"F0",x"21",x"0F",x"21", -- 0x2B48
    x"0F",x"FF",x"FF",x"00",x"FF",x"FF",x"EB",x"03", -- 0x2B50
    x"53",x"73",x"F0",x"52",x"FF",x"27",x"0F",x"0F", -- 0x2B58
    x"0F",x"0F",x"37",x"45",x"00",x"5F",x"D5",x"FF", -- 0x2B60
    x"18",x"2B",x"F7",x"2A",x"54",x"2B",x"46",x"2B", -- 0x2B68
    x"3E",x"2B",x"20",x"2B",x"65",x"2B",x"58",x"2B", -- 0x2B70
    x"52",x"31",x"51",x"61",x"F0",x"F0",x"61",x"51", -- 0x2B78
    x"31",x"52",x"00",x"FF",x"5F",x"05",x"53",x"21", -- 0x2B80
    x"52",x"F0",x"52",x"21",x"53",x"F0",x"52",x"21", -- 0x2B88
    x"53",x"00",x"FF",x"55",x"15",x"12",x"23",x"FF", -- 0x2B90
    x"21",x"41",x"F0",x"F0",x"41",x"21",x"FF",x"23", -- 0x2B98
    x"12",x"25",x"13",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x2BA0
    x"FF",x"FF",x"FF",x"0F",x"FF",x"FF",x"12",x"12", -- 0x2BA8
    x"FF",x"21",x"F0",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x2BB0
    x"FF",x"0F",x"83",x"2B",x"78",x"2B",x"92",x"2B", -- 0x2BB8
    x"86",x"2B",x"83",x"2B",x"78",x"2B",x"92",x"2B", -- 0x2BC0
    x"86",x"2B",x"A7",x"2B",x"95",x"2B",x"B7",x"2B", -- 0x2BC8
    x"AC",x"2B",x"A7",x"2B",x"95",x"2B",x"B7",x"2B", -- 0x2BD0
    x"AC",x"2B",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE0
    x"00",x"7E",x"00",x"FC",x"01",x"F8",x"03",x"F1", -- 0x2BE8
    x"1F",x"F3",x"3F",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x2BF0
    x"1F",x"F3",x"03",x"F1",x"01",x"F8",x"00",x"FC", -- 0x2BF8
    x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C10
    x"2C",x"2C",x"3C",x"2C",x"24",x"2C",x"44",x"2C", -- 0x2C18
    x"4C",x"2C",x"34",x"2C",x"76",x"7F",x"7F",x"FE", -- 0x2C20
    x"FE",x"FF",x"7F",x"3A",x"00",x"00",x"1C",x"1E", -- 0x2C28
    x"3F",x"3F",x"3E",x"1E",x"38",x"7C",x"7C",x"FC", -- 0x2C30
    x"FC",x"78",x"00",x"00",x"40",x"E0",x"E0",x"60", -- 0x2C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38", -- 0x2C40
    x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C48
    x"02",x"07",x"07",x"02",x"00",x"00",x"00",x"2E", -- 0x2C50
    x"0C",x"2E",x"40",x"0C",x"2F",x"00",x"00",x"00", -- 0x2C58
    x"18",x"0C",x"2E",x"26",x"03",x"44",x"10",x"03", -- 0x2C60
    x"44",x"2A",x"0C",x"2F",x"22",x"03",x"44",x"10", -- 0x2C68
    x"03",x"44",x"2E",x"03",x"44",x"14",x"03",x"44", -- 0x2C70
    x"0C",x"03",x"44",x"02",x"03",x"44",x"04",x"03", -- 0x2C78
    x"44",x"0E",x"03",x"44",x"18",x"03",x"44",x"06", -- 0x2C80
    x"03",x"44",x"08",x"03",x"44",x"12",x"03",x"44", -- 0x2C88
    x"30",x"03",x"44",x"16",x"03",x"44",x"24",x"03", -- 0x2C90
    x"44",x"26",x"03",x"44",x"2C",x"0C",x"2C",x"0E", -- 0x2C98
    x"03",x"44",x"2C",x"03",x"44",x"40",x"0C",x"2D", -- 0x2CA0
    x"00",x"00",x"00",x"32",x"0C",x"2C",x"30",x"0C", -- 0x2CA8
    x"2D",x"00",x"00",x"00",x"38",x"7C",x"7C",x"FC", -- 0x2CB0
    x"FC",x"78",x"00",x"00",x"40",x"E0",x"E0",x"60", -- 0x2CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38", -- 0x2CC0
    x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC8
    x"02",x"07",x"07",x"02",x"00",x"00",x"00",x"2E", -- 0x2CD0
    x"0C",x"2E",x"40",x"0C",x"2F",x"00",x"00",x"00", -- 0x2CD8
    x"18",x"0C",x"2E",x"26",x"03",x"44",x"10",x"03", -- 0x2CE0
    x"44",x"2A",x"0C",x"2F",x"22",x"03",x"44",x"10", -- 0x2CE8
    x"03",x"44",x"2E",x"03",x"44",x"14",x"03",x"44", -- 0x2CF0
    x"0C",x"03",x"44",x"02",x"03",x"44",x"04",x"03", -- 0x2CF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF8
    x"5F",x"E6",x"1F",x"C6",x"08",x"DD",x"77",x"0B", -- 0x3000
    x"C9",x"E5",x"2A",x"8C",x"40",x"23",x"7C",x"E6", -- 0x3008
    x"1F",x"67",x"22",x"8C",x"40",x"7E",x"E1",x"C9", -- 0x3010
    x"D9",x"4F",x"3A",x"00",x"40",x"FE",x"04",x"CA", -- 0x3018
    x"48",x"28",x"79",x"2A",x"0E",x"41",x"23",x"86", -- 0x3020
    x"C3",x"40",x"28",x"D9",x"4F",x"3A",x"00",x"40", -- 0x3028
    x"FE",x"04",x"79",x"CA",x"48",x"28",x"2A",x"0E", -- 0x3030
    x"41",x"86",x"27",x"77",x"23",x"7E",x"CE",x"00", -- 0x3038
    x"27",x"77",x"23",x"7E",x"CE",x"00",x"27",x"77", -- 0x3040
    x"D9",x"C9",x"3A",x"21",x"41",x"A7",x"C8",x"3A", -- 0x3048
    x"00",x"40",x"FE",x"04",x"C8",x"2A",x"0E",x"41", -- 0x3050
    x"23",x"23",x"7E",x"A7",x"C2",x"66",x"28",x"2B", -- 0x3058
    x"7E",x"21",x"68",x"40",x"BE",x"D8",x"3A",x"00", -- 0x3060
    x"40",x"FE",x"18",x"21",x"60",x"50",x"CA",x"74", -- 0x3068
    x"28",x"21",x"A0",x"53",x"34",x"21",x"10",x"41", -- 0x3070
    x"34",x"AF",x"32",x"21",x"41",x"11",x"CB",x"2A", -- 0x3078
    x"CD",x"1F",x"27",x"C9",x"C9",x"8F",x"28",x"BB", -- 0x3080
    x"28",x"E7",x"28",x"13",x"29",x"3F",x"29",x"B2", -- 0x3088
    x"10",x"F7",x"10",x"72",x"11",x"31",x"11",x"4B", -- 0x3090
    x"12",x"4B",x"12",x"4B",x"12",x"4F",x"13",x"4F", -- 0x3098
    x"13",x"4F",x"13",x"72",x"11",x"72",x"11",x"72", -- 0x30A0
    x"11",x"83",x"13",x"83",x"13",x"83",x"13",x"D3", -- 0x30A8
    x"13",x"D3",x"13",x"D3",x"13",x"02",x"14",x"02", -- 0x30B0
    x"14",x"02",x"14",x"00",x"00",x"00",x"00",x"00", -- 0x30B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C0
    x"00",x"B3",x"14",x"B3",x"14",x"B3",x"14",x"27", -- 0x30C8
    x"15",x"27",x"15",x"27",x"15",x"83",x"13",x"83", -- 0x30D0
    x"13",x"83",x"13",x"00",x"00",x"00",x"00",x"00", -- 0x30D8
    x"00",x"02",x"14",x"02",x"14",x"02",x"14",x"B2", -- 0x30E0
    x"10",x"F7",x"10",x"73",x"17",x"31",x"11",x"4B", -- 0x30E8
    x"12",x"4B",x"12",x"4B",x"12",x"6F",x"15",x"6F", -- 0x30F0
    x"15",x"6F",x"15",x"73",x"17",x"73",x"17",x"73", -- 0x30F8
    x"17",x"83",x"13",x"83",x"13",x"83",x"13",x"DE", -- 0x3100
    x"13",x"DE",x"13",x"DE",x"13",x"02",x"14",x"02", -- 0x3108
    x"14",x"02",x"14",x"B2",x"10",x"F7",x"10",x"72", -- 0x3110
    x"11",x"31",x"11",x"4B",x"12",x"4B",x"12",x"4B", -- 0x3118
    x"12",x"81",x"16",x"81",x"16",x"81",x"16",x"C2", -- 0x3120
    x"17",x"C2",x"17",x"C2",x"17",x"83",x"13",x"83", -- 0x3128
    x"13",x"83",x"13",x"4B",x"17",x"4B",x"17",x"4B", -- 0x3130
    x"17",x"02",x"14",x"02",x"14",x"02",x"14",x"B2", -- 0x3138
    x"10",x"F7",x"10",x"72",x"11",x"31",x"11",x"4B", -- 0x3140
    x"12",x"4B",x"12",x"4B",x"12",x"A4",x"15",x"A4", -- 0x3148
    x"15",x"A4",x"15",x"2F",x"16",x"2F",x"16",x"2F", -- 0x3150
    x"16",x"83",x"13",x"83",x"13",x"83",x"13",x"FF", -- 0x3158
    x"15",x"FF",x"15",x"FF",x"15",x"02",x"14",x"02", -- 0x3160
    x"14",x"02",x"14",x"5E",x"4D",x"7C",x"88",x"5E", -- 0x3168
    x"88",x"4A",x"7A",x"4A",x"72",x"4A",x"60",x"7C", -- 0x3170
    x"A6",x"5E",x"88",x"4A",x"7A",x"4A",x"72",x"4A", -- 0x3178
    x"60",x"7C",x"A6",x"5E",x"88",x"4A",x"7A",x"4A", -- 0x3180
    x"72",x"4A",x"7A",x"7C",x"60",x"4F",x"11",x"47", -- 0x3188
    x"FF",x"47",x"11",x"7C",x"4D",x"7C",x"4D",x"00", -- 0x3190
    x"FE",x"41",x"8F",x"41",x"A1",x"41",x"8F",x"41", -- 0x3198
    x"A1",x"41",x"8F",x"41",x"A1",x"05",x"FF",x"41", -- 0x31A0
    x"8F",x"41",x"A1",x"41",x"8F",x"41",x"A1",x"41", -- 0x31A8
    x"8F",x"41",x"A1",x"05",x"FF",x"41",x"8F",x"41", -- 0x31B0
    x"A1",x"41",x"8F",x"41",x"A1",x"41",x"8F",x"41", -- 0x31B8
    x"A1",x"41",x"FD",x"8F",x"A1",x"41",x"FC",x"01", -- 0x31C0
    x"A6",x"41",x"FC",x"FF",x"00",x"00",x"FE",x"C4", -- 0x31C8
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C2",x"FF",x"C4", -- 0x31D0
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C2",x"FF",x"C4", -- 0x31D8
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C1",x"FD",x"E5", -- 0x31E0
    x"D8",x"C1",x"FC",x"FF",x"30",x"00",x"FE",x"C2", -- 0x31E8
    x"1E",x"C2",x"57",x"C2",x"81",x"C2",x"2B",x"C2", -- 0x31F0
    x"60",x"C2",x"88",x"C2",x"37",x"C2",x"69",x"C2", -- 0x31F8
    x"8F",x"00",x"FE",x"C4",x"DC",x"C3",x"D6",x"C2", -- 0x3200
    x"E5",x"C1",x"E1",x"00",x"FE",x"C2",x"A6",x"C4", -- 0x3208
    x"B9",x"C2",x"A6",x"C4",x"1E",x"C2",x"A6",x"C4", -- 0x3210
    x"B9",x"C2",x"A6",x"00",x"FE",x"43",x"11",x"42", -- 0x3218
    x"1E",x"42",x"11",x"C3",x"4D",x"41",x"37",x"42", -- 0x3220
    x"81",x"42",x"11",x"C2",x"60",x"43",x"1E",x"00", -- 0x3228
    x"FE",x"44",x"FB",x"1E",x"11",x"44",x"FA",x"42", -- 0x3230
    x"4D",x"42",x"7A",x"6C",x"95",x"56",x"95",x"42", -- 0x3238
    x"69",x"42",x"7A",x"56",x"95",x"42",x"60",x"42", -- 0x3240
    x"7A",x"56",x"9B",x"42",x"60",x"42",x"7A",x"6C", -- 0x3248
    x"9B",x"42",x"4D",x"42",x"7A",x"56",x"95",x"42", -- 0x3250
    x"60",x"42",x"7A",x"61",x"9B",x"42",x"7A",x"4B", -- 0x3258
    x"95",x"42",x"72",x"56",x"88",x"42",x"60",x"56", -- 0x3260
    x"7A",x"42",x"4D",x"6C",x"72",x"56",x"72",x"42", -- 0x3268
    x"72",x"56",x"88",x"42",x"7A",x"42",x"95",x"6C", -- 0x3270
    x"A6",x"42",x"4D",x"42",x"72",x"6C",x"9B",x"42", -- 0x3278
    x"7A",x"4B",x"95",x"4B",x"7A",x"42",x"72",x"4B", -- 0x3280
    x"9B",x"4B",x"88",x"42",x"7A",x"42",x"95",x"56", -- 0x3288
    x"A6",x"42",x"60",x"42",x"7A",x"56",x"9B",x"42", -- 0x3290
    x"4D",x"42",x"7A",x"6C",x"95",x"42",x"4D",x"42", -- 0x3298
    x"72",x"6C",x"88",x"6C",x"7A",x"6C",x"7A",x"00", -- 0x32A0
    x"FE",x"41",x"FD",x"69",x"72",x"41",x"FC",x"FF", -- 0x32A8
    x"57",x"41",x"FD",x"42",x"57",x"41",x"FC",x"01", -- 0x32B0
    x"88",x"41",x"FD",x"95",x"88",x"41",x"FC",x"FF", -- 0x32B8
    x"1E",x"41",x"FD",x"1E",x"11",x"41",x"FC",x"01", -- 0x32C0
    x"E5",x"00",x"FE",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x32C8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x32D0
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x32D8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x32E0
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x32E8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"00",x"FE",x"F0", -- 0x32F0
    x"41",x"41",x"53",x"53",x"FF",x"53",x"31",x"F0", -- 0x32F8
    x"43",x"35",x"0F",x"12",x"12",x"12",x"54",x"52", -- 0x3300
    x"51",x"F0",x"41",x"35",x"0F",x"15",x"35",x"FF", -- 0x3308
    x"53",x"53",x"52",x"F0",x"52",x"53",x"41",x"00", -- 0x3310
    x"FF",x"FF",x"57",x"00",x"80",x"FA",x"FF",x"57", -- 0x3318
    x"32",x"32",x"32",x"32",x"32",x"32",x"F0",x"21", -- 0x3320
    x"FF",x"12",x"0F",x"12",x"FF",x"21",x"F0",x"21", -- 0x3328
    x"FF",x"12",x"0F",x"12",x"FF",x"21",x"F0",x"32", -- 0x3330
    x"32",x"32",x"32",x"32",x"32",x"00",x"FF",x"7F", -- 0x3338
    x"15",x"80",x"EA",x"7F",x"55",x"01",x"FF",x"FF", -- 0x3340
    x"FF",x"21",x"21",x"F0",x"F0",x"21",x"0F",x"21", -- 0x3348
    x"0F",x"FF",x"FF",x"00",x"FF",x"FF",x"EB",x"03", -- 0x3350
    x"53",x"73",x"F0",x"52",x"FF",x"27",x"0F",x"0F", -- 0x3358
    x"0F",x"0F",x"37",x"45",x"00",x"5F",x"D5",x"FF", -- 0x3360
    x"18",x"2B",x"F7",x"2A",x"54",x"2B",x"46",x"2B", -- 0x3368
    x"3E",x"2B",x"20",x"2B",x"65",x"2B",x"58",x"2B", -- 0x3370
    x"52",x"31",x"51",x"61",x"F0",x"F0",x"61",x"51", -- 0x3378
    x"31",x"52",x"00",x"FF",x"5F",x"05",x"53",x"21", -- 0x3380
    x"52",x"F0",x"52",x"21",x"53",x"F0",x"52",x"21", -- 0x3388
    x"53",x"00",x"FF",x"55",x"15",x"12",x"23",x"FF", -- 0x3390
    x"21",x"41",x"F0",x"F0",x"41",x"21",x"FF",x"23", -- 0x3398
    x"12",x"25",x"13",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x33A0
    x"FF",x"FF",x"FF",x"0F",x"FF",x"FF",x"12",x"12", -- 0x33A8
    x"FF",x"21",x"F0",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x33B0
    x"FF",x"0F",x"83",x"2B",x"78",x"2B",x"92",x"2B", -- 0x33B8
    x"86",x"2B",x"83",x"2B",x"78",x"2B",x"92",x"2B", -- 0x33C0
    x"86",x"2B",x"A7",x"2B",x"95",x"2B",x"B7",x"2B", -- 0x33C8
    x"AC",x"2B",x"A7",x"2B",x"95",x"2B",x"B7",x"2B", -- 0x33D0
    x"AC",x"2B",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E0
    x"00",x"7E",x"00",x"FC",x"01",x"F8",x"03",x"F1", -- 0x33E8
    x"1F",x"F3",x"3F",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x33F0
    x"1F",x"F3",x"03",x"F1",x"01",x"F8",x"00",x"FC", -- 0x33F8
    x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3410
    x"2C",x"2C",x"3C",x"2C",x"24",x"2C",x"44",x"2C", -- 0x3418
    x"4C",x"2C",x"34",x"2C",x"76",x"7F",x"7F",x"FE", -- 0x3420
    x"FE",x"FF",x"7F",x"3A",x"00",x"00",x"1C",x"1E", -- 0x3428
    x"3F",x"3F",x"3E",x"1E",x"38",x"7C",x"7C",x"FC", -- 0x3430
    x"FC",x"78",x"00",x"00",x"40",x"E0",x"E0",x"60", -- 0x3438
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38", -- 0x3440
    x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3448
    x"02",x"07",x"07",x"02",x"00",x"00",x"00",x"2E", -- 0x3450
    x"0C",x"2E",x"40",x"0C",x"2F",x"00",x"00",x"00", -- 0x3458
    x"18",x"0C",x"2E",x"26",x"03",x"44",x"10",x"03", -- 0x3460
    x"44",x"2A",x"0C",x"2F",x"22",x"03",x"44",x"10", -- 0x3468
    x"03",x"44",x"2E",x"03",x"44",x"14",x"03",x"44", -- 0x3470
    x"0C",x"03",x"44",x"02",x"03",x"44",x"04",x"03", -- 0x3478
    x"44",x"0E",x"03",x"44",x"18",x"03",x"44",x"06", -- 0x3480
    x"03",x"44",x"08",x"03",x"44",x"12",x"03",x"44", -- 0x3488
    x"30",x"03",x"44",x"16",x"03",x"44",x"24",x"03", -- 0x3490
    x"44",x"26",x"03",x"44",x"2C",x"0C",x"2C",x"0E", -- 0x3498
    x"03",x"44",x"2C",x"03",x"44",x"40",x"0C",x"2D", -- 0x34A0
    x"00",x"00",x"00",x"32",x"0C",x"2C",x"30",x"0C", -- 0x34A8
    x"2D",x"00",x"00",x"00",x"38",x"7C",x"7C",x"FC", -- 0x34B0
    x"FC",x"78",x"00",x"00",x"40",x"E0",x"E0",x"60", -- 0x34B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38", -- 0x34C0
    x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C8
    x"02",x"07",x"07",x"02",x"00",x"00",x"00",x"2E", -- 0x34D0
    x"0C",x"2E",x"40",x"0C",x"2F",x"00",x"00",x"00", -- 0x34D8
    x"18",x"0C",x"2E",x"26",x"03",x"44",x"10",x"03", -- 0x34E0
    x"44",x"2A",x"0C",x"2F",x"22",x"03",x"44",x"10", -- 0x34E8
    x"03",x"44",x"2E",x"03",x"44",x"14",x"03",x"44", -- 0x34F0
    x"0C",x"03",x"44",x"02",x"03",x"44",x"04",x"03", -- 0x34F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37F8
    x"5F",x"E6",x"1F",x"C6",x"08",x"DD",x"77",x"0B", -- 0x3800
    x"C9",x"E5",x"2A",x"8C",x"40",x"23",x"7C",x"E6", -- 0x3808
    x"1F",x"67",x"22",x"8C",x"40",x"7E",x"E1",x"C9", -- 0x3810
    x"D9",x"4F",x"3A",x"00",x"40",x"FE",x"04",x"CA", -- 0x3818
    x"48",x"28",x"79",x"2A",x"0E",x"41",x"23",x"86", -- 0x3820
    x"C3",x"40",x"28",x"D9",x"4F",x"3A",x"00",x"40", -- 0x3828
    x"FE",x"04",x"79",x"CA",x"48",x"28",x"2A",x"0E", -- 0x3830
    x"41",x"86",x"27",x"77",x"23",x"7E",x"CE",x"00", -- 0x3838
    x"27",x"77",x"23",x"7E",x"CE",x"00",x"27",x"77", -- 0x3840
    x"D9",x"C9",x"3A",x"21",x"41",x"A7",x"C8",x"3A", -- 0x3848
    x"00",x"40",x"FE",x"04",x"C8",x"2A",x"0E",x"41", -- 0x3850
    x"23",x"23",x"7E",x"A7",x"C2",x"66",x"28",x"2B", -- 0x3858
    x"7E",x"21",x"68",x"40",x"BE",x"D8",x"3A",x"00", -- 0x3860
    x"40",x"FE",x"18",x"21",x"60",x"50",x"CA",x"74", -- 0x3868
    x"28",x"21",x"A0",x"53",x"34",x"21",x"10",x"41", -- 0x3870
    x"34",x"AF",x"32",x"21",x"41",x"11",x"CB",x"2A", -- 0x3878
    x"CD",x"1F",x"27",x"C9",x"C9",x"8F",x"28",x"BB", -- 0x3880
    x"28",x"E7",x"28",x"13",x"29",x"3F",x"29",x"B2", -- 0x3888
    x"10",x"F7",x"10",x"72",x"11",x"31",x"11",x"4B", -- 0x3890
    x"12",x"4B",x"12",x"4B",x"12",x"4F",x"13",x"4F", -- 0x3898
    x"13",x"4F",x"13",x"72",x"11",x"72",x"11",x"72", -- 0x38A0
    x"11",x"83",x"13",x"83",x"13",x"83",x"13",x"D3", -- 0x38A8
    x"13",x"D3",x"13",x"D3",x"13",x"02",x"14",x"02", -- 0x38B0
    x"14",x"02",x"14",x"00",x"00",x"00",x"00",x"00", -- 0x38B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C0
    x"00",x"B3",x"14",x"B3",x"14",x"B3",x"14",x"27", -- 0x38C8
    x"15",x"27",x"15",x"27",x"15",x"83",x"13",x"83", -- 0x38D0
    x"13",x"83",x"13",x"00",x"00",x"00",x"00",x"00", -- 0x38D8
    x"00",x"02",x"14",x"02",x"14",x"02",x"14",x"B2", -- 0x38E0
    x"10",x"F7",x"10",x"73",x"17",x"31",x"11",x"4B", -- 0x38E8
    x"12",x"4B",x"12",x"4B",x"12",x"6F",x"15",x"6F", -- 0x38F0
    x"15",x"6F",x"15",x"73",x"17",x"73",x"17",x"73", -- 0x38F8
    x"17",x"83",x"13",x"83",x"13",x"83",x"13",x"DE", -- 0x3900
    x"13",x"DE",x"13",x"DE",x"13",x"02",x"14",x"02", -- 0x3908
    x"14",x"02",x"14",x"B2",x"10",x"F7",x"10",x"72", -- 0x3910
    x"11",x"31",x"11",x"4B",x"12",x"4B",x"12",x"4B", -- 0x3918
    x"12",x"81",x"16",x"81",x"16",x"81",x"16",x"C2", -- 0x3920
    x"17",x"C2",x"17",x"C2",x"17",x"83",x"13",x"83", -- 0x3928
    x"13",x"83",x"13",x"4B",x"17",x"4B",x"17",x"4B", -- 0x3930
    x"17",x"02",x"14",x"02",x"14",x"02",x"14",x"B2", -- 0x3938
    x"10",x"F7",x"10",x"72",x"11",x"31",x"11",x"4B", -- 0x3940
    x"12",x"4B",x"12",x"4B",x"12",x"A4",x"15",x"A4", -- 0x3948
    x"15",x"A4",x"15",x"2F",x"16",x"2F",x"16",x"2F", -- 0x3950
    x"16",x"83",x"13",x"83",x"13",x"83",x"13",x"FF", -- 0x3958
    x"15",x"FF",x"15",x"FF",x"15",x"02",x"14",x"02", -- 0x3960
    x"14",x"02",x"14",x"5E",x"4D",x"7C",x"88",x"5E", -- 0x3968
    x"88",x"4A",x"7A",x"4A",x"72",x"4A",x"60",x"7C", -- 0x3970
    x"A6",x"5E",x"88",x"4A",x"7A",x"4A",x"72",x"4A", -- 0x3978
    x"60",x"7C",x"A6",x"5E",x"88",x"4A",x"7A",x"4A", -- 0x3980
    x"72",x"4A",x"7A",x"7C",x"60",x"4F",x"11",x"47", -- 0x3988
    x"FF",x"47",x"11",x"7C",x"4D",x"7C",x"4D",x"00", -- 0x3990
    x"FE",x"41",x"8F",x"41",x"A1",x"41",x"8F",x"41", -- 0x3998
    x"A1",x"41",x"8F",x"41",x"A1",x"05",x"FF",x"41", -- 0x39A0
    x"8F",x"41",x"A1",x"41",x"8F",x"41",x"A1",x"41", -- 0x39A8
    x"8F",x"41",x"A1",x"05",x"FF",x"41",x"8F",x"41", -- 0x39B0
    x"A1",x"41",x"8F",x"41",x"A1",x"41",x"8F",x"41", -- 0x39B8
    x"A1",x"41",x"FD",x"8F",x"A1",x"41",x"FC",x"01", -- 0x39C0
    x"A6",x"41",x"FC",x"FF",x"00",x"00",x"FE",x"C4", -- 0x39C8
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C2",x"FF",x"C4", -- 0x39D0
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C2",x"FF",x"C4", -- 0x39D8
    x"E5",x"C2",x"FF",x"C4",x"E5",x"C1",x"FD",x"E5", -- 0x39E0
    x"D8",x"C1",x"FC",x"FF",x"30",x"00",x"FE",x"C2", -- 0x39E8
    x"1E",x"C2",x"57",x"C2",x"81",x"C2",x"2B",x"C2", -- 0x39F0
    x"60",x"C2",x"88",x"C2",x"37",x"C2",x"69",x"C2", -- 0x39F8
    x"8F",x"00",x"FE",x"C4",x"DC",x"C3",x"D6",x"C2", -- 0x3A00
    x"E5",x"C1",x"E1",x"00",x"FE",x"C2",x"A6",x"C4", -- 0x3A08
    x"B9",x"C2",x"A6",x"C4",x"1E",x"C2",x"A6",x"C4", -- 0x3A10
    x"B9",x"C2",x"A6",x"00",x"FE",x"43",x"11",x"42", -- 0x3A18
    x"1E",x"42",x"11",x"C3",x"4D",x"41",x"37",x"42", -- 0x3A20
    x"81",x"42",x"11",x"C2",x"60",x"43",x"1E",x"00", -- 0x3A28
    x"FE",x"44",x"FB",x"1E",x"11",x"44",x"FA",x"42", -- 0x3A30
    x"4D",x"42",x"7A",x"6C",x"95",x"56",x"95",x"42", -- 0x3A38
    x"69",x"42",x"7A",x"56",x"95",x"42",x"60",x"42", -- 0x3A40
    x"7A",x"56",x"9B",x"42",x"60",x"42",x"7A",x"6C", -- 0x3A48
    x"9B",x"42",x"4D",x"42",x"7A",x"56",x"95",x"42", -- 0x3A50
    x"60",x"42",x"7A",x"61",x"9B",x"42",x"7A",x"4B", -- 0x3A58
    x"95",x"42",x"72",x"56",x"88",x"42",x"60",x"56", -- 0x3A60
    x"7A",x"42",x"4D",x"6C",x"72",x"56",x"72",x"42", -- 0x3A68
    x"72",x"56",x"88",x"42",x"7A",x"42",x"95",x"6C", -- 0x3A70
    x"A6",x"42",x"4D",x"42",x"72",x"6C",x"9B",x"42", -- 0x3A78
    x"7A",x"4B",x"95",x"4B",x"7A",x"42",x"72",x"4B", -- 0x3A80
    x"9B",x"4B",x"88",x"42",x"7A",x"42",x"95",x"56", -- 0x3A88
    x"A6",x"42",x"60",x"42",x"7A",x"56",x"9B",x"42", -- 0x3A90
    x"4D",x"42",x"7A",x"6C",x"95",x"42",x"4D",x"42", -- 0x3A98
    x"72",x"6C",x"88",x"6C",x"7A",x"6C",x"7A",x"00", -- 0x3AA0
    x"FE",x"41",x"FD",x"69",x"72",x"41",x"FC",x"FF", -- 0x3AA8
    x"57",x"41",x"FD",x"42",x"57",x"41",x"FC",x"01", -- 0x3AB0
    x"88",x"41",x"FD",x"95",x"88",x"41",x"FC",x"FF", -- 0x3AB8
    x"1E",x"41",x"FD",x"1E",x"11",x"41",x"FC",x"01", -- 0x3AC0
    x"E5",x"00",x"FE",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x3AC8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x3AD0
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x3AD8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x3AE0
    x"1E",x"C2",x"FF",x"C4",x"1E",x"C2",x"FF",x"C4", -- 0x3AE8
    x"1E",x"C2",x"FF",x"C4",x"1E",x"00",x"FE",x"F0", -- 0x3AF0
    x"41",x"41",x"53",x"53",x"FF",x"53",x"31",x"F0", -- 0x3AF8
    x"43",x"35",x"0F",x"12",x"12",x"12",x"54",x"52", -- 0x3B00
    x"51",x"F0",x"41",x"35",x"0F",x"15",x"35",x"FF", -- 0x3B08
    x"53",x"53",x"52",x"F0",x"52",x"53",x"41",x"00", -- 0x3B10
    x"FF",x"FF",x"57",x"00",x"80",x"FA",x"FF",x"57", -- 0x3B18
    x"32",x"32",x"32",x"32",x"32",x"32",x"F0",x"21", -- 0x3B20
    x"FF",x"12",x"0F",x"12",x"FF",x"21",x"F0",x"21", -- 0x3B28
    x"FF",x"12",x"0F",x"12",x"FF",x"21",x"F0",x"32", -- 0x3B30
    x"32",x"32",x"32",x"32",x"32",x"00",x"FF",x"7F", -- 0x3B38
    x"15",x"80",x"EA",x"7F",x"55",x"01",x"FF",x"FF", -- 0x3B40
    x"FF",x"21",x"21",x"F0",x"F0",x"21",x"0F",x"21", -- 0x3B48
    x"0F",x"FF",x"FF",x"00",x"FF",x"FF",x"EB",x"03", -- 0x3B50
    x"53",x"73",x"F0",x"52",x"FF",x"27",x"0F",x"0F", -- 0x3B58
    x"0F",x"0F",x"37",x"45",x"00",x"5F",x"D5",x"FF", -- 0x3B60
    x"18",x"2B",x"F7",x"2A",x"54",x"2B",x"46",x"2B", -- 0x3B68
    x"3E",x"2B",x"20",x"2B",x"65",x"2B",x"58",x"2B", -- 0x3B70
    x"52",x"31",x"51",x"61",x"F0",x"F0",x"61",x"51", -- 0x3B78
    x"31",x"52",x"00",x"FF",x"5F",x"05",x"53",x"21", -- 0x3B80
    x"52",x"F0",x"52",x"21",x"53",x"F0",x"52",x"21", -- 0x3B88
    x"53",x"00",x"FF",x"55",x"15",x"12",x"23",x"FF", -- 0x3B90
    x"21",x"41",x"F0",x"F0",x"41",x"21",x"FF",x"23", -- 0x3B98
    x"12",x"25",x"13",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x3BA0
    x"FF",x"FF",x"FF",x"0F",x"FF",x"FF",x"12",x"12", -- 0x3BA8
    x"FF",x"21",x"F0",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x3BB0
    x"FF",x"0F",x"83",x"2B",x"78",x"2B",x"92",x"2B", -- 0x3BB8
    x"86",x"2B",x"83",x"2B",x"78",x"2B",x"92",x"2B", -- 0x3BC0
    x"86",x"2B",x"A7",x"2B",x"95",x"2B",x"B7",x"2B", -- 0x3BC8
    x"AC",x"2B",x"A7",x"2B",x"95",x"2B",x"B7",x"2B", -- 0x3BD0
    x"AC",x"2B",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE0
    x"00",x"7E",x"00",x"FC",x"01",x"F8",x"03",x"F1", -- 0x3BE8
    x"1F",x"F3",x"3F",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x3BF0
    x"1F",x"F3",x"03",x"F1",x"01",x"F8",x"00",x"FC", -- 0x3BF8
    x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C10
    x"2C",x"2C",x"3C",x"2C",x"24",x"2C",x"44",x"2C", -- 0x3C18
    x"4C",x"2C",x"34",x"2C",x"76",x"7F",x"7F",x"FE", -- 0x3C20
    x"FE",x"FF",x"7F",x"3A",x"00",x"00",x"1C",x"1E", -- 0x3C28
    x"3F",x"3F",x"3E",x"1E",x"38",x"7C",x"7C",x"FC", -- 0x3C30
    x"FC",x"78",x"00",x"00",x"40",x"E0",x"E0",x"60", -- 0x3C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38", -- 0x3C40
    x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C48
    x"02",x"07",x"07",x"02",x"00",x"00",x"00",x"2E", -- 0x3C50
    x"0C",x"2E",x"40",x"0C",x"2F",x"00",x"00",x"00", -- 0x3C58
    x"18",x"0C",x"2E",x"26",x"03",x"44",x"10",x"03", -- 0x3C60
    x"44",x"2A",x"0C",x"2F",x"22",x"03",x"44",x"10", -- 0x3C68
    x"03",x"44",x"2E",x"03",x"44",x"14",x"03",x"44", -- 0x3C70
    x"0C",x"03",x"44",x"02",x"03",x"44",x"04",x"03", -- 0x3C78
    x"44",x"0E",x"03",x"44",x"18",x"03",x"44",x"06", -- 0x3C80
    x"03",x"44",x"08",x"03",x"44",x"12",x"03",x"44", -- 0x3C88
    x"30",x"03",x"44",x"16",x"03",x"44",x"24",x"03", -- 0x3C90
    x"44",x"26",x"03",x"44",x"2C",x"0C",x"2C",x"0E", -- 0x3C98
    x"03",x"44",x"2C",x"03",x"44",x"40",x"0C",x"2D", -- 0x3CA0
    x"00",x"00",x"00",x"32",x"0C",x"2C",x"30",x"0C", -- 0x3CA8
    x"2D",x"00",x"00",x"00",x"38",x"7C",x"7C",x"FC", -- 0x3CB0
    x"FC",x"78",x"00",x"00",x"40",x"E0",x"E0",x"60", -- 0x3CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38", -- 0x3CC0
    x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC8
    x"02",x"07",x"07",x"02",x"00",x"00",x"00",x"2E", -- 0x3CD0
    x"0C",x"2E",x"40",x"0C",x"2F",x"00",x"00",x"00", -- 0x3CD8
    x"18",x"0C",x"2E",x"26",x"03",x"44",x"10",x"03", -- 0x3CE0
    x"44",x"2A",x"0C",x"2F",x"22",x"03",x"44",x"10", -- 0x3CE8
    x"03",x"44",x"2E",x"03",x"44",x"14",x"03",x"44", -- 0x3CF0
    x"0C",x"03",x"44",x"02",x"03",x"44",x"04",x"03", -- 0x3CF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
       DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
