library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity hector1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of hector1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"40",X"32",X"02",X"28",X"C3",X"0C",X"00",X"F3",X"C3",X"04",X"08",X"3E",X"38",X"32",X"00",
		X"30",X"AF",X"32",X"00",X"10",X"32",X"00",X"18",X"06",X"3E",X"21",X"C0",X"5F",X"F9",X"77",X"23",
		X"05",X"C2",X"1E",X"00",X"3A",X"00",X"08",X"B7",X"CA",X"00",X"08",X"3A",X"00",X"30",X"77",X"3E",
		X"80",X"32",X"DB",X"5F",X"C3",X"8C",X"01",X"FF",X"E5",X"D5",X"C5",X"F5",X"3A",X"F5",X"5F",X"B7",
		X"C2",X"6A",X"00",X"21",X"C0",X"5F",X"7E",X"1F",X"1F",X"1F",X"E6",X"07",X"F5",X"11",X"F6",X"5F",
		X"83",X"5F",X"3A",X"00",X"30",X"12",X"F1",X"3D",X"C2",X"5D",X"00",X"3E",X"06",X"87",X"87",X"87",
		X"AE",X"E6",X"F8",X"AE",X"F6",X"40",X"77",X"32",X"00",X"30",X"2A",X"EF",X"5F",X"23",X"22",X"EF",
		X"5F",X"11",X"06",X"38",X"21",X"C8",X"5F",X"01",X"CF",X"5F",X"1A",X"2F",X"A6",X"C2",X"89",X"00",
		X"2B",X"0B",X"1D",X"F2",X"7A",X"00",X"C3",X"24",X"01",X"F5",X"0A",X"2F",X"E3",X"A4",X"E1",X"CA",
		X"80",X"00",X"11",X"02",X"07",X"F5",X"21",X"C9",X"5F",X"7E",X"87",X"D2",X"9F",X"00",X"1D",X"C2",
		X"9A",X"00",X"23",X"15",X"C2",X"99",X"00",X"F1",X"1D",X"FA",X"24",X"01",X"16",X"08",X"0F",X"D2",
		X"B5",X"00",X"5A",X"3E",X"80",X"15",X"C2",X"AE",X"00",X"57",X"0A",X"B2",X"02",X"79",X"D6",X"C9",
		X"87",X"87",X"87",X"83",X"3D",X"FE",X"02",X"21",X"D2",X"5F",X"C2",X"D3",X"00",X"7E",X"2F",X"77",
		X"C3",X"24",X"01",X"FE",X"07",X"DA",X"E9",X"00",X"57",X"3A",X"00",X"38",X"2F",X"E6",X"80",X"B6",
		X"7A",X"CA",X"F5",X"00",X"FE",X"17",X"D2",X"F0",X"00",X"21",X"75",X"01",X"85",X"6F",X"7E",X"11",
		X"C6",X"23",X"C3",X"03",X"01",X"C6",X"23",X"FE",X"41",X"DA",X"03",X"01",X"FE",X"5B",X"D2",X"03",
		X"01",X"C6",X"20",X"57",X"3A",X"00",X"38",X"E6",X"C0",X"EE",X"80",X"7A",X"C2",X"16",X"01",X"FE",
		X"60",X"DA",X"16",X"01",X"D6",X"60",X"32",X"D1",X"5F",X"21",X"D0",X"5F",X"7E",X"B7",X"CA",X"23",
		X"01",X"36",X"80",X"34",X"01",X"00",X"38",X"11",X"C2",X"5F",X"21",X"C9",X"5F",X"0A",X"F6",X"C0",
		X"FE",X"0A",X"2F",X"12",X"A6",X"77",X"03",X"13",X"23",X"3E",X"07",X"B9",X"C2",X"31",X"01",X"21",
		X"C1",X"5F",X"46",X"3A",X"07",X"38",X"2F",X"77",X"A0",X"47",X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",
		X"21",X"F2",X"5F",X"77",X"2B",X"78",X"E6",X"0F",X"77",X"3A",X"F5",X"5F",X"B7",X"C2",X"6A",X"01",
		X"21",X"C0",X"5F",X"7E",X"EE",X"C0",X"77",X"32",X"00",X"30",X"2A",X"F3",X"5F",X"7D",X"B4",X"E5",
		X"C0",X"E1",X"F1",X"C1",X"D1",X"E1",X"FB",X"C9",X"08",X"09",X"0D",X"20",X"2A",X"5E",X"23",X"5F",
		X"26",X"40",X"3C",X"3E",X"22",X"27",X"24",X"25",X"21",X"3A",X"28",X"29",X"FB",X"CD",X"73",X"05",
		X"01",X"E8",X"01",X"CD",X"D3",X"01",X"3A",X"00",X"4C",X"FE",X"31",X"F5",X"03",X"01",X"EB",X"0F",
		X"CC",X"D3",X"01",X"01",X"17",X"02",X"CD",X"36",X"06",X"CD",X"E0",X"07",X"47",X"F1",X"78",X"20",
		X"05",X"FE",X"72",X"CA",X"00",X"4C",X"D6",X"6D",X"CA",X"57",X"08",X"3C",X"20",X"D8",X"01",X"01",
		X"01",X"11",X"00",X"00",X"CD",X"1C",X"02",X"B7",X"20",X"08",X"3A",X"00",X"4C",X"FE",X"31",X"CA",
		X"00",X"4C",X"C7",X"0A",X"FE",X"FF",X"C8",X"CD",X"2F",X"06",X"03",X"0A",X"5F",X"03",X"0A",X"57",
		X"03",X"CD",X"4F",X"05",X"03",X"C3",X"D3",X"01",X"03",X"0C",X"0A",X"54",X"41",X"50",X"45",X"5A",
		X"00",X"02",X"1C",X"0A",X"4C",X"3A",X"4C",X"45",X"43",X"54",X"55",X"52",X"45",X"20",X"4B",X"37",
		X"00",X"02",X"26",X"0A",X"4D",X"3A",X"4D",X"4F",X"4E",X"49",X"54",X"45",X"55",X"52",X"00",X"FF",
		X"4C",X"41",X"4E",X"43",X"45",X"00",X"FF",X"04",X"01",X"02",X"07",X"00",X"F3",X"AF",X"32",X"D3",
		X"5F",X"D5",X"C5",X"CD",X"CA",X"02",X"CD",X"DD",X"02",X"01",X"1D",X"00",X"CD",X"F6",X"07",X"01",
		X"64",X"01",X"1E",X"00",X"CD",X"B1",X"03",X"C1",X"C5",X"01",X"05",X"00",X"11",X"D4",X"5F",X"CD",
		X"1A",X"03",X"C1",X"B7",X"CA",X"5D",X"02",X"32",X"D3",X"5F",X"78",X"B7",X"C2",X"38",X"02",X"D1",
		X"7A",X"B7",X"C2",X"58",X"02",X"CD",X"E3",X"02",X"3A",X"D3",X"5F",X"FB",X"C9",X"C5",X"2A",X"DD",
		X"5F",X"7C",X"B5",X"CA",X"6F",X"02",X"22",X"D4",X"5F",X"2A",X"DF",X"5F",X"22",X"D6",X"5F",X"3A",
		X"D8",X"5F",X"FE",X"FD",X"C2",X"7B",X"02",X"C1",X"C3",X"4F",X"02",X"FE",X"FE",X"C2",X"AE",X"02",
		X"21",X"D9",X"5F",X"01",X"01",X"00",X"CD",X"1A",X"03",X"C1",X"B7",X"CA",X"99",X"02",X"32",X"D3",
		X"5F",X"78",X"B7",X"C2",X"38",X"02",X"C3",X"4F",X"02",X"2A",X"D6",X"5F",X"EB",X"2A",X"D4",X"5F",
		X"3A",X"D9",X"5F",X"77",X"23",X"1B",X"7A",X"B3",X"C2",X"A0",X"02",X"C3",X"38",X"02",X"2A",X"D4",
		X"5F",X"EB",X"2A",X"D6",X"5F",X"44",X"4D",X"CD",X"00",X"03",X"C1",X"B7",X"CA",X"38",X"02",X"32",
		X"D3",X"5F",X"78",X"B7",X"C2",X"38",X"02",X"C3",X"4F",X"02",X"0F",X"2F",X"E6",X"40",X"32",X"02",
		X"28",X"3A",X"C0",X"5F",X"F6",X"07",X"32",X"C0",X"5F",X"32",X"00",X"30",X"C9",X"F5",X"3E",X"FF",
		X"C3",X"E5",X"02",X"F5",X"AF",X"E5",X"21",X"DB",X"5F",X"AE",X"E6",X"40",X"AE",X"77",X"32",X"00",
		X"10",X"21",X"C0",X"5F",X"7E",X"E6",X"07",X"F6",X"38",X"77",X"32",X"00",X"30",X"E1",X"F1",X"C9",
		X"E5",X"CD",X"DD",X"02",X"AF",X"32",X"D3",X"5F",X"CD",X"1A",X"03",X"21",X"D3",X"5F",X"B6",X"77",
		X"78",X"B1",X"C2",X"08",X"03",X"E1",X"3A",X"D3",X"5F",X"C9",X"E5",X"C5",X"CD",X"4F",X"03",X"C1",
		X"67",X"D2",X"36",X"03",X"6F",X"7B",X"84",X"5F",X"7A",X"CE",X"00",X"57",X"79",X"94",X"4F",X"7A",
		X"DE",X"00",X"47",X"7D",X"E1",X"C9",X"CD",X"9A",X"03",X"DA",X"24",X"03",X"12",X"13",X"0B",X"25",
		X"CA",X"4C",X"03",X"78",X"B1",X"C2",X"36",X"03",X"3E",X"04",X"E1",X"C9",X"E1",X"AF",X"C9",X"CD",
		X"D0",X"03",X"FE",X"15",X"DA",X"4F",X"03",X"CD",X"D0",X"03",X"FE",X"21",X"D2",X"4F",X"03",X"FE",
		X"15",X"D2",X"57",X"03",X"C5",X"FE",X"0E",X"3F",X"0E",X"80",X"DA",X"A8",X"03",X"CD",X"D0",X"03",
		X"FE",X"21",X"D2",X"95",X"03",X"FE",X"15",X"0E",X"40",X"DA",X"A5",X"03",X"CD",X"D0",X"03",X"FE",
		X"0E",X"D2",X"95",X"03",X"CD",X"D0",X"03",X"FE",X"21",X"D2",X"95",X"03",X"FE",X"15",X"DA",X"95",
		X"03",X"00",X"3E",X"01",X"01",X"3E",X"02",X"C1",X"37",X"C9",X"C5",X"0E",X"80",X"CD",X"D0",X"03",
		X"FE",X"15",X"D2",X"95",X"03",X"FE",X"0E",X"3F",X"79",X"1F",X"4F",X"D2",X"9D",X"03",X"B7",X"C1",
		X"C9",X"C5",X"CD",X"D0",X"03",X"FE",X"21",X"D2",X"CC",X"03",X"FE",X"15",X"DA",X"CC",X"03",X"0B",
		X"78",X"B1",X"C2",X"B2",X"03",X"7B",X"B7",X"C4",X"CA",X"02",X"C1",X"C9",X"C1",X"C3",X"B1",X"03",
		X"E5",X"2A",X"DA",X"5F",X"3A",X"00",X"30",X"AD",X"F2",X"D4",X"03",X"AD",X"32",X"DA",X"5F",X"95",
		X"E1",X"E6",X"7F",X"C9",X"C5",X"06",X"08",X"79",X"0F",X"4F",X"9F",X"E6",X"08",X"C6",X"08",X"CD",
		X"F8",X"03",X"05",X"C2",X"E7",X"03",X"C1",X"C9",X"D6",X"02",X"CD",X"FF",X"03",X"3E",X"02",X"E5",
		X"2A",X"DA",X"5F",X"85",X"E6",X"7F",X"6F",X"3A",X"00",X"30",X"E6",X"7F",X"BD",X"C2",X"07",X"04",
		X"7C",X"EE",X"80",X"32",X"00",X"10",X"67",X"22",X"DA",X"5F",X"E1",X"C9",X"3A",X"00",X"30",X"E6",
		X"7F",X"32",X"DA",X"5F",X"78",X"B1",X"C8",X"3E",X"1B",X"CD",X"F8",X"03",X"0B",X"C3",X"24",X"04",
		X"CD",X"33",X"04",X"3E",X"08",X"CD",X"F8",X"03",X"01",X"01",X"00",X"C3",X"24",X"04",X"79",X"B7",
		X"C8",X"E5",X"D5",X"57",X"2A",X"E1",X"5F",X"7C",X"B5",X"C2",X"4F",X"04",X"21",X"7A",X"06",X"7A",
		X"FE",X"61",X"DA",X"5A",X"04",X"D6",X"43",X"C3",X"6F",X"04",X"FE",X"1E",X"3D",X"DA",X"6F",X"04",
		X"D6",X"1D",X"57",X"2A",X"E3",X"5F",X"7C",X"B5",X"7A",X"C2",X"6F",X"04",X"21",X"6E",X"06",X"5E",
		X"23",X"56",X"23",X"E5",X"D5",X"CD",X"18",X"05",X"D1",X"7A",X"C6",X"07",X"1F",X"1F",X"1F",X"E6",
		X"1F",X"EB",X"E3",X"CD",X"1D",X"05",X"22",X"E5",X"5F",X"E1",X"D1",X"D5",X"C5",X"01",X"00",X"00",
		X"CD",X"9D",X"04",X"C1",X"D1",X"E1",X"C9",X"CD",X"F7",X"05",X"CD",X"B3",X"05",X"E5",X"21",X"DB",
		X"04",X"22",X"EB",X"5F",X"E1",X"7C",X"B7",X"C8",X"7D",X"B7",X"C8",X"C5",X"D5",X"E5",X"22",X"E9",
		X"5F",X"E5",X"C5",X"D5",X"E5",X"2A",X"EB",X"5F",X"CD",X"DA",X"04",X"E1",X"D1",X"C1",X"0C",X"1C",
		X"2D",X"C2",X"B2",X"04",X"E3",X"7D",X"E3",X"6F",X"79",X"95",X"4F",X"7B",X"95",X"5F",X"04",X"14",
		X"25",X"C2",X"B2",X"04",X"E1",X"E1",X"D1",X"C1",X"37",X"C9",X"E9",X"CD",X"ED",X"04",X"C8",X"3A",
		X"EE",X"5F",X"4F",X"CD",X"2D",X"05",X"47",X"79",X"AE",X"A0",X"AE",X"77",X"C9",X"3A",X"EA",X"5F",
		X"C6",X"07",X"1F",X"1F",X"1F",X"E6",X"1F",X"D5",X"59",X"16",X"00",X"2A",X"E5",X"5F",X"CD",X"1D",
		X"05",X"78",X"1F",X"1F",X"1F",X"E6",X"1F",X"5F",X"16",X"00",X"19",X"78",X"E6",X"07",X"5F",X"7E",
		X"87",X"1D",X"F2",X"10",X"05",X"9F",X"D1",X"C9",X"16",X"00",X"21",X"00",X"00",X"D5",X"B7",X"1F",
		X"D2",X"24",X"05",X"19",X"EB",X"29",X"EB",X"B7",X"C2",X"1F",X"05",X"D1",X"C9",X"6B",X"26",X"00",
		X"29",X"29",X"29",X"29",X"29",X"7A",X"1F",X"1F",X"E6",X"3F",X"B5",X"6F",X"7A",X"EB",X"E6",X"03",
		X"21",X"4B",X"05",X"85",X"6F",X"7E",X"2A",X"E7",X"5F",X"19",X"C9",X"03",X"0C",X"30",X"C0",X"CD",
		X"F7",X"05",X"0A",X"CD",X"5C",X"05",X"D0",X"03",X"C3",X"52",X"05",X"79",X"CD",X"3F",X"04",X"D0",
		X"3A",X"EA",X"5F",X"3C",X"82",X"FE",X"67",X"57",X"D8",X"3A",X"E9",X"5F",X"3C",X"83",X"5F",X"16",
		X"06",X"37",X"C9",X"0E",X"00",X"E5",X"D5",X"79",X"CD",X"E8",X"05",X"4F",X"21",X"00",X"40",X"11",
		X"A0",X"09",X"71",X"23",X"1B",X"7A",X"B3",X"C2",X"82",X"05",X"D1",X"E1",X"C9",X"CD",X"F7",X"05",
		X"21",X"D2",X"05",X"22",X"EB",X"5F",X"CD",X"B3",X"05",X"CD",X"E8",X"05",X"32",X"ED",X"5F",X"C3",
		X"A5",X"04",X"CD",X"F7",X"05",X"21",X"DF",X"04",X"22",X"EB",X"5F",X"60",X"69",X"CD",X"BE",X"05",
		X"C3",X"A5",X"04",X"60",X"69",X"5E",X"23",X"56",X"23",X"EB",X"22",X"E5",X"5F",X"EB",X"5E",X"23",
		X"56",X"23",X"D5",X"7E",X"23",X"CD",X"2F",X"06",X"5E",X"23",X"56",X"23",X"7E",X"E1",X"01",X"00",
		X"00",X"C9",X"CD",X"ED",X"04",X"C8",X"CD",X"2D",X"05",X"47",X"A6",X"4F",X"3A",X"EE",X"5F",X"A0",
		X"B9",X"C0",X"3A",X"ED",X"5F",X"C3",X"E8",X"04",X"E6",X"03",X"C5",X"4F",X"87",X"87",X"81",X"87",
		X"87",X"81",X"87",X"87",X"81",X"C1",X"C9",X"E5",X"21",X"00",X"40",X"22",X"E7",X"5F",X"E1",X"C9",
		X"E5",X"D5",X"C5",X"CD",X"F7",X"05",X"79",X"CD",X"E8",X"05",X"CD",X"E2",X"04",X"C1",X"D1",X"E1",
		X"CD",X"F7",X"05",X"E5",X"D5",X"C5",X"50",X"59",X"78",X"E6",X"03",X"47",X"CD",X"2D",X"05",X"7E",
		X"0F",X"0F",X"05",X"F2",X"20",X"06",X"07",X"07",X"E6",X"03",X"C1",X"D1",X"E1",X"C9",X"79",X"CD",
		X"E8",X"05",X"32",X"EE",X"5F",X"C9",X"D5",X"3A",X"DB",X"5F",X"E6",X"C0",X"CD",X"5E",X"06",X"32",
		X"00",X"10",X"32",X"DB",X"5F",X"0B",X"3A",X"DC",X"5F",X"E6",X"80",X"CD",X"5E",X"06",X"57",X"03",
		X"0A",X"0F",X"0F",X"E6",X"40",X"B2",X"32",X"00",X"18",X"32",X"DC",X"5F",X"D1",X"C9",X"57",X"0A",
		X"03",X"E6",X"07",X"B2",X"57",X"03",X"0A",X"E6",X"07",X"17",X"17",X"17",X"B2",X"C9",X"05",X"05",
		X"00",X"50",X"20",X"50",X"00",X"C0",X"60",X"30",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"20",
		X"20",X"20",X"00",X"20",X"50",X"50",X"00",X"00",X"00",X"50",X"F8",X"50",X"F8",X"50",X"70",X"A0",
		X"70",X"28",X"70",X"C8",X"D0",X"20",X"58",X"98",X"20",X"50",X"20",X"50",X"28",X"20",X"40",X"00",
		X"00",X"00",X"20",X"40",X"40",X"40",X"20",X"20",X"10",X"10",X"10",X"20",X"A8",X"70",X"F8",X"70",
		X"A8",X"00",X"20",X"70",X"20",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"08",X"10",X"20",X"40",X"80",X"70",X"88",X"88",X"88",X"70",X"20",
		X"60",X"20",X"20",X"70",X"F8",X"08",X"F8",X"80",X"F8",X"F8",X"08",X"38",X"08",X"F8",X"90",X"90",
		X"F8",X"10",X"10",X"F0",X"80",X"F0",X"08",X"F0",X"F8",X"80",X"F8",X"88",X"F8",X"F8",X"08",X"10",
		X"20",X"20",X"F8",X"88",X"F8",X"88",X"F8",X"F8",X"88",X"F8",X"08",X"F8",X"00",X"20",X"00",X"20",
		X"00",X"00",X"20",X"00",X"20",X"40",X"10",X"20",X"40",X"20",X"10",X"00",X"70",X"00",X"70",X"00",
		X"40",X"20",X"10",X"20",X"40",X"F8",X"88",X"38",X"00",X"20",X"30",X"48",X"50",X"40",X"38",X"70",
		X"88",X"F8",X"88",X"88",X"F8",X"88",X"F0",X"88",X"F8",X"F8",X"80",X"80",X"80",X"F8",X"F0",X"88",
		X"88",X"88",X"F0",X"F8",X"80",X"E0",X"80",X"F8",X"F8",X"80",X"E0",X"80",X"80",X"F8",X"80",X"98",
		X"88",X"F8",X"88",X"88",X"F8",X"88",X"88",X"70",X"20",X"20",X"20",X"70",X"08",X"08",X"08",X"88",
		X"F8",X"88",X"90",X"E0",X"90",X"88",X"80",X"80",X"80",X"80",X"F8",X"88",X"D8",X"A8",X"88",X"88",
		X"88",X"C8",X"A8",X"98",X"88",X"F8",X"88",X"88",X"88",X"F8",X"F8",X"88",X"F8",X"80",X"80",X"F8",
		X"88",X"A8",X"90",X"E8",X"F8",X"88",X"F8",X"90",X"88",X"F8",X"80",X"F8",X"08",X"F8",X"F8",X"20",
		X"20",X"20",X"20",X"88",X"88",X"88",X"88",X"F8",X"88",X"88",X"50",X"70",X"20",X"88",X"88",X"A8",
		X"D8",X"88",X"88",X"50",X"20",X"50",X"88",X"88",X"50",X"20",X"20",X"20",X"F8",X"10",X"20",X"40",
		X"F8",X"30",X"20",X"20",X"20",X"30",X"80",X"40",X"20",X"10",X"08",X"60",X"20",X"20",X"20",X"60",
		X"20",X"50",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"20",X"10",X"00",X"00",X"00",X"21",
		X"DC",X"5F",X"7E",X"EE",X"80",X"77",X"32",X"00",X"18",X"F5",X"C5",X"60",X"69",X"01",X"FF",X"FF",
		X"09",X"DA",X"D0",X"07",X"C1",X"F1",X"FA",X"BF",X"07",X"1B",X"7A",X"B3",X"C2",X"BF",X"07",X"C9",
		X"3A",X"D0",X"5F",X"B7",X"CA",X"E0",X"07",X"3A",X"D0",X"5F",X"B7",X"C8",X"07",X"3E",X"00",X"32",
		X"D0",X"5F",X"3A",X"D1",X"5F",X"C9",X"C5",X"0B",X"78",X"B1",X"C2",X"F7",X"07",X"C1",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"22",X"B5",X"49",X"E1",X"22",X"B3",X"49",X"F5",X"E1",X"22",X"AB",X"49",
		X"21",X"00",X"00",X"39",X"31",X"B3",X"49",X"E5",X"D5",X"C5",X"31",X"C0",X"5F",X"3A",X"A0",X"49",
		X"3C",X"3C",X"BD",X"CA",X"49",X"08",X"0E",X"40",X"3A",X"A5",X"49",X"B7",X"C2",X"3D",X"08",X"23",
		X"23",X"22",X"B1",X"49",X"2A",X"B3",X"49",X"2B",X"22",X"B3",X"49",X"0E",X"2A",X"2A",X"B3",X"49",
		X"CD",X"74",X"0B",X"CD",X"67",X"0C",X"C3",X"A7",X"08",X"2B",X"2B",X"22",X"B1",X"49",X"21",X"00",
		X"00",X"22",X"B3",X"49",X"C3",X"A7",X"08",X"CD",X"73",X"05",X"01",X"CC",X"0F",X"CD",X"36",X"06",
		X"01",X"D1",X"0F",X"CD",X"D3",X"01",X"FB",X"CD",X"56",X"09",X"FE",X"03",X"20",X"11",X"F3",X"21",
		X"E0",X"48",X"F9",X"11",X"FF",X"7F",X"0E",X"00",X"CD",X"46",X"09",X"D2",X"57",X"08",X"76",X"3E",
		X"C3",X"32",X"03",X"4C",X"21",X"57",X"08",X"22",X"04",X"4C",X"00",X"00",X"00",X"21",X"00",X"4A",
		X"22",X"B1",X"49",X"CD",X"BC",X"09",X"21",X"DF",X"0F",X"22",X"E1",X"5F",X"3A",X"DB",X"5F",X"F6",
		X"80",X"32",X"DB",X"5F",X"CD",X"73",X"05",X"31",X"C0",X"5F",X"21",X"A7",X"08",X"E5",X"FB",X"AF",
		X"32",X"FF",X"5F",X"32",X"A5",X"49",X"CD",X"E3",X"02",X"3E",X"01",X"CD",X"2F",X"06",X"21",X"DE",
		X"08",X"3E",X"1F",X"CD",X"93",X"0C",X"CD",X"2F",X"06",X"CD",X"CC",X"0C",X"D6",X"41",X"F8",X"FE",
		X"1A",X"F0",X"0E",X"02",X"87",X"16",X"00",X"5F",X"19",X"CD",X"B4",X"0C",X"EB",X"E9",X"28",X"09",
		X"2B",X"00",X"A4",X"08",X"12",X"09",X"75",X"0F",X"40",X"09",X"6B",X"09",X"91",X"09",X"F7",X"4B",
		X"FA",X"4B",X"FD",X"4B",X"AF",X"0D",X"C2",X"09",X"03",X"0A",X"29",X"0A",X"AA",X"09",X"00",X"08",
		X"53",X"09",X"59",X"0A",X"C2",X"0E",X"2C",X"0B",X"5D",X"0B",X"F5",X"0D",X"8C",X"0A",X"7B",X"0D",
		X"00",X"4C",X"CD",X"F0",X"0B",X"CD",X"74",X"0B",X"CD",X"8B",X"0C",X"7D",X"E6",X"03",X"C2",X"18",
		X"09",X"CD",X"3E",X"0C",X"D8",X"C3",X"15",X"09",X"CD",X"F0",X"0B",X"CD",X"74",X"0B",X"7E",X"CD",
		X"2B",X"0C",X"23",X"7D",X"E6",X"07",X"C2",X"2E",X"09",X"CD",X"3E",X"0C",X"D8",X"C3",X"2B",X"09",
		X"CD",X"C0",X"0B",X"C1",X"D1",X"E1",X"71",X"CD",X"AA",X"0B",X"D8",X"CD",X"7F",X"0B",X"3F",X"DA",
		X"46",X"09",X"C9",X"CD",X"DD",X"02",X"CD",X"E0",X"07",X"F5",X"C5",X"D5",X"E5",X"01",X"18",X"00",
		X"11",X"35",X"00",X"F3",X"CD",X"BF",X"07",X"FB",X"C3",X"86",X"0C",X"CD",X"99",X"0C",X"CA",X"7A",
		X"09",X"CD",X"A9",X"0C",X"CD",X"F0",X"0B",X"22",X"B3",X"49",X"31",X"AB",X"49",X"F1",X"C1",X"D1",
		X"E1",X"22",X"A0",X"49",X"F9",X"21",X"08",X"00",X"E5",X"2A",X"B3",X"49",X"E5",X"2A",X"B5",X"49",
		X"C9",X"CD",X"C4",X"0B",X"D1",X"E1",X"E5",X"19",X"CD",X"74",X"0B",X"E1",X"E5",X"CD",X"BA",X"0C",
		X"CD",X"77",X"0B",X"E1",X"CD",X"B9",X"0C",X"C3",X"53",X"0C",X"CD",X"F0",X"0B",X"7D",X"B7",X"CA",
		X"ED",X"0D",X"87",X"85",X"87",X"C6",X"05",X"FE",X"4D",X"DA",X"BE",X"09",X"3E",X"4D",X"32",X"A4",
		X"49",X"C9",X"CD",X"C0",X"0B",X"C1",X"D1",X"E1",X"79",X"95",X"78",X"9C",X"D2",X"E8",X"09",X"CD",
		X"DB",X"09",X"D8",X"03",X"CD",X"7F",X"0B",X"D2",X"CF",X"09",X"C9",X"7E",X"02",X"E5",X"C5",X"60",
		X"69",X"4F",X"CD",X"AA",X"0B",X"C1",X"E1",X"C9",X"D5",X"C5",X"CD",X"B9",X"0C",X"EB",X"DA",X"ED",
		X"0D",X"E1",X"19",X"E5",X"C1",X"E1",X"CD",X"DB",X"09",X"D8",X"2B",X"0B",X"7B",X"B2",X"1B",X"C2",
		X"F6",X"09",X"C9",X"21",X"00",X"00",X"CD",X"99",X"0C",X"CA",X"23",X"0A",X"D6",X"30",X"DA",X"ED",
		X"0D",X"FE",X"0A",X"D2",X"ED",X"0D",X"E5",X"D1",X"29",X"29",X"19",X"29",X"5F",X"16",X"00",X"19",
		X"C3",X"06",X"0A",X"CD",X"7A",X"0B",X"C3",X"77",X"0B",X"CD",X"F0",X"0B",X"CD",X"7A",X"0B",X"11",
		X"F0",X"D8",X"CD",X"4A",X"0A",X"11",X"18",X"FC",X"CD",X"4A",X"0A",X"11",X"9C",X"FF",X"CD",X"4A",
		X"0A",X"11",X"F6",X"FF",X"CD",X"4A",X"0A",X"11",X"FF",X"FF",X"AF",X"E5",X"19",X"D2",X"55",X"0A",
		X"C1",X"3C",X"C3",X"4B",X"0A",X"E1",X"C3",X"61",X"0C",X"CD",X"F0",X"0B",X"CD",X"74",X"0B",X"7E",
		X"CD",X"58",X"0C",X"CD",X"89",X"0B",X"DA",X"79",X"0A",X"CA",X"79",X"0A",X"E5",X"CD",X"C2",X"0B",
		X"50",X"C1",X"E1",X"71",X"CD",X"AA",X"0B",X"D8",X"7A",X"FE",X"2E",X"C8",X"FE",X"0D",X"23",X"CA",
		X"5C",X"0A",X"FE",X"08",X"2B",X"2B",X"CA",X"5C",X"0A",X"C3",X"ED",X"0D",X"CD",X"99",X"0C",X"21",
		X"9F",X"0F",X"CA",X"F3",X"0A",X"BE",X"CA",X"B4",X"0A",X"57",X"7E",X"B7",X"FA",X"ED",X"0D",X"23",
		X"23",X"23",X"23",X"7A",X"C3",X"95",X"0A",X"FE",X"4D",X"C0",X"E3",X"23",X"E3",X"E5",X"2A",X"B5",
		X"49",X"7E",X"E1",X"C9",X"7E",X"F5",X"CD",X"19",X"0B",X"F1",X"CD",X"A7",X"0A",X"1A",X"CD",X"58",
		X"0C",X"05",X"CA",X"CA",X"0A",X"1B",X"1A",X"CD",X"58",X"0C",X"04",X"CD",X"89",X"0B",X"4F",X"DA",
		X"E9",X"0A",X"CA",X"E9",X"0A",X"E5",X"D5",X"C5",X"CD",X"F0",X"0B",X"78",X"C1",X"D1",X"4F",X"7D",
		X"12",X"05",X"CA",X"E8",X"0A",X"13",X"7C",X"12",X"E1",X"7E",X"B7",X"F8",X"79",X"FE",X"0D",X"CA",
		X"B4",X"0A",X"C9",X"CD",X"19",X"0B",X"F8",X"CD",X"A7",X"0A",X"1A",X"CD",X"58",X"0C",X"05",X"CA",
		X"0A",X"0B",X"1B",X"1A",X"CD",X"58",X"0C",X"C3",X"F3",X"0A",X"CD",X"7A",X"0B",X"CD",X"1C",X"0B",
		X"F8",X"FE",X"50",X"CA",X"FA",X"0A",X"C3",X"03",X"0B",X"CD",X"31",X"0D",X"7E",X"B7",X"F8",X"CD",
		X"B3",X"0C",X"46",X"23",X"CD",X"37",X"0C",X"0E",X"3D",X"C3",X"67",X"0C",X"CD",X"F5",X"0B",X"C2",
		X"35",X"0B",X"21",X"00",X"00",X"46",X"23",X"7C",X"B5",X"C8",X"7E",X"BB",X"C2",X"35",X"0B",X"23",
		X"7E",X"2B",X"BA",X"C2",X"35",X"0B",X"3E",X"02",X"CD",X"93",X"0C",X"CD",X"77",X"0B",X"78",X"CD",
		X"8D",X"0C",X"CD",X"52",X"0C",X"EB",X"CD",X"3E",X"0C",X"D8",X"C3",X"35",X"0B",X"CD",X"C4",X"0B",
		X"D1",X"E1",X"01",X"00",X"00",X"7E",X"81",X"4F",X"D2",X"6C",X"0B",X"04",X"CD",X"7F",X"0B",X"D2",
		X"65",X"0B",X"60",X"69",X"CD",X"31",X"0D",X"CD",X"53",X"0C",X"3E",X"20",X"C3",X"37",X"0C",X"23",
		X"7C",X"B5",X"37",X"C8",X"7B",X"95",X"7A",X"9C",X"C9",X"3E",X"2D",X"CD",X"37",X"0C",X"CD",X"CC",
		X"0C",X"CD",X"A9",X"0C",X"FE",X"20",X"C8",X"FE",X"2C",X"C8",X"FE",X"2E",X"C8",X"FE",X"3F",X"C8",
		X"FE",X"08",X"C8",X"FE",X"0D",X"37",X"3F",X"C0",X"37",X"C9",X"7E",X"47",X"B9",X"C8",X"3E",X"3F",
		X"CD",X"93",X"0C",X"CD",X"23",X"0A",X"79",X"CD",X"8D",X"0C",X"78",X"CD",X"58",X"0C",X"37",X"C9",
		X"0C",X"21",X"0E",X"01",X"21",X"00",X"00",X"CD",X"99",X"0C",X"47",X"CD",X"02",X"0C",X"DA",X"DA",
		X"0B",X"29",X"29",X"29",X"29",X"B5",X"6F",X"C3",X"C7",X"0B",X"E3",X"E5",X"78",X"CD",X"94",X"0B",
		X"D2",X"E8",X"0B",X"0D",X"C2",X"ED",X"0D",X"C9",X"C2",X"ED",X"0D",X"0D",X"C2",X"C4",X"0B",X"C9",
		X"CD",X"C2",X"0B",X"E1",X"C9",X"CD",X"C2",X"0B",X"D1",X"78",X"FE",X"0D",X"C8",X"CD",X"F0",X"0B",
		X"0D",X"C9",X"D6",X"30",X"D8",X"C6",X"E9",X"D8",X"C6",X"06",X"F2",X"10",X"0C",X"C6",X"07",X"D8",
		X"C6",X"0A",X"B7",X"C9",X"E6",X"0F",X"FE",X"0A",X"FA",X"1D",X"0C",X"C6",X"07",X"C6",X"30",X"C9",
		X"CD",X"56",X"09",X"FE",X"08",X"DA",X"37",X"0C",X"FE",X"1F",X"D8",X"FE",X"61",X"FA",X"37",X"0C",
		X"FE",X"7B",X"F2",X"37",X"0C",X"D6",X"20",X"C5",X"4F",X"CD",X"67",X"0C",X"C1",X"C9",X"CD",X"E7",
		X"07",X"C8",X"CD",X"59",X"09",X"FE",X"0D",X"37",X"C8",X"CD",X"56",X"09",X"FE",X"0D",X"37",X"C8",
		X"B7",X"C9",X"EB",X"7C",X"CD",X"58",X"0C",X"7D",X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",X"61",X"0C",
		X"F1",X"CD",X"14",X"0C",X"C3",X"37",X"0C",X"F5",X"C5",X"D5",X"E5",X"2A",X"A6",X"49",X"3E",X"44",
		X"BD",X"DC",X"31",X"0D",X"3A",X"FF",X"5F",X"B7",X"C4",X"A8",X"49",X"2A",X"A6",X"49",X"EB",X"CD",
		X"5B",X"05",X"EB",X"22",X"A6",X"49",X"E1",X"D1",X"C1",X"F1",X"C9",X"7E",X"23",X"CD",X"58",X"0C",
		X"C3",X"7A",X"0B",X"CD",X"31",X"0D",X"C3",X"37",X"0C",X"E5",X"2A",X"B9",X"49",X"7E",X"23",X"FE",
		X"20",X"CA",X"9D",X"0C",X"FE",X"0D",X"C3",X"AE",X"0C",X"E5",X"2A",X"B9",X"49",X"2B",X"22",X"B9",
		X"49",X"E1",X"C9",X"23",X"5E",X"23",X"56",X"23",X"C9",X"EB",X"7D",X"93",X"6F",X"7C",X"9A",X"67",
		X"C9",X"23",X"4E",X"23",X"46",X"23",X"78",X"B1",X"C9",X"37",X"3F",X"C9",X"E5",X"D5",X"C5",X"06",
		X"00",X"21",X"BB",X"49",X"22",X"B9",X"49",X"CD",X"20",X"0C",X"FE",X"18",X"CA",X"A7",X"08",X"FE",
		X"0D",X"CA",X"2A",X"0D",X"FE",X"08",X"CA",X"FA",X"0C",X"DA",X"F1",X"0C",X"FE",X"1F",X"DA",X"D7",
		X"0C",X"77",X"23",X"04",X"78",X"FE",X"1A",X"DA",X"D7",X"0C",X"05",X"FA",X"2A",X"0D",X"2B",X"E5",
		X"2A",X"A6",X"49",X"7C",X"FE",X"07",X"D2",X"12",X"0D",X"26",X"66",X"7D",X"D6",X"06",X"6F",X"C3",
		X"15",X"0D",X"D6",X"06",X"67",X"22",X"A6",X"49",X"AF",X"32",X"EE",X"5F",X"EB",X"3C",X"CD",X"5C",
		X"05",X"0E",X"03",X"CD",X"2E",X"06",X"E1",X"C3",X"D7",X"0C",X"77",X"CD",X"99",X"0C",X"C3",X"93",
		X"04",X"F5",X"C5",X"D5",X"E5",X"21",X"E0",X"48",X"3E",X"C0",X"36",X"00",X"23",X"3D",X"C2",X"3A",
		X"0D",X"21",X"A4",X"49",X"7E",X"B7",X"CC",X"BC",X"09",X"CD",X"B7",X"09",X"7E",X"D6",X"06",X"4F",
		X"3E",X"4D",X"96",X"6F",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"11",X"00",X"40",X"19",X"EB",
		X"21",X"C0",X"00",X"19",X"06",X"20",X"7E",X"12",X"23",X"13",X"05",X"C2",X"66",X"0D",X"0D",X"C2",
		X"64",X"0D",X"21",X"42",X"06",X"22",X"A6",X"49",X"C3",X"86",X"0C",X"CD",X"99",X"0C",X"C2",X"D4",
		X"0D",X"21",X"88",X"0D",X"22",X"F3",X"5F",X"C9",X"21",X"D0",X"5F",X"7E",X"B7",X"CA",X"72",X"01",
		X"23",X"7E",X"2B",X"FE",X"11",X"C2",X"9D",X"0D",X"AF",X"77",X"C3",X"A7",X"08",X"FE",X"10",X"C2",
		X"72",X"01",X"AF",X"77",X"3C",X"32",X"A5",X"49",X"F1",X"C1",X"D1",X"E1",X"C3",X"04",X"08",X"21",
		X"00",X"00",X"22",X"DD",X"5F",X"CD",X"99",X"0C",X"CA",X"C9",X"0D",X"CD",X"A9",X"0C",X"CD",X"C4",
		X"0B",X"E1",X"22",X"DF",X"5F",X"E1",X"22",X"DD",X"5F",X"01",X"01",X"01",X"11",X"00",X"00",X"CD",
		X"1C",X"02",X"F3",X"06",X"AF",X"B7",X"F5",X"2A",X"F3",X"5F",X"7C",X"B5",X"CA",X"EB",X"0D",X"22",
		X"A2",X"49",X"CD",X"74",X"0B",X"21",X"00",X"00",X"22",X"F3",X"5F",X"F1",X"C8",X"3E",X"3F",X"CD",
		X"93",X"0C",X"C3",X"A7",X"08",X"CD",X"99",X"0C",X"CA",X"20",X"0E",X"CD",X"A9",X"0C",X"CD",X"C4",
		X"0B",X"21",X"D5",X"49",X"11",X"07",X"00",X"72",X"19",X"36",X"FF",X"19",X"36",X"FD",X"D1",X"E1",
		X"22",X"DD",X"49",X"22",X"E1",X"49",X"CD",X"B9",X"0C",X"DA",X"ED",X"0D",X"23",X"22",X"DF",X"49",
		X"01",X"D5",X"49",X"F3",X"E5",X"D5",X"C5",X"60",X"69",X"CD",X"DD",X"02",X"01",X"00",X"06",X"CD",
		X"24",X"04",X"7E",X"FE",X"FC",X"CA",X"61",X"0E",X"32",X"D8",X"5F",X"CD",X"B3",X"0C",X"EB",X"22",
		X"D4",X"5F",X"EB",X"CD",X"B4",X"0C",X"EB",X"22",X"D6",X"5F",X"EB",X"CD",X"B4",X"0C",X"B7",X"CA",
		X"2C",X"0E",X"F5",X"D5",X"CD",X"A1",X"0E",X"D1",X"F1",X"FE",X"FD",X"C2",X"6E",X"0E",X"CD",X"30",
		X"04",X"01",X"FF",X"7F",X"CD",X"F6",X"07",X"CD",X"E3",X"02",X"FB",X"C3",X"93",X"04",X"FE",X"FE",
		X"C2",X"82",X"0E",X"0E",X"01",X"CD",X"E4",X"03",X"4B",X"CD",X"E4",X"03",X"01",X"80",X"00",X"C3",
		X"2F",X"0E",X"E5",X"2A",X"D6",X"5F",X"4D",X"44",X"E1",X"78",X"B7",X"C2",X"95",X"0E",X"B1",X"C4",
		X"A7",X"0E",X"C3",X"32",X"0E",X"C5",X"0E",X"00",X"CD",X"A7",X"0E",X"C1",X"05",X"14",X"C3",X"89",
		X"0E",X"01",X"05",X"00",X"11",X"D4",X"5F",X"E5",X"D5",X"C5",X"CD",X"E4",X"03",X"EB",X"C5",X"4E",
		X"CD",X"E4",X"03",X"C1",X"23",X"0D",X"C2",X"AE",X"0E",X"01",X"04",X"00",X"CD",X"24",X"04",X"C3",
		X"93",X"04",X"CD",X"F5",X"0B",X"CA",X"CB",X"0E",X"22",X"B7",X"49",X"EB",X"CD",X"3E",X"0C",X"D8",
		X"CD",X"74",X"0B",X"5E",X"23",X"CD",X"00",X"0F",X"CD",X"23",X"0F",X"FE",X"03",X"C2",X"E9",X"0E",
		X"CD",X"B4",X"0C",X"CD",X"52",X"0C",X"C3",X"CB",X"0E",X"FE",X"02",X"C2",X"CC",X"0E",X"56",X"CD",
		X"8B",X"0C",X"3E",X"3B",X"CD",X"37",X"0C",X"7A",X"E6",X"7F",X"CD",X"2B",X"0C",X"C3",X"CC",X"0E",
		X"E5",X"D5",X"2A",X"B7",X"49",X"7C",X"B5",X"CA",X"ED",X"0D",X"1C",X"7E",X"23",X"B7",X"F2",X"0B",
		X"0F",X"1D",X"C2",X"0B",X"0F",X"E6",X"7F",X"CD",X"37",X"0C",X"7E",X"23",X"B7",X"F2",X"17",X"0F",
		X"D1",X"E1",X"C9",X"E5",X"D5",X"16",X"01",X"3E",X"F3",X"BB",X"CA",X"44",X"0F",X"21",X"47",X"0F",
		X"14",X"23",X"7E",X"BB",X"CA",X"44",X"0F",X"FE",X"F3",X"C2",X"31",X"0F",X"3E",X"03",X"BA",X"C2",
		X"30",X"0F",X"16",X"01",X"7A",X"D1",X"E1",X"C9",X"06",X"0E",X"16",X"1E",X"26",X"2E",X"36",X"3E",
		X"C6",X"CE",X"D3",X"D6",X"DB",X"DE",X"E6",X"EE",X"F6",X"FE",X"F3",X"01",X"11",X"21",X"22",X"2A",
		X"31",X"32",X"3A",X"C2",X"C3",X"C4",X"CA",X"CC",X"CD",X"D2",X"D4",X"DA",X"DC",X"E2",X"E4",X"EA",
		X"EC",X"F2",X"F4",X"FA",X"FC",X"F3",X"06",X"00",X"21",X"00",X"40",X"7D",X"AC",X"A8",X"77",X"23",
		X"7C",X"FE",X"80",X"C2",X"7B",X"0F",X"21",X"00",X"40",X"7D",X"AC",X"A8",X"BE",X"C2",X"9B",X"0F",
		X"23",X"7C",X"FE",X"80",X"C2",X"89",X"0F",X"04",X"C3",X"78",X"0F",X"22",X"A2",X"49",X"C7",X"41",
		X"AC",X"49",X"01",X"46",X"AB",X"49",X"01",X"42",X"AE",X"49",X"01",X"43",X"AD",X"49",X"01",X"44",
		X"B0",X"49",X"01",X"45",X"AF",X"49",X"01",X"48",X"B6",X"49",X"01",X"4C",X"B5",X"49",X"01",X"4D",
		X"00",X"00",X"01",X"50",X"B4",X"49",X"02",X"53",X"B2",X"49",X"02",X"FF",X"00",X"07",X"06",X"03",
		X"00",X"02",X"26",X"1D",X"4D",X"4F",X"4E",X"49",X"54",X"45",X"55",X"52",X"00",X"FF",X"00",X"05",
		X"05",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"08",X"10",X"A0",X"40",X"02",X"30",X"0A",X"52",X"3A",
		X"52",X"45",X"44",X"45",X"4D",X"41",X"52",X"52",X"41",X"47",X"45",X"00",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
