library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu1_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu1_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7F",X"30",X"00",X"8E",X"00",X"00",X"4F",X"B7",X"30",X"00",X"B7",X"20",X"00",X"30",X"01",X"26",
		X"F5",X"86",X"44",X"1F",X"8B",X"8E",X"50",X"00",X"CC",X"00",X"00",X"ED",X"81",X"ED",X"81",X"8C",
		X"58",X"00",X"25",X"F7",X"B7",X"20",X"00",X"10",X"CE",X"50",X"00",X"B7",X"20",X"00",X"8E",X"40",
		X"00",X"CC",X"00",X"00",X"ED",X"81",X"ED",X"81",X"B7",X"20",X"00",X"8C",X"50",X"00",X"25",X"F4",
		X"B7",X"20",X"00",X"8E",X"57",X"40",X"BF",X"52",X"3A",X"BF",X"52",X"38",X"CC",X"FF",X"FF",X"ED",
		X"81",X"8C",X"57",X"7F",X"23",X"F9",X"B7",X"20",X"00",X"8E",X"57",X"80",X"BF",X"52",X"3C",X"BF",
		X"52",X"3E",X"B6",X"28",X"60",X"43",X"B7",X"57",X"33",X"43",X"C6",X"01",X"85",X"0F",X"27",X"06",
		X"5C",X"85",X"F0",X"27",X"01",X"5F",X"D7",X"8C",X"B6",X"30",X"00",X"43",X"B7",X"57",X"34",X"48",
		X"48",X"09",X"AB",X"48",X"09",X"AB",X"97",X"F6",X"CE",X"BC",X"00",X"D6",X"AB",X"58",X"EC",X"C5",
		X"97",X"B7",X"F7",X"57",X"CF",X"96",X"F6",X"48",X"09",X"AC",X"48",X"09",X"AC",X"48",X"09",X"AE",
		X"48",X"49",X"49",X"CE",X"BC",X"08",X"A6",X"C6",X"97",X"AA",X"B6",X"57",X"33",X"84",X"0F",X"48",
		X"8E",X"BC",X"0C",X"EC",X"86",X"DD",X"8D",X"B6",X"57",X"33",X"84",X"F0",X"12",X"44",X"44",X"44",
		X"8E",X"BC",X"0C",X"EC",X"86",X"DD",X"8F",X"B7",X"20",X"00",X"8E",X"57",X"A0",X"CE",X"BC",X"2C",
		X"EC",X"C1",X"ED",X"81",X"8C",X"57",X"BE",X"25",X"F7",X"7F",X"57",X"36",X"FC",X"BC",X"2D",X"FD",
		X"57",X"37",X"B7",X"20",X"00",X"4F",X"B7",X"3A",X"00",X"B7",X"38",X"00",X"97",X"00",X"B7",X"3C",
		X"00",X"97",X"02",X"B7",X"3E",X"00",X"B7",X"45",X"06",X"B7",X"28",X"00",X"BD",X"8F",X"C5",X"B7",
		X"20",X"00",X"B6",X"28",X"00",X"84",X"18",X"27",X"2F",X"7C",X"57",X"C5",X"8D",X"34",X"86",X"03",
		X"97",X"F6",X"8E",X"00",X"00",X"3D",X"B7",X"20",X"00",X"30",X"1F",X"26",X"F8",X"0A",X"F6",X"26",
		X"F1",X"BD",X"8F",X"C5",X"BD",X"8F",X"ED",X"4F",X"5F",X"BD",X"8F",X"0C",X"C6",X"02",X"BD",X"8F",
		X"0C",X"D6",X"8C",X"CB",X"03",X"BD",X"8F",X"0C",X"86",X"01",X"B7",X"30",X"00",X"1C",X"EF",X"7E",
		X"83",X"AF",X"8E",X"40",X"22",X"86",X"0F",X"97",X"F6",X"30",X"88",X"20",X"86",X"0D",X"97",X"F7",
		X"B7",X"20",X"00",X"1F",X"13",X"86",X"05",X"C6",X"0F",X"A7",X"C0",X"E7",X"C9",X"07",X"FF",X"4C",
		X"A7",X"C4",X"E7",X"C9",X"08",X"00",X"33",X"C8",X"1F",X"4C",X"A7",X"C0",X"E7",X"C9",X"07",X"FF",
		X"4C",X"A7",X"C4",X"E7",X"C9",X"08",X"00",X"30",X"02",X"0A",X"F7",X"26",X"D3",X"30",X"06",X"0A",
		X"F6",X"26",X"C6",X"8E",X"40",X"5C",X"CC",X"20",X"0F",X"A7",X"84",X"A7",X"01",X"E7",X"89",X"08",
		X"00",X"E7",X"89",X"08",X"01",X"30",X"88",X"20",X"8C",X"44",X"1C",X"25",X"EC",X"39",X"B7",X"20",
		X"00",X"4F",X"B7",X"30",X"00",X"B6",X"52",X"37",X"88",X"01",X"B7",X"52",X"37",X"8E",X"50",X"00",
		X"CE",X"51",X"78",X"86",X"2F",X"97",X"F6",X"B6",X"52",X"37",X"26",X"04",X"30",X"89",X"00",X"BC",
		X"B6",X"57",X"C8",X"26",X"14",X"EC",X"C4",X"ED",X"84",X"EC",X"42",X"C0",X"07",X"ED",X"02",X"30",
		X"04",X"33",X"44",X"0A",X"F6",X"26",X"EE",X"20",X"18",X"EC",X"C4",X"43",X"80",X"12",X"ED",X"84",
		X"EC",X"42",X"88",X"C0",X"53",X"C0",X"06",X"ED",X"02",X"30",X"04",X"33",X"44",X"0A",X"F6",X"26",
		X"E8",X"7C",X"57",X"C7",X"96",X"02",X"B7",X"3E",X"00",X"96",X"00",X"B7",X"3C",X"00",X"B6",X"45",
		X"06",X"B7",X"28",X"00",X"B6",X"57",X"C8",X"84",X"01",X"B7",X"30",X"04",X"B7",X"30",X"05",X"B6",
		X"28",X"00",X"43",X"B7",X"57",X"30",X"B6",X"28",X"40",X"43",X"B7",X"57",X"32",X"FC",X"57",X"C5",
		X"4A",X"27",X"07",X"81",X"03",X"26",X"09",X"7E",X"83",X"27",X"C0",X"02",X"C1",X"01",X"23",X"09",
		X"B6",X"28",X"20",X"43",X"B7",X"57",X"31",X"20",X"36",X"BE",X"57",X"CA",X"7A",X"57",X"CC",X"26",
		X"0D",X"30",X"02",X"BF",X"57",X"CA",X"EC",X"84",X"B7",X"57",X"31",X"F7",X"57",X"CC",X"B6",X"57",
		X"31",X"84",X"CF",X"F6",X"57",X"C7",X"C4",X"0F",X"26",X"02",X"8A",X"10",X"F6",X"52",X"B9",X"C1",
		X"30",X"27",X"07",X"F6",X"52",X"C9",X"C1",X"38",X"26",X"02",X"8A",X"20",X"B7",X"57",X"31",X"96",
		X"8C",X"10",X"26",X"00",X"B2",X"5F",X"B6",X"57",X"30",X"44",X"09",X"83",X"44",X"09",X"84",X"44",
		X"09",X"8B",X"BD",X"82",X"AF",X"BD",X"82",X"DA",X"BD",X"82",X"94",X"BD",X"82",X"FA",X"BD",X"83",
		X"02",X"7E",X"83",X"27",X"96",X"8B",X"84",X"07",X"81",X"01",X"26",X"3D",X"BD",X"91",X"FA",X"96",
		X"82",X"81",X"99",X"27",X"34",X"8B",X"01",X"19",X"97",X"82",X"86",X"05",X"7E",X"8F",X"0C",X"96",
		X"83",X"84",X"07",X"81",X"01",X"26",X"22",X"BD",X"91",X"FA",X"0C",X"87",X"0C",X"85",X"96",X"85",
		X"91",X"8D",X"26",X"15",X"86",X"05",X"BD",X"8F",X"0C",X"0F",X"85",X"96",X"8E",X"9B",X"82",X"19",
		X"25",X"03",X"97",X"82",X"39",X"86",X"99",X"97",X"82",X"39",X"96",X"84",X"84",X"07",X"81",X"01",
		X"26",X"F7",X"BD",X"91",X"FA",X"0C",X"89",X"0C",X"86",X"96",X"86",X"91",X"8F",X"26",X"EA",X"86",
		X"05",X"BD",X"8F",X"0C",X"0F",X"86",X"96",X"90",X"20",X"D3",X"8E",X"44",X"87",X"CE",X"30",X"02",
		X"20",X"06",X"8E",X"44",X"89",X"CE",X"30",X"01",X"6D",X"84",X"27",X"12",X"6A",X"01",X"A6",X"01",
		X"84",X"1F",X"27",X"0B",X"81",X"1F",X"27",X"0A",X"81",X"10",X"26",X"02",X"6F",X"C4",X"39",X"6A",
		X"84",X"39",X"86",X"01",X"A7",X"C4",X"39",X"BE",X"52",X"3E",X"BC",X"52",X"3C",X"27",X"13",X"A6",
		X"80",X"B7",X"3A",X"00",X"B7",X"38",X"00",X"8C",X"57",X"A0",X"25",X"03",X"8E",X"57",X"80",X"BF",
		X"52",X"3E",X"B6",X"57",X"C5",X"48",X"8E",X"BC",X"4A",X"AD",X"96",X"FC",X"52",X"35",X"10",X"83",
		X"FF",X"FF",X"26",X"1C",X"8E",X"BD",X"5E",X"C6",X"06",X"A6",X"80",X"AB",X"80",X"5A",X"26",X"FB",
		X"81",X"1B",X"27",X"0C",X"CC",X"00",X"52",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"20",X"22",
		X"B6",X"94",X"FA",X"81",X"35",X"27",X"0C",X"CC",X"00",X"52",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",
		X"0C",X"20",X"0F",X"B6",X"A8",X"FC",X"81",X"34",X"27",X"08",X"B6",X"57",X"C8",X"88",X"01",X"B7",
		X"57",X"C8",X"86",X"01",X"B7",X"30",X"00",X"3B",X"84",X"7F",X"CE",X"FF",X"FF",X"EF",X"81",X"8C",
		X"57",X"80",X"25",X"03",X"8E",X"57",X"40",X"BF",X"52",X"3A",X"8E",X"BC",X"54",X"AD",X"96",X"4F",
		X"BE",X"52",X"3A",X"EC",X"84",X"48",X"24",X"E0",X"20",X"F5",X"CC",X"20",X"20",X"8E",X"40",X"40",
		X"ED",X"81",X"8C",X"43",X"C0",X"26",X"F9",X"39",X"4F",X"8E",X"BC",X"6E",X"58",X"EE",X"8B",X"AE",
		X"C1",X"E6",X"C0",X"A6",X"C0",X"81",X"40",X"27",X"0B",X"A7",X"84",X"E7",X"89",X"08",X"00",X"30",
		X"88",X"E0",X"20",X"EF",X"39",X"4F",X"8E",X"BC",X"6E",X"58",X"EE",X"8B",X"AE",X"C1",X"33",X"41",
		X"A6",X"C0",X"81",X"40",X"27",X"0E",X"CC",X"20",X"0F",X"A7",X"84",X"E7",X"89",X"08",X"00",X"30",
		X"88",X"E0",X"20",X"EC",X"39",X"8E",X"57",X"36",X"CE",X"46",X"61",X"86",X"0F",X"97",X"F0",X"7E",
		X"8F",X"7E",X"B6",X"57",X"C5",X"81",X"03",X"26",X"1E",X"96",X"AF",X"26",X"0D",X"8E",X"57",X"39",
		X"CE",X"47",X"81",X"86",X"0F",X"97",X"F0",X"7E",X"8F",X"7E",X"8E",X"57",X"3C",X"CE",X"45",X"41",
		X"86",X"0F",X"97",X"F0",X"7E",X"8F",X"7E",X"39",X"86",X"0F",X"97",X"F0",X"8E",X"44",X"82",X"CE",
		X"44",X"7F",X"7E",X"8F",X"B4",X"B6",X"57",X"C5",X"81",X"03",X"26",X"52",X"CE",X"C2",X"7A",X"E6",
		X"C5",X"D7",X"91",X"CE",X"57",X"39",X"96",X"AF",X"27",X"02",X"33",X"43",X"A6",X"42",X"9B",X"91",
		X"19",X"A7",X"42",X"24",X"10",X"A6",X"41",X"8B",X"01",X"19",X"A7",X"41",X"24",X"07",X"A6",X"C4",
		X"8B",X"01",X"19",X"A7",X"C4",X"EC",X"C4",X"10",X"B3",X"57",X"36",X"27",X"0F",X"25",X"93",X"FD",
		X"57",X"36",X"A6",X"42",X"B7",X"57",X"38",X"BD",X"84",X"05",X"20",X"86",X"A6",X"42",X"B1",X"57",
		X"38",X"10",X"23",X"FF",X"7D",X"B7",X"57",X"38",X"BD",X"84",X"05",X"7E",X"84",X"12",X"39",X"8E",
		X"47",X"BE",X"4F",X"5A",X"26",X"02",X"86",X"20",X"A7",X"84",X"30",X"88",X"E0",X"8C",X"46",X"3E",
		X"24",X"F1",X"39",X"86",X"0F",X"97",X"F0",X"8E",X"44",X"E2",X"CE",X"46",X"FF",X"7E",X"8F",X"B4",
		X"8E",X"45",X"FE",X"CC",X"01",X"8F",X"A7",X"84",X"E7",X"89",X"08",X"00",X"CB",X"40",X"A7",X"01",
		X"E7",X"89",X"08",X"01",X"CB",X"40",X"A7",X"88",X"20",X"E7",X"89",X"08",X"20",X"CB",X"40",X"A7",
		X"88",X"21",X"E7",X"89",X"08",X"21",X"39",X"CE",X"C2",X"84",X"8E",X"C2",X"98",X"4F",X"B7",X"45",
		X"0B",X"48",X"EC",X"C6",X"B7",X"45",X"0C",X"86",X"21",X"58",X"49",X"FB",X"45",X"0B",X"CB",X"03",
		X"1F",X"02",X"A6",X"89",X"00",X"8B",X"A7",X"A9",X"08",X"00",X"A6",X"80",X"A7",X"A4",X"31",X"A8",
		X"E0",X"7A",X"45",X"0C",X"26",X"EC",X"7C",X"45",X"0B",X"B6",X"45",X"0B",X"81",X"0A",X"25",X"D1",
		X"39",X"7C",X"57",X"C9",X"39",X"B6",X"57",X"C9",X"8E",X"C3",X"AE",X"48",X"6E",X"96",X"B6",X"57",
		X"C8",X"26",X"04",X"B6",X"57",X"31",X"39",X"B6",X"57",X"32",X"39",X"0F",X"AF",X"5F",X"B6",X"57",
		X"C5",X"4A",X"26",X"05",X"F6",X"57",X"CD",X"58",X"5C",X"4F",X"FD",X"57",X"E1",X"5F",X"DD",X"1A",
		X"DD",X"1C",X"FD",X"57",X"39",X"FD",X"57",X"3B",X"FD",X"57",X"3D",X"97",X"DD",X"97",X"E5",X"B7",
		X"57",X"E4",X"FD",X"57",X"E5",X"FD",X"57",X"E7",X"FD",X"57",X"E9",X"FD",X"57",X"EB",X"FD",X"57",
		X"ED",X"DD",X"36",X"DD",X"38",X"FD",X"52",X"35",X"8E",X"00",X"00",X"CE",X"44",X"42",X"C6",X"0C",
		X"BD",X"8C",X"DA",X"B6",X"57",X"CF",X"B7",X"57",X"E3",X"96",X"AA",X"B7",X"57",X"E0",X"86",X"10",
		X"B7",X"57",X"EF",X"CE",X"C3",X"D2",X"96",X"AC",X"97",X"F6",X"48",X"9B",X"F6",X"33",X"C6",X"A6",
		X"C4",X"97",X"B1",X"EC",X"41",X"DD",X"B2",X"4F",X"5F",X"BD",X"8F",X"0C",X"86",X"04",X"BD",X"8F",
		X"0C",X"B6",X"57",X"C5",X"4A",X"27",X"77",X"96",X"B0",X"27",X"3F",X"CC",X"00",X"01",X"BD",X"8F",
		X"0C",X"0C",X"AF",X"86",X"04",X"BD",X"8F",X"0C",X"0F",X"AF",X"CC",X"30",X"0F",X"97",X"61",X"97",
		X"81",X"F7",X"4C",X"61",X"F7",X"4C",X"81",X"8E",X"57",X"E0",X"CE",X"57",X"F0",X"C6",X"10",X"BD",
		X"8C",X"E0",X"8E",X"00",X"00",X"CE",X"44",X"62",X"C6",X"0C",X"BD",X"8C",X"DA",X"96",X"B1",X"97",
		X"B4",X"DC",X"B2",X"DD",X"B5",X"CC",X"20",X"0F",X"20",X"13",X"CC",X"01",X"01",X"BD",X"8F",X"0C",
		X"CC",X"20",X"0F",X"97",X"61",X"97",X"81",X"F7",X"4C",X"61",X"F7",X"4C",X"81",X"97",X"A1",X"97",
		X"C1",X"97",X"E1",X"B7",X"45",X"01",X"B7",X"45",X"21",X"B7",X"45",X"41",X"F7",X"4C",X"A1",X"F7",
		X"4C",X"C1",X"F7",X"4C",X"E1",X"F7",X"4D",X"01",X"F7",X"4D",X"21",X"F7",X"4D",X"41",X"B6",X"57",
		X"C5",X"4A",X"10",X"26",X"FE",X"EB",X"86",X"01",X"B7",X"57",X"E0",X"B6",X"57",X"CD",X"26",X"1C",
		X"CC",X"03",X"04",X"97",X"48",X"D7",X"4A",X"CC",X"05",X"03",X"B7",X"57",X"E6",X"F7",X"57",X"E2",
		X"CC",X"0D",X"19",X"B7",X"57",X"E3",X"F7",X"57",X"EE",X"7E",X"85",X"21",X"CC",X"01",X"0B",X"97",
		X"48",X"F7",X"57",X"E3",X"CC",X"06",X"05",X"B7",X"57",X"E1",X"F7",X"57",X"E2",X"CC",X"10",X"08",
		X"FD",X"57",X"EB",X"CC",X"00",X"01",X"DD",X"42",X"97",X"E7",X"B7",X"57",X"3F",X"C3",X"02",X"02",
		X"DD",X"44",X"C3",X"02",X"02",X"DD",X"46",X"7E",X"85",X"21",X"4F",X"97",X"DA",X"97",X"DD",X"97",
		X"E5",X"B7",X"4C",X"00",X"97",X"E7",X"86",X"0A",X"BD",X"8F",X"0C",X"BD",X"90",X"35",X"7E",X"85",
		X"21",X"4F",X"5F",X"DD",X"E9",X"DD",X"D8",X"DD",X"EB",X"97",X"F5",X"CE",X"57",X"D0",X"8E",X"57",
		X"E0",X"96",X"AF",X"27",X"03",X"8E",X"57",X"F0",X"C6",X"10",X"BD",X"8C",X"E0",X"CE",X"44",X"14",
		X"8E",X"44",X"42",X"96",X"AF",X"27",X"03",X"8E",X"44",X"62",X"C6",X"18",X"BD",X"8C",X"E0",X"B6",
		X"57",X"D1",X"8B",X"01",X"19",X"97",X"E2",X"B6",X"57",X"C5",X"4A",X"27",X"0B",X"CC",X"00",X"19",
		X"BD",X"8F",X"0C",X"86",X"09",X"BD",X"8F",X"0C",X"7E",X"85",X"21",X"7F",X"57",X"C8",X"96",X"AE",
		X"26",X"07",X"96",X"AF",X"27",X"03",X"7C",X"57",X"C8",X"CC",X"04",X"00",X"FD",X"57",X"C2",X"4F",
		X"FD",X"57",X"C0",X"BD",X"92",X"99",X"BD",X"A9",X"4E",X"CC",X"A5",X"08",X"8E",X"4E",X"80",X"CE",
		X"51",X"B8",X"36",X"16",X"80",X"03",X"81",X"78",X"24",X"F8",X"BD",X"92",X"6C",X"86",X"40",X"B7",
		X"57",X"CE",X"F6",X"57",X"D0",X"5C",X"86",X"07",X"BD",X"8F",X"0C",X"BD",X"8C",X"6A",X"7E",X"85",
		X"21",X"BD",X"93",X"0D",X"BD",X"A9",X"D9",X"7A",X"57",X"CE",X"27",X"1A",X"B6",X"57",X"CE",X"85",
		X"0F",X"26",X"12",X"44",X"44",X"44",X"44",X"8B",X"3F",X"8E",X"51",X"7A",X"A7",X"84",X"30",X"04",
		X"8C",X"51",X"B8",X"25",X"F7",X"39",X"86",X"01",X"B7",X"57",X"C2",X"86",X"10",X"B7",X"57",X"CE",
		X"BD",X"95",X"F8",X"86",X"01",X"97",X"99",X"96",X"9B",X"97",X"9C",X"B6",X"57",X"C5",X"4A",X"26",
		X"09",X"B6",X"57",X"D6",X"26",X"04",X"86",X"04",X"97",X"97",X"7E",X"85",X"21",X"BD",X"93",X"0D",
		X"BD",X"A9",X"D9",X"7A",X"57",X"CE",X"27",X"0B",X"B6",X"57",X"CE",X"48",X"48",X"8E",X"51",X"7B",
		X"6F",X"86",X"39",X"F6",X"57",X"D0",X"86",X"07",X"BD",X"8F",X"0C",X"BD",X"AD",X"31",X"BD",X"91",
		X"F2",X"86",X"30",X"B7",X"57",X"CE",X"7E",X"85",X"21",X"BD",X"AD",X"57",X"BD",X"93",X"0D",X"0F",
		X"EF",X"BD",X"AE",X"5F",X"BD",X"A9",X"D9",X"7A",X"57",X"CE",X"27",X"01",X"39",X"BD",X"90",X"78",
		X"7A",X"57",X"CE",X"CC",X"02",X"00",X"DD",X"2C",X"F7",X"52",X"34",X"7E",X"85",X"21",X"BD",X"B1",
		X"15",X"BD",X"94",X"F2",X"BD",X"AD",X"57",X"BD",X"93",X"0D",X"BD",X"A8",X"E6",X"BD",X"96",X"45",
		X"BD",X"9A",X"A1",X"BD",X"A0",X"A9",X"BD",X"AE",X"5F",X"BD",X"A9",X"D9",X"BD",X"A7",X"C6",X"BD",
		X"A7",X"7C",X"BD",X"90",X"86",X"B6",X"52",X"40",X"4C",X"10",X"27",X"00",X"C6",X"4A",X"26",X"BC",
		X"BD",X"91",X"F6",X"4F",X"5F",X"DD",X"E9",X"97",X"CC",X"B7",X"52",X"34",X"B7",X"4C",X"00",X"7A",
		X"57",X"D3",X"B6",X"57",X"C4",X"27",X"54",X"96",X"AF",X"26",X"06",X"D7",X"36",X"D7",X"38",X"20",
		X"04",X"D7",X"37",X"D7",X"39",X"4F",X"FD",X"57",X"D9",X"FD",X"57",X"DB",X"FD",X"57",X"DD",X"B7",
		X"57",X"D4",X"B7",X"57",X"C4",X"B6",X"57",X"D2",X"4C",X"81",X"06",X"25",X"01",X"4F",X"B7",X"57",
		X"D2",X"86",X"01",X"F6",X"57",X"D5",X"54",X"24",X"01",X"40",X"BB",X"57",X"D6",X"B7",X"57",X"D6",
		X"27",X"04",X"81",X"05",X"26",X"03",X"7C",X"57",X"D5",X"B6",X"57",X"D1",X"81",X"99",X"25",X"02",
		X"86",X"98",X"8B",X"01",X"19",X"B7",X"57",X"D1",X"BD",X"91",X"30",X"7A",X"57",X"D0",X"8E",X"57",
		X"D0",X"CE",X"57",X"E0",X"96",X"AF",X"27",X"03",X"CE",X"57",X"F0",X"C6",X"10",X"BD",X"8C",X"E0",
		X"8E",X"44",X"14",X"CE",X"44",X"42",X"96",X"AF",X"27",X"03",X"CE",X"44",X"62",X"C6",X"18",X"BD",
		X"8C",X"E0",X"B6",X"57",X"D0",X"27",X"21",X"96",X"AF",X"26",X"07",X"B6",X"57",X"F0",X"27",X"0D",
		X"20",X"05",X"B6",X"57",X"E0",X"27",X"06",X"96",X"AF",X"88",X"01",X"97",X"AF",X"4F",X"5F",X"DD",
		X"00",X"DD",X"02",X"4C",X"B7",X"57",X"C9",X"39",X"BD",X"90",X"35",X"86",X"28",X"B7",X"57",X"CE",
		X"7E",X"85",X"21",X"B6",X"57",X"C4",X"27",X"39",X"CC",X"00",X"00",X"97",X"EF",X"DD",X"E9",X"B7",
		X"52",X"34",X"B7",X"57",X"C4",X"FD",X"57",X"D9",X"FD",X"57",X"DB",X"FD",X"57",X"DD",X"B7",X"57",
		X"D4",X"B7",X"4C",X"00",X"BD",X"91",X"F6",X"8E",X"57",X"D0",X"CE",X"57",X"E0",X"96",X"AF",X"27",
		X"03",X"CE",X"57",X"F0",X"C6",X"10",X"BD",X"8C",X"E0",X"7F",X"57",X"CE",X"86",X"0E",X"B7",X"57",
		X"C9",X"39",X"BD",X"93",X"0D",X"7A",X"57",X"CE",X"26",X"08",X"86",X"0A",X"BD",X"8F",X"0C",X"7E",
		X"85",X"21",X"39",X"BD",X"91",X"EF",X"4F",X"5F",X"DD",X"00",X"DD",X"02",X"B7",X"3C",X"00",X"B7",
		X"3E",X"00",X"F6",X"57",X"C5",X"5A",X"27",X"1E",X"C6",X"0F",X"F7",X"45",X"06",X"C6",X"18",X"BD",
		X"8F",X"0C",X"C6",X"27",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"BD",X"92",X"85",X"86",X"80",
		X"B7",X"57",X"CE",X"7E",X"85",X"21",X"86",X"0D",X"B7",X"57",X"C9",X"39",X"96",X"82",X"27",X"2B",
		X"96",X"AF",X"26",X"07",X"B6",X"57",X"F0",X"26",X"22",X"20",X"05",X"B6",X"57",X"E0",X"26",X"1B",
		X"96",X"82",X"4A",X"26",X"09",X"B6",X"57",X"30",X"84",X"08",X"27",X"0F",X"20",X"07",X"B6",X"57",
		X"30",X"84",X"18",X"27",X"06",X"86",X"0D",X"B7",X"57",X"C9",X"39",X"7A",X"57",X"CE",X"27",X"22",
		X"B6",X"57",X"CE",X"81",X"60",X"25",X"1A",X"85",X"07",X"26",X"16",X"12",X"44",X"44",X"44",X"40",
		X"8B",X"2A",X"1F",X"89",X"8E",X"4B",X"34",X"ED",X"84",X"30",X"88",X"E0",X"8C",X"48",X"D4",X"24",
		X"F6",X"39",X"CC",X"01",X"18",X"BD",X"8F",X"0C",X"C6",X"27",X"BD",X"83",X"E5",X"C6",X"28",X"BD",
		X"83",X"E5",X"BD",X"90",X"BA",X"96",X"B9",X"26",X"08",X"86",X"0C",X"B7",X"57",X"C9",X"7E",X"8A",
		X"CC",X"BD",X"92",X"71",X"BD",X"8F",X"20",X"7E",X"85",X"21",X"96",X"82",X"27",X"2B",X"96",X"AF",
		X"26",X"07",X"B6",X"57",X"F0",X"26",X"22",X"20",X"05",X"B6",X"57",X"E0",X"26",X"1B",X"96",X"82",
		X"4A",X"26",X"09",X"B6",X"57",X"30",X"84",X"08",X"27",X"0F",X"20",X"07",X"B6",X"57",X"30",X"84",
		X"18",X"27",X"06",X"86",X"0D",X"B7",X"57",X"C9",X"39",X"96",X"C3",X"84",X"0F",X"44",X"8B",X"0A",
		X"97",X"F6",X"9E",X"C2",X"DE",X"C4",X"96",X"BC",X"4C",X"26",X"08",X"86",X"41",X"A7",X"C4",X"86",
		X"01",X"97",X"BC",X"B6",X"57",X"C7",X"44",X"24",X"29",X"0C",X"BD",X"D6",X"BD",X"86",X"0F",X"C4",
		X"04",X"26",X"02",X"96",X"F6",X"C6",X"08",X"A7",X"89",X"08",X"00",X"30",X"88",X"E0",X"5A",X"26",
		X"F6",X"A7",X"C9",X"08",X"00",X"B6",X"57",X"C7",X"4C",X"26",X"06",X"0A",X"BB",X"10",X"27",X"00",
		X"85",X"39",X"BD",X"85",X"2E",X"44",X"09",X"C8",X"44",X"09",X"C9",X"44",X"44",X"44",X"09",X"CA",
		X"10",X"8E",X"C3",X"DE",X"96",X"CA",X"84",X"07",X"4A",X"27",X"40",X"96",X"C9",X"81",X"FF",X"26",
		X"04",X"0F",X"C9",X"20",X"05",X"84",X"07",X"4A",X"27",X"1B",X"96",X"C8",X"81",X"FF",X"26",X"04",
		X"0F",X"C8",X"20",X"C1",X"84",X"07",X"4A",X"26",X"BC",X"0A",X"BC",X"D6",X"BC",X"2A",X"11",X"C6",
		X"1B",X"D7",X"BC",X"20",X"0B",X"0C",X"BC",X"D6",X"BC",X"C1",X"1B",X"23",X"03",X"5F",X"D7",X"BC",
		X"A6",X"A5",X"A7",X"C4",X"C6",X"0F",X"E7",X"C9",X"08",X"00",X"39",X"BD",X"92",X"7B",X"9E",X"C6",
		X"D6",X"BC",X"A6",X"A5",X"A7",X"80",X"D6",X"F6",X"E7",X"C9",X"08",X"00",X"33",X"C8",X"E0",X"11",
		X"83",X"40",X"F0",X"25",X"11",X"86",X"41",X"A7",X"C4",X"86",X"08",X"97",X"BB",X"86",X"01",X"97",
		X"BC",X"9F",X"C6",X"DF",X"C4",X"39",X"BD",X"92",X"76",X"7E",X"85",X"21",X"96",X"AF",X"26",X"08",
		X"B6",X"57",X"F0",X"27",X"0B",X"7E",X"88",X"A7",X"B6",X"57",X"E0",X"27",X"03",X"7E",X"88",X"A7",
		X"7E",X"85",X"21",X"39",X"4F",X"B7",X"57",X"C8",X"B7",X"57",X"C6",X"97",X"AF",X"86",X"01",X"B7",
		X"57",X"C5",X"7E",X"8F",X"ED",X"FC",X"51",X"79",X"DD",X"94",X"BD",X"90",X"35",X"DC",X"1A",X"FD",
		X"45",X"07",X"DC",X"1C",X"FD",X"45",X"09",X"FC",X"57",X"C0",X"FD",X"45",X"02",X"FC",X"57",X"C2",
		X"FD",X"45",X"04",X"BD",X"92",X"67",X"5F",X"96",X"AF",X"26",X"06",X"D7",X"36",X"D7",X"38",X"20",
		X"04",X"D7",X"37",X"D7",X"39",X"7E",X"85",X"21",X"BD",X"93",X"0D",X"B6",X"57",X"CE",X"81",X"F0",
		X"22",X"7E",X"25",X"0E",X"4F",X"5F",X"8E",X"51",X"78",X"ED",X"81",X"8C",X"51",X"B8",X"25",X"F9",
		X"20",X"6E",X"8E",X"51",X"78",X"B6",X"57",X"CE",X"44",X"25",X"1A",X"D6",X"95",X"C4",X"F0",X"96",
		X"D6",X"CE",X"C3",X"FA",X"EB",X"C6",X"D7",X"95",X"CC",X"80",X"78",X"A7",X"03",X"0F",X"F6",X"E7",
		X"84",X"0F",X"F7",X"20",X"26",X"CC",X"80",X"00",X"B3",X"57",X"C0",X"B3",X"57",X"C0",X"B3",X"57",
		X"C0",X"B3",X"57",X"C0",X"A7",X"03",X"D7",X"F6",X"CC",X"78",X"00",X"B3",X"57",X"C2",X"B3",X"57",
		X"C2",X"B3",X"57",X"C2",X"B3",X"57",X"C2",X"A7",X"84",X"D7",X"F7",X"DC",X"94",X"ED",X"01",X"A6",
		X"03",X"D6",X"F6",X"F3",X"57",X"C0",X"A7",X"07",X"D7",X"F6",X"A6",X"84",X"D6",X"F7",X"F3",X"57",
		X"C2",X"A7",X"04",X"D7",X"F7",X"DC",X"94",X"ED",X"05",X"30",X"04",X"8C",X"51",X"B4",X"25",X"DF",
		X"7C",X"57",X"CE",X"26",X"12",X"FC",X"45",X"07",X"DD",X"1A",X"FC",X"45",X"09",X"DD",X"1C",X"86",
		X"0A",X"BD",X"8F",X"0C",X"7E",X"85",X"21",X"39",X"96",X"AF",X"26",X"49",X"B6",X"57",X"E1",X"81",
		X"99",X"25",X"02",X"86",X"98",X"8B",X"01",X"19",X"B7",X"57",X"E1",X"B6",X"57",X"E2",X"4C",X"81",
		X"06",X"25",X"01",X"4F",X"B7",X"57",X"E2",X"B6",X"57",X"E1",X"B7",X"57",X"D1",X"BD",X"91",X"30",
		X"8E",X"44",X"14",X"CE",X"44",X"42",X"C6",X"18",X"BD",X"8C",X"E0",X"86",X"01",X"F6",X"57",X"E5",
		X"54",X"24",X"01",X"40",X"BB",X"57",X"E6",X"B7",X"57",X"E6",X"27",X"04",X"81",X"05",X"26",X"4C",
		X"7C",X"57",X"E5",X"20",X"47",X"B6",X"57",X"F1",X"81",X"99",X"25",X"02",X"86",X"98",X"8B",X"01",
		X"19",X"B7",X"57",X"F1",X"B6",X"57",X"F2",X"4C",X"81",X"06",X"25",X"01",X"4F",X"B7",X"57",X"F2",
		X"B6",X"57",X"F1",X"B7",X"57",X"D1",X"BD",X"91",X"30",X"8E",X"44",X"14",X"CE",X"44",X"62",X"C6",
		X"18",X"BD",X"8C",X"E0",X"86",X"01",X"F6",X"57",X"F5",X"54",X"24",X"01",X"40",X"BB",X"57",X"F6",
		X"B7",X"57",X"F6",X"27",X"04",X"81",X"05",X"26",X"03",X"7C",X"57",X"F5",X"CC",X"00",X"00",X"FD",
		X"57",X"C0",X"4C",X"FD",X"57",X"C2",X"B7",X"57",X"C9",X"39",X"CE",X"51",X"EC",X"86",X"03",X"97",
		X"F6",X"CC",X"4A",X"43",X"DD",X"F7",X"CC",X"60",X"90",X"DD",X"F9",X"8D",X"44",X"CC",X"4A",X"44",
		X"DD",X"F7",X"CC",X"73",X"98",X"DD",X"F9",X"86",X"03",X"97",X"F6",X"8D",X"34",X"86",X"02",X"97",
		X"F6",X"CC",X"4D",X"43",X"DD",X"F7",X"86",X"98",X"97",X"F9",X"86",X"90",X"D6",X"AF",X"27",X"04",
		X"86",X"88",X"0C",X"F8",X"97",X"FA",X"8D",X"19",X"B6",X"57",X"C5",X"4A",X"27",X"04",X"96",X"B0",
		X"26",X"0E",X"CE",X"51",X"ED",X"86",X"FF",X"C6",X"08",X"A7",X"C4",X"33",X"44",X"5A",X"26",X"F9",
		X"39",X"DC",X"F9",X"A7",X"43",X"E7",X"C4",X"DC",X"F7",X"ED",X"41",X"0C",X"F7",X"86",X"10",X"9B",
		X"F9",X"97",X"F9",X"33",X"44",X"0A",X"F6",X"26",X"E8",X"39",X"AF",X"C1",X"5A",X"26",X"FB",X"39",
		X"A6",X"80",X"A7",X"C0",X"5A",X"26",X"F9",X"39",X"7C",X"57",X"C5",X"7F",X"57",X"C6",X"39",X"7C",
		X"57",X"C6",X"39",X"B6",X"57",X"C6",X"8E",X"C4",X"02",X"48",X"AD",X"96",X"96",X"8C",X"27",X"06",
		X"4A",X"26",X"07",X"7E",X"8E",X"C9",X"96",X"82",X"26",X"DE",X"39",X"86",X"0E",X"B7",X"45",X"06",
		X"86",X"0C",X"BD",X"8F",X"0C",X"8E",X"C4",X"0E",X"CE",X"51",X"78",X"10",X"8E",X"52",X"40",X"CC",
		X"FF",X"40",X"ED",X"41",X"EC",X"81",X"A7",X"43",X"E7",X"C4",X"A6",X"80",X"A7",X"A0",X"33",X"44",
		X"11",X"83",X"51",X"AC",X"25",X"E9",X"CC",X"00",X"20",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",
		X"C6",X"06",X"BD",X"8F",X"0C",X"86",X"03",X"BD",X"8F",X"0C",X"4C",X"BD",X"8F",X"0C",X"D6",X"8C",
		X"26",X"04",X"4C",X"BD",X"8F",X"0C",X"CC",X"30",X"0F",X"B7",X"45",X"81",X"B7",X"45",X"A1",X"B7",
		X"46",X"A1",X"B7",X"46",X"C1",X"F7",X"4D",X"81",X"F7",X"4D",X"A1",X"F7",X"4E",X"A1",X"F7",X"4E",
		X"C1",X"BD",X"8F",X"20",X"7F",X"57",X"CE",X"7E",X"8E",X"9B",X"7A",X"57",X"CE",X"27",X"5B",X"B6",
		X"57",X"CE",X"81",X"A0",X"26",X"1A",X"CC",X"00",X"1A",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",
		X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",
		X"8E",X"52",X"40",X"CE",X"51",X"78",X"A6",X"80",X"2B",X"27",X"4A",X"A7",X"1F",X"81",X"30",X"22",
		X"20",X"26",X"10",X"11",X"83",X"51",X"8C",X"25",X"05",X"BD",X"92",X"16",X"20",X"03",X"BD",X"92",
		X"1A",X"86",X"30",X"85",X"07",X"26",X"0A",X"44",X"44",X"44",X"27",X"02",X"8B",X"55",X"4A",X"A7",
		X"41",X"33",X"44",X"11",X"83",X"51",X"AC",X"25",X"CD",X"39",X"7F",X"57",X"C7",X"0F",X"D8",X"BD",
		X"A0",X"98",X"7F",X"57",X"C9",X"8E",X"C4",X"47",X"B6",X"57",X"CD",X"88",X"01",X"B7",X"57",X"CD",
		X"27",X"03",X"8E",X"C5",X"C1",X"BF",X"57",X"CA",X"EC",X"84",X"B7",X"57",X"31",X"F7",X"57",X"CC",
		X"7E",X"8C",X"EF",X"BD",X"85",X"25",X"B6",X"57",X"C9",X"4A",X"10",X"27",X"FE",X"E1",X"F6",X"57",
		X"C7",X"C4",X"04",X"27",X"02",X"C6",X"09",X"8E",X"C4",X"35",X"3A",X"CE",X"45",X"5E",X"A6",X"80",
		X"A7",X"C4",X"33",X"C8",X"E0",X"11",X"83",X"44",X"5E",X"24",X"F3",X"39",X"86",X"0A",X"BD",X"8F",
		X"0C",X"BD",X"90",X"35",X"7E",X"8C",X"EF",X"7F",X"57",X"C6",X"39",X"B6",X"57",X"C6",X"48",X"8E",
		X"C7",X"75",X"6E",X"96",X"BD",X"91",X"EF",X"BD",X"91",X"FA",X"86",X"0A",X"BD",X"8F",X"0C",X"BD",
		X"90",X"35",X"86",X"0E",X"B7",X"45",X"06",X"86",X"0C",X"BD",X"8F",X"0C",X"CC",X"00",X"1A",X"BD",
		X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",
		X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"4F",X"5F",X"DD",X"00",X"DD",X"02",X"C6",X"54",X"BD",X"8F",
		X"0C",X"5C",X"BD",X"8F",X"0C",X"C6",X"0D",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"D6",X"AC",
		X"58",X"CB",X"10",X"4F",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"BD",X"8C",X"EF",X"8E",X"45",
		X"5E",X"CC",X"20",X"0F",X"A7",X"84",X"E7",X"89",X"08",X"00",X"30",X"88",X"E0",X"8C",X"44",X"5E",
		X"24",X"F2",X"39",X"B6",X"57",X"30",X"84",X"08",X"26",X"1A",X"96",X"82",X"4A",X"26",X"01",X"39",
		X"CC",X"00",X"0F",X"BD",X"8F",X"0C",X"7E",X"8C",X"EF",X"B6",X"57",X"30",X"84",X"18",X"27",X"EF",
		X"81",X"08",X"26",X"14",X"96",X"8C",X"4A",X"27",X"21",X"96",X"82",X"8B",X"99",X"19",X"97",X"82",
		X"86",X"05",X"BD",X"8F",X"0C",X"4F",X"20",X"12",X"96",X"8C",X"26",X"0E",X"96",X"82",X"8B",X"98",
		X"19",X"97",X"82",X"86",X"05",X"BD",X"8F",X"0C",X"86",X"01",X"97",X"B0",X"86",X"03",X"B7",X"57",
		X"C5",X"7F",X"57",X"C9",X"BD",X"91",X"EF",X"BD",X"92",X"8A",X"20",X"92",X"34",X"10",X"BE",X"52",
		X"38",X"ED",X"81",X"8C",X"57",X"80",X"25",X"03",X"8E",X"57",X"40",X"BF",X"52",X"38",X"35",X"90",
		X"86",X"0E",X"B7",X"45",X"06",X"CC",X"00",X"07",X"BD",X"8F",X"0C",X"5C",X"8E",X"41",X"B0",X"4F",
		X"BD",X"8F",X"0C",X"86",X"30",X"A7",X"84",X"A7",X"88",X"E0",X"CB",X"02",X"E7",X"89",X"08",X"00",
		X"E7",X"89",X"07",X"E0",X"C0",X"02",X"30",X"02",X"5C",X"C1",X"0C",X"23",X"E2",X"8E",X"57",X"A0",
		X"86",X"0A",X"97",X"F0",X"CE",X"42",X"70",X"8D",X"25",X"33",X"C8",X"80",X"86",X"03",X"97",X"F6",
		X"A6",X"80",X"A7",X"C4",X"96",X"F0",X"A7",X"C9",X"08",X"00",X"33",X"C8",X"E0",X"0A",X"F6",X"26",
		X"EF",X"33",X"C9",X"01",X"A2",X"0C",X"F0",X"96",X"F0",X"81",X"0E",X"23",X"DA",X"39",X"8D",X"02",
		X"8D",X"00",X"A6",X"80",X"1F",X"89",X"44",X"44",X"44",X"44",X"8D",X"02",X"1F",X"98",X"84",X"0F",
		X"26",X"10",X"A6",X"C8",X"20",X"81",X"20",X"26",X"08",X"86",X"20",X"A7",X"C4",X"33",X"C8",X"E0",
		X"39",X"4F",X"10",X"8E",X"C7",X"7B",X"A6",X"A6",X"A7",X"C4",X"96",X"F0",X"A7",X"C9",X"08",X"00",
		X"33",X"C8",X"E0",X"39",X"A6",X"84",X"E6",X"84",X"44",X"44",X"44",X"44",X"8D",X"02",X"1F",X"98",
		X"84",X"0F",X"7E",X"8F",X"A2",X"CE",X"44",X"40",X"BD",X"8F",X"DA",X"CE",X"44",X"41",X"BD",X"8F",
		X"DA",X"CE",X"44",X"5E",X"BD",X"8F",X"DA",X"CE",X"44",X"5F",X"C6",X"1C",X"86",X"20",X"A7",X"C4",
		X"86",X"0F",X"A7",X"C9",X"08",X"00",X"33",X"C8",X"20",X"5A",X"26",X"F0",X"39",X"C6",X"20",X"D7",
		X"E3",X"CE",X"40",X"00",X"86",X"20",X"34",X"40",X"C6",X"20",X"D7",X"E4",X"C6",X"0F",X"A7",X"C4",
		X"E7",X"C9",X"08",X"00",X"33",X"C8",X"20",X"0A",X"E4",X"26",X"F3",X"35",X"40",X"33",X"41",X"0A",
		X"E3",X"26",X"E3",X"86",X"20",X"C6",X"0F",X"8E",X"45",X"FE",X"A7",X"84",X"E7",X"89",X"08",X"00",
		X"A7",X"01",X"E7",X"89",X"08",X"01",X"A7",X"88",X"20",X"E7",X"89",X"08",X"20",X"A7",X"88",X"21",
		X"E7",X"89",X"08",X"21",X"39",X"CE",X"50",X"03",X"CC",X"00",X"8D",X"A7",X"C4",X"33",X"44",X"5A",
		X"26",X"F9",X"8E",X"52",X"40",X"86",X"2F",X"97",X"F6",X"4F",X"ED",X"84",X"ED",X"02",X"ED",X"04",
		X"ED",X"06",X"ED",X"08",X"ED",X"0A",X"ED",X"0C",X"ED",X"0E",X"30",X"88",X"10",X"0A",X"F6",X"26",
		X"E9",X"39",X"CE",X"51",X"A7",X"8E",X"52",X"F0",X"CC",X"08",X"00",X"E7",X"C4",X"E7",X"84",X"33",
		X"44",X"30",X"88",X"10",X"4A",X"26",X"F4",X"39",X"CE",X"51",X"EF",X"CC",X"08",X"00",X"E7",X"C4",
		X"33",X"44",X"4A",X"26",X"F9",X"39",X"CE",X"57",X"39",X"8E",X"44",X"B1",X"0D",X"AF",X"27",X"06",
		X"CE",X"57",X"3C",X"8E",X"44",X"B4",X"EC",X"C4",X"10",X"A3",X"01",X"25",X"1C",X"7C",X"57",X"D0",
		X"F6",X"57",X"D0",X"86",X"07",X"BD",X"8F",X"0C",X"BD",X"92",X"58",X"A6",X"84",X"AB",X"02",X"19",
		X"A7",X"02",X"86",X"00",X"A9",X"01",X"19",X"A7",X"01",X"39",X"8E",X"57",X"39",X"CE",X"57",X"B8",
		X"0F",X"B9",X"86",X"05",X"97",X"BA",X"96",X"AF",X"27",X"02",X"30",X"03",X"A6",X"84",X"A1",X"C4",
		X"25",X"30",X"26",X"07",X"EC",X"01",X"10",X"A3",X"41",X"25",X"27",X"0C",X"B9",X"0A",X"BA",X"27",
		X"24",X"33",X"5A",X"A6",X"84",X"A1",X"C4",X"25",X"1A",X"26",X"07",X"EC",X"01",X"10",X"A3",X"41",
		X"25",X"11",X"31",X"46",X"EC",X"C4",X"ED",X"A1",X"EC",X"42",X"ED",X"A1",X"EC",X"44",X"ED",X"A4",
		X"20",X"DB",X"39",X"33",X"46",X"A6",X"80",X"A7",X"C0",X"EC",X"84",X"ED",X"C1",X"DF",X"C6",X"CC",
		X"20",X"20",X"A7",X"C0",X"ED",X"C4",X"8E",X"C7",X"85",X"96",X"BA",X"48",X"48",X"30",X"86",X"EC",
		X"81",X"DD",X"C2",X"EC",X"84",X"DD",X"C4",X"86",X"08",X"97",X"BB",X"86",X"FF",X"97",X"BC",X"39",
		X"B6",X"57",X"D1",X"81",X"06",X"25",X"1F",X"81",X"21",X"25",X"1C",X"81",X"41",X"25",X"1F",X"81",
		X"56",X"25",X"38",X"81",X"62",X"25",X"5D",X"CC",X"00",X"01",X"DD",X"14",X"CC",X"02",X"03",X"DD",
		X"16",X"CC",X"04",X"05",X"DD",X"18",X"39",X"86",X"06",X"97",X"F6",X"7E",X"91",X"BE",X"96",X"16",
		X"26",X"0A",X"CC",X"00",X"01",X"DD",X"14",X"86",X"02",X"97",X"16",X"39",X"4C",X"81",X"06",X"25",
		X"09",X"86",X"05",X"97",X"F6",X"8D",X"47",X"4C",X"97",X"16",X"39",X"96",X"17",X"26",X"0B",X"CC",
		X"00",X"01",X"DD",X"14",X"CC",X"02",X"03",X"DD",X"16",X"39",X"4C",X"81",X"06",X"25",X"EB",X"0C",
		X"16",X"96",X"16",X"81",X"05",X"25",X"09",X"86",X"04",X"97",X"F6",X"8D",X"21",X"4C",X"97",X"16",
		X"4C",X"97",X"17",X"39",X"80",X"38",X"97",X"F6",X"48",X"48",X"9B",X"F6",X"8E",X"C7",X"99",X"30",
		X"86",X"EC",X"84",X"DD",X"14",X"EC",X"02",X"DD",X"16",X"A6",X"04",X"97",X"18",X"39",X"0C",X"15",
		X"96",X"15",X"81",X"06",X"25",X"07",X"0C",X"14",X"96",X"14",X"4C",X"97",X"15",X"39",X"F6",X"57",
		X"34",X"58",X"25",X"07",X"F6",X"57",X"C5",X"5A",X"26",X"01",X"39",X"34",X"10",X"BE",X"52",X"3C",
		X"A7",X"80",X"8C",X"57",X"A0",X"25",X"03",X"8E",X"57",X"80",X"BF",X"52",X"3C",X"35",X"90",X"4F",
		X"20",X"E9",X"86",X"01",X"20",X"DE",X"86",X"81",X"20",X"E1",X"86",X"02",X"20",X"DD",X"86",X"03",
		X"20",X"CC",X"86",X"04",X"20",X"CE",X"86",X"05",X"20",X"CA",X"86",X"06",X"20",X"C0",X"86",X"07",
		X"20",X"C2",X"86",X"08",X"20",X"B8",X"86",X"09",X"20",X"B4",X"86",X"0A",X"20",X"B0",X"86",X"0B",
		X"20",X"AC",X"86",X"0C",X"20",X"A8",X"86",X"81",X"8D",X"B1",X"86",X"0D",X"20",X"A6",X"86",X"8D",
		X"20",X"A9",X"86",X"81",X"8D",X"A5",X"86",X"0E",X"20",X"9A",X"86",X"8E",X"20",X"9D",X"86",X"0F",
		X"20",X"8C",X"86",X"10",X"20",X"88",X"86",X"11",X"8D",X"84",X"86",X"9F",X"8D",X"80",X"86",X"1A",
		X"BD",X"91",X"CE",X"86",X"19",X"7E",X"91",X"CE",X"86",X"12",X"7E",X"91",X"D4",X"86",X"13",X"BD",
		X"91",X"CE",X"86",X"14",X"7E",X"91",X"CE",X"86",X"15",X"7E",X"91",X"D4",X"86",X"16",X"7E",X"91",
		X"CE",X"86",X"17",X"7E",X"91",X"D4",X"86",X"97",X"7E",X"91",X"DB",X"86",X"18",X"7E",X"91",X"D4",
		X"86",X"1B",X"7E",X"91",X"CE",X"86",X"1C",X"7E",X"91",X"D4",X"86",X"1D",X"7E",X"91",X"D4",X"86",
		X"1F",X"7E",X"91",X"CE",X"86",X"20",X"7E",X"91",X"CE",X"8E",X"40",X"00",X"CC",X"0A",X"0A",X"ED",
		X"81",X"8C",X"44",X"00",X"25",X"F9",X"4F",X"5F",X"DD",X"0A",X"DD",X"0C",X"DD",X"0E",X"DD",X"06",
		X"DD",X"08",X"DD",X"00",X"DD",X"02",X"8E",X"C7",X"B7",X"B6",X"57",X"D6",X"A6",X"86",X"B7",X"45",
		X"06",X"DC",X"1A",X"C3",X"00",X"80",X"84",X"07",X"5F",X"DD",X"1A",X"DD",X"1E",X"DC",X"1C",X"C3",
		X"01",X"90",X"84",X"07",X"5F",X"DD",X"1C",X"DD",X"20",X"39",X"96",X"11",X"5F",X"44",X"56",X"44",
		X"56",X"44",X"56",X"DB",X"10",X"58",X"49",X"C3",X"C7",X"C5",X"1F",X"02",X"10",X"AE",X"A4",X"96",
		X"13",X"48",X"48",X"48",X"9B",X"12",X"E6",X"A6",X"8B",X"82",X"44",X"A6",X"A6",X"25",X"08",X"44",
		X"44",X"44",X"44",X"AB",X"A8",X"40",X"39",X"84",X"0F",X"AB",X"A8",X"40",X"39",X"96",X"01",X"97",
		X"00",X"96",X"03",X"97",X"02",X"B6",X"57",X"C9",X"81",X"0F",X"26",X"47",X"B6",X"57",X"CE",X"80",
		X"F0",X"25",X"1F",X"27",X"17",X"81",X"01",X"22",X"12",X"CC",X"20",X"0F",X"8E",X"40",X"00",X"CE",
		X"48",X"00",X"A7",X"80",X"E7",X"C0",X"8C",X"44",X"00",X"25",X"F7",X"39",X"5F",X"DD",X"02",X"DD",
		X"00",X"39",X"FC",X"45",X"02",X"DD",X"3A",X"FC",X"45",X"04",X"DD",X"3C",X"4F",X"F6",X"57",X"CE",
		X"58",X"49",X"58",X"49",X"58",X"49",X"BD",X"A6",X"6F",X"DC",X"3A",X"FD",X"57",X"C0",X"DC",X"3C",
		X"FD",X"57",X"C2",X"DC",X"06",X"34",X"02",X"F3",X"57",X"C0",X"DD",X"06",X"35",X"02",X"0F",X"F6",
		X"F6",X"57",X"DD",X"27",X"16",X"F6",X"54",X"6D",X"26",X"11",X"F6",X"54",X"60",X"5A",X"2B",X"0B",
		X"54",X"C4",X"03",X"5C",X"D7",X"F6",X"8E",X"C7",X"BC",X"AB",X"85",X"90",X"06",X"27",X"3E",X"1F",
		X"89",X"40",X"9B",X"03",X"97",X"03",X"1D",X"2A",X"18",X"D3",X"1A",X"84",X"07",X"DD",X"1A",X"CB",
		X"07",X"D1",X"1F",X"2A",X"28",X"DC",X"1E",X"83",X"00",X"08",X"84",X"07",X"DD",X"1E",X"5F",X"20",
		X"17",X"D3",X"1A",X"84",X"07",X"DD",X"1A",X"C0",X"08",X"D1",X"1F",X"2B",X"10",X"DC",X"1E",X"C3",
		X"00",X"08",X"84",X"07",X"DD",X"1E",X"C6",X"01",X"86",X"08",X"BD",X"8F",X"0C",X"DC",X"08",X"34",
		X"02",X"F3",X"57",X"C2",X"DD",X"08",X"35",X"02",X"D6",X"F6",X"27",X"04",X"CB",X"04",X"AB",X"85",
		X"90",X"08",X"27",X"3E",X"1F",X"89",X"9B",X"01",X"97",X"01",X"1D",X"2A",X"19",X"D3",X"1C",X"84",
		X"07",X"DD",X"1C",X"CB",X"07",X"D1",X"21",X"2A",X"29",X"DC",X"20",X"83",X"00",X"08",X"84",X"07",
		X"DD",X"20",X"C6",X"02",X"20",X"17",X"D3",X"1C",X"84",X"07",X"DD",X"1C",X"C0",X"08",X"D1",X"21",
		X"2B",X"10",X"DC",X"20",X"C3",X"00",X"08",X"84",X"07",X"DD",X"20",X"C6",X"03",X"86",X"08",X"7E",
		X"8F",X"0C",X"39",X"D7",X"22",X"96",X"22",X"4A",X"27",X"02",X"86",X"F8",X"90",X"1F",X"44",X"44",
		X"44",X"C1",X"03",X"D6",X"21",X"25",X"02",X"C0",X"08",X"44",X"56",X"44",X"56",X"44",X"56",X"C3",
		X"40",X"00",X"DD",X"04",X"D6",X"1F",X"96",X"22",X"81",X"01",X"26",X"02",X"CB",X"F8",X"54",X"54",
		X"54",X"C4",X"07",X"D7",X"12",X"96",X"22",X"40",X"81",X"FF",X"DC",X"1E",X"25",X"03",X"C3",X"00",
		X"F8",X"58",X"49",X"58",X"49",X"84",X"1F",X"97",X"10",X"D6",X"21",X"96",X"22",X"81",X"03",X"25",
		X"02",X"CB",X"F8",X"54",X"54",X"54",X"C4",X"07",X"D7",X"13",X"96",X"22",X"81",X"03",X"DC",X"20",
		X"25",X"03",X"C3",X"00",X"F8",X"58",X"49",X"58",X"49",X"84",X"1F",X"97",X"11",X"86",X"20",X"97",
		X"2F",X"96",X"22",X"84",X"02",X"26",X"2D",X"BD",X"92",X"DA",X"9E",X"04",X"E7",X"84",X"A7",X"89",
		X"08",X"00",X"0A",X"2F",X"27",X"4B",X"1F",X"10",X"5C",X"C5",X"1F",X"26",X"02",X"C0",X"20",X"DD",
		X"04",X"0C",X"13",X"96",X"13",X"84",X"07",X"26",X"DE",X"97",X"13",X"96",X"11",X"4C",X"84",X"1F",
		X"97",X"11",X"20",X"D3",X"BD",X"92",X"DA",X"9E",X"04",X"E7",X"84",X"A7",X"89",X"08",X"00",X"0A",
		X"2F",X"27",X"1E",X"1F",X"10",X"83",X"40",X"20",X"84",X"03",X"8B",X"40",X"DD",X"04",X"0C",X"12",
		X"96",X"12",X"84",X"07",X"26",X"DE",X"97",X"12",X"96",X"10",X"4C",X"84",X"1F",X"97",X"10",X"20",
		X"D3",X"39",X"FC",X"52",X"35",X"C3",X"00",X"01",X"FD",X"52",X"35",X"10",X"83",X"FF",X"FF",X"26",
		X"2E",X"B6",X"52",X"36",X"8E",X"BD",X"5E",X"C6",X"06",X"A6",X"80",X"AB",X"80",X"5A",X"26",X"FB",
		X"81",X"1B",X"27",X"0C",X"CC",X"00",X"52",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"20",X"0F",
		X"B6",X"A8",X"FC",X"81",X"34",X"27",X"08",X"B6",X"57",X"C8",X"88",X"01",X"B7",X"57",X"C8",X"B6",
		X"57",X"DD",X"10",X"26",X"00",X"83",X"B6",X"57",X"D1",X"81",X"06",X"25",X"07",X"CC",X"40",X"3D",
		X"DD",X"F6",X"20",X"05",X"CC",X"30",X"2D",X"DD",X"F6",X"B6",X"57",X"DB",X"91",X"F6",X"24",X"55",
		X"91",X"F7",X"25",X"04",X"86",X"FF",X"97",X"F5",X"B6",X"57",X"DC",X"B1",X"57",X"DF",X"24",X"45",
		X"8B",X"03",X"B1",X"57",X"DF",X"25",X"04",X"86",X"FF",X"97",X"F5",X"DC",X"E9",X"C3",X"00",X"01",
		X"DD",X"E9",X"10",X"83",X"02",X"80",X"26",X"32",X"96",X"EB",X"44",X"91",X"EC",X"25",X"0E",X"96",
		X"EC",X"81",X"03",X"24",X"08",X"0F",X"EB",X"0F",X"EC",X"0F",X"E9",X"0F",X"EA",X"7C",X"57",X"DF",
		X"B6",X"57",X"DF",X"81",X"21",X"25",X"05",X"86",X"20",X"B7",X"57",X"DF",X"CC",X"00",X"00",X"DD",
		X"E9",X"DD",X"EB",X"20",X"05",X"86",X"FF",X"B7",X"57",X"DD",X"96",X"F5",X"27",X"1C",X"B6",X"4C",
		X"00",X"26",X"06",X"7A",X"4C",X"00",X"BD",X"92",X"80",X"8E",X"45",X"FE",X"B6",X"57",X"C7",X"44",
		X"44",X"84",X"03",X"8B",X"01",X"C6",X"8F",X"BD",X"84",X"C6",X"0D",X"9C",X"27",X"02",X"0A",X"9C",
		X"B6",X"57",X"C7",X"84",X"1F",X"26",X"06",X"0A",X"B8",X"10",X"27",X"00",X"1B",X"0D",X"A7",X"27",
		X"0C",X"0A",X"A4",X"26",X"12",X"0F",X"A7",X"96",X"A5",X"97",X"A6",X"20",X"0A",X"0A",X"A6",X"26",
		X"06",X"0C",X"A7",X"96",X"A3",X"97",X"A4",X"39",X"96",X"B7",X"97",X"B8",X"F6",X"57",X"D3",X"7C",
		X"57",X"D3",X"C1",X"17",X"25",X"06",X"C6",X"17",X"F7",X"57",X"D3",X"39",X"4F",X"DD",X"F6",X"58",
		X"46",X"58",X"46",X"58",X"46",X"D3",X"F6",X"C3",X"F3",X"C4",X"1F",X"03",X"A6",X"C4",X"97",X"98",
		X"A6",X"41",X"97",X"9B",X"A6",X"42",X"97",X"A3",X"A6",X"43",X"97",X"A5",X"97",X"A6",X"A6",X"44",
		X"97",X"96",X"A6",X"45",X"97",X"9A",X"A6",X"46",X"97",X"97",X"A6",X"47",X"97",X"9D",X"A6",X"48",
		X"97",X"A2",X"0F",X"A7",X"39",X"B6",X"57",X"D2",X"81",X"02",X"27",X"04",X"81",X"05",X"26",X"08",
		X"9E",X"2C",X"27",X"04",X"30",X"1F",X"9F",X"2C",X"8E",X"54",X"60",X"CE",X"52",X"00",X"A6",X"84",
		X"27",X"1A",X"4C",X"10",X"27",X"00",X"DB",X"10",X"2A",X"01",X"F7",X"F6",X"52",X"40",X"5C",X"FA",
		X"57",X"C4",X"EA",X"0D",X"10",X"26",X"02",X"9F",X"A7",X"84",X"20",X"51",X"B6",X"52",X"40",X"4C",
		X"BA",X"52",X"34",X"BA",X"57",X"C4",X"26",X"0A",X"B6",X"57",X"DD",X"27",X"06",X"BD",X"92",X"26",
		X"20",X"1F",X"39",X"DC",X"2C",X"26",X"FB",X"4A",X"F6",X"57",X"D2",X"C1",X"02",X"27",X"05",X"40",
		X"C1",X"05",X"26",X"EE",X"A7",X"0D",X"BD",X"92",X"32",X"A6",X"0D",X"2B",X"04",X"C6",X"68",X"20",
		X"02",X"C6",X"30",X"6A",X"84",X"E7",X"0A",X"E7",X"0B",X"10",X"8E",X"53",X"A0",X"86",X"FE",X"A7",
		X"A4",X"31",X"30",X"10",X"8C",X"53",X"50",X"24",X"F6",X"A6",X"0D",X"26",X"67",X"86",X"FD",X"F6",
		X"52",X"41",X"E7",X"01",X"CB",X"A0",X"D7",X"F6",X"C4",X"3F",X"58",X"CB",X"40",X"08",X"F6",X"25",
		X"09",X"08",X"F6",X"24",X"0E",X"1E",X"89",X"40",X"20",X"09",X"40",X"50",X"08",X"F6",X"24",X"03",
		X"1E",X"89",X"40",X"80",X"08",X"A7",X"43",X"A7",X"4B",X"8B",X"10",X"A7",X"47",X"A7",X"4F",X"E7",
		X"48",X"E7",X"4C",X"C0",X"10",X"E7",X"C4",X"E7",X"44",X"6F",X"02",X"6F",X"03",X"6F",X"08",X"6F",
		X"09",X"C6",X"40",X"A6",X"0D",X"27",X"0D",X"B6",X"57",X"D2",X"81",X"05",X"86",X"F5",X"25",X"06",
		X"86",X"F9",X"20",X"02",X"86",X"A1",X"ED",X"41",X"4C",X"ED",X"45",X"4C",X"ED",X"49",X"4C",X"ED",
		X"4D",X"7E",X"99",X"17",X"4F",X"5F",X"ED",X"04",X"CC",X"FE",X"E8",X"ED",X"06",X"CC",X"80",X"FD",
		X"20",X"B1",X"A6",X"0D",X"26",X"63",X"FC",X"57",X"C2",X"58",X"49",X"58",X"49",X"58",X"49",X"58",
		X"49",X"DD",X"F7",X"58",X"49",X"D3",X"F7",X"8B",X"78",X"97",X"F6",X"FC",X"57",X"C0",X"58",X"49",
		X"58",X"49",X"58",X"49",X"58",X"49",X"DD",X"F7",X"58",X"49",X"D3",X"F7",X"8B",X"80",X"E6",X"43",
		X"CB",X"08",X"E7",X"43",X"E6",X"C4",X"CB",X"08",X"E7",X"C4",X"D6",X"F6",X"BD",X"A5",X"E0",X"A6",
		X"43",X"80",X"08",X"A7",X"43",X"A6",X"C4",X"80",X"08",X"A7",X"C4",X"1F",X"98",X"C6",X"01",X"A0",
		X"01",X"2A",X"01",X"50",X"EB",X"01",X"E7",X"01",X"BD",X"A6",X"21",X"CC",X"01",X"60",X"BD",X"A6",
		X"6F",X"DC",X"3A",X"ED",X"04",X"DC",X"3C",X"ED",X"06",X"A6",X"43",X"E6",X"02",X"E3",X"04",X"F3",
		X"57",X"C0",X"A7",X"43",X"E7",X"02",X"A7",X"4B",X"8B",X"10",X"A7",X"47",X"A7",X"4F",X"8B",X"F9",
		X"81",X"02",X"23",X"6B",X"A6",X"C4",X"E6",X"03",X"E3",X"06",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",
		X"03",X"A7",X"44",X"8B",X"10",X"A7",X"48",X"A7",X"4C",X"8B",X"02",X"81",X"02",X"23",X"50",X"A6",
		X"84",X"10",X"2A",X"01",X"32",X"A6",X"0D",X"10",X"26",X"01",X"2C",X"EC",X"08",X"4C",X"81",X"03",
		X"26",X"38",X"5C",X"C1",X"03",X"26",X"01",X"5F",X"E7",X"09",X"58",X"58",X"CB",X"A1",X"E7",X"41",
		X"5C",X"E7",X"45",X"5C",X"E7",X"49",X"5C",X"E7",X"4D",X"B6",X"28",X"20",X"84",X"0F",X"26",X"19",
		X"34",X"50",X"8E",X"F4",X"9C",X"CE",X"46",X"A0",X"A6",X"80",X"88",X"56",X"A7",X"C4",X"33",X"C8",
		X"E0",X"11",X"83",X"44",X"E0",X"22",X"F1",X"35",X"50",X"4F",X"A7",X"08",X"7E",X"99",X"17",X"6F",
		X"43",X"6F",X"47",X"6F",X"4B",X"6F",X"4F",X"A6",X"0D",X"27",X"0D",X"86",X"FE",X"A7",X"84",X"BD",
		X"92",X"3A",X"BD",X"91",X"F2",X"7E",X"99",X"17",X"A6",X"84",X"2A",X"07",X"86",X"FE",X"A7",X"84",
		X"7E",X"99",X"17",X"86",X"C0",X"B7",X"57",X"CE",X"86",X"FF",X"B7",X"57",X"C4",X"6F",X"84",X"7E",
		X"99",X"17",X"81",X"78",X"10",X"23",X"00",X"8B",X"86",X"06",X"A7",X"84",X"4F",X"5F",X"ED",X"04",
		X"ED",X"06",X"A6",X"0D",X"26",X"54",X"86",X"0D",X"A7",X"0E",X"C6",X"78",X"8E",X"53",X"A0",X"86",
		X"0C",X"97",X"F6",X"8D",X"37",X"8E",X"54",X"30",X"86",X"09",X"97",X"F6",X"8D",X"2E",X"8E",X"55",
		X"10",X"86",X"08",X"97",X"F6",X"8D",X"25",X"CC",X"E9",X"40",X"ED",X"41",X"4C",X"ED",X"45",X"4C",
		X"ED",X"49",X"4C",X"ED",X"4D",X"C6",X"03",X"BD",X"A5",X"AB",X"CC",X"06",X"08",X"BD",X"8F",X"0C",
		X"BD",X"92",X"2E",X"BD",X"92",X"4A",X"8E",X"54",X"60",X"7E",X"97",X"A9",X"A6",X"84",X"4C",X"26",
		X"02",X"E7",X"84",X"30",X"10",X"0A",X"F6",X"26",X"F3",X"39",X"4C",X"48",X"8B",X"ED",X"A7",X"41",
		X"4C",X"A7",X"45",X"4C",X"A7",X"49",X"4C",X"A7",X"4D",X"86",X"0C",X"A7",X"0E",X"5F",X"BD",X"A5",
		X"AB",X"CC",X"06",X"05",X"BD",X"8F",X"0C",X"BD",X"92",X"3A",X"BD",X"92",X"46",X"BD",X"91",X"F2",
		X"7E",X"97",X"A9",X"6A",X"84",X"10",X"26",X"FE",X"B0",X"6A",X"0E",X"10",X"2B",X"FF",X"30",X"86",
		X"06",X"A7",X"84",X"E6",X"0E",X"58",X"58",X"CB",X"B5",X"E7",X"41",X"5C",X"E7",X"45",X"5C",X"E7",
		X"49",X"5C",X"E7",X"4D",X"7E",X"97",X"A9",X"10",X"8E",X"F4",X"AA",X"A6",X"84",X"4C",X"26",X"75",
		X"6A",X"0B",X"26",X"71",X"B6",X"57",X"D3",X"48",X"40",X"8B",X"18",X"AB",X"0A",X"A7",X"0B",X"8E",
		X"53",X"A0",X"CE",X"51",X"D0",X"A6",X"84",X"81",X"FE",X"26",X"51",X"B6",X"52",X"03",X"8B",X"08",
		X"A7",X"43",X"B6",X"52",X"00",X"8B",X"08",X"A7",X"C4",X"F6",X"54",X"6C",X"CB",X"2B",X"F7",X"54",
		X"6C",X"E7",X"01",X"6F",X"08",X"B6",X"54",X"6D",X"2A",X"1D",X"BD",X"A6",X"21",X"B6",X"57",X"D3",
		X"C6",X"0C",X"3D",X"C3",X"00",X"10",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"04",X"DC",X"3C",X"ED",
		X"06",X"6F",X"09",X"C6",X"20",X"20",X"07",X"CB",X"08",X"C4",X"F0",X"54",X"54",X"54",X"EC",X"A5",
		X"ED",X"41",X"6C",X"84",X"BD",X"92",X"22",X"B6",X"54",X"6D",X"27",X"09",X"30",X"10",X"33",X"5C",
		X"8C",X"53",X"50",X"24",X"A0",X"8E",X"53",X"A0",X"CE",X"51",X"D0",X"A6",X"84",X"10",X"27",X"00",
		X"88",X"4C",X"10",X"2B",X"00",X"83",X"10",X"26",X"00",X"CD",X"B6",X"54",X"6D",X"2A",X"15",X"6C",
		X"09",X"A6",X"09",X"85",X"07",X"26",X"45",X"44",X"44",X"44",X"84",X"07",X"8B",X"22",X"A6",X"A6",
		X"A7",X"42",X"20",X"38",X"CC",X"80",X"78",X"BD",X"A5",X"E0",X"1F",X"98",X"C6",X"01",X"A0",X"01",
		X"2A",X"01",X"50",X"EB",X"01",X"E7",X"01",X"BD",X"A6",X"21",X"F6",X"57",X"D3",X"58",X"58",X"58",
		X"4F",X"C3",X"01",X"40",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"04",X"DC",X"3C",X"ED",X"06",X"A6",
		X"01",X"8B",X"08",X"84",X"F0",X"44",X"44",X"44",X"EC",X"A6",X"ED",X"41",X"6A",X"08",X"26",X"04",
		X"86",X"78",X"A7",X"84",X"A6",X"43",X"E6",X"02",X"E3",X"04",X"F3",X"57",X"C0",X"A7",X"43",X"E7",
		X"02",X"8B",X"08",X"81",X"10",X"23",X"58",X"A6",X"C4",X"E6",X"03",X"E3",X"06",X"F3",X"57",X"C2",
		X"A7",X"C4",X"E7",X"03",X"40",X"81",X"10",X"23",X"46",X"30",X"10",X"33",X"5C",X"8C",X"53",X"50",
		X"10",X"24",X"FF",X"67",X"B6",X"54",X"6D",X"27",X"35",X"B6",X"54",X"60",X"81",X"FE",X"26",X"2E",
		X"A6",X"47",X"AA",X"4B",X"AA",X"4F",X"AA",X"C8",X"13",X"AA",X"C8",X"17",X"AA",X"C8",X"1B",X"26",
		X"1D",X"4F",X"B7",X"54",X"60",X"B7",X"54",X"6D",X"A7",X"88",X"10",X"A7",X"88",X"20",X"A7",X"88",
		X"30",X"A7",X"88",X"40",X"A7",X"88",X"50",X"A7",X"88",X"60",X"86",X"02",X"97",X"2C",X"39",X"6F",
		X"43",X"86",X"FE",X"A7",X"84",X"20",X"B2",X"81",X"78",X"23",X"0D",X"4F",X"5F",X"ED",X"04",X"ED",
		X"06",X"BD",X"92",X"0E",X"86",X"11",X"A7",X"84",X"6A",X"84",X"27",X"E3",X"A6",X"84",X"85",X"03",
		X"26",X"97",X"44",X"44",X"8B",X"29",X"A6",X"A6",X"E6",X"42",X"C4",X"C0",X"ED",X"41",X"7E",X"9A",
		X"04",X"DC",X"D8",X"C3",X"00",X"01",X"DD",X"D8",X"B6",X"57",X"DD",X"26",X"68",X"B6",X"57",X"C7",
		X"2B",X"64",X"B6",X"54",X"60",X"26",X"5E",X"B6",X"57",X"CE",X"27",X"05",X"7A",X"57",X"CE",X"26",
		X"25",X"B6",X"57",X"D2",X"81",X"02",X"27",X"1E",X"81",X"05",X"27",X"1A",X"10",X"8E",X"F4",X"D8",
		X"48",X"A6",X"B6",X"26",X"11",X"B6",X"52",X"34",X"81",X"02",X"24",X"3A",X"10",X"8E",X"F4",X"E2",
		X"B6",X"57",X"D2",X"48",X"AD",X"B6",X"B6",X"57",X"C5",X"4A",X"26",X"05",X"B6",X"57",X"D6",X"27",
		X"25",X"DC",X"2C",X"27",X"21",X"86",X"10",X"F6",X"57",X"DE",X"3D",X"DD",X"F6",X"CC",X"02",X"80",
		X"93",X"F6",X"10",X"93",X"D8",X"24",X"0F",X"B6",X"52",X"34",X"81",X"02",X"24",X"08",X"96",X"DA",
		X"26",X"04",X"7E",X"9E",X"2C",X"39",X"96",X"99",X"27",X"04",X"0A",X"99",X"26",X"F7",X"96",X"98",
		X"97",X"99",X"96",X"97",X"97",X"D4",X"B6",X"57",X"C7",X"2A",X"06",X"96",X"E5",X"81",X"03",X"24",
		X"1C",X"8E",X"52",X"F0",X"CE",X"51",X"A4",X"A6",X"84",X"26",X"07",X"BD",X"9D",X"69",X"0A",X"D4",
		X"27",X"D3",X"30",X"88",X"10",X"33",X"44",X"8C",X"53",X"50",X"25",X"EB",X"39",X"0F",X"E5",X"B6",
		X"57",X"C5",X"4A",X"26",X"05",X"B6",X"57",X"D6",X"26",X"BB",X"96",X"DA",X"26",X"B7",X"DC",X"2C",
		X"27",X"B3",X"B6",X"52",X"34",X"81",X"06",X"24",X"AC",X"8E",X"53",X"50",X"CE",X"51",X"BC",X"A6",
		X"84",X"26",X"34",X"7C",X"52",X"34",X"B6",X"57",X"D1",X"81",X"06",X"25",X"1D",X"96",X"E7",X"26",
		X"04",X"96",X"14",X"20",X"15",X"96",X"E7",X"81",X"06",X"25",X"03",X"4F",X"97",X"E7",X"10",X"8E",
		X"44",X"14",X"A6",X"A6",X"26",X"04",X"0F",X"E7",X"96",X"14",X"0C",X"E7",X"48",X"10",X"8E",X"F4",
		X"EC",X"AD",X"B6",X"0A",X"D4",X"27",X"0A",X"30",X"88",X"10",X"33",X"44",X"8C",X"53",X"B0",X"25",
		X"BE",X"39",X"BD",X"A0",X"9E",X"84",X"1F",X"9B",X"D4",X"85",X"01",X"27",X"01",X"40",X"BB",X"52",
		X"41",X"97",X"D2",X"BD",X"9D",X"C7",X"CC",X"FF",X"00",X"A7",X"84",X"E7",X"03",X"BD",X"A0",X"9E",
		X"84",X"0F",X"85",X"01",X"27",X"01",X"40",X"A7",X"01",X"BD",X"A5",X"DE",X"EB",X"01",X"E7",X"01",
		X"BD",X"A6",X"21",X"CC",X"01",X"10",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"06",X"DC",X"3C",X"ED",
		X"08",X"86",X"40",X"A7",X"42",X"CC",X"00",X"00",X"A7",X"04",X"ED",X"0C",X"39",X"CC",X"FF",X"01",
		X"A7",X"84",X"E7",X"03",X"6F",X"04",X"BD",X"A0",X"9E",X"84",X"1F",X"BB",X"57",X"C7",X"A7",X"05",
		X"BD",X"A0",X"9E",X"84",X"F8",X"8B",X"80",X"A7",X"43",X"F6",X"52",X"41",X"CB",X"04",X"2A",X"1B",
		X"86",X"EF",X"A7",X"C4",X"86",X"C0",X"A7",X"01",X"86",X"40",X"A7",X"41",X"86",X"40",X"A7",X"42",
		X"CC",X"FE",X"A0",X"ED",X"06",X"86",X"C0",X"A7",X"02",X"20",X"15",X"CC",X"01",X"40",X"A7",X"C4",
		X"E7",X"01",X"CC",X"40",X"00",X"ED",X"41",X"CC",X"01",X"60",X"ED",X"06",X"86",X"40",X"A7",X"02",
		X"CC",X"00",X"00",X"ED",X"08",X"ED",X"0C",X"39",X"6A",X"84",X"CC",X"02",X"00",X"ED",X"03",X"BD",
		X"A0",X"9E",X"84",X"3F",X"8B",X"40",X"A7",X"05",X"CC",X"40",X"30",X"A7",X"42",X"E7",X"0B",X"BD",
		X"A0",X"9E",X"BB",X"57",X"C7",X"A7",X"43",X"CC",X"00",X"00",X"ED",X"06",X"ED",X"0C",X"B6",X"52",
		X"41",X"2A",X"0D",X"CC",X"FE",X"80",X"ED",X"08",X"CC",X"C0",X"EF",X"A7",X"01",X"E7",X"C4",X"39",
		X"CC",X"01",X"80",X"ED",X"08",X"CC",X"40",X"01",X"A7",X"01",X"E7",X"C4",X"39",X"6A",X"84",X"CC",
		X"00",X"00",X"ED",X"04",X"ED",X"06",X"ED",X"08",X"CC",X"24",X"40",X"ED",X"41",X"CC",X"00",X"03",
		X"A7",X"01",X"E7",X"03",X"BD",X"A0",X"9E",X"84",X"1F",X"BB",X"57",X"C7",X"A7",X"02",X"BD",X"A0",
		X"9E",X"A7",X"43",X"B6",X"52",X"41",X"2B",X"0A",X"86",X"01",X"A7",X"C4",X"CC",X"01",X"48",X"ED",
		X"0A",X"39",X"86",X"EF",X"A7",X"C4",X"CC",X"FE",X"B8",X"ED",X"0A",X"39",X"BD",X"A0",X"9E",X"84",
		X"1F",X"9B",X"D4",X"85",X"01",X"27",X"01",X"40",X"BB",X"52",X"41",X"97",X"D2",X"BD",X"9D",X"C7",
		X"CC",X"FF",X"04",X"A7",X"84",X"E7",X"03",X"CC",X"40",X"20",X"A7",X"42",X"E7",X"41",X"BD",X"A0",
		X"9E",X"1F",X"89",X"C4",X"0F",X"85",X"01",X"27",X"01",X"50",X"FB",X"52",X"41",X"C0",X"80",X"E7",
		X"01",X"BD",X"A6",X"21",X"CC",X"01",X"50",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"06",X"DC",X"3C",
		X"ED",X"08",X"86",X"20",X"A7",X"04",X"A7",X"05",X"CC",X"00",X"00",X"ED",X"0C",X"39",X"B6",X"57",
		X"3F",X"7C",X"57",X"3F",X"F6",X"57",X"3F",X"C1",X"0B",X"25",X"03",X"7F",X"57",X"3F",X"10",X"8E",
		X"F4",X"F8",X"48",X"EC",X"A6",X"A7",X"43",X"E7",X"C4",X"86",X"40",X"A7",X"42",X"CC",X"FF",X"05",
		X"A7",X"84",X"E7",X"03",X"BD",X"A5",X"DE",X"BD",X"A6",X"21",X"CC",X"01",X"80",X"BD",X"A6",X"6F",
		X"DC",X"3A",X"ED",X"06",X"DC",X"3C",X"ED",X"08",X"39",X"0C",X"E5",X"BD",X"A0",X"9E",X"84",X"1F",
		X"9B",X"D4",X"85",X"01",X"27",X"01",X"40",X"BB",X"52",X"41",X"97",X"D2",X"8D",X"49",X"CC",X"FF",
		X"06",X"A7",X"84",X"E7",X"03",X"BD",X"A0",X"9E",X"84",X"0F",X"85",X"01",X"27",X"01",X"40",X"BB",
		X"52",X"41",X"80",X"80",X"A7",X"01",X"E6",X"01",X"BD",X"A6",X"21",X"CC",X"00",X"C4",X"BD",X"A6",
		X"6F",X"DC",X"3A",X"ED",X"06",X"DC",X"3C",X"ED",X"08",X"96",X"96",X"A7",X"0A",X"BD",X"A0",X"9E",
		X"84",X"3F",X"85",X"20",X"27",X"01",X"40",X"9B",X"9A",X"A7",X"0B",X"86",X"11",X"A7",X"04",X"CC",
		X"00",X"00",X"A7",X"05",X"ED",X"0C",X"39",X"34",X"20",X"8B",X"20",X"84",X"C0",X"48",X"49",X"49",
		X"48",X"10",X"8E",X"F5",X"90",X"EC",X"A6",X"4C",X"26",X"29",X"59",X"25",X"13",X"96",X"D2",X"80",
		X"A0",X"48",X"48",X"4D",X"26",X"02",X"86",X"04",X"A7",X"43",X"86",X"01",X"A7",X"C4",X"35",X"A0",
		X"86",X"60",X"90",X"D2",X"48",X"48",X"4D",X"26",X"02",X"86",X"FC",X"A7",X"43",X"86",X"EF",X"A7",
		X"C4",X"35",X"A0",X"49",X"25",X"13",X"C6",X"A0",X"D0",X"D2",X"58",X"58",X"5D",X"26",X"02",X"C6",
		X"EF",X"E7",X"C4",X"86",X"04",X"A7",X"43",X"35",X"A0",X"D6",X"D2",X"C0",X"E0",X"58",X"58",X"5D",
		X"26",X"02",X"C6",X"01",X"E7",X"C4",X"86",X"FC",X"A7",X"43",X"35",X"A0",X"B6",X"57",X"DE",X"81",
		X"28",X"25",X"01",X"39",X"BD",X"92",X"42",X"CC",X"00",X"00",X"DD",X"D8",X"97",X"D5",X"F6",X"52",
		X"41",X"C0",X"80",X"BD",X"A6",X"21",X"CC",X"01",X"04",X"BD",X"A6",X"6F",X"8E",X"53",X"50",X"CE",
		X"51",X"BC",X"B6",X"57",X"C7",X"84",X"03",X"85",X"01",X"27",X"01",X"40",X"BB",X"52",X"41",X"97",
		X"D3",X"BD",X"A0",X"9E",X"84",X"03",X"48",X"10",X"8E",X"F5",X"0C",X"10",X"AE",X"A6",X"A6",X"A0",
		X"97",X"3E",X"A6",X"84",X"26",X"2D",X"0C",X"D5",X"7C",X"52",X"34",X"EC",X"A1",X"E7",X"0E",X"9B",
		X"D3",X"97",X"D2",X"BD",X"9D",X"C7",X"CC",X"FE",X"07",X"A7",X"84",X"E7",X"03",X"CC",X"FF",X"40",
		X"ED",X"41",X"DC",X"3A",X"ED",X"06",X"DC",X"3C",X"ED",X"08",X"CC",X"00",X"00",X"ED",X"0C",X"0A",
		X"3E",X"27",X"0A",X"30",X"88",X"10",X"33",X"44",X"8C",X"53",X"B0",X"25",X"C5",X"39",X"39",X"DC",
		X"1A",X"10",X"83",X"01",X"70",X"25",X"F7",X"10",X"83",X"02",X"61",X"24",X"F1",X"B6",X"52",X"41",
		X"80",X"20",X"84",X"40",X"26",X"E8",X"7C",X"57",X"D9",X"20",X"1A",X"DC",X"1C",X"10",X"83",X"04",
		X"70",X"25",X"DB",X"10",X"83",X"05",X"61",X"24",X"D5",X"B6",X"52",X"41",X"8B",X"20",X"84",X"40",
		X"26",X"CC",X"7C",X"57",X"DA",X"0F",X"E8",X"8E",X"53",X"50",X"CE",X"51",X"BC",X"86",X"05",X"97",
		X"F6",X"B6",X"52",X"41",X"8B",X"20",X"84",X"C0",X"27",X"08",X"48",X"24",X"1A",X"48",X"24",X"2C",
		X"20",X"3F",X"10",X"8E",X"F5",X"40",X"CC",X"AE",X"40",X"DD",X"F8",X"CC",X"04",X"96",X"DD",X"FA",
		X"CC",X"00",X"0A",X"DD",X"FC",X"20",X"3D",X"10",X"8E",X"F5",X"54",X"CC",X"AD",X"00",X"DD",X"F8",
		X"CC",X"9E",X"01",X"DD",X"FA",X"CC",X"0A",X"00",X"DD",X"FC",X"20",X"28",X"10",X"8E",X"F5",X"68",
		X"CC",X"AE",X"C0",X"DD",X"F8",X"CC",X"FC",X"96",X"DD",X"FA",X"CC",X"00",X"0A",X"DD",X"FC",X"20",
		X"13",X"10",X"8E",X"F5",X"7C",X"CC",X"AD",X"40",X"DD",X"F8",X"CC",X"9E",X"EF",X"DD",X"FA",X"CC",
		X"0A",X"00",X"DD",X"FC",X"A6",X"84",X"26",X"2F",X"7C",X"52",X"34",X"0C",X"E8",X"EC",X"A1",X"ED",
		X"06",X"EC",X"A1",X"ED",X"08",X"DC",X"F8",X"ED",X"41",X"DC",X"FA",X"93",X"FC",X"DD",X"FA",X"A7",
		X"43",X"E7",X"C4",X"CC",X"00",X"00",X"ED",X"0C",X"86",X"54",X"A7",X"01",X"CC",X"FF",X"08",X"A7",
		X"84",X"E7",X"03",X"0A",X"F6",X"27",X"0A",X"30",X"88",X"10",X"33",X"44",X"8C",X"53",X"B0",X"25",
		X"C3",X"39",X"96",X"AF",X"26",X"05",X"96",X"36",X"27",X"05",X"39",X"96",X"37",X"26",X"FB",X"DC",
		X"1A",X"10",X"83",X"03",X"80",X"25",X"F3",X"10",X"83",X"04",X"81",X"24",X"ED",X"DC",X"1C",X"10",
		X"83",X"02",X"80",X"25",X"E5",X"10",X"83",X"03",X"81",X"24",X"DF",X"96",X"AF",X"26",X"04",X"0C",
		X"36",X"20",X"02",X"0C",X"37",X"8E",X"53",X"50",X"CE",X"51",X"BC",X"A6",X"84",X"26",X"3A",X"6A",
		X"84",X"7C",X"52",X"34",X"86",X"09",X"A7",X"03",X"B6",X"52",X"41",X"2B",X"16",X"CC",X"80",X"EF",
		X"A7",X"43",X"E7",X"C4",X"CC",X"00",X"00",X"ED",X"06",X"CC",X"FF",X"18",X"ED",X"08",X"86",X"40",
		X"A7",X"42",X"39",X"CC",X"80",X"01",X"A7",X"43",X"E7",X"C4",X"CC",X"00",X"00",X"ED",X"06",X"CC");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
