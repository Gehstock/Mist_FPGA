library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"5E",X"23",X"56",X"D5",X"C9",X"15",X"08",X"2F",X"08",X"45",X"08",X"62",X"08",X"62",X"08",X"62",
		X"08",X"62",X"08",X"62",X"08",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"CB",X"21",X"06",X"00",
		X"21",X"B3",X"08",X"09",X"5E",X"23",X"56",X"DD",X"73",X"04",X"DD",X"72",X"05",X"18",X"23",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"4E",X"06",X"00",X"21",X"4B",X"09",X"09",X"7E",X"32",X"A2",X"42",
		X"DD",X"77",X"01",X"18",X"0D",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"06",X"DD",
		X"77",X"07",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",
		X"D9",X"07",X"06",X"00",X"DF",X"DD",X"36",X"00",X"FF",X"C9",X"CD",X"72",X"08",X"06",X"00",X"DF",
		X"18",X"33",X"78",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"01",X"10",X"04",X"DD",X"77",X"00",
		X"C9",X"07",X"18",X"F7",X"C5",X"CD",X"72",X"08",X"C1",X"78",X"E6",X"1F",X"3D",X"07",X"4F",X"06",
		X"00",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",X"EF",X"DD",X"46",X"06",
		X"78",X"DD",X"77",X"07",X"DF",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",
		X"74",X"03",X"C9",X"D3",X"08",X"D7",X"08",X"DB",X"08",X"DF",X"08",X"E3",X"08",X"E7",X"08",X"EB",
		X"08",X"EF",X"08",X"F3",X"08",X"F7",X"08",X"FB",X"08",X"FF",X"08",X"03",X"09",X"07",X"09",X"0B",
		X"09",X"0F",X"09",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",X"06",X"F3",
		X"05",X"9E",X"05",X"4E",X"05",X"01",X"05",X"B9",X"04",X"76",X"04",X"36",X"04",X"F9",X"03",X"C0",
		X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",
		X"02",X"3B",X"02",X"1B",X"02",X"FD",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",X"01",X"7D",
		X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",
		X"00",X"E3",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",
		X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",
		X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"04",X"08",X"34",X"2C",X"25",
		X"21",X"1D",X"1A",X"18",X"16",X"14",X"13",X"11",X"10",X"0F",X"0A",X"21",X"A5",X"42",X"7E",X"A7",
		X"C0",X"21",X"93",X"09",X"11",X"80",X"42",X"01",X"18",X"00",X"ED",X"B0",X"3A",X"A3",X"42",X"87",
		X"4F",X"87",X"81",X"4F",X"06",X"00",X"21",X"AB",X"09",X"09",X"11",X"82",X"42",X"CD",X"89",X"09",
		X"11",X"8A",X"42",X"CD",X"89",X"09",X"11",X"92",X"42",X"7E",X"12",X"CD",X"90",X"09",X"7E",X"12",
		X"23",X"13",X"C9",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"0A",X"6A",X"0A",X"8D",
		X"0A",X"CE",X"0A",X"E7",X"0A",X"3A",X"0B",X"FB",X"0A",X"19",X"0B",X"3A",X"0B",X"15",X"0C",X"3A",
		X"0B",X"3A",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"B5",X"0B",X"E6",X"0B",X"3A",X"0B",X"2A",
		X"0C",X"55",X"0C",X"3A",X"0B",X"7E",X"0C",X"BA",X"0C",X"3A",X"0B",X"EE",X"0C",X"1A",X"0D",X"3A",
		X"0B",X"43",X"0D",X"7B",X"0D",X"3A",X"0B",X"9F",X"0D",X"D2",X"0D",X"3A",X"0B",X"03",X"0E",X"5C",
		X"0E",X"3A",X"0B",X"81",X"0E",X"B0",X"0E",X"3A",X"0B",X"DD",X"0E",X"13",X"0F",X"3A",X"0B",X"47",
		X"0F",X"78",X"0F",X"3A",X"0B",X"A7",X"0F",X"E2",X"0F",X"3A",X"0B",X"74",X"11",X"C7",X"11",X"3A",
		X"0B",X"F1",X"11",X"17",X"12",X"3A",X"0B",X"18",X"12",X"40",X"12",X"3A",X"0B",X"66",X"12",X"92",
		X"12",X"3A",X"0B",X"BE",X"12",X"DD",X"12",X"3A",X"0B",X"F6",X"12",X"19",X"13",X"3A",X"0B",X"3A",
		X"13",X"7A",X"13",X"3A",X"0B",X"B8",X"13",X"EC",X"13",X"3A",X"0B",X"1E",X"14",X"48",X"14",X"3A",
		X"0B",X"34",X"10",X"CA",X"10",X"3A",X"0B",X"1F",X"0B",X"3F",X"0A",X"5F",X"07",X"91",X"8D",X"8D",
		X"8D",X"91",X"8D",X"8D",X"8D",X"92",X"92",X"91",X"91",X"AF",X"A0",X"92",X"92",X"91",X"91",X"8F",
		X"8F",X"96",X"96",X"94",X"92",X"91",X"8F",X"AD",X"A0",X"FF",X"1F",X"05",X"5F",X"07",X"8D",X"91",
		X"88",X"91",X"8D",X"91",X"88",X"91",X"8F",X"92",X"88",X"92",X"8F",X"92",X"88",X"92",X"8F",X"92",
		X"88",X"92",X"8F",X"92",X"88",X"92",X"8F",X"92",X"88",X"92",X"B1",X"A0",X"FF",X"1F",X"05",X"5F",
		X"07",X"80",X"8D",X"80",X"8D",X"80",X"8D",X"80",X"8D",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",
		X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"AD",X"A0",X"FF",
		X"E7",X"3E",X"01",X"32",X"A3",X"42",X"32",X"A6",X"42",X"F7",X"C3",X"61",X"09",X"DD",X"21",X"80",
		X"42",X"C3",X"A1",X"07",X"E7",X"F7",X"C9",X"DD",X"21",X"88",X"42",X"C3",X"A1",X"07",X"1F",X"0C",
		X"3F",X"0F",X"5F",X"07",X"AD",X"80",X"8A",X"B2",X"B2",X"B6",X"74",X"72",X"71",X"6F",X"CD",X"AB",
		X"AD",X"A8",X"AD",X"AA",X"AD",X"C6",X"FF",X"1F",X"06",X"5F",X"07",X"AA",X"AD",X"AA",X"AD",X"A6",
		X"AD",X"AA",X"AD",X"A8",X"AD",X"AB",X"AD",X"A6",X"AD",X"CA",X"FF",X"1F",X"0B",X"3F",X"0C",X"5F",
		X"07",X"8D",X"8F",X"91",X"92",X"B4",X"B1",X"8D",X"8F",X"91",X"8F",X"AD",X"AD",X"8D",X"8F",X"91",
		X"92",X"B4",X"B1",X"94",X"92",X"91",X"8F",X"CD",X"FF",X"1F",X"0B",X"5F",X"07",X"85",X"88",X"85",
		X"88",X"85",X"88",X"85",X"88",X"85",X"88",X"85",X"88",X"85",X"88",X"85",X"88",X"85",X"88",X"85",
		X"88",X"85",X"88",X"85",X"88",X"86",X"88",X"86",X"88",X"C5",X"FF",X"E7",X"AF",X"32",X"C8",X"42",
		X"3E",X"02",X"32",X"A3",X"42",X"32",X"A6",X"42",X"F7",X"C3",X"61",X"09",X"DD",X"21",X"80",X"42",
		X"C3",X"A1",X"07",X"E7",X"F7",X"C9",X"DD",X"21",X"88",X"42",X"C3",X"A1",X"07",X"E7",X"F7",X"C9",
		X"DD",X"21",X"90",X"42",X"C3",X"A1",X"07",X"E7",X"21",X"A7",X"42",X"34",X"7E",X"FE",X"01",X"28",
		X"10",X"FE",X"18",X"28",X"11",X"32",X"A3",X"42",X"F7",X"3E",X"01",X"32",X"A5",X"42",X"C3",X"61",
		X"09",X"36",X"05",X"7E",X"18",X"EF",X"36",X"04",X"3E",X"18",X"18",X"E9",X"E7",X"F7",X"C9",X"DD",
		X"21",X"80",X"42",X"C3",X"A1",X"07",X"DD",X"21",X"88",X"42",X"C3",X"A1",X"07",X"E7",X"3E",X"03",
		X"32",X"A3",X"42",X"F7",X"C3",X"5B",X"09",X"3A",X"A5",X"42",X"A7",X"C2",X"B4",X"07",X"DD",X"21",
		X"80",X"42",X"C3",X"A1",X"07",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"9B",X"60",X"7D",X"BB",X"A6",
		X"9B",X"60",X"7D",X"BB",X"B8",X"9B",X"60",X"7B",X"BD",X"80",X"9B",X"99",X"93",X"B8",X"A0",X"8F",
		X"60",X"6F",X"8F",X"93",X"B6",X"8F",X"60",X"6F",X"8F",X"94",X"B8",X"9B",X"60",X"7B",X"BD",X"80",
		X"9B",X"99",X"93",X"B4",X"A0",X"FF",X"1F",X"0B",X"5F",X"06",X"98",X"60",X"77",X"B8",X"B4",X"98",
		X"60",X"77",X"B8",X"B4",X"98",X"60",X"76",X"B5",X"80",X"95",X"96",X"97",X"B4",X"A0",X"8F",X"60",
		X"6F",X"8F",X"93",X"B6",X"8F",X"60",X"6D",X"8C",X"8F",X"B4",X"98",X"60",X"76",X"B4",X"80",X"93",
		X"8F",X"8D",X"AC",X"A0",X"FF",X"1F",X"0B",X"3F",X"0E",X"5F",X"06",X"8F",X"60",X"6F",X"93",X"96",
		X"BB",X"A0",X"98",X"60",X"78",X"9B",X"98",X"B6",X"A0",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",
		X"8D",X"96",X"B6",X"80",X"97",X"B6",X"94",X"8D",X"B4",X"8D",X"97",X"B7",X"80",X"99",X"B7",X"96",
		X"8D",X"B6",X"96",X"99",X"B9",X"80",X"9B",X"B9",X"97",X"96",X"94",X"92",X"91",X"94",X"9B",X"99",
		X"97",X"91",X"D2",X"A0",X"FF",X"1F",X"0B",X"5F",X"06",X"8D",X"92",X"B2",X"80",X"91",X"B2",X"91",
		X"8D",X"B1",X"8D",X"94",X"B4",X"80",X"96",X"B4",X"92",X"8D",X"B2",X"92",X"96",X"B6",X"80",X"97",
		X"B6",X"94",X"92",X"91",X"8F",X"8D",X"91",X"97",X"96",X"94",X"8D",X"D2",X"A0",X"FF",X"1F",X"0B",
		X"3F",X"0D",X"5F",X"06",X"C0",X"A0",X"94",X"60",X"75",X"96",X"9E",X"96",X"9E",X"B6",X"96",X"60",
		X"75",X"94",X"9D",X"94",X"9D",X"B4",X"9D",X"60",X"73",X"B2",X"BB",X"B9",X"B8",X"B9",X"BB",X"BD",
		X"94",X"60",X"75",X"96",X"92",X"96",X"92",X"B6",X"96",X"60",X"79",X"94",X"99",X"94",X"99",X"BD",
		X"94",X"60",X"74",X"B4",X"BB",X"B9",X"B8",X"D9",X"C0",X"FF",X"1F",X"05",X"5F",X"06",X"E0",X"B2",
		X"80",X"8D",X"92",X"AD",X"92",X"AD",X"80",X"88",X"8D",X"A8",X"8D",X"A8",X"80",X"88",X"88",X"A8",
		X"88",X"AD",X"80",X"88",X"8D",X"94",X"91",X"8D",X"B2",X"80",X"8D",X"92",X"AD",X"92",X"AD",X"80",
		X"88",X"8D",X"A8",X"8D",X"88",X"94",X"83",X"94",X"88",X"94",X"88",X"94",X"E0",X"FF",X"1F",X"0B",
		X"3F",X"0D",X"5F",X"06",X"B8",X"80",X"96",X"96",X"94",X"B3",X"B1",X"80",X"AF",X"8D",X"AC",X"CA",
		X"AF",X"B6",X"DB",X"9B",X"80",X"8C",X"8D",X"AF",X"B8",X"94",X"80",X"8C",X"8D",X"AF",X"B8",X"94",
		X"80",X"98",X"99",X"B8",X"B6",X"B8",X"B6",X"D4",X"A0",X"FF",X"1F",X"05",X"5F",X"06",X"A3",X"80",
		X"AF",X"8F",X"AF",X"A3",X"80",X"AF",X"8F",X"AF",X"A3",X"AF",X"AF",X"AF",X"A3",X"AF",X"8F",X"8F",
		X"83",X"83",X"A8",X"B4",X"A8",X"B4",X"A8",X"B4",X"A8",X"B4",X"AA",X"B3",X"AF",X"B3",X"B4",X"AF",
		X"88",X"80",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"98",X"98",X"98",X"98",X"98",X"98",X"96",
		X"98",X"99",X"B1",X"80",X"B1",X"B1",X"96",X"96",X"96",X"96",X"B6",X"94",X"96",X"98",X"AF",X"80",
		X"AF",X"AF",X"98",X"98",X"98",X"98",X"98",X"98",X"96",X"98",X"99",X"99",X"99",X"99",X"B1",X"91",
		X"94",X"93",X"B3",X"80",X"8F",X"8F",X"98",X"96",X"D4",X"A0",X"FF",X"1F",X"05",X"5F",X"06",X"A8",
		X"80",X"88",X"C8",X"AA",X"80",X"8A",X"CA",X"AF",X"80",X"8F",X"CF",X"B4",X"80",X"8F",X"AF",X"AC",
		X"A8",X"80",X"88",X"C8",X"AA",X"80",X"8A",X"CA",X"A3",X"80",X"83",X"C3",X"A8",X"C0",X"FF",X"1F",
		X"0B",X"3F",X"0D",X"5F",X"06",X"94",X"60",X"72",X"91",X"94",X"B9",X"9B",X"99",X"96",X"99",X"AF",
		X"9B",X"60",X"79",X"98",X"60",X"76",X"94",X"94",X"96",X"94",X"D4",X"94",X"60",X"72",X"91",X"94",
		X"B9",X"9B",X"99",X"96",X"99",X"AF",X"9B",X"60",X"79",X"98",X"60",X"76",X"94",X"94",X"96",X"98",
		X"D9",X"FF",X"1F",X"0B",X"5F",X"06",X"94",X"60",X"72",X"91",X"94",X"B9",X"98",X"94",X"92",X"91",
		X"B2",X"92",X"60",X"76",X"94",X"60",X"74",X"92",X"92",X"92",X"92",X"D1",X"94",X"60",X"72",X"91",
		X"94",X"B9",X"98",X"94",X"92",X"91",X"B2",X"92",X"60",X"76",X"94",X"60",X"74",X"92",X"92",X"92",
		X"92",X"D1",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"88",X"86",X"65",X"68",X"6D",X"71",X"B4",
		X"80",X"92",X"71",X"74",X"6D",X"71",X"A8",X"80",X"91",X"6F",X"72",X"6C",X"6F",X"A8",X"80",X"92",
		X"71",X"74",X"6D",X"71",X"A8",X"88",X"60",X"66",X"65",X"68",X"6D",X"71",X"B4",X"8D",X"60",X"6B",
		X"6A",X"6D",X"72",X"76",X"B9",X"98",X"96",X"94",X"60",X"71",X"96",X"60",X"71",X"94",X"60",X"71",
		X"72",X"68",X"6C",X"6F",X"B4",X"80",X"92",X"71",X"68",X"6D",X"71",X"B4",X"80",X"91",X"6F",X"68",
		X"71",X"60",X"6F",X"68",X"71",X"60",X"6F",X"68",X"74",X"60",X"D9",X"FF",X"1F",X"0B",X"5F",X"06",
		X"A0",X"AD",X"AC",X"A0",X"AA",X"A8",X"A0",X"A6",X"A5",X"A0",X"A8",X"A6",X"A0",X"AD",X"A7",X"A0",
		X"AA",X"A8",X"A0",X"A5",X"A6",X"A5",X"A8",X"A6",X"A0",X"A8",X"A5",X"A0",X"A6",X"A8",X"A6",X"C5",
		X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"94",X"99",X"99",X"9B",X"9B",X"9D",X"9D",X"98",X"9B",
		X"B9",X"B6",X"B4",X"80",X"92",X"91",X"8F",X"91",X"92",X"94",X"B4",X"99",X"98",X"94",X"96",X"98",
		X"B9",X"80",X"92",X"91",X"8F",X"91",X"92",X"94",X"B4",X"99",X"98",X"94",X"96",X"98",X"B9",X"FF",
		X"1F",X"0B",X"5F",X"06",X"94",X"94",X"94",X"94",X"94",X"94",X"94",X"92",X"92",X"B1",X"B3",X"B4",
		X"80",X"8F",X"8D",X"8C",X"8D",X"8F",X"8F",X"8F",X"B4",X"92",X"92",X"92",X"92",X"B1",X"80",X"8F",
		X"8D",X"8C",X"8D",X"8F",X"8F",X"8F",X"B4",X"92",X"92",X"92",X"92",X"B1",X"FF",X"1F",X"0B",X"3F",
		X"0D",X"5F",X"06",X"87",X"60",X"68",X"AA",X"80",X"8F",X"8E",X"60",X"6C",X"CA",X"8F",X"60",X"6F",
		X"6E",X"71",X"94",X"9A",X"60",X"78",X"96",X"8E",X"8F",X"93",X"8A",X"80",X"87",X"60",X"68",X"AA",
		X"80",X"8F",X"8E",X"60",X"6C",X"CA",X"8F",X"60",X"6F",X"6E",X"71",X"94",X"9A",X"60",X"78",X"96",
		X"8E",X"CF",X"FF",X"1F",X"0B",X"5F",X"06",X"87",X"60",X"68",X"AA",X"80",X"8F",X"8E",X"60",X"6C",
		X"CA",X"8F",X"60",X"6F",X"6E",X"6E",X"91",X"96",X"60",X"74",X"91",X"88",X"87",X"88",X"87",X"80",
		X"87",X"60",X"68",X"AA",X"80",X"87",X"88",X"60",X"68",X"C7",X"8F",X"60",X"6F",X"6E",X"6E",X"91",
		X"96",X"60",X"74",X"91",X"88",X"C7",X"FF",X"1F",X"0B",X"3F",X"0D",X"5F",X"06",X"8A",X"8F",X"8E",
		X"91",X"AA",X"8C",X"8E",X"8F",X"93",X"AA",X"8A",X"8F",X"8E",X"91",X"AA",X"8C",X"8E",X"8F",X"93",
		X"AA",X"87",X"60",X"68",X"AA",X"80",X"8F",X"8E",X"60",X"6C",X"CA",X"8F",X"60",X"6F",X"6E",X"71",
		X"94",X"9A",X"60",X"78",X"96",X"8E",X"CF",X"FF",X"1F",X"0B",X"5F",X"06",X"8A",X"87",X"88",X"88",
		X"A8",X"88",X"88",X"87",X"8A",X"A7",X"87",X"87",X"88",X"88",X"A8",X"88",X"88",X"87",X"8A",X"A7",
		X"87",X"60",X"68",X"AA",X"80",X"87",X"88",X"60",X"68",X"C7",X"8F",X"60",X"6F",X"6E",X"6E",X"91",
		X"96",X"60",X"74",X"91",X"88",X"C7",X"FF",X"1F",X"0B",X"3F",X"0C",X"5F",X"06",X"B4",X"91",X"8D",
		X"B9",X"98",X"96",X"B4",X"99",X"91",X"8F",X"B4",X"80",X"94",X"94",X"94",X"94",X"96",X"94",X"91",
		X"8D",X"99",X"99",X"99",X"99",X"9B",X"99",X"96",X"92",X"94",X"94",X"94",X"94",X"96",X"94",X"91",
		X"8D",X"99",X"99",X"99",X"99",X"9B",X"99",X"96",X"92",X"94",X"91",X"80",X"91",X"B9",X"B1",X"94",
		X"CF",X"FF",X"1F",X"05",X"5F",X"06",X"D9",X"D6",X"D9",X"D8",X"8D",X"91",X"88",X"91",X"8D",X"91",
		X"88",X"91",X"8D",X"92",X"8A",X"92",X"8D",X"92",X"8A",X"92",X"8D",X"91",X"88",X"91",X"8D",X"91");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
