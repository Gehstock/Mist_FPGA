library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity satans_hollow_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of satans_hollow_sp_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"77",X"7E",
		X"00",X"00",X"76",X"7E",X"00",X"00",X"76",X"7D",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"D7",X"00",X"DD",X"DD",X"66",X"DD",X"66",X"DD",
		X"66",X"77",X"66",X"DD",X"77",X"00",X"77",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"77",X"00",X"00",X"77",X"70",X"00",X"00",X"76",X"7E",X"00",X"00",X"76",X"7E",
		X"00",X"00",X"77",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"77",X"7E",
		X"00",X"00",X"76",X"7E",X"00",X"60",X"76",X"7D",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"00",X"D0",X"DD",X"DD",X"66",X"7D",X"66",X"DD",
		X"66",X"77",X"66",X"DD",X"00",X"70",X"77",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"77",X"00",X"00",X"77",X"70",X"00",X"00",X"76",X"7E",X"00",X"00",X"76",X"7E",
		X"00",X"00",X"77",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"77",X"77",X"7E",
		X"00",X"67",X"76",X"7E",X"00",X"67",X"76",X"7D",X"00",X"77",X"77",X"70",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"D7",X"00",X"DD",X"DD",X"66",X"DD",X"66",X"DD",
		X"66",X"77",X"66",X"DD",X"77",X"00",X"77",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"77",X"00",X"00",X"77",X"70",X"00",X"00",X"76",X"7E",X"00",X"00",X"76",X"7E",
		X"00",X"00",X"77",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"DD",X"00",X"77",X"7E",
		X"00",X"DD",X"76",X"7E",X"00",X"77",X"76",X"7D",X"77",X"00",X"77",X"70",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"00",X"DD",X"DD",X"DD",X"66",X"0D",X"66",X"DD",
		X"66",X"07",X"66",X"DD",X"00",X"77",X"77",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"77",X"00",X"00",X"77",X"70",X"00",X"00",X"76",X"7E",X"00",X"00",X"76",X"7E",
		X"00",X"00",X"77",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"77",X"77",X"7E",
		X"00",X"67",X"76",X"7E",X"00",X"67",X"76",X"7D",X"00",X"77",X"77",X"70",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"D7",X"00",X"DD",X"DD",X"66",X"DD",X"66",X"DD",
		X"66",X"77",X"66",X"DD",X"77",X"00",X"77",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"77",X"00",X"77",X"77",X"70",X"00",X"67",X"76",X"7E",X"00",X"67",X"76",X"7E",
		X"00",X"77",X"77",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"DD",X"00",X"77",X"7E",
		X"00",X"DD",X"76",X"7E",X"00",X"77",X"76",X"7D",X"77",X"00",X"77",X"70",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"00",X"DD",X"DD",X"DD",X"66",X"07",X"66",X"DD",
		X"66",X"07",X"66",X"DD",X"00",X"77",X"77",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D7",
		X"00",X"00",X"00",X"77",X"DD",X"00",X"77",X"70",X"00",X"DD",X"76",X"7E",X"00",X"77",X"76",X"7E",
		X"77",X"00",X"77",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",
		X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"41",X"00",X"00",X"00",X"33",X"00",X"00",X"01",X"13",X"00",X"00",X"14",X"13",X"11",
		X"00",X"01",X"01",X"44",X"01",X"00",X"00",X"32",X"00",X"10",X"10",X"32",X"00",X"F1",X"10",X"32",
		X"00",X"6F",X"41",X"32",X"00",X"11",X"41",X"11",X"00",X"33",X"33",X"00",X"00",X"11",X"43",X"00",
		X"00",X"1F",X"41",X"00",X"00",X"F1",X"41",X"00",X"00",X"11",X"11",X"11",X"01",X"13",X"14",X"43",
		X"00",X"43",X"14",X"14",X"00",X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"1C",X"14",X"00",X"00",X"CC",X"42",X"00",X"00",X"CC",X"23",X"00",X"00",X"1C",X"31",X"00",X"00",
		X"1C",X"10",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"C9",
		X"00",X"00",X"9C",X"CC",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"CC",X"0F",X"00",X"00",X"CC",X"0F",X"00",X"00",X"C9",X"0F",X"00",X"00",X"90",X"0F",
		X"00",X"00",X"90",X"0F",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"FC",X"00",X"00",X"99",X"F9",
		X"00",X"00",X"99",X"0F",X"00",X"00",X"FF",X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"0C",X"00",X"00",X"99",X"FF",X"00",X"00",X"CC",X"F0",X"00",X"0F",X"99",X"00",
		X"00",X"99",X"FF",X"00",X"00",X"99",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"90",X"99",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9B",X"99",X"0F",X"99",X"9B",X"99",X"FF",X"90",X"9B",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"00",X"CC",X"C0",
		X"00",X"00",X"CF",X"CC",X"00",X"00",X"CF",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"CC",X"C0",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"90",X"00",
		X"00",X"05",X"06",X"60",X"00",X"90",X"06",X"66",X"00",X"9F",X"F6",X"C6",X"00",X"95",X"F6",X"CC",
		X"00",X"9F",X"66",X"CC",X"00",X"55",X"6F",X"CC",X"00",X"09",X"60",X"CC",X"00",X"F9",X"66",X"CC",
		X"00",X"90",X"C6",X"CC",X"00",X"00",X"66",X"C6",X"00",X"00",X"C6",X"C6",X"00",X"00",X"CC",X"C6",
		X"00",X"00",X"CC",X"66",X"00",X"00",X"CC",X"60",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",
		X"00",X"BC",X"BB",X"00",X"00",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"9C",X"C0",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"09",X"99",X"09",X"22",X"00",X"00",X"99",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"09",X"90",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"11",X"11",X"00",X"00",X"1C",X"B1",X"00",X"0C",X"1C",X"99",X"00",X"00",X"11",X"BB",X"B0",
		X"00",X"11",X"B9",X"B9",X"09",X"11",X"B1",X"91",X"0B",X"11",X"9B",X"11",X"B9",X"11",X"BB",X"A1",
		X"9B",X"91",X"11",X"9A",X"9B",X"B9",X"11",X"11",X"9B",X"BB",X"99",X"A1",X"9B",X"BB",X"BB",X"A1",
		X"9B",X"BB",X"BB",X"11",X"9B",X"B9",X"B1",X"9A",X"99",X"91",X"BB",X"A1",X"9B",X"91",X"BB",X"11",
		X"9B",X"11",X"BB",X"91",X"09",X"11",X"BB",X"B9",X"09",X"11",X"B9",X"00",X"00",X"1C",X"91",X"00",
		X"0C",X"1C",X"11",X"00",X"00",X"11",X"1B",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"09",X"00",X"00",X"00",X"91",X"00",
		X"00",X"00",X"91",X"00",X"0C",X"77",X"77",X"77",X"CC",X"FF",X"FF",X"FF",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"B9",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"91",X"00",X"00",X"BB",X"11",
		X"00",X"00",X"9B",X"11",X"00",X"00",X"99",X"1A",X"00",X"00",X"9B",X"1C",X"00",X"00",X"0A",X"1C",
		X"00",X"00",X"AA",X"1C",X"00",X"00",X"A0",X"CC",X"00",X"00",X"00",X"C1",X"00",X"00",X"00",X"1B",
		X"00",X"00",X"09",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"A1",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"BB",X"1A",X"00",X"00",
		X"BB",X"A1",X"00",X"00",X"BB",X"11",X"00",X"00",X"9B",X"B0",X"00",X"00",X"B1",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"F9",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"99",
		X"88",X"88",X"88",X"79",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"F9",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"77",X"88",X"88",X"88",X"99",
		X"88",X"88",X"8F",X"99",X"88",X"88",X"F9",X"99",X"88",X"88",X"99",X"79",X"88",X"88",X"99",X"99",
		X"88",X"88",X"FF",X"97",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"97",X"88",X"88",X"88",X"99",
		X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"97",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"99",
		X"88",X"88",X"88",X"77",X"88",X"88",X"88",X"97",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"F9",
		X"88",X"88",X"F8",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"09",X"BB",X"B1",X"00",X"09",X"BB",X"B1",X"00",X"09",X"BB",X"91",X"00",X"09",X"BB",X"91",
		X"00",X"00",X"BB",X"1C",X"00",X"00",X"BB",X"CA",X"00",X"00",X"BB",X"CA",X"00",X"00",X"BB",X"AA",
		X"00",X"00",X"AB",X"CA",X"00",X"00",X"AB",X"CA",X"00",X"00",X"BB",X"C1",X"00",X"00",X"BB",X"1B",
		X"00",X"00",X"B9",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"0C",X"BB",X"BB",X"00",X"0C",X"BB",X"BB",
		X"00",X"C0",X"BB",X"9B",X"00",X"00",X"11",X"99",X"00",X"00",X"19",X"09",X"00",X"00",X"19",X"00",
		X"00",X"09",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"19",X"1C",X"00",X"11",X"B9",X"11",X"00",X"11",X"B9",X"11",X"00",X"BB",X"B9",X"1C",X"00",
		X"BB",X"B9",X"19",X"00",X"1B",X"BB",X"B9",X"00",X"9B",X"B1",X"91",X"00",X"BB",X"BB",X"11",X"00",
		X"B9",X"BB",X"B0",X"00",X"BB",X"9B",X"00",X"00",X"99",X"11",X"00",X"00",X"9B",X"11",X"00",X"00",
		X"99",X"10",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"0D",X"0D",X"00",X"00",X"0D",X"DD",X"00",
		X"00",X"0D",X"DD",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"03",X"90",X"22",
		X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"22",X"00",X"32",X"03",X"33",X"00",X"23",X"33",X"33",
		X"00",X"02",X"33",X"22",X"00",X"00",X"22",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"02",X"33",
		X"00",X"00",X"02",X"30",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",
		X"00",X"55",X"CC",X"00",X"00",X"55",X"CC",X"00",X"00",X"55",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"55",X"00",
		X"00",X"09",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"05",X"55",X"00",X"00",X"00",X"C5",X"00",X"00",X"00",X"C5",X"99",X"00",X"00",X"CC",X"99",
		X"00",X"5C",X"CC",X"50",X"00",X"5C",X"C5",X"00",X"00",X"00",X"C5",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"9C",X"00",
		X"D9",X"55",X"99",X"CC",X"D9",X"55",X"99",X"5C",X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",X"95",
		X"90",X"55",X"CC",X"55",X"90",X"55",X"CC",X"55",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"55",X"99",X"55",X"00",X"55",X"99",X"95",X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",X"99",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"55",X"CC",X"CC",X"00",X"55",X"CC",X"CC",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"55",
		X"CC",X"55",X"99",X"99",X"CC",X"55",X"99",X"59",X"CC",X"55",X"99",X"99",X"CC",X"55",X"99",X"55",
		X"65",X"55",X"99",X"55",X"65",X"55",X"99",X"55",X"CC",X"99",X"9F",X"55",X"CC",X"99",X"FF",X"55",
		X"00",X"99",X"9F",X"99",X"00",X"99",X"9F",X"99",X"00",X"99",X"FF",X"55",X"00",X"99",X"FF",X"55",
		X"00",X"55",X"99",X"CC",X"00",X"55",X"99",X"CC",X"CC",X"55",X"99",X"55",X"CC",X"55",X"99",X"55",
		X"CC",X"55",X"55",X"99",X"CC",X"55",X"55",X"99",X"00",X"99",X"CC",X"55",X"00",X"99",X"CC",X"55",
		X"00",X"55",X"CC",X"CC",X"00",X"55",X"CC",X"CC",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"09",X"00",X"00",X"9F",X"99",X"90",X"99",X"FF",X"99",
		X"99",X"99",X"FF",X"99",X"9C",X"CC",X"FF",X"99",X"9C",X"CC",X"FF",X"C9",X"9F",X"C9",X"CC",X"99",
		X"9F",X"CF",X"99",X"99",X"9F",X"9C",X"9C",X"F9",X"09",X"99",X"FF",X"99",X"00",X"F9",X"FC",X"99",
		X"00",X"FF",X"CC",X"99",X"00",X"9F",X"CC",X"99",X"00",X"F9",X"F9",X"99",X"00",X"F9",X"99",X"99",
		X"00",X"F9",X"99",X"99",X"00",X"FF",X"00",X"99",X"00",X"9F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"00",X"99",X"00",X"F9",X"99",X"99",
		X"00",X"F9",X"99",X"99",X"00",X"F9",X"F9",X"99",X"00",X"9F",X"CC",X"99",X"00",X"FF",X"99",X"99",
		X"00",X"99",X"FC",X"99",X"09",X"99",X"FF",X"99",X"9F",X"9C",X"9C",X"F9",X"9F",X"CF",X"99",X"99",
		X"99",X"C9",X"CC",X"99",X"9C",X"CC",X"FF",X"C9",X"9C",X"CC",X"99",X"99",X"99",X"99",X"99",X"99",
		X"90",X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"99",X"09",X"00",
		X"00",X"99",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"CC",X"00",X"09",X"09",X"0C",X"00",X"99",X"00",X"0C",X"09",X"99",X"99",
		X"0C",X"00",X"09",X"00",X"00",X"99",X"09",X"90",X"00",X"09",X"00",X"C0",X"00",X"00",X"00",X"CC",
		X"00",X"CC",X"99",X"99",X"00",X"CC",X"99",X"99",X"00",X"0C",X"00",X"99",X"00",X"00",X"C0",X"99",
		X"00",X"00",X"C0",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"09",X"33",X"03",X"22",X"00",X"00",X"33",X"33",
		X"00",X"00",X"22",X"33",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"32",X"00",X"30",
		X"00",X"33",X"00",X"30",X"00",X"03",X"20",X"33",X"00",X"00",X"22",X"33",X"00",X"00",X"33",X"33",
		X"00",X"00",X"33",X"33",X"00",X"00",X"03",X"33",X"00",X"00",X"22",X"33",X"00",X"00",X"32",X"33",
		X"00",X"02",X"33",X"33",X"00",X"22",X"22",X"33",X"00",X"33",X"22",X"00",X"00",X"33",X"32",X"00",
		X"00",X"33",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"99",X"00",X"00",X"03",X"30",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"30",X"00",X"00",X"20",X"30",X"00",X"00",X"22",X"30",X"00",X"00",X"33",X"33",
		X"00",X"22",X"33",X"33",X"00",X"33",X"03",X"33",X"00",X"33",X"22",X"33",X"00",X"33",X"22",X"33",
		X"00",X"03",X"33",X"33",X"00",X"00",X"32",X"33",X"00",X"00",X"22",X"33",X"00",X"00",X"22",X"33",
		X"00",X"00",X"32",X"03",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"33",X"49",X"00",X"00",X"32",X"41",
		X"00",X"20",X"20",X"49",X"00",X"32",X"20",X"44",X"00",X"03",X"20",X"00",X"00",X"03",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"06",X"33",X"00",X"00",X"06",X"33",X"00",
		X"00",X"06",X"23",X"00",X"00",X"06",X"23",X"00",X"00",X"06",X"22",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"20",X"00",X"00",X"02",X"22",X"00",
		X"00",X"02",X"22",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"30",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"20",X"20",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"03",X"30",X"00",
		X"00",X"03",X"06",X"00",X"00",X"03",X"06",X"00",X"00",X"03",X"66",X"00",X"00",X"03",X"66",X"00",
		X"00",X"03",X"06",X"00",X"00",X"03",X"06",X"00",X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"03",X"00",X"04",X"00",X"33",X"00",X"34",X"00",X"33",X"00",X"44",X"00",X"33",X"00",X"24",
		X"00",X"33",X"00",X"04",X"00",X"33",X"00",X"00",X"00",X"33",X"03",X"00",X"00",X"33",X"32",X"00",
		X"00",X"32",X"32",X"00",X"00",X"32",X"20",X"00",X"00",X"32",X"20",X"00",X"00",X"32",X"00",X"22",
		X"00",X"33",X"00",X"23",X"00",X"33",X"00",X"33",X"00",X"33",X"22",X"30",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"32",X"00",X"00",X"33",X"23",X"00",X"00",X"30",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"49",X"00",X"03",X"00",X"41",
		X"00",X"03",X"00",X"49",X"00",X"33",X"00",X"44",X"00",X"32",X"00",X"00",X"00",X"32",X"03",X"00",
		X"00",X"32",X"32",X"00",X"00",X"32",X"32",X"00",X"00",X"32",X"22",X"00",X"00",X"33",X"20",X"00",
		X"00",X"33",X"20",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"23",X"22",X"00",
		X"00",X"23",X"33",X"00",X"00",X"33",X"33",X"22",X"00",X"00",X"22",X"32",X"00",X"00",X"33",X"33",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"9C",X"00",X"00",X"99",X"9C",X"00",X"00",X"90",X"9C",
		X"00",X"00",X"90",X"9C",X"00",X"0C",X"00",X"9C",X"00",X"CC",X"99",X"9C",X"00",X"99",X"99",X"9C",
		X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"90",X"00",X"99",X"09",X"90",X"0C",X"00",X"09",X"00",
		X"0C",X"09",X"9F",X"FF",X"0C",X"99",X"00",X"00",X"CC",X"FF",X"99",X"00",X"CC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"88",X"80",X"00",X"00",X"88",X"88",X"00",
		X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",
		X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"80",X"08",X"88",X"88",X"88",X"08",X"C8",X"58",X"88",
		X"08",X"89",X"88",X"88",X"08",X"95",X"88",X"88",X"88",X"C9",X"CC",X"88",X"08",X"99",X"98",X"88",
		X"08",X"C5",X"9C",X"88",X"08",X"95",X"58",X"88",X"08",X"9C",X"85",X"88",X"08",X"89",X"88",X"88",
		X"08",X"88",X"88",X"88",X"08",X"88",X"88",X"88",X"00",X"88",X"88",X"80",X"00",X"88",X"88",X"00",
		X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",
		X"00",X"88",X"88",X"00",X"00",X"88",X"80",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"90",X"99",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9B",X"99",X"0F",X"99",X"9B",X"99",X"FF",X"90",X"9B",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"09",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"C9",X"00",
		X"00",X"CC",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"0C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"55",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"92",X"00",X"90",
		X"00",X"99",X"00",X"90",X"00",X"09",X"20",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",
		X"00",X"02",X"99",X"99",X"00",X"22",X"22",X"99",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EF",
		X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"99",X"99",X"99",X"EE",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"FE",
		X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"30",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"20",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"99",
		X"00",X"22",X"99",X"99",X"00",X"99",X"09",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",
		X"00",X"09",X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"92",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"99",X"49",X"00",X"00",X"92",X"41",
		X"00",X"20",X"20",X"49",X"00",X"92",X"20",X"44",X"00",X"09",X"20",X"00",X"00",X"09",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"06",X"99",X"00",X"00",X"06",X"99",X"00",
		X"00",X"06",X"29",X"00",X"00",X"06",X"29",X"00",X"00",X"06",X"22",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"20",X"00",X"00",X"02",X"22",X"00",
		X"00",X"02",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"30",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"20",X"20",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"90",X"00",
		X"00",X"09",X"06",X"00",X"00",X"09",X"06",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",
		X"00",X"09",X"06",X"00",X"00",X"09",X"06",X"00",X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"09",X"00",X"04",X"00",X"99",X"00",X"34",X"00",X"99",X"00",X"44",X"00",X"99",X"00",X"24",
		X"00",X"99",X"00",X"04",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"92",X"00",
		X"00",X"92",X"92",X"00",X"00",X"92",X"20",X"00",X"00",X"92",X"20",X"00",X"00",X"92",X"00",X"22",
		X"00",X"99",X"00",X"29",X"00",X"99",X"00",X"99",X"00",X"99",X"22",X"90",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"49",X"00",X"09",X"00",X"41",
		X"00",X"09",X"00",X"49",X"00",X"99",X"00",X"44",X"00",X"92",X"00",X"00",X"00",X"92",X"09",X"00",
		X"00",X"92",X"92",X"00",X"00",X"92",X"92",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"20",X"00",
		X"00",X"99",X"20",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"29",X"22",X"00",
		X"00",X"29",X"99",X"00",X"00",X"99",X"99",X"22",X"00",X"00",X"22",X"92",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
