library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity nrx_nchr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of nrx_nchr_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"66",X"33",X"33",X"33",X"22",X"CC",X"00",X"11",X"22",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"00",
		X"EE",X"33",X"77",X"EE",X"CC",X"00",X"FF",X"00",X"33",X"66",X"00",X"11",X"33",X"77",X"77",X"00",
		X"FF",X"66",X"CC",X"EE",X"33",X"33",X"EE",X"00",X"33",X"00",X"00",X"11",X"00",X"66",X"33",X"00",
		X"EE",X"EE",X"66",X"66",X"FF",X"66",X"66",X"00",X"00",X"11",X"33",X"66",X"77",X"00",X"00",X"00",
		X"EE",X"00",X"EE",X"33",X"33",X"33",X"EE",X"00",X"77",X"66",X"77",X"00",X"00",X"66",X"33",X"00",
		X"EE",X"00",X"00",X"EE",X"33",X"33",X"EE",X"00",X"11",X"33",X"66",X"77",X"66",X"66",X"33",X"00",
		X"FF",X"33",X"66",X"CC",X"88",X"88",X"88",X"00",X"77",X"66",X"00",X"00",X"11",X"11",X"11",X"00",
		X"CC",X"22",X"22",X"CC",X"FF",X"33",X"EE",X"00",X"33",X"66",X"77",X"33",X"44",X"44",X"33",X"00",
		X"EE",X"33",X"33",X"FF",X"33",X"66",X"CC",X"00",X"33",X"66",X"66",X"33",X"00",X"00",X"33",X"00",
		X"CC",X"66",X"33",X"33",X"FF",X"33",X"33",X"00",X"11",X"33",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"EE",X"33",X"33",X"EE",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"77",X"00",
		X"EE",X"33",X"00",X"00",X"00",X"33",X"EE",X"00",X"11",X"33",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"66",X"33",X"33",X"33",X"66",X"CC",X"00",X"77",X"66",X"66",X"66",X"66",X"66",X"77",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"99",X"11",X"11",X"99",X"22",X"CC",X"33",X"44",X"99",X"AA",X"AA",X"99",X"44",X"33",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"07",X"07",X"00",X"0F",X"0F",X"0C",X"0F",X"0F",X"08",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"01",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"0F",X"0F",X"01",X"0F",X"0F",X"01",X"0F",X"0F",
		X"0F",X"0F",X"09",X"09",X"09",X"09",X"09",X"09",X"0F",X"0F",X"09",X"09",X"09",X"09",X"09",X"09",
		X"0F",X"0F",X"08",X"08",X"08",X"08",X"0F",X"0F",X"00",X"09",X"09",X"09",X"09",X"09",X"09",X"08",
		X"03",X"07",X"06",X"06",X"06",X"06",X"07",X"03",X"0E",X"0E",X"00",X"00",X"00",X"00",X"0E",X"0E",
		X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"0F",X"0F",X"01",X"01",X"01",X"01",X"0F",X"0F",
		X"EE",X"11",X"DD",X"55",X"FF",X"00",X"EE",X"00",X"33",X"44",X"55",X"55",X"55",X"44",X"33",X"00",
		X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"00",X"33",X"33",
		X"66",X"66",X"22",X"44",X"00",X"00",X"00",X"00",X"33",X"33",X"11",X"22",X"00",X"00",X"00",X"00",
		X"66",X"66",X"FF",X"66",X"FF",X"66",X"66",X"00",X"33",X"33",X"77",X"33",X"77",X"33",X"33",X"00",
		X"88",X"EE",X"88",X"EE",X"BB",X"EE",X"88",X"00",X"00",X"33",X"66",X"33",X"00",X"33",X"00",X"00",
		X"11",X"22",X"44",X"88",X"33",X"55",X"77",X"00",X"77",X"55",X"66",X"00",X"11",X"22",X"44",X"00",
		X"00",X"88",X"88",X"33",X"AA",X"44",X"BB",X"00",X"33",X"44",X"55",X"33",X"66",X"44",X"33",X"00",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"11",X"00",X"00",X"00",X"00",
		X"CC",X"88",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"11",X"33",X"33",X"33",X"11",X"00",X"00",
		X"88",X"CC",X"66",X"66",X"66",X"CC",X"88",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"88",X"AA",X"CC",X"88",X"CC",X"AA",X"88",X"00",X"00",X"22",X"11",X"00",X"11",X"22",X"00",X"00",
		X"00",X"88",X"88",X"EE",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"22",X"00",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"66",X"33",X"33",X"33",X"22",X"CC",X"00",X"11",X"22",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"00",
		X"EE",X"33",X"77",X"EE",X"CC",X"00",X"FF",X"00",X"33",X"66",X"00",X"11",X"33",X"77",X"77",X"00",
		X"FF",X"66",X"CC",X"EE",X"33",X"33",X"EE",X"00",X"33",X"00",X"00",X"11",X"00",X"66",X"33",X"00",
		X"EE",X"EE",X"66",X"66",X"FF",X"66",X"66",X"00",X"00",X"11",X"33",X"66",X"77",X"00",X"00",X"00",
		X"EE",X"00",X"EE",X"33",X"33",X"33",X"EE",X"00",X"77",X"66",X"77",X"00",X"00",X"66",X"33",X"00",
		X"EE",X"00",X"00",X"EE",X"33",X"33",X"EE",X"00",X"11",X"33",X"66",X"77",X"66",X"66",X"33",X"00",
		X"FF",X"33",X"66",X"CC",X"88",X"88",X"88",X"00",X"77",X"66",X"00",X"00",X"11",X"11",X"11",X"00",
		X"CC",X"22",X"22",X"CC",X"FF",X"33",X"EE",X"00",X"33",X"66",X"77",X"33",X"44",X"44",X"33",X"00",
		X"EE",X"33",X"33",X"FF",X"33",X"66",X"CC",X"00",X"33",X"66",X"66",X"33",X"00",X"00",X"33",X"00",
		X"00",X"88",X"88",X"00",X"88",X"88",X"00",X"00",X"00",X"11",X"11",X"00",X"11",X"11",X"00",X"00",
		X"00",X"88",X"88",X"00",X"88",X"88",X"00",X"00",X"00",X"11",X"11",X"00",X"11",X"00",X"11",X"00",
		X"66",X"CC",X"88",X"00",X"88",X"CC",X"66",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"77",X"77",X"00",X"77",X"77",X"00",X"00",
		X"00",X"88",X"CC",X"66",X"CC",X"88",X"00",X"00",X"33",X"11",X"00",X"00",X"00",X"11",X"33",X"00",
		X"EE",X"33",X"33",X"66",X"CC",X"00",X"CC",X"CC",X"33",X"66",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"66",X"33",X"33",X"FF",X"33",X"33",X"00",X"11",X"33",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"EE",X"33",X"33",X"EE",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"77",X"00",
		X"EE",X"33",X"00",X"00",X"00",X"33",X"EE",X"00",X"11",X"33",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"66",X"33",X"33",X"33",X"66",X"CC",X"00",X"77",X"66",X"66",X"66",X"66",X"66",X"77",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"FF",X"00",X"00",X"77",X"33",X"33",X"FF",X"00",X"11",X"33",X"66",X"66",X"66",X"33",X"11",X"00",
		X"33",X"33",X"33",X"FF",X"33",X"33",X"33",X"00",X"66",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"33",X"00",
		X"33",X"66",X"CC",X"88",X"CC",X"EE",X"77",X"00",X"66",X"66",X"66",X"77",X"77",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"33",X"77",X"FF",X"FF",X"BB",X"33",X"33",X"00",X"66",X"77",X"77",X"77",X"66",X"66",X"66",X"00",
		X"33",X"33",X"BB",X"FF",X"FF",X"77",X"33",X"00",X"66",X"77",X"77",X"77",X"66",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"33",X"EE",X"00",X"00",X"00",X"77",X"66",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"33",X"FF",X"66",X"DD",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"77",X"CC",X"EE",X"77",X"00",X"77",X"66",X"66",X"66",X"77",X"66",X"66",X"00",
		X"CC",X"66",X"00",X"EE",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"33",X"00",X"66",X"33",X"00",
		X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"33",X"33",X"33",X"77",X"EE",X"CC",X"88",X"00",X"66",X"66",X"66",X"77",X"33",X"11",X"00",X"00",
		X"33",X"33",X"BB",X"FF",X"FF",X"77",X"33",X"00",X"66",X"66",X"66",X"77",X"77",X"77",X"66",X"00",
		X"33",X"77",X"EE",X"CC",X"EE",X"77",X"33",X"00",X"66",X"77",X"33",X"11",X"33",X"77",X"66",X"00",
		X"33",X"33",X"33",X"EE",X"CC",X"CC",X"CC",X"00",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"77",X"EE",X"CC",X"88",X"00",X"FF",X"00",X"77",X"00",X"00",X"11",X"33",X"77",X"77",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0F",X"0F",X"3F",X"BF",X"DB",X"FF",X"F6",X"FF",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"0F",X"3F",
		X"0F",X"EF",X"7F",X"96",X"F3",X"FF",X"F9",X"FF",X"0F",X"4F",X"FF",X"F3",X"FF",X"F7",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"87",X"8F",X"0F",X"4F",X"0F",X"0F",X"CF",X"87",X"FC",X"FF",X"BF",X"EF",
		X"FA",X"FB",X"FD",X"FF",X"B6",X"DB",X"EF",X"F6",X"7F",X"7E",X"3D",X"5F",X"7D",X"7D",X"3F",X"7E",
		X"F9",X"F7",X"FE",X"7F",X"FF",X"F9",X"EF",X"F7",X"F7",X"F7",X"9F",X"EF",X"FE",X"F5",X"7F",X"FF",
		X"EB",X"EB",X"CF",X"2F",X"EB",X"E7",X"EF",X"6F",X"FD",X"F3",X"FC",X"FF",X"F5",X"FB",X"EF",X"FB",
		X"7E",X"FF",X"FB",X"FD",X"7B",X"1F",X"0F",X"0F",X"3F",X"2F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"F9",X"EF",X"0F",X"CC",X"FF",X"FD",X"FD",X"17",X"E9",X"6F",X"0F",
		X"0F",X"CF",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"F7",X"FF",X"FA",X"F7",X"7F",X"0F",X"0F",X"0F",
		X"FF",X"5F",X"0F",X"8F",X"C3",X"F3",X"9F",X"3F",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"CF",X"FF",
		X"FF",X"EF",X"CF",X"CF",X"8F",X"FF",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"3F",X"1F",X"1F",X"1F",X"1F",X"3F",X"FF",X"3F",X"2F",X"2F",X"2F",X"79",X"F8",X"78",
		X"7F",X"FF",X"FF",X"DF",X"1F",X"3F",X"3C",X"FC",X"FF",X"FF",X"FF",X"FF",X"EF",X"CF",X"CF",X"EF",
		X"0F",X"0F",X"DF",X"6F",X"2F",X"0F",X"3F",X"3F",X"FF",X"BF",X"1F",X"0F",X"1F",X"9F",X"EF",X"C7",
		X"5F",X"9F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"78",X"F8",X"1E",X"1F",X"1F",X"3F",X"FF",X"FF",
		X"3C",X"3F",X"1F",X"1F",X"2F",X"6F",X"FF",X"FF",X"FF",X"EF",X"CF",X"CF",X"CF",X"EF",X"FF",X"FF",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"97",X"0F",X"0F",X"0F",X"1F",X"3F",X"FF",
		X"FF",X"7F",X"7F",X"9F",X"9F",X"1F",X"3F",X"FF",X"FF",X"CF",X"CF",X"3C",X"3C",X"1F",X"EF",X"FF",
		X"EE",X"7F",X"1D",X"9F",X"97",X"9F",X"3F",X"7F",X"EC",X"CF",X"8F",X"3E",X"38",X"3E",X"8F",X"CF",
		X"DD",X"7F",X"3F",X"9F",X"95",X"9F",X"3F",X"7F",X"FF",X"CF",X"8F",X"3E",X"34",X"3E",X"8F",X"CF",
		X"1D",X"1F",X"C7",X"C3",X"C7",X"1F",X"3F",X"FF",X"CD",X"CF",X"17",X"9E",X"9B",X"CF",X"EF",X"FF",
		X"EF",X"3F",X"1F",X"C7",X"C3",X"C7",X"1F",X"3F",X"33",X"EF",X"CF",X"9F",X"9E",X"9F",X"CF",X"EB",
		X"8B",X"7F",X"3F",X"9F",X"97",X"9F",X"3F",X"6F",X"6E",X"CF",X"8F",X"3E",X"3C",X"3E",X"8F",X"4F",
		X"7F",X"3F",X"9F",X"97",X"9F",X"3F",X"7F",X"FF",X"E6",X"8F",X"3E",X"3C",X"3E",X"8F",X"CF",X"FF",
		X"3F",X"1F",X"C7",X"C3",X"C7",X"1F",X"3E",X"FF",X"EF",X"CF",X"9F",X"9E",X"9F",X"CF",X"AF",X"FF",
		X"FF",X"7F",X"3F",X"9F",X"97",X"9F",X"3F",X"7F",X"FF",X"CF",X"8F",X"3E",X"3C",X"3E",X"8F",X"CF",
		X"7F",X"3F",X"9F",X"97",X"9F",X"3F",X"5D",X"FF",X"CF",X"8F",X"3E",X"3C",X"3E",X"8F",X"0B",X"FF",
		X"FF",X"FE",X"FE",X"FF",X"EF",X"FE",X"FC",X"ED",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F3",X"FF",X"FF",X"F7",X"F7",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"F7",X"FF",X"DF",X"CF",X"F8",X"BC",X"E8",X"BC",X"3C",
		X"E9",X"DF",X"F8",X"F8",X"F8",X"78",X"78",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FE",X"EF",X"D6",X"FF",X"FF",X"F3",X"B3",X"F1",X"B1",X"10",X"91",X"91",X"11",
		X"77",X"11",X"7F",X"77",X"31",X"75",X"FA",X"FF",X"78",X"E0",X"E3",X"E8",X"E0",X"E0",X"C0",X"EC",
		X"68",X"D2",X"F2",X"F6",X"FE",X"FE",X"FE",X"FF",X"FE",X"EF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"FB",X"FF",X"FE",X"FF",X"FF",X"31",X"90",X"B1",X"FC",X"77",X"77",X"77",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"EC",X"EC",X"FF",X"FF",X"F2",X"F0",X"FF",X"79",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"10",X"10",X"00",X"00",X"00",X"00",X"10",X"10",
		X"F0",X"F0",X"F0",X"F0",X"30",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"78",X"1E",X"78",X"F0",X"F0",X"F0",X"78",X"1E",X"0F",X"0F",X"0F",X"1E",X"78",
		X"F0",X"F0",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"3C",X"3C",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"FC",X"F6",X"F0",X"FC",X"F6",X"F6",X"FC",X"F0",X"F3",X"F6",X"F6",X"F3",X"F0",X"F6",X"F3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F2",X"FE",X"F0",X"F0",X"F6",X"F6",X"F6",X"F6",X"F6",X"F7",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F3",X"F7",X"EF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"60",X"40",X"F0",X"70",X"70",X"C0",X"B3",X"F0",X"E0",X"F0",X"C0",X"83",X"C1",X"E0",X"D0",
		X"F0",X"F0",X"30",X"DC",X"9C",X"0E",X"0F",X"0F",X"F0",X"F0",X"C0",X"B3",X"33",X"67",X"67",X"67",
		X"F0",X"F0",X"F0",X"F0",X"D0",X"70",X"38",X"38",X"F0",X"F0",X"90",X"F0",X"B0",X"C0",X"41",X"60",
		X"67",X"67",X"67",X"67",X"47",X"47",X"00",X"0D",X"F0",X"F0",X"F0",X"C0",X"83",X"83",X"81",X"C1",
		X"0F",X"0C",X"1F",X"2F",X"2F",X"4F",X"4F",X"0F",X"09",X"0D",X"0D",X"0D",X"0D",X"09",X"0D",X"0E",
		X"70",X"F0",X"70",X"38",X"38",X"1C",X"18",X"1C",X"60",X"70",X"88",X"0F",X"0F",X"0B",X"0D",X"0D",
		X"0D",X"0D",X"0D",X"0D",X"07",X"83",X"C0",X"F0",X"83",X"83",X"C0",X"E0",X"F0",X"90",X"90",X"F0",
		X"0F",X"0F",X"0F",X"0E",X"0F",X"0E",X"10",X"F0",X"0E",X"08",X"0B",X"0B",X"0F",X"0E",X"10",X"F0",
		X"18",X"70",X"70",X"F0",X"F0",X"50",X"70",X"F0",X"0D",X"0F",X"00",X"70",X"60",X"C1",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"D0",X"D0",X"D0",X"D0",X"D0",X"60",X"F0",X"E0",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",
		X"F0",X"E0",X"50",X"50",X"D0",X"D0",X"D0",X"60",X"F0",X"C0",X"B0",X"B0",X"E0",X"D0",X"B0",X"80",
		X"F0",X"E0",X"50",X"50",X"D0",X"50",X"50",X"E0",X"F0",X"C0",X"B0",X"F0",X"E0",X"F0",X"B0",X"C0",
		X"F0",X"E0",X"D0",X"D0",X"D0",X"50",X"D0",X"E0",X"F0",X"A0",X"A0",X"A0",X"A0",X"80",X"E0",X"E0",
		X"F0",X"60",X"D0",X"D0",X"50",X"50",X"50",X"E0",X"F0",X"80",X"B0",X"80",X"F0",X"F0",X"B0",X"C0",
		X"F0",X"E0",X"50",X"D0",X"D0",X"50",X"50",X"E0",X"F0",X"C0",X"B0",X"B0",X"80",X"B0",X"B0",X"C0",
		X"F0",X"60",X"50",X"D0",X"D0",X"D0",X"D0",X"E0",X"F0",X"80",X"F0",X"E0",X"E0",X"D0",X"D0",X"D0",
		X"F0",X"E0",X"50",X"50",X"D0",X"50",X"50",X"E0",X"F0",X"C0",X"B0",X"B0",X"C0",X"B0",X"B0",X"C0",
		X"F0",X"E0",X"50",X"50",X"50",X"50",X"50",X"E0",X"F0",X"C0",X"B0",X"B0",X"C0",X"F0",X"B0",X"C0",
		X"00",X"10",X"B0",X"F0",X"B0",X"10",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"30",X"D0",X"D0",X"D0",X"D0",X"D0",X"30",X"F0",X"70",X"A0",X"A0",X"A0",X"A0",X"A0",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"90",X"60",X"60",X"60",X"60",X"60",X"90",
		X"F0",X"90",X"60",X"E0",X"D0",X"B0",X"00",X"F0",X"F0",X"F0",X"F0",X"50",X"B0",X"50",X"F0",X"F0",
		X"F0",X"00",X"D0",X"90",X"E0",X"60",X"90",X"F0",X"F0",X"F0",X"F0",X"50",X"B0",X"50",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"B0",X"F0",X"B0",X"10",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"D0",X"F0",X"D0",X"80",X"80",X"C0",
		X"B0",X"F0",X"90",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"D0",X"F0",X"90",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E1",X"69",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"96",X"87",X"C3",X"C3",X"E1",X"E1",
		X"F0",X"C3",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"B4",X"3C",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"96",X"1E",X"1E",X"3C",X"3C",X"3C",X"78",X"78",X"78",X"2D",X"0F",X"0F",X"0F",X"0F",
		X"8F",X"5F",X"5F",X"9F",X"5F",X"5F",X"9F",X"0F",X"F3",X"E3",X"E3",X"3F",X"A7",X"E3",X"F3",X"E1",
		X"8F",X"8F",X"CF",X"AF",X"9F",X"8F",X"8F",X"0F",X"CF",X"2F",X"2F",X"EF",X"2F",X"2F",X"2F",X"0F",
		X"F8",X"7C",X"78",X"FC",X"7C",X"5E",X"DE",X"1E",X"9F",X"AF",X"AF",X"AF",X"AF",X"AF",X"9F",X"0F",
		X"0F",X"0F",X"0F",X"1E",X"78",X"F0",X"F0",X"F0",X"E1",X"C3",X"C3",X"87",X"87",X"1E",X"78",X"F0",
		X"0F",X"0F",X"0F",X"69",X"78",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"96",X"D2",
		X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"1E",X"1E",X"1E",X"96",X"D2",X"D2",
		X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"CC",X"BB",X"F0",X"E0",X"D1",X"B3",X"B3",X"B3",X"91",X"FF",
		X"F7",X"FF",X"77",X"BB",X"BB",X"BB",X"33",X"CC",X"F0",X"70",X"00",X"77",X"77",X"FF",X"33",X"DD",
		X"F0",X"70",X"B8",X"DC",X"DC",X"DC",X"DC",X"30",X"F8",X"EC",X"DD",X"DD",X"FF",X"FF",X"FF",X"FF",
		X"77",X"77",X"55",X"BB",X"33",X"BB",X"CC",X"66",X"FF",X"FF",X"FF",X"FF",X"44",X"D9",X"D1",X"C0",
		X"33",X"BB",X"BB",X"22",X"AA",X"DD",X"FF",X"FF",X"CC",X"FF",X"FF",X"EE",X"DD",X"DD",X"BB",X"77",
		X"CC",X"EE",X"EE",X"EE",X"FF",X"10",X"F0",X"F0",X"FF",X"FF",X"FF",X"33",X"DD",X"DD",X"EE",X"EE",
		X"DD",X"DD",X"EE",X"FF",X"EE",X"EE",X"00",X"F0",X"B3",X"B3",X"B3",X"77",X"77",X"91",X"E0",X"F0",
		X"EE",X"99",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"77",X"99",X"EE",X"DD",X"DD",X"30",
		X"70",X"B8",X"B8",X"DC",X"DC",X"30",X"F0",X"F0",X"CC",X"FF",X"FF",X"FF",X"FF",X"BB",X"88",X"70",
		X"0F",X"69",X"69",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"87",X"87",X"87",X"87",X"87",X"87",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"00",
		X"00",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"00",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"00",
		X"00",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"00",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"00",
		X"00",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"00",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"EE",X"00",X"CC",X"00",X"00",X"00",X"00",X"08",X"77",X"66",X"77",X"66",X"66",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"CC",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"33",X"00",X"00",X"02",
		X"EE",X"00",X"CC",X"00",X"EE",X"00",X"00",X"02",X"77",X"66",X"77",X"66",X"77",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"08",X"66",X"66",X"66",X"66",X"77",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"66",X"33",X"33",X"FF",X"33",X"33",X"00",X"11",X"33",X"66",X"66",X"66",X"33",X"11",X"00",
		X"FF",X"00",X"00",X"77",X"33",X"33",X"FF",X"00",X"11",X"33",X"66",X"66",X"77",X"66",X"66",X"00",
		X"33",X"33",X"33",X"77",X"EE",X"CC",X"88",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"66",X"66",X"66",X"77",X"33",X"11",X"00",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"66",X"77",X"77",X"77",X"66",X"66",X"66",X"00",
		X"33",X"77",X"FF",X"FF",X"BB",X"33",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"EE",X"33",X"33",X"77",X"CC",X"EE",X"77",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"77",X"66",X"66",X"66",X"77",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"08",X"00",X"33",X"33",X"33",X"00",X"00",X"01",X"03",
		X"03",X"8B",X"CF",X"8B",X"07",X"07",X"0F",X"1E",X"08",X"3B",X"7F",X"3B",X"0C",X"0C",X"0F",X"0F",
		X"08",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"03",X"00",X"EE",X"EE",X"FF",X"EE",X"EE",X"00",
		X"3C",X"3C",X"3C",X"3C",X"2F",X"6F",X"6F",X"66",X"87",X"86",X"86",X"86",X"9F",X"CE",X"CE",X"CC",
		X"0C",X"0C",X"3B",X"7F",X"77",X"66",X"08",X"0C",X"00",X"00",X"00",X"00",X"01",X"00",X"66",X"FF",
		X"11",X"33",X"11",X"00",X"0F",X"0F",X"0F",X"16",X"CD",X"8B",X"8B",X"07",X"0F",X"0F",X"4B",X"E1",
		X"0C",X"0E",X"06",X"88",X"CC",X"EE",X"CC",X"88",X"EE",X"FF",X"45",X"01",X"00",X"11",X"11",X"00",
		X"1E",X"3C",X"3E",X"7E",X"DD",X"DD",X"BB",X"33",X"E1",X"C3",X"86",X"8E",X"BF",X"9D",X"33",X"11",
		X"CC",X"CC",X"8B",X"8F",X"0F",X"0E",X"19",X"77",X"00",X"33",X"77",X"FF",X"77",X"11",X"03",X"77",
		X"00",X"07",X"8F",X"8F",X"07",X"1E",X"3C",X"F8",X"11",X"33",X"3B",X"0C",X"0F",X"87",X"C3",X"87",
		X"77",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",X"33",X"77",X"66",X"00",X"00",X"00",
		X"F0",X"ED",X"8F",X"0F",X"2E",X"33",X"77",X"33",X"87",X"0F",X"0F",X"07",X"88",X"CC",X"88",X"00",
		X"00",X"00",X"EE",X"EE",X"EE",X"44",X"0F",X"0F",X"77",X"77",X"77",X"11",X"07",X"EF",X"FF",X"07",
		X"CC",X"CC",X"CD",X"01",X"0F",X"0F",X"F0",X"F0",X"00",X"00",X"08",X"0C",X"0C",X"0F",X"0F",X"87",
		X"0F",X"44",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"FF",X"EF",X"07",X"11",X"77",X"77",X"77",X"00",
		X"F0",X"0F",X"0F",X"01",X"CD",X"CC",X"CC",X"00",X"0F",X"0F",X"0C",X"0C",X"08",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
