library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity popeye_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of popeye_sp_bits_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FC",X"00",X"FC",X"C0",X"1E",X"E0",X"1E",X"F0",X"0E",X"F8",X"06",X"FC",X"00",X"F8",X"00",X"F0",
		X"0F",X"00",X"07",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"39",X"98",X"CC",X"CE",X"E6",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"F0",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"1E",X"1F",X"3F",X"3F",
		X"1F",X"1F",X"0F",X"43",X"28",X"04",X"10",X"20",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"83",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"FC",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",X"E1",X"C1",X"07",X"0E",X"3F",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"1F",X"1F",X"0F",X"0E",X"A6",X"A6",X"47",X"87",X"8F",X"4F",
		X"5F",X"BF",X"FF",X"FC",X"C0",X"00",X"00",X"00",X"00",X"0F",X"08",X"08",X"10",X"20",X"00",X"00",
		X"0F",X"0F",X"07",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"12",X"07",X"03",X"00",X"00",X"10",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",
		X"00",X"10",X"00",X"00",X"7F",X"FE",X"1C",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"03",X"01",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"7F",X"87",X"E0",X"F8",X"F0",X"00",X"80",X"01",X"0F",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",
		X"40",X"70",X"30",X"10",X"00",X"04",X"00",X"00",X"60",X"70",X"19",X"00",X"00",X"00",X"00",X"00",
		X"70",X"FC",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"08",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"50",X"78",X"70",X"30",X"10",X"01",X"03",X"03",X"05",X"0F",X"0F",X"47",X"63",X"71",X"BC",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"06",X"07",X"03",X"10",X"B8",X"DD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"8F",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"7F",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",
		X"00",X"00",X"00",X"08",X"0C",X"0E",X"02",X"00",X"00",X"06",X"0F",X"2F",X"7F",X"7F",X"7F",X"7F",
		X"BF",X"DF",X"DF",X"7F",X"7F",X"3F",X"1F",X"2F",X"3F",X"1F",X"1F",X"0F",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"02",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7C",X"FF",X"FF",X"7F",X"EF",X"CF",X"9F",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"81",X"C1",X"47",X"E9",X"73",X"A2",
		X"40",X"80",X"80",X"E0",X"80",X"00",X"00",X"60",X"84",X"04",X"18",X"00",X"81",X"4F",X"83",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"02",X"02",X"01",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"00",X"0F",X"03",X"0F",X"03",X"1F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"81",X"81",X"E3",X"25",X"F9",X"31",X"93",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"00",X"2A",X"49",X"84",X"00",
		X"02",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"20",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"87",X"83",X"C1",X"E0",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"F0",X"C1",X"C1",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"C0",X"80",X"00",X"00",
		X"FF",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"07",X"07",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",
		X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"38",X"0E",X"07",X"0F",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"07",X"03",X"00",X"00",X"00",
		X"00",X"0E",X"3C",X"78",X"F0",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"EF",X"EE",X"C7",X"87",X"83",X"01",X"83",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"87",X"C7",X"8F",X"0D",X"09",X"08",X"98",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"04",X"0E",X"1C",X"38",X"31",X"3B",X"1F",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"F8",X"FC",X"FA",X"FA",X"FA",X"F6",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"06",X"00",X"00",X"0C",X"18",X"38",X"30",X"70",X"70",X"60",X"60",X"00",X"00",
		X"00",X"00",X"33",X"33",X"30",X"30",X"30",X"F0",X"F0",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"FE",X"FE",X"06",X"06",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"38",
		X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"00",
		X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"1E",X"1F",X"1F",X"1F",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1E",X"1C",X"1C",X"1E",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"CF",X"CF",X"C3",X"C3",X"C3",X"CF",X"CF",X"C3",X"C3",X"C3",X"CF",X"CF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"8F",X"DF",X"FF",X"FF",X"FF",X"FF",X"F1",X"E1",X"E1",X"C1",X"81",X"81",X"8F",X"FE",
		X"FF",X"FF",X"FF",X"E3",X"D8",X"FC",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"07",X"01",X"00",X"00",
		X"E3",X"C3",X"83",X"07",X"06",X"0E",X"9C",X"F8",X"70",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"1F",X"1F",X"03",X"03",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FC",X"00",X"FC",X"00",
		X"FC",X"00",X"FC",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FE",X"00",X"FC",X"00",X"FC",X"00",
		X"3F",X"3F",X"00",X"3F",X"2E",X"2C",X"2A",X"28",X"3F",X"3F",X"3F",X"60",X"E9",X"F5",X"7E",X"3E",
		X"00",X"41",X"33",X"07",X"03",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"FE",X"FE",X"FF",X"6F",X"31",
		X"00",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",X"78",X"71",X"39",X"0F",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FE",X"FE",X"FF",X"6F",X"30",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"30",X"30",X"38",X"7C",X"1E",X"1E",X"3F",X"1F",X"1F",X"1F",X"0F",X"07",
		X"03",X"03",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"F0",X"F2",X"FD",X"FD",X"FD",X"FB",X"FB",
		X"F7",X"F7",X"6E",X"2C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"C3",X"E7",X"1F",X"03",X"C3",X"7F",X"3F",
		X"3F",X"1D",X"1B",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"F0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",
		X"CF",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"03",X"03",X"0F",X"0F",
		X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"7E",X"7C",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"47",X"C3",X"F9",X"7F",X"3E",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"01",X"01",X"00",X"88",X"C9",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EE",
		X"EC",X"F0",X"F9",X"F7",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7C",X"78",X"20",
		X"30",X"78",X"F8",X"F8",X"F1",X"6D",X"07",X"07",X"1F",X"FE",X"F4",X"C8",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"3F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"0F",X"1F",X"3F",X"7F",X"E7",X"C7",X"07",X"27",X"E6",X"E0",X"F0",X"E3",X"D1",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"C0",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"02",X"00",X"00",
		X"01",X"01",X"00",X"40",X"28",X"04",X"10",X"20",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"01",X"01",X"01",X"03",X"02",X"02",X"02",X"01",X"06",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"0E",X"06",X"66",X"64",X"CC",X"38",X"F0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"F0",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FE",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"F8",X"FC",X"FC",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"FF",X"FB",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"00",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7E",
		X"00",X"00",X"03",X"01",X"20",X"2C",X"2D",X"2D",X"0D",X"2D",X"21",X"2C",X"2D",X"2D",X"0D",X"2D",
		X"21",X"2C",X"2D",X"2D",X"0D",X"05",X"00",X"08",X"08",X"08",X"04",X"04",X"06",X"02",X"01",X"00",
		X"FD",X"FE",X"FF",X"7F",X"1F",X"8F",X"26",X"C6",X"D4",X"E4",X"F0",X"E6",X"A4",X"94",X"10",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"03",X"7B",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"18",X"18",X"1C",X"DF",X"EF",X"3F",X"1B",X"1D",X"9E",X"1F",X"9F",X"FF",X"DF",X"9F",X"DF",X"DF",
		X"00",X"00",X"80",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"83",X"FF",
		X"FF",X"F7",X"3F",X"C0",X"FF",X"3F",X"1F",X"1F",X"9F",X"1F",X"9F",X"FF",X"DF",X"9F",X"DF",X"DF",
		X"BF",X"BF",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"12",X"14",X"04",X"49",X"40",X"A0",X"98",X"81",X"C3",X"FF",X"FF",X"7F",X"7C",X"3E",X"06",
		X"3F",X"3D",X"1E",X"1C",X"1C",X"0E",X"0F",X"17",X"07",X"0B",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"C1",X"E2",X"E0",X"70",X"3A",X"B8",X"B8",X"F4",X"78",X"F0",X"90",X"C8",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C7",X"8F",X"FF",X"FF",X"FF",X"E7",X"C3",X"FF",X"FF",X"FF",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"90",
		X"F8",X"BD",X"BF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"F3",X"F2",X"FD",X"FD",X"FD",X"3B",X"27",X"DF",X"EF",X"DF",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FB",X"FB",X"FB",X"FB",X"7B",X"8F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",
		X"07",X"07",X"07",X"07",X"07",X"4F",X"8F",X"8F",X"CF",X"5F",X"7F",X"7F",X"7F",X"FF",X"DF",X"C7",
		X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"01",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"FF",X"FF",X"FB",X"F7",X"7F",X"EF",X"DF",X"BF",X"7F",X"7F",
		X"78",X"70",X"E0",X"E9",X"FE",X"C6",X"B3",X"B9",X"9C",X"EE",X"F7",X"FB",X"9C",X"0C",X"8F",X"5F",
		X"82",X"A4",X"C8",X"10",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0F",X"0F",X"07",X"03",X"04",X"07",X"03",X"03",X"01",X"01",
		X"01",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"01",X"01",X"01",X"02",X"04",X"08",X"0A",X"0B",
		X"0B",X"09",X"1C",X"1E",X"27",X"03",X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"3F",X"3F",X"FE",X"FF",X"FE",X"4C",X"CC",X"FC",X"FF",X"DE",X"F6",X"F7",
		X"79",X"78",X"BC",X"DC",X"DE",X"EF",X"F7",X"FB",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0B",X"09",X"07",X"03",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",
		X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",
		X"34",X"02",X"09",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"1F",X"1E",X"1E",X"0C",X"00",X"00",X"01",
		X"1F",X"1F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"70",X"38",X"B8",X"B8",X"F4",X"78",X"F0",X"90",X"C8",X"00",
		X"03",X"07",X"16",X"0D",X"0D",X"0D",X"1E",X"0F",X"0E",X"17",X"01",X"02",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"05",X"00",X"D0",X"DE",X"DE",X"DE",X"DE",X"06",X"D8",
		X"DE",X"DE",X"DE",X"DE",X"06",X"D8",X"DE",X"DE",X"DE",X"DE",X"02",X"00",X"F8",X"FF",X"00",X"00",
		X"BE",X"BE",X"1F",X"1F",X"17",X"17",X"37",X"77",X"FF",X"FE",X"F0",X"00",X"02",X"02",X"02",X"02",
		X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",
		X"07",X"05",X"04",X"03",X"00",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"BF",X"DF",X"EF",X"FF",X"FF",X"FF",X"FE",X"FD",X"3E",
		X"4F",X"33",X"82",X"FF",X"3A",X"10",X"00",X"28",X"50",X"F8",X"68",X"00",X"80",X"F8",X"F4",X"08",
		X"F7",X"FF",X"FF",X"FF",X"7F",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"1E",
		X"FF",X"7F",X"FC",X"FC",X"4F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3E",X"7F",X"7F",
		X"BE",X"BE",X"1F",X"1F",X"17",X"17",X"37",X"77",X"FB",X"FB",X"FB",X"73",X"07",X"0F",X"07",X"07",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",
		X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FE",X"FC",X"F8",
		X"F8",X"F0",X"F0",X"B0",X"B1",X"B2",X"B2",X"B4",X"DC",X"D8",X"E8",X"F8",X"F0",X"E0",X"C0",X"88",
		X"08",X"10",X"20",X"00",X"00",X"20",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"FF",X"BF",X"9F",X"8F",X"87",X"C3",X"61",X"F0",X"B0",X"F8",X"FA",X"FB",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"08",X"01",X"02",X"04",X"00",X"01",
		X"01",X"01",X"01",X"07",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FC",X"FC",X"F8",X"F8",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"F0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"FF",X"FF",X"FF",X"FC",X"00",
		X"FE",X"FF",X"FF",X"FF",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",X"1F",X"3F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"9F",X"9F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",
		X"3F",X"1F",X"1F",X"5F",X"8F",X"CF",X"7F",X"6F",X"4F",X"EF",X"EF",X"CF",X"DF",X"BF",X"79",X"FE",
		X"09",X"0A",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"81",X"47",X"7F",X"7F",X"3F",X"3F",X"01",X"0F",X"0F",X"06",X"06",X"02",X"02",
		X"03",X"03",X"03",X"01",X"05",X"03",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"01",X"00",X"04",
		X"03",X"07",X"0B",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FC",X"DE",X"DE",X"BE",X"BE",X"BE",X"7C",X"78",X"79",
		X"F2",X"E0",X"00",X"00",X"7C",X"F6",X"F6",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"F7",X"77",X"0E",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"3F",X"7F",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"FC",X"F7",X"F3",X"F9",X"FE",X"FF",X"7F",X"1F",X"DC",X"BA",X"F7",
		X"F7",X"E1",X"5C",X"5F",X"7F",X"2E",X"04",X"00",X"0C",X"05",X"0B",X"19",X"00",X"03",X"05",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"3F",X"3F",X"36",X"26",
		X"CF",X"07",X"03",X"19",X"3C",X"3F",X"3F",X"3F",X"0E",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"FF",X"FF",X"7F",X"FF",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"1F",X"37",X"33",X"1F",X"01",X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"70",X"30",X"7F",
		X"00",X"00",X"00",X"00",X"0F",X"17",X"1F",X"1F",X"0F",X"0F",X"3F",X"3F",X"3F",X"30",X"30",X"7F",
		X"80",X"E0",X"F0",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",
		X"FC",X"FF",X"FF",X"FB",X"FB",X"FB",X"FD",X"FE",X"FF",X"FF",X"FE",X"FC",X"F0",X"E0",X"60",X"C0",
		X"00",X"00",X"00",X"00",X"03",X"07",X"05",X"0E",X"1F",X"1F",X"3F",X"3F",X"3F",X"30",X"30",X"7F",
		X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7D",X"35",X"1D",X"3F",X"17",X"02",X"00",X"05",X"02",X"07",X"05",X"04",X"02",X"03",X"05",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"01",X"09",X"02",X"04",X"09",X"02",X"00",X"00",X"00",
		X"00",X"00",X"3E",X"37",X"13",X"0F",X"C7",X"E7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"7F",X"FF",X"DE",X"CD",X"7F",X"07",X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"30",X"30",X"7F",
		X"FE",X"7F",X"3F",X"FF",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"BF",X"BF",X"BF",X"DF",X"EF",X"F0",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"60",X"C0",
		X"E0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"70",X"7F",
		X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"F3",X"E4",X"48",X"40",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"3F",X"3F",X"FF",X"FF",X"DF",X"CF",X"C7",X"63",X"E1",X"B0",X"F8",X"3C",X"1E",X"0B",X"2F",X"1F",
		X"7F",X"3E",X"10",X"3F",X"17",X"02",X"00",X"05",X"02",X"07",X"05",X"00",X"03",X"07",X"09",X"02",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"F0",X"F9",X"FB",X"FB",X"FB",X"FF",X"FF",X"7F",X"7E",X"7E",X"7E",X"7C",X"3C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"F0",X"FC",X"FE",X"0E",X"FC",X"F0",X"FE",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"D0",X"F8",
		X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"04",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"0F",X"0F",X"0F",X"3F",X"3F",
		X"1F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"A0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"08",X"0C",X"5C",X"7F",X"3F",X"0F",X"03",X"03",X"01",X"01",X"18",X"18",X"10",X"88",
		X"3C",X"22",X"02",X"22",X"62",X"86",X"10",X"41",X"C0",X"E0",X"C0",X"E0",X"E0",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"2F",X"1E",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",
		X"07",X"0F",X"0C",X"0C",X"0F",X"07",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"78",X"30",X"00",X"00",
		X"03",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"02",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"FF",X"FF",X"FF",X"7F",X"FF",X"BF",X"9B",X"01",
		X"01",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"06",X"03",X"01",
		X"00",X"00",X"00",X"08",X"1C",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",
		X"03",X"07",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"1F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"3F",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"07",X"00",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"1F",X"0F",X"0F",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E3",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",
		X"81",X"E3",X"FB",X"FC",X"FF",X"FF",X"FF",X"FE",X"7E",X"3D",X"3B",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FB",X"F9",X"F1",X"F1",X"E1",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"F3",X"C3",X"83",X"03",X"03",X"03",X"03",X"83",
		X"03",X"03",X"03",X"0F",X"0F",X"03",X"03",X"07",X"0E",X"0C",X"0C",X"0D",X"0D",X"07",X"03",X"01",
		X"01",X"03",X"07",X"0D",X"0D",X"0C",X"0C",X"0D",X"0D",X"07",X"03",X"01",X"01",X"03",X"07",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1E",X"1E",X"0F",X"06",
		X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"7F",X"3F",X"1E",X"4C",X"8C",X"18",X"00",X"21",X"61",X"00",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",X"F0",X"F0",X"F0",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"FB",X"F9",X"F0",X"F0",X"F1",X"FF",X"7F",X"3F",X"7C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"FB",X"F9",X"F0",X"F0",X"F1",X"FF",X"7F",X"3F",X"7C",X"00",
		X"00",X"00",X"80",X"FC",X"FE",X"CE",X"C4",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"07",X"0E",X"0C",X"1C",X"18",X"18",X"18",X"11",X"10",X"D2",X"F4",X"F1",X"6A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"C0",X"E0",X"F8",X"FC",X"FE",X"FF",
		X"FE",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"06",X"1D",X"33",X"77",X"6F",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"77",X"77",X"77",X"3B",
		X"3B",X"1B",X"1D",X"0D",X"06",X"02",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FD",
		X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"9E",X"8E",X"07",X"CB",
		X"0E",X"1F",X"3F",X"3F",X"3F",X"3F",X"15",X"04",X"04",X"44",X"44",X"88",X"30",X"60",X"60",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"1F",X"7F",X"FF",X"FB",X"FB",
		X"F6",X"A6",X"4F",X"0F",X"1F",X"1C",X"18",X"00",X"01",X"00",X"00",X"00",X"01",X"01",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"1F",X"0F",X"06",X"02",X"10",X"08",X"00",X"00",X"00",X"00",
		X"FC",X"BC",X"5E",X"EC",X"FC",X"FC",X"FC",X"BE",X"DE",X"FF",X"FF",X"FF",X"87",X"83",X"CE",X"00",
		X"00",X"33",X"3F",X"7F",X"7D",X"7C",X"3C",X"06",X"86",X"86",X"0E",X"1E",X"FC",X"F8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"07",X"06",X"06",X"06",X"04",X"04",X"35",X"3D",X"3C",X"1A",X"00",X"00",X"00",
		X"7C",X"FE",X"D4",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"02",X"07",X"07",X"01",X"00",X"00",
		X"07",X"0F",X"0F",X"0C",X"00",X"00",X"08",X"3F",X"7F",X"7F",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",
		X"00",X"00",X"01",X"03",X"03",X"07",X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",
		X"FC",X"3C",X"DE",X"EC",X"F4",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"87",X"03",X"01",X"CE",X"00",
		X"00",X"32",X"7F",X"7F",X"7D",X"3C",X"0C",X"8C",X"9C",X"3C",X"78",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1F",X"1E",X"34",X"34",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"8E",X"0C",X"1C",X"18",X"38",X"70",X"F8",X"00",X"00",X"FC",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"3F",X"7B",X"73",X"C1",X"81",X"63",X"03",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FB",X"C3",X"07",X"06",X"0E",X"8E",X"CC",X"9E",X"9E",X"00",X"00",X"E0",X"FC",X"FE",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FE",X"FC",X"FC",X"EC",X"D4",X"BC",X"BC",X"FE",X"FF",X"FF",X"C7",X"83",X"86",X"80",
		X"00",X"32",X"7F",X"7F",X"79",X"3C",X"0C",X"0C",X"9C",X"3C",X"78",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"C6",X"83",X"01",X"87",X"03",
		X"07",X"33",X"7F",X"7F",X"79",X"3C",X"0C",X"8C",X"9C",X"3C",X"78",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"07",X"02",X"12",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"F9",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"87",X"01",X"00",X"00",
		X"00",X"03",X"1F",X"3F",X"7F",X"FF",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"01",X"00",
		X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"00",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3E",X"1C",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"FF",X"FF",X"C0",X"60",X"60",X"10",X"18",X"18",X"04",X"04",X"06",X"01",X"03",X"07",X"03",X"01",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"07",X"07",X"06",X"06",X"07",X"07",
		X"00",X"01",X"03",X"06",X"06",X"07",X"07",X"06",X"06",X"06",X"07",X"07",X"06",X"06",X"07",X"07",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"FE",X"FE",X"06",X"06",X"FE",X"FE",
		X"00",X"01",X"03",X"06",X"06",X"07",X"07",X"06",X"06",X"06",X"FE",X"FE",X"06",X"06",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"01",X"09",X"0D",X"0D",X"09",X"01",X"43",X"67",X"7F",X"3F",X"3F",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"E3",X"FB",X"FC",X"FF",X"FF",X"FF",X"FE",X"7E",X"3D",X"3B",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",
		X"C4",X"C8",X"D0",X"F0",X"F0",X"FA",X"FE",X"FC",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"40",X"F0",X"E0",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",
		X"F8",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"FC",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"79",X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"02",
		X"07",X"0B",X"01",X"01",X"0D",X"0F",X"1F",X"1F",X"1F",X"1F",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"00",X"00",X"03",X"04",X"08",X"08",X"08",X"08",X"1C",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"04",X"1C",X"04",X"0E",X"38",X"10",X"10",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"0E",
		X"1E",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"C7",X"83",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"F8",X"FC",X"3E",X"0F",X"07",
		X"0F",X"1E",X"3E",X"3C",X"7C",X"7E",X"7F",X"7F",X"3F",X"FF",X"3F",X"0F",X"87",X"C3",X"83",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"03",X"52",X"90",X"00",
		X"40",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"04",X"06",X"05",X"10",X"38",X"3C",X"0E",X"03",
		X"2C",X"26",X"1F",X"07",X"03",X"03",X"07",X"0F",X"3E",X"3C",X"98",X"D0",X"C0",X"E0",X"E0",X"F0",
		X"F0",X"FA",X"FB",X"FB",X"FB",X"FA",X"F8",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"87",X"4F",X"1F",
		X"3E",X"3C",X"BE",X"FE",X"7F",X"FF",X"BF",X"BF",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"01",X"43",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"04",
		X"00",X"18",X"38",X"1C",X"1F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"1C",X"20",X"41",X"41",X"40",X"40",X"40",X"E0",X"E1",X"00",
		X"F0",X"F0",X"F9",X"FB",X"FF",X"FF",X"FF",X"FF",X"7C",X"18",X"C0",X"20",X"A0",X"80",X"90",X"08",
		X"00",X"80",X"00",X"00",X"B2",X"7E",X"7C",X"F8",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"7B",X"03",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"05",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"03",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"0E",
		X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"3E",X"7C",X"FC",X"F8",X"FE",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"00",X"00",X"40",X"00",
		X"40",X"00",X"00",X"00",X"34",X"3C",X"7C",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"07",
		X"07",X"03",X"03",X"01",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"08",X"03",X"04",X"08",X"08",X"10",X"10",X"10",X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"7C",X"7E",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",
		X"F8",X"F8",X"F0",X"F8",X"F8",X"FC",X"0C",X"00",X"00",X"20",X"14",X"0C",X"88",X"C0",X"E0",X"FE",
		X"FE",X"FA",X"F2",X"F2",X"E2",X"02",X"02",X"12",X"8E",X"87",X"07",X"47",X"87",X"0F",X"03",X"0B",
		X"13",X"07",X"87",X"C3",X"E3",X"E1",X"E0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"1D",X"3B",X"7B",X"77",X"F7",
		X"EF",X"EF",X"1F",X"F7",X"6F",X"0F",X"1F",X"1E",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"5C",X"6E",X"76",X"36",X"16",X"D6",X"F6",X"F4",X"F2",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"09",X"11",X"11",X"20",X"60",X"30",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"11",X"1E",X"0F",X"03",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3F",X"1F",X"5F",X"3F",X"3F",X"BF",X"5E",X"1E",X"9C",X"9C",X"1C",X"3C",X"38",
		X"38",X"3E",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"01",X"01",X"01",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"DF",X"1F",X"3E",X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",
		X"F8",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"FD",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F1",X"E3",X"E2",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"FC",X"F8",X"78",X"30",X"60",X"00",X"00",X"00",X"80",X"84",X"D2",
		X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"07",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"05",X"06",X"03",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"3E",X"1C",X"1C",X"98",X"08",X"18",X"98",X"98",
		X"FC",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"78",X"30",X"60",X"00",X"00",X"40",X"20",X"A4",
		X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"7F",X"1E",X"1E",X"1E",X"BF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"C7",X"0F",X"0F",X"17",X"02",X"32",X"60",X"50",X"88",X"C0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"1C",X"BE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FD",X"78",X"30",X"60",X"00",X"00",X"00",X"80",X"84",X"D2",
		X"50",X"12",X"20",X"00",X"00",X"20",X"A6",X"7E",X"FF",X"FF",X"FE",X"7C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"05",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"04",X"50",X"28",X"20",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"FC",X"F8",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F9",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F8",X"78",X"30",X"60",X"00",X"00",X"40",X"20",X"A4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"1F",X"3E",X"3C",X"3C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"0C",X"10",X"10",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"16",X"09",
		X"00",X"00",X"00",X"00",X"7C",X"FF",X"FF",X"7F",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"C7",X"0F",X"0F",X"17",X"02",X"32",X"60",X"50",X"88",X"C0",X"F0",X"F8",
		X"F0",X"F8",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F8",X"78",X"30",X"60",X"00",X"00",X"40",X"A4",
		X"22",X"40",X"02",X"00",X"80",X"80",X"20",X"A6",X"7E",X"FF",X"FF",X"FE",X"7C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"16",X"09",
		X"08",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
