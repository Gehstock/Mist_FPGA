library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity skyskip_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of skyskip_sp_bits_2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"C8",X"7C",X"FC",
		X"F6",X"F7",X"EB",X"CD",X"0E",X"96",X"D8",X"B8",X"CC",X"CC",X"8C",X"8E",X"86",X"06",X"06",X"00",
		X"F1",X"FF",X"FF",X"FE",X"FF",X"FF",X"3F",X"C0",X"FF",X"0F",X"00",X"00",X"80",X"F8",X"0F",X"00",
		X"00",X"00",X"01",X"03",X"C7",X"EE",X"FC",X"F8",X"F8",X"EC",X"CC",X"04",X"C6",X"66",X"22",X"33",
		X"93",X"11",X"C1",X"F1",X"F9",X"FC",X"FC",X"37",X"CF",X"F7",X"F7",X"FF",X"C1",X"FE",X"FF",X"97",
		X"8B",X"CD",X"C7",X"8F",X"9F",X"FE",X"FC",X"FE",X"FF",X"F0",X"88",X"1C",X"0D",X"06",X"8C",X"78",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"03",X"FF",X"FC",X"00",X"00",X"00",X"01",X"07",
		X"76",X"77",X"BB",X"FD",X"FE",X"FF",X"7F",X"BE",X"BE",X"1C",X"00",X"00",X"C0",X"FC",X"FF",X"00",
		X"FF",X"FC",X"00",X"17",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",X"9F",X"FF",X"F0",X"E4",X"E6",X"E3",X"61",X"30",X"1C",X"07",
		X"F0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"F0",X"FC",X"FE",X"FF",X"CF",X"BF",X"BF",X"7F",X"7F",X"FF",X"FE",X"EC",X"C2",X"C2",X"C4",X"E4",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"07",X"07",X"0E",X"0C",X"0C",X"08",X"08",X"18",X"3C",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"7E",X"FD",X"EC",X"C8",X"8C",X"08",X"00",X"80",X"80",X"80",X"C0",X"C0",
		X"FC",X"FC",X"7D",X"FF",X"FE",X"FC",X"EE",X"47",X"82",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"33",
		X"23",X"23",X"37",X"1F",X"0F",X"0E",X"06",X"00",X"00",X"00",X"00",X"1C",X"FC",X"E0",X"00",X"00",
		X"23",X"23",X"37",X"1F",X"0F",X"0E",X"06",X"00",X"E0",X"E0",X"00",X"00",X"02",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"4C",X"84",X"08",X"CC",X"00",X"00",X"40",X"00",X"00",X"40",
		X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"03",X"01",X"03",X"07",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"21",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"70",X"38",X"18",X"00",X"00",X"00",
		X"FF",X"FF",X"3C",X"0E",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C0",X"E0",X"70",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"1F",X"0C",X"00",X"00",X"00",X"00",X"00",X"01",X"F9",X"F8",X"00",X"04",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"F4",X"DC",X"CC",X"C0",X"C0",X"C0",X"C0",X"E0",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"3C",X"1C",X"0C",X"0C",X"0C",X"6C",X"7C",X"F8",X"F0",X"C0",
		X"FF",X"FE",X"78",X"00",X"00",X"01",X"3E",X"00",X"7C",X"FE",X"FF",X"FF",X"FF",X"FF",X"9F",X"EF",
		X"EF",X"F6",X"F7",X"FB",X"FF",X"F7",X"EF",X"1F",X"F9",X"69",X"E9",X"A9",X"A9",X"AF",X"BF",X"FF",
		X"EF",X"F6",X"F7",X"F7",X"F7",X"F7",X"EF",X"1F",X"FF",X"7F",X"3F",X"3F",X"3F",X"3F",X"BF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"EF",X"1F",X"FF",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"CF",X"46",X"46",X"47",X"07",X"83",X"E3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"A7",X"46",X"46",X"47",X"47",X"27",X"83",X"E3",
		X"F1",X"F1",X"78",X"78",X"F8",X"B8",X"10",X"00",X"80",X"C0",X"80",X"80",X"C0",X"E0",X"30",X"98",
		X"F1",X"F1",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"C0",X"E0",X"30",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",
		X"2E",X"7E",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"0C",X"0C",X"1C",X"3C",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"3E",X"3C",X"1C",X"18",
		X"00",X"18",X"0C",X"04",X"06",X"02",X"82",X"82",X"82",X"C2",X"C2",X"C2",X"C4",X"C4",X"88",X"88",
		X"98",X"10",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"BF",X"3F",X"FF",X"FE",X"FE",X"7E",X"7F",X"FF",X"FE",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FE",X"FE",
		X"FF",X"7F",X"7E",X"3E",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"DE",X"FE",X"FE",X"FC",X"B8",X"48",X"40",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"8F",X"0F",X"07",X"07",X"07",X"07",X"0F",X"9F",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"3F",X"0F",X"0F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"80",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"81",X"80",X"00",X"80",
		X"80",X"80",X"80",X"90",X"91",X"91",X"81",X"00",X"01",X"01",X"01",X"07",X"0F",X"1F",X"1F",X"3F",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"81",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",X"FB",X"FB",X"F3",X"F3",X"F3",X"F3",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"FB",X"F9",X"FC",X"7E",X"6E",X"6C",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"1F",X"7F",X"FE",X"FC",X"F0",X"C0",X"01",X"02",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",
		X"00",X"00",X"00",X"80",X"C0",X"E3",X"FF",X"7F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",
		X"E1",X"C0",X"C0",X"81",X"03",X"0F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"E1",X"C0",X"C0",X"81",X"03",X"0F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",
		X"FF",X"7F",X"7F",X"3F",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"3F",X"3F",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"7C",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"8F",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"3F",X"3F",X"7F",X"7F",X"FC",X"FA",X"F4",X"F4",X"F4",X"F2",X"78",X"7C",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FA",X"F4",X"F4",X"F4",X"72",X"78",X"FC",
		X"FC",X"F7",X"F7",X"F7",X"F7",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"40",X"20",X"20",X"20",X"20",X"10",X"18",X"08",X"08",X"08",X"18",X"10",
		X"E0",X"F0",X"18",X"04",X"02",X"22",X"C1",X"01",X"01",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"60",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"F8",X"FC",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",
		X"1E",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"7C",X"7C",X"7F",X"7F",X"7E",X"7E",X"7F",X"7F",X"7C",X"7C",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E0",X"C0",X"C0",X"C0",X"CE",X"CE",X"CE",X"CE",X"CE",X"CE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E7",X"E7",X"E7",X"07",X"07",X"E7",X"E7",X"C7",X"07",X"07",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3C",X"38",X"30",X"20",X"00",X"00",X"00",X"00",
		X"00",X"18",X"D4",X"F8",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"FA",X"FF",X"FE",X"FC",
		X"F8",X"FC",X"FC",X"C0",X"5C",X"28",X"E0",X"E2",X"E2",X"E2",X"42",X"46",X"44",X"6C",X"38",X"10",
		X"00",X"3F",X"FF",X"E6",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"FA",X"FB",X"FF",X"FE",X"FC",
		X"F8",X"FC",X"FC",X"C0",X"5C",X"28",X"E0",X"E0",X"E0",X"E0",X"60",X"42",X"43",X"47",X"7E",X"38",
		X"00",X"0F",X"1F",X"FF",X"0F",X"05",X"F5",X"E2",X"5A",X"FE",X"FE",X"FE",X"5A",X"E4",X"F4",X"F4",
		X"E4",X"04",X"00",X"80",X"FE",X"FC",X"FE",X"F6",X"F6",X"E6",X"E6",X"CF",X"27",X"AA",X"A2",X"C0",
		X"3F",X"3E",X"38",X"F8",X"0C",X"04",X"F4",X"E2",X"5A",X"FD",X"FD",X"FF",X"5B",X"E2",X"F0",X"F0",
		X"E0",X"00",X"00",X"80",X"FE",X"FC",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"A0",X"A0",X"20",X"C0",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FF",X"7D",X"3F",X"7B",X"3F",X"BF",X"E6",X"C6",X"C6",X"C4",X"E8",X"A0",X"80",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"7C",X"3C",X"78",X"38",X"F0",X"C0",X"C0",X"C0",X"E0",X"A0",X"80",
		X"C0",X"80",X"00",X"00",X"FF",X"FC",X"DC",X"8C",X"8C",X"AC",X"AC",X"DC",X"FC",X"FC",X"F8",X"F0",
		X"7E",X"7E",X"7C",X"30",X"00",X"00",X"E0",X"C0",X"86",X"F3",X"FB",X"FB",X"FB",X"FB",X"F3",X"E2",
		X"C0",X"FF",X"FC",X"DC",X"8C",X"8C",X"AC",X"AC",X"DC",X"FC",X"FC",X"F8",X"F0",X"00",X"00",X"00",
		X"38",X"7C",X"7C",X"78",X"30",X"00",X"00",X"E0",X"C0",X"80",X"F0",X"F8",X"FA",X"FA",X"FB",X"F3",
		X"E3",X"C7",X"83",X"00",X"FF",X"FC",X"DC",X"8C",X"8C",X"AC",X"AC",X"DC",X"FC",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"07",X"3F",X"37",X"33",X"31",X"71",X"E0",X"91",X"D1",X"FB",X"FB",X"7F",X"1F",
		X"00",X"00",X"00",X"07",X"3F",X"77",X"33",X"31",X"71",X"60",X"11",X"91",X"FB",X"FB",X"FF",X"7F",
		X"3F",X"79",X"F7",X"EF",X"7B",X"75",X"3B",X"3F",X"3F",X"1F",X"1B",X"1B",X"1F",X"0F",X"06",X"00",
		X"00",X"00",X"0C",X"1F",X"1B",X"3B",X"71",X"71",X"31",X"80",X"91",X"91",X"FB",X"FB",X"FF",X"3F",
		X"3F",X"79",X"F7",X"EF",X"7B",X"75",X"3B",X"3F",X"3B",X"1B",X"D1",X"F9",X"FB",X"7F",X"3E",X"1C",
		X"38",X"FE",X"FF",X"C7",X"EE",X"7C",X"FF",X"FF",X"FF",X"38",X"07",X"06",X"0E",X"1F",X"7F",X"7F",
		X"38",X"F2",X"F3",X"E3",X"E3",X"E3",X"E7",X"FF",X"FF",X"F8",X"3F",X"06",X"0E",X"1F",X"7F",X"7F",
		X"BE",X"9C",X"99",X"91",X"10",X"30",X"36",X"72",X"15",X"0F",X"0F",X"0F",X"0B",X"01",X"00",X"00",
		X"00",X"00",X"7B",X"8F",X"DE",X"FC",X"FF",X"FF",X"FF",X"30",X"17",X"06",X"8E",X"CF",X"FF",X"FF",
		X"8F",X"FF",X"FF",X"C7",X"EE",X"7C",X"FF",X"FF",X"FF",X"F8",X"C7",X"E6",X"6E",X"6F",X"7F",X"7F",
		X"FE",X"FC",X"F9",X"F0",X"F0",X"F2",X"76",X"32",X"15",X"0F",X"0F",X"0F",X"0B",X"01",X"00",X"00",
		X"FC",X"3C",X"FC",X"FE",X"7E",X"BF",X"BF",X"BF",X"7F",X"DF",X"88",X"1E",X"3C",X"3D",X"7F",X"7F",
		X"00",X"00",X"60",X"E0",X"E0",X"F8",X"FC",X"FF",X"FF",X"7F",X"00",X"3E",X"BC",X"F9",X"F3",X"F7",
		X"90",X"F0",X"F0",X"F0",X"F8",X"FE",X"FF",X"FF",X"7F",X"3F",X"00",X"3E",X"BC",X"F9",X"F3",X"77",
		X"AB",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"FF",X"00",X"29",X"21",X"00",X"00",X"C1",X"C1",X"00",
		X"82",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"82",X"C3",X"E6",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"D8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"1E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"FC",X"1E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"1E",X"0F",
		X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"83",X"83",X"C1",X"C0",X"C0",X"E0",X"E0",X"E0",X"60",X"60",X"60",X"30",X"30",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"F0",X"E0",X"E0",X"F0",X"F8",X"FF",X"FF",X"FF",X"7F",X"0F",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"E0",X"E0",X"E0",X"70",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"48",X"7C",X"7F",X"3F",X"1F",X"1F",X"0F",X"06",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FC",X"1E",X"02",X"02",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"10",X"18",X"0F",X"07",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"3F",X"77",X"33",X"31",X"71",X"60",X"11",X"91",X"FB",X"FB",X"FF",X"7F",
		X"00",X"00",X"0C",X"1F",X"1B",X"3B",X"71",X"F1",X"31",X"80",X"D1",X"F1",X"FB",X"FB",X"7F",X"1F",
		X"3F",X"79",X"F7",X"EF",X"7B",X"75",X"3B",X"3F",X"3F",X"1F",X"1B",X"1B",X"1F",X"0F",X"06",X"00",
		X"3F",X"79",X"F7",X"EF",X"7B",X"75",X"3B",X"3F",X"3B",X"1B",X"D1",X"F1",X"FB",X"7F",X"3E",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CE",X"7F",X"38",X"07",X"06",X"0E",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"44",X"EF",X"FF",X"FF",X"FF",X"F8",X"C7",X"E6",X"6E",X"6F",X"7F",X"7F",
		X"FE",X"FC",X"F9",X"F0",X"F0",X"F2",X"76",X"32",X"15",X"0F",X"0F",X"0F",X"0B",X"01",X"00",X"FF",
		X"FF",X"F0",X"F0",X"F0",X"F8",X"FE",X"FF",X"FF",X"7F",X"3F",X"00",X"3E",X"BC",X"F9",X"F3",X"77",
		X"FF",X"00",X"60",X"E0",X"E0",X"F8",X"FC",X"FF",X"FF",X"7F",X"00",X"3E",X"BC",X"F9",X"F3",X"F7",
		X"AB",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"FF",X"00",X"28",X"21",X"00",X"00",X"00",X"00",X"FF",
		X"AB",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"FF",X"00",X"28",X"21",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"60",X"00",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"F0",X"F8",X"FC",X"FA",X"F6",X"EF",X"EF",X"EF",X"EF",X"F6",X"FA",X"FC",X"F8",X"F0",X"C0",
		X"C0",X"F0",X"E8",X"DC",X"3E",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"3E",X"DC",X"E8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"40",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"40",
		X"01",X"EB",X"C3",X"00",X"00",X"00",X"0F",X"01",X"07",X"1F",X"7E",X"F8",X"E0",X"80",X"00",X"00",
		X"11",X"1B",X"0B",X"00",X"00",X"00",X"0F",X"01",X"07",X"1F",X"7E",X"F8",X"E0",X"80",X"00",X"00",
		X"7B",X"7B",X"FB",X"F9",X"0E",X"0F",X"07",X"07",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"80",X"80",X"80",X"FF",X"FF",X"FF",X"80",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"3C",X"3D",X"3B",X"3B",X"3D",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"DF",X"EF",X"F7",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"30",X"70",X"28",X"00",X"82",X"C3",X"61",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"30",X"70",X"20",X"04",X"81",X"C0",X"60",X"A0",
		X"00",X"00",X"00",X"00",X"08",X"1C",X"36",X"7B",X"6D",X"76",X"78",X"3F",X"1F",X"3C",X"7C",X"FE",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F7",X"E9",X"C0",X"C8",X"D9",X"FF",X"EF",X"C7",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"0D",X"1D",X"1D",X"3C",X"FE",X"FE",
		X"00",X"30",X"30",X"10",X"10",X"10",X"08",X"18",X"08",X"88",X"80",X"8C",X"CC",X"CC",X"C8",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"10",X"88",X"80",X"8C",X"CC",X"CC",X"C8",X"C4",
		X"C4",X"E2",X"E2",X"E2",X"C1",X"01",X"03",X"03",X"80",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"C2",X"E1",X"E2",X"E3",X"C0",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"F0",X"CF",X"DE",X"C0",X"D0",X"D0",X"F8",X"EF",X"BF",X"9F",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"01",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"07",X"07",X"0C",X"09",X"FB",X"FB",X"FB",X"FB",
		X"F8",X"FF",X"0B",X"FB",X"93",X"83",X"83",X"9B",X"FF",X"0F",X"00",X"00",X"00",X"C3",X"EB",X"01",
		X"F8",X"FF",X"0B",X"FB",X"93",X"83",X"83",X"9B",X"FF",X"0F",X"00",X"00",X"00",X"0B",X"1D",X"11",
		X"01",X"03",X"03",X"03",X"01",X"01",X"03",X"03",X"E4",X"FA",X"F7",X"EF",X"EE",X"F2",X"DD",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"3F",X"7E",X"78",X"FD",X"FD",X"7B",X"3B",X"1F",X"06",X"00",X"C0",X"E0",X"50",X"06",X"03",X"01",
		X"3F",X"7E",X"78",X"FD",X"FD",X"7B",X"3B",X"1F",X"06",X"00",X"C0",X"E0",X"50",X"04",X"08",X"00",
		X"80",X"00",X"00",X"80",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"1F",X"3F",X"3F",X"BD",X"DE",X"FF",X"7F",X"EF",X"CF",X"87",
		X"80",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"8C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"FF",X"7F",X"3F",X"1F",X"0F",X"87",X"07",X"80",X"80",X"00",X"20",X"30",X"18",X"00",X"00",
		X"87",X"FF",X"7F",X"3F",X"1F",X"0F",X"80",X"07",X"80",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"FB",
		X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"FB",
		X"00",X"60",X"60",X"C0",X"80",X"F8",X"FC",X"FE",X"FE",X"FC",X"EC",X"EC",X"EE",X"F6",X"F6",X"F7",
		X"F7",X"7B",X"3A",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"F6",X"F6",X"F4",X"F0",X"66",X"76",X"76",X"76",X"37",X"37",X"3F",X"3F",X"1F",X"1F",X"0E",
		X"FA",X"F6",X"F6",X"F4",X"F0",X"66",X"76",X"76",X"76",X"37",X"37",X"3F",X"3F",X"1F",X"1F",X"0E",
		X"30",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",
		X"30",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"30",X"E0",X"F0",X"FC",X"FF",
		X"FF",X"FE",X"F6",X"F6",X"F6",X"F6",X"F6",X"76",X"76",X"36",X"3E",X"1C",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"DE",X"DE",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"DE",X"DE",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
