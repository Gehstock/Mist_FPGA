library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_sp_bits is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"22",
		X"00",X"66",X"77",X"00",X"00",X"66",X"77",X"00",X"00",X"66",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"66",X"00",
		X"00",X"02",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"27",X"00",
		X"72",X"66",X"22",X"77",X"72",X"66",X"22",X"67",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"26",
		X"20",X"66",X"77",X"66",X"20",X"66",X"77",X"66",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"66",X"22",X"66",X"00",X"66",X"22",X"26",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"20",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"27",X"00",
		X"72",X"66",X"22",X"77",X"72",X"66",X"22",X"67",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"26",
		X"20",X"66",X"77",X"66",X"20",X"66",X"77",X"66",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"66",X"22",X"66",X"00",X"66",X"22",X"26",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"CC",X"00",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"77",
		X"CC",X"77",X"22",X"22",X"CC",X"77",X"22",X"72",X"CC",X"77",X"22",X"22",X"CC",X"77",X"22",X"77",
		X"67",X"77",X"22",X"77",X"67",X"77",X"22",X"77",X"CC",X"22",X"27",X"77",X"CC",X"22",X"77",X"77",
		X"00",X"22",X"27",X"22",X"00",X"22",X"27",X"22",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"77",
		X"00",X"77",X"22",X"CC",X"00",X"77",X"22",X"00",X"CC",X"77",X"22",X"77",X"CC",X"77",X"22",X"77",
		X"CC",X"77",X"77",X"22",X"CC",X"77",X"77",X"22",X"00",X"22",X"CC",X"77",X"00",X"22",X"CC",X"77",
		X"00",X"77",X"CC",X"CC",X"00",X"77",X"CC",X"CC",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"01",X"00",X"22",X"01",X"11",X"00",X"C1",X"11",
		X"1D",X"10",X"1A",X"13",X"1D",X"10",X"00",X"33",X"1D",X"10",X"00",X"33",X"1D",X"11",X"A1",X"33",
		X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"AD",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"DD",X"33",
		X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"D2",X"33",
		X"1D",X"1D",X"22",X"33",X"1D",X"1D",X"2D",X"33",X"1D",X"1D",X"3D",X"23",X"1D",X"1D",X"33",X"23",
		X"1D",X"1D",X"33",X"23",X"1D",X"1D",X"3D",X"23",X"1D",X"1D",X"2D",X"33",X"1D",X"1D",X"22",X"33",
		X"1D",X"1D",X"D2",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"11",X"11",X"33",X"1D",X"10",X"00",X"13",
		X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"00",X"DD",X"DD",X"DD",X"01",X"33",X"33",X"33",X"11",X"11",X"11",X"11",
		X"11",X"22",X"A2",X"2A",X"01",X"11",X"11",X"11",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"11",X"12",X"11",X"00",X"DD",X"22",X"DD",X"00",X"DD",X"2D",X"2D",X"00",X"DD",X"3D",X"2D",
		X"00",X"DD",X"33",X"2D",X"00",X"DD",X"3D",X"2D",X"00",X"DD",X"2D",X"2D",X"02",X"DD",X"22",X"DD",
		X"22",X"12",X"12",X"AD",X"A3",X"33",X"33",X"1A",X"A3",X"33",X"33",X"32",X"22",X"12",X"12",X"1D",
		X"02",X"DD",X"DD",X"AD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"11",X"11",X"11",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"01",X"11",X"11",X"11",X"11",X"22",X"A2",X"2A",
		X"11",X"11",X"11",X"11",X"01",X"33",X"33",X"33",X"00",X"DD",X"DD",X"DD",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"05",X"55",X"00",X"00",X"55",X"C2",X"00",X"00",X"5C",
		X"CC",X"50",X"00",X"5C",X"C2",X"50",X"00",X"C6",X"55",X"50",X"02",X"CA",X"55",X"50",X"5C",X"C6",
		X"C2",X"50",X"7C",X"C6",X"CC",X"52",X"C7",X"C6",X"C2",X"52",X"7C",X"C6",X"55",X"52",X"7C",X"CA",
		X"55",X"52",X"C7",X"C6",X"C2",X"52",X"77",X"C6",X"CC",X"CC",X"55",X"C6",X"C2",X"C7",X"55",X"C6",
		X"55",X"C7",X"55",X"CA",X"55",X"C7",X"55",X"C6",X"C2",X"C7",X"55",X"C6",X"CC",X"C7",X"55",X"C6",
		X"C2",X"C7",X"55",X"C6",X"55",X"C7",X"55",X"CA",X"55",X"C7",X"55",X"C6",X"C2",X"CC",X"55",X"C6",
		X"CC",X"57",X"77",X"C6",X"C2",X"55",X"CC",X"C6",X"55",X"50",X"22",X"CA",X"55",X"50",X"22",X"CC",
		X"05",X"00",X"77",X"5C",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"52",X"25",X"2C",X"00",X"52",X"25",X"2C",X"05",X"CC",X"55",X"CC",X"55",X"55",X"5A",X"55",
		X"56",X"CC",X"CC",X"C6",X"5C",X"CC",X"CC",X"CC",X"55",X"66",X"6A",X"66",X"00",X"CC",X"CC",X"CC",
		X"00",X"55",X"CC",X"C5",X"00",X"00",X"77",X"C7",X"00",X"00",X"77",X"CC",X"00",X"05",X"75",X"77",
		X"00",X"05",X"55",X"77",X"00",X"55",X"55",X"57",X"00",X"CC",X"55",X"57",X"00",X"57",X"55",X"57",
		X"00",X"57",X"55",X"57",X"00",X"CC",X"55",X"57",X"00",X"55",X"55",X"57",X"00",X"05",X"55",X"77",
		X"00",X"05",X"75",X"77",X"00",X"00",X"77",X"CC",X"00",X"00",X"77",X"C7",X"00",X"55",X"CC",X"C5",
		X"00",X"CC",X"CC",X"CC",X"55",X"66",X"6A",X"66",X"5C",X"CC",X"CC",X"CC",X"56",X"CC",X"CC",X"C6",
		X"55",X"55",X"5A",X"55",X"05",X"CC",X"55",X"CC",X"00",X"52",X"25",X"2C",X"00",X"5C",X"C5",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"33",X"00",
		X"00",X"0F",X"93",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"55",X"99",X"00",X"55",X"55",X"99",
		X"00",X"0F",X"AA",X"90",X"00",X"FF",X"AA",X"00",X"00",X"F3",X"AA",X"F0",X"00",X"33",X"A5",X"3F",
		X"00",X"55",X"F5",X"55",X"00",X"39",X"99",X"3F",X"00",X"F3",X"9A",X"F0",X"00",X"FF",X"9A",X"00",
		X"00",X"0F",X"9A",X"50",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"00",
		X"00",X"0F",X"93",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"3F",X"00",X"00",X"03",X"F0",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"05",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"22",X"00",X"00",X"BE",X"22",X"00",X"00",X"BB",X"22",
		X"22",X"22",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"02",X"00",X"22",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"7E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"23",X"00",X"00",X"02",X"22",X"00",X"00",X"72",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"33",X"00",X"00",X"A6",X"3B",
		X"00",X"00",X"A6",X"AA",X"00",X"00",X"A7",X"3A",X"00",X"00",X"AA",X"3A",X"00",X"00",X"0A",X"AA",
		X"00",X"00",X"00",X"3B",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"72",X"02",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"D0",X"20",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"DD",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"DD",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C7",
		X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"0F",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"0F",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"07",X"FF",X"FF",X"00",X"00",X"FF",X"CC",
		X"00",X"00",X"FF",X"77",X"00",X"00",X"FF",X"CC",X"00",X"00",X"0F",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"2C",X"00",X"00",X"FF",X"2C",X"77",X"00",X"FF",
		X"00",X"77",X"FF",X"CC",X"00",X"07",X"FF",X"77",X"00",X"00",X"FF",X"CC",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F7",
		X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"7C",X"00",X"00",X"FF",X"C7",X"02",X"77",X"FF",X"C7",
		X"02",X"77",X"FF",X"C7",X"00",X"00",X"FF",X"C7",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"CF",
		X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"33",X"00",X"EE",X"33",X"99",X"00",X"EE",X"EE",X"99",
		X"33",X"E9",X"EE",X"99",X"3E",X"99",X"EE",X"EE",X"9E",X"99",X"9E",X"99",X"99",X"9E",X"9E",X"E9",
		X"99",X"9E",X"EE",X"33",X"9E",X"E9",X"EE",X"EE",X"33",X"EE",X"E3",X"99",X"00",X"EE",X"30",X"99",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"EE",X"00",X"00",X"99",X"99",X"30",X"00",X"9E",X"93",X"30",X"00",
		X"EE",X"3E",X"30",X"00",X"33",X"E9",X"30",X"00",X"EE",X"33",X"30",X"00",X"33",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"33",X"00",X"EE",X"33",X"99",X"00",X"EE",X"EE",X"99",
		X"33",X"E9",X"EE",X"EE",X"3E",X"99",X"EE",X"99",X"9E",X"99",X"9E",X"99",X"99",X"9E",X"9E",X"E9",
		X"99",X"9E",X"EE",X"33",X"3E",X"E9",X"EE",X"99",X"03",X"EE",X"E3",X"EE",X"00",X"EE",X"30",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"33",X"00",X"00",X"33",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"99",
		X"00",X"44",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"44",X"00",
		X"00",X"99",X"94",X"00",X"00",X"9E",X"94",X"00",X"00",X"9E",X"44",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"CC",X"CC",X"EE",
		X"0E",X"EE",X"EE",X"CC",X"EE",X"CC",X"CC",X"CC",X"EE",X"CC",X"CC",X"CF",X"EE",X"CC",X"CC",X"CF",
		X"EE",X"CC",X"CC",X"CF",X"EE",X"CC",X"CC",X"CF",X"1E",X"CC",X"CC",X"CC",X"0E",X"EE",X"EE",X"CC",
		X"00",X"CC",X"CC",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"0F",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"CC",X"CC",X"77",
		X"07",X"77",X"77",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CF",X"77",X"CC",X"CC",X"CF",
		X"77",X"CC",X"CC",X"CF",X"77",X"CC",X"CC",X"CF",X"77",X"CC",X"CC",X"CC",X"07",X"77",X"77",X"CC",
		X"00",X"CC",X"CC",X"77",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"0F",X"CC",X"00",
		X"00",X"0F",X"CC",X"00",X"00",X"04",X"CC",X"00",X"00",X"04",X"CC",X"00",X"00",X"07",X"CC",X"00",
		X"00",X"07",X"CC",X"00",X"00",X"07",X"CC",X"00",X"00",X"07",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"10",
		X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"03",X"13",X"13",X"13",X"01",X"31",X"31",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"D0",X"FD",X"FD",X"FD",X"F0",X"0F",X"DF",X"DF",X"DF",X"0D",X"FD",X"FD",X"FD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"10",
		X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",
		X"60",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"55",X"55",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"40",
		X"60",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FA",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"50",X"00",X"00",X"0A",X"AF",X"7F",X"00",X"A0",X"A0",X"00",
		X"0A",X"00",X"07",X"0F",X"A5",X"00",X"70",X"00",X"50",X"00",X"00",X"0F",X"00",X"00",X"50",X"F0",
		X"90",X"0E",X"0E",X"0E",X"0E",X"90",X"A0",X"E0",X"20",X"09",X"0A",X"0B",X"0E",X"E0",X"E0",X"A0",
		X"00",X"0E",X"4B",X"09",X"00",X"E0",X"A0",X"2A",X"00",X"0A",X"0B",X"00",X"00",X"00",X"EA",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"02",X"00",X"00",
		X"2E",X"A0",X"00",X"00",X"90",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"7B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"20",X"00",X"00",
		X"02",X"0B",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"79",X"00",X"00",
		X"00",X"79",X"07",X"00",X"00",X"79",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"97",X"00",X"00",
		X"00",X"97",X"00",X"07",X"00",X"97",X"00",X"00",X"00",X"47",X"40",X"00",X"70",X"44",X"00",X"00",
		X"03",X"44",X"00",X"00",X"70",X"47",X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"97",X"00",X"07",
		X"00",X"97",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"07",X"00",
		X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"55",X"00",X"55",
		X"00",X"C5",X"00",X"CC",X"00",X"50",X"00",X"CC",X"00",X"00",X"00",X"5C",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"55",X"05",X"00",X"00",X"CC",X"00",
		X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"00",X"05",X"05",X"05",
		X"00",X"5C",X"00",X"05",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"75",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"55",X"55",X"55",X"00",X"CC",X"CC",X"C5",
		X"00",X"CC",X"CC",X"C5",X"00",X"CC",X"CC",X"C5",X"00",X"CC",X"55",X"55",X"00",X"CC",X"00",X"05",
		X"00",X"C5",X"00",X"55",X"00",X"50",X"00",X"C5",X"00",X"00",X"00",X"C5",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"C5",X"00",X"50",X"00",X"C5",X"00",X"C5",X"00",X"55",
		X"00",X"CC",X"00",X"05",X"00",X"CC",X"55",X"55",X"00",X"CC",X"CC",X"C5",X"00",X"CC",X"CC",X"C5",
		X"00",X"CC",X"CC",X"C5",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"77",X"22",X"00",X"00",X"77",X"22",X"00",X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"77",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"77",X"00",X"66",X"00",X"77",X"00",X"66",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"77",X"00",
		X"22",X"66",X"22",X"77",X"22",X"66",X"22",X"77",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"77",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"77",X"00",X"66",X"00",X"77",X"00",X"66",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"77",X"00",
		X"22",X"66",X"22",X"77",X"22",X"66",X"22",X"77",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"CC",X"77",X"00",X"00",X"CC",X"77",X"CC",X"00",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"77",
		X"CC",X"22",X"77",X"77",X"CC",X"22",X"77",X"77",X"77",X"22",X"22",X"77",X"77",X"22",X"22",X"27",
		X"72",X"22",X"22",X"0C",X"22",X"22",X"22",X"CC",X"77",X"22",X"72",X"77",X"77",X"22",X"77",X"77",
		X"CC",X"22",X"27",X"22",X"CC",X"22",X"77",X"27",X"CC",X"22",X"27",X"77",X"CC",X"22",X"22",X"77",
		X"77",X"77",X"22",X"CC",X"77",X"77",X"22",X"00",X"77",X"22",X"22",X"77",X"77",X"22",X"22",X"77",
		X"CC",X"22",X"77",X"22",X"CC",X"22",X"77",X"22",X"00",X"27",X"77",X"77",X"00",X"77",X"77",X"77",
		X"00",X"CC",X"77",X"CC",X"00",X"CC",X"77",X"CC",X"CC",X"00",X"55",X"00",X"CC",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",X"00",X"0C",X"BB",X"00",X"00",X"0C",X"BB",X"00",
		X"00",X"0C",X"BB",X"00",X"00",X"0C",X"BB",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",
		X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"01",X"11",X"02",X"00",X"11",X"11",X"22",X"00",X"12",X"31",X"1C",X"00",X"1A",
		X"31",X"A1",X"00",X"12",X"31",X"00",X"00",X"12",X"31",X"00",X"00",X"12",X"31",X"11",X"11",X"1A",
		X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"1A",
		X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"22",X"12",
		X"31",X"DD",X"33",X"1A",X"31",X"DD",X"D3",X"12",X"31",X"DD",X"D3",X"12",X"31",X"DD",X"33",X"12",
		X"31",X"DD",X"33",X"12",X"31",X"DD",X"D3",X"1A",X"31",X"DD",X"D3",X"12",X"31",X"DD",X"33",X"12",
		X"31",X"DA",X"22",X"12",X"31",X"DD",X"DD",X"1A",X"31",X"11",X"11",X"12",X"31",X"00",X"00",X"12",
		X"31",X"00",X"00",X"1A",X"11",X"00",X"00",X"12",X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"01",
		X"01",X"11",X"11",X"11",X"11",X"DD",X"DD",X"DD",X"13",X"33",X"33",X"33",X"11",X"11",X"11",X"11",
		X"2A",X"2A",X"22",X"22",X"11",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"01",X"33",X"22",X"31",
		X"00",X"11",X"23",X"11",X"00",X"DD",X"33",X"D0",X"00",X"DD",X"D3",X"10",X"00",X"DD",X"D3",X"10",
		X"00",X"DD",X"33",X"10",X"00",X"DD",X"D3",X"10",X"21",X"DD",X"D3",X"10",X"2C",X"DD",X"33",X"10",
		X"33",X"11",X"23",X"10",X"33",X"33",X"22",X"10",X"33",X"33",X"33",X"10",X"33",X"1A",X"1A",X"10",
		X"2C",X"DD",X"DD",X"10",X"21",X"DD",X"DD",X"10",X"00",X"DD",X"DD",X"10",X"00",X"11",X"11",X"11",
		X"01",X"33",X"33",X"31",X"11",X"33",X"33",X"33",X"11",X"11",X"11",X"11",X"2A",X"2A",X"22",X"22",
		X"11",X"11",X"11",X"11",X"13",X"33",X"33",X"33",X"11",X"DD",X"DD",X"DD",X"01",X"11",X"11",X"11",
		X"55",X"00",X"00",X"55",X"5A",X"00",X"00",X"CC",X"C5",X"00",X"00",X"CC",X"C5",X"00",X"00",X"CC",
		X"C5",X"00",X"00",X"C6",X"55",X"00",X"00",X"CC",X"5A",X"00",X"00",X"CC",X"C5",X"00",X"22",X"CC",
		X"C5",X"22",X"22",X"CC",X"C5",X"22",X"C2",X"C6",X"55",X"22",X"7C",X"CC",X"5A",X"22",X"7C",X"CC",
		X"C5",X"2C",X"77",X"CC",X"C5",X"C7",X"77",X"CC",X"C5",X"77",X"57",X"C6",X"55",X"77",X"55",X"CC",
		X"5A",X"75",X"55",X"CC",X"C5",X"55",X"55",X"CC",X"C5",X"55",X"55",X"CC",X"C5",X"55",X"55",X"C6",
		X"55",X"55",X"55",X"CC",X"5A",X"75",X"55",X"CC",X"C5",X"77",X"55",X"CC",X"C5",X"C7",X"57",X"CC",
		X"C5",X"C7",X"77",X"C6",X"55",X"CC",X"CC",X"CC",X"5A",X"07",X"22",X"CC",X"C5",X"07",X"22",X"CC",
		X"55",X"07",X"77",X"CC",X"55",X"07",X"0C",X"5C",X"05",X"07",X"00",X"55",X"05",X"07",X"00",X"05",
		X"55",X"C2",X"52",X"25",X"55",X"C2",X"52",X"25",X"5C",X"C5",X"CC",X"55",X"A5",X"55",X"55",X"5A",
		X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"55",X"66",X"66",X"6A",X"05",X"CC",X"CC",X"CC",
		X"00",X"55",X"CC",X"55",X"00",X"55",X"77",X"50",X"00",X"55",X"55",X"C0",X"00",X"55",X"55",X"C7",
		X"00",X"5C",X"55",X"C2",X"00",X"C7",X"55",X"C2",X"00",X"7C",X"55",X"C2",X"00",X"C7",X"55",X"C2",
		X"00",X"C7",X"55",X"C2",X"00",X"7C",X"55",X"C2",X"00",X"C7",X"55",X"C2",X"00",X"5C",X"55",X"C2",
		X"00",X"55",X"55",X"C7",X"00",X"55",X"55",X"C0",X"00",X"55",X"77",X"50",X"00",X"55",X"CC",X"55",
		X"05",X"CC",X"CC",X"CC",X"55",X"66",X"66",X"6A",X"CC",X"CC",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",
		X"A5",X"55",X"55",X"5A",X"5C",X"C5",X"CC",X"55",X"55",X"C2",X"52",X"25",X"55",X"CC",X"5C",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"F0",X"00",
		X"00",X"FA",X"3F",X"00",X"00",X"59",X"33",X"00",X"00",X"55",X"93",X"90",X"00",X"55",X"59",X"00",
		X"00",X"53",X"AA",X"00",X"00",X"33",X"A5",X"00",X"00",X"39",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"55",X"55",X"F0",X"00",X"33",X"99",X"00",X"00",X"93",X"99",X"00",X"00",X"39",X"A9",X"00",
		X"00",X"93",X"AA",X"00",X"00",X"93",X"53",X"00",X"00",X"33",X"33",X"50",X"00",X"33",X"3A",X"00",
		X"00",X"33",X"3F",X"00",X"00",X"33",X"F0",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"02",X"00",X"EE",X"22",X"23",X"0E",X"EE",X"22",
		X"32",X"2E",X"EE",X"00",X"23",X"00",X"E0",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"02",X"E2",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"20",X"00",X"00",X"22",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"33",X"00",X"00",X"2A",X"B3",
		X"00",X"00",X"22",X"B3",X"00",X"00",X"22",X"B3",X"00",X"00",X"72",X"B3",X"00",X"00",X"A7",X"B3",
		X"00",X"00",X"AA",X"B3",X"00",X"00",X"0A",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"02",X"20",X"00",X"00",X"22",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"20",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"02",X"20",X"00",
		X"00",X"02",X"00",X"00",X"DD",X"20",X"00",X"00",X"D6",X"20",X"00",X"00",X"D6",X"00",X"00",X"00",
		X"D6",X"DD",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"20",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"07",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"07",X"CF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"0F",X"C7",X"00",X"00",X"07",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",
		X"00",X"00",X"0F",X"CF",X"00",X"00",X"0F",X"7C",X"00",X"00",X"7F",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0F",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"7F",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"2C",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0F",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"7F",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"F7",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"7C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",
		X"00",X"00",X"07",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",
		X"00",X"00",X"07",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"07",X"FF",X"F7",
		X"00",X"00",X"FF",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"7C",X"00",X"00",X"F0",X"CC",X"70",X"0F",X"F7",
		X"7C",X"77",X"FF",X"FF",X"07",X"77",X"FF",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"FF",X"07",X"00",X"FC",X"CF",X"CC",X"77",X"FC",X"CF",
		X"CC",X"77",X"FC",X"CF",X"07",X"00",X"FC",X"CF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"EE",X"39",X"93",X"33",X"EE",X"E9",X"99",
		X"E9",X"99",X"99",X"99",X"9E",X"9E",X"99",X"EE",X"9C",X"E9",X"99",X"99",X"EC",X"99",X"99",X"99",
		X"EC",X"99",X"99",X"33",X"9C",X"E9",X"E9",X"EE",X"93",X"EE",X"E9",X"99",X"30",X"EE",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"3E",X"33",X"00",X"00",
		X"9E",X"99",X"00",X"00",X"EE",X"EE",X"00",X"00",X"E9",X"99",X"00",X"00",X"E9",X"33",X"00",X"00",
		X"33",X"EE",X"00",X"00",X"EE",X"99",X"00",X"00",X"E9",X"33",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"EE",X"39",X"9E",X"33",X"EE",X"E9",X"9E",
		X"E9",X"99",X"99",X"EE",X"9E",X"9E",X"99",X"99",X"9C",X"E9",X"99",X"99",X"EC",X"99",X"99",X"93",
		X"EC",X"99",X"99",X"33",X"9C",X"E9",X"E9",X"99",X"93",X"EE",X"E9",X"EE",X"30",X"EE",X"33",X"9E",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"33",X"00",X"00",X"99",X"E9",X"00",X"00",
		X"33",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"4E",X"E0",X"00",X"00",X"44",X"EE",X"00",
		X"00",X"04",X"E9",X"99",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"04",X"EE",X"00",
		X"00",X"44",X"EE",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"40",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"EE",X"40",X"00",X"00",X"E9",X"40",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"E0",X"00",X"99",X"0F",X"E9",X"00",X"EE",X"CC",X"CC",X"E0",
		X"EE",X"EE",X"CC",X"E0",X"EE",X"CC",X"CC",X"E0",X"EC",X"CC",X"CC",X"FF",X"EC",X"CC",X"CC",X"FF",
		X"EC",X"CC",X"CC",X"FF",X"EC",X"CC",X"CC",X"FF",X"EE",X"CC",X"CC",X"E0",X"EE",X"EE",X"CC",X"E0",
		X"EE",X"CC",X"CC",X"E0",X"99",X"0F",X"E9",X"00",X"00",X"09",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"9E",X"EE",X"00",X"00",X"9E",X"EE",X"00",
		X"00",X"9E",X"CE",X"00",X"00",X"9E",X"CE",X"00",X"00",X"9E",X"CE",X"00",X"00",X"9E",X"CE",X"00",
		X"00",X"0C",X"CE",X"00",X"00",X"0C",X"CE",X"00",X"00",X"0C",X"CE",X"00",X"00",X"FC",X"CE",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"EC",X"CC",X"00",X"00",X"E9",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"0E",X"1C",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"70",X"00",X"FF",X"0F",X"74",X"00",X"77",X"CC",X"CC",X"70",
		X"77",X"77",X"CC",X"70",X"77",X"CC",X"CC",X"70",X"7C",X"CC",X"CC",X"FF",X"7C",X"CC",X"CC",X"FF",
		X"7C",X"CC",X"CC",X"FF",X"7C",X"CC",X"CC",X"FF",X"77",X"CC",X"CC",X"70",X"77",X"77",X"CC",X"70",
		X"77",X"CC",X"CC",X"70",X"FF",X"0F",X"74",X"00",X"00",X"0F",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"F7",X"77",X"00",X"00",X"F7",X"77",X"00",
		X"00",X"F7",X"C7",X"00",X"00",X"F7",X"C7",X"00",X"00",X"F7",X"C7",X"00",X"00",X"F7",X"C7",X"00",
		X"00",X"0C",X"C7",X"00",X"00",X"0C",X"C7",X"00",X"00",X"0C",X"C7",X"00",X"00",X"FC",X"C7",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"CC",X"00",X"00",X"4C",X"CC",X"00",
		X"00",X"7C",X"CC",X"00",X"00",X"74",X"CC",X"00",X"00",X"04",X"CC",X"00",X"00",X"07",X"4C",X"00",
		X"00",X"07",X"CC",X"00",X"00",X"07",X"CC",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"10",
		X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",
		X"13",X"13",X"13",X"10",X"31",X"31",X"31",X"30",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"05",X"35",X"35",X"35",
		X"0B",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",
		X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",
		X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",
		X"06",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",
		X"06",X"60",X"60",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"7F",X"00",X"00",X"00",X"A0",X"00",X"02",X"00",X"00",X"A0",X"79",X"00",X"B0",X"7F",X"00",
		X"00",X"00",X"00",X"09",X"00",X"A0",X"00",X"0A",X"00",X"00",X"00",X"50",X"00",X"F0",X"90",X"00",
		X"A0",X"07",X"09",X"00",X"0A",X"A0",X"90",X"A0",X"79",X"09",X"09",X"02",X"00",X"E0",X"20",X"90",
		X"00",X"00",X"0B",X"05",X"00",X"A0",X"A0",X"E0",X"00",X"09",X"00",X"02",X"00",X"E0",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"07",X"00",X"00",X"00",X"90",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"07",X"11",X"00",X"00",
		X"03",X"99",X"00",X"00",X"03",X"99",X"00",X"00",X"03",X"99",X"00",X"00",X"03",X"79",X"00",X"00",
		X"03",X"79",X"00",X"00",X"03",X"79",X"07",X"00",X"03",X"79",X"00",X"00",X"03",X"93",X"00",X"00",
		X"03",X"93",X"00",X"00",X"03",X"93",X"00",X"07",X"04",X"93",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"43",X"00",X"00",X"44",X"93",X"00",X"00",X"04",X"93",X"00",X"07",X"03",X"93",X"00",X"00",
		X"03",X"93",X"00",X"00",X"03",X"79",X"00",X"00",X"07",X"79",X"07",X"00",X"00",X"79",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"70",X"00",X"77",X"55",X"50",X"00",X"55",
		X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",
		X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",
		X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"55",X"00",X"50",X"55",X"00",X"00",X"C5",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"5C",X"CC",X"55",X"CC",
		X"5C",X"C5",X"00",X"CC",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"CC",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"C5",X"50",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"05",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",
		X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"05",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"50",X"00",X"00",X"00",X"C5",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"22",X"77",X"00",
		X"00",X"22",X"77",X"00",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"77",X"77",X"00",X"22",X"77",X"77",X"00",X"22",
		X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"77",X"66",X"66",X"00",X"77",X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"22",X"62",X"66",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"22",X"66",X"22",X"22",X"22",X"66",
		X"00",X"77",X"77",X"22",X"00",X"72",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",
		X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"77",X"77",X"00",X"22",X"77",X"77",X"00",X"22",
		X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"77",X"66",X"66",X"00",X"77",X"66",X"66",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"22",X"62",X"66",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"22",X"66",X"22",X"22",X"22",X"66",
		X"00",X"77",X"77",X"22",X"00",X"72",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",
		X"77",X"66",X"00",X"00",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"CC",X"77",X"00",X"00",X"0C",
		X"77",X"00",X"00",X"00",X"77",X"CC",X"00",X"00",X"C7",X"77",X"CC",X"00",X"CC",X"77",X"CC",X"00",
		X"00",X"22",X"77",X"C0",X"00",X"22",X"77",X"C0",X"CC",X"22",X"77",X"C0",X"CC",X"22",X"77",X"C0",
		X"77",X"22",X"22",X"00",X"77",X"22",X"22",X"00",X"22",X"22",X"22",X"C0",X"22",X"72",X"77",X"C0",
		X"77",X"77",X"72",X"77",X"77",X"77",X"22",X"77",X"77",X"22",X"22",X"CC",X"77",X"22",X"22",X"CC",
		X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"77",X"22",X"22",X"CC",X"77",X"72",X"22",X"CC",
		X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"55",X"00",X"CC",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"AA",X"A0",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"BB",X"C0",X"00",X"00",X"BB",X"C0",X"00",
		X"00",X"BB",X"C0",X"00",X"00",X"BB",X"C0",X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"2A",X"00",X"10",X"11",X"23",X"00",X"11",X"21",X"33",X"00",X"11",X"A1",X"33",X"00",X"13",
		X"21",X"13",X"00",X"13",X"21",X"23",X"00",X"13",X"21",X"13",X"00",X"13",X"A1",X"A3",X"11",X"13",
		X"21",X"13",X"DD",X"13",X"21",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"A1",X"A3",X"DD",X"13",
		X"21",X"13",X"DD",X"13",X"21",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"21",X"A3",X"22",X"13",
		X"A1",X"13",X"32",X"13",X"21",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"21",X"A3",X"33",X"13",
		X"21",X"13",X"33",X"13",X"A1",X"23",X"DD",X"13",X"21",X"13",X"DD",X"13",X"21",X"13",X"32",X"13",
		X"21",X"13",X"22",X"13",X"A1",X"D2",X"DD",X"13",X"21",X"11",X"11",X"13",X"21",X"00",X"00",X"13",
		X"A1",X"00",X"00",X"13",X"21",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"10",
		X"11",X"11",X"11",X"10",X"DD",X"DD",X"DD",X"11",X"33",X"33",X"33",X"31",X"11",X"11",X"11",X"11",
		X"22",X"22",X"2A",X"A2",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"11",X"13",X"33",X"22",X"10",
		X"11",X"11",X"32",X"00",X"00",X"DD",X"33",X"00",X"00",X"DD",X"3D",X"00",X"00",X"DD",X"3D",X"00",
		X"00",X"DD",X"33",X"00",X"00",X"DD",X"3D",X"00",X"A0",X"DD",X"3D",X"00",X"10",X"DD",X"33",X"00",
		X"12",X"12",X"32",X"00",X"33",X"33",X"22",X"00",X"33",X"33",X"33",X"00",X"12",X"12",X"12",X"00",
		X"10",X"DD",X"DD",X"00",X"A0",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"11",X"11",X"11",X"00",
		X"13",X"33",X"33",X"10",X"33",X"33",X"33",X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"2A",X"A2",
		X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"31",X"DD",X"DD",X"DD",X"11",X"11",X"11",X"11",X"10",
		X"55",X"00",X"00",X"55",X"CC",X"00",X"00",X"A5",X"CC",X"00",X"00",X"5C",X"CC",X"00",X"00",X"5C",
		X"6C",X"00",X"00",X"5C",X"CC",X"00",X"00",X"55",X"CC",X"00",X"00",X"A5",X"CC",X"22",X"00",X"5C",
		X"CC",X"22",X"22",X"5C",X"6C",X"2C",X"22",X"5C",X"CC",X"C7",X"22",X"55",X"CC",X"C7",X"22",X"A5",
		X"CC",X"77",X"C2",X"5C",X"CC",X"77",X"7C",X"5C",X"6C",X"75",X"77",X"5C",X"CC",X"55",X"77",X"55",
		X"CC",X"55",X"57",X"A5",X"CC",X"55",X"55",X"5C",X"CC",X"55",X"55",X"5C",X"6C",X"55",X"55",X"5C",
		X"CC",X"55",X"55",X"55",X"CC",X"55",X"57",X"A5",X"CC",X"55",X"77",X"5C",X"CC",X"75",X"7C",X"5C",
		X"6C",X"77",X"7C",X"5C",X"CC",X"CC",X"CC",X"55",X"CC",X"22",X"70",X"A5",X"CC",X"22",X"70",X"5C",
		X"CC",X"77",X"70",X"55",X"C5",X"C0",X"70",X"55",X"55",X"00",X"70",X"50",X"55",X"00",X"70",X"05",
		X"2C",X"55",X"C2",X"55",X"2C",X"55",X"C2",X"55",X"CC",X"5C",X"C5",X"25",X"55",X"A5",X"55",X"55",
		X"C6",X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"A6",X"66",X"6C",X"5C",X"CC",X"CC",X"C5",
		X"55",X"55",X"CC",X"50",X"00",X"55",X"77",X"00",X"00",X"55",X"55",X"00",X"00",X"5C",X"55",X"77",
		X"00",X"C7",X"55",X"27",X"00",X"77",X"55",X"27",X"00",X"C7",X"55",X"27",X"00",X"7C",X"55",X"27",
		X"00",X"7C",X"55",X"27",X"00",X"C7",X"55",X"27",X"00",X"77",X"55",X"27",X"00",X"C7",X"55",X"27",
		X"00",X"5C",X"55",X"77",X"00",X"55",X"55",X"00",X"00",X"55",X"77",X"00",X"05",X"55",X"CC",X"50",
		X"55",X"CC",X"CC",X"C5",X"CC",X"A6",X"66",X"6C",X"CC",X"CC",X"CC",X"CC",X"C6",X"CC",X"6C",X"CC",
		X"55",X"A5",X"55",X"55",X"CC",X"5C",X"C5",X"25",X"2C",X"55",X"C2",X"55",X"CC",X"55",X"CC",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"A0",X"33",X"00",
		X"00",X"AF",X"33",X"00",X"00",X"AA",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"35",X"39",X"00",
		X"00",X"3A",X"93",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"93",X"00",
		X"00",X"99",X"33",X"00",X"00",X"39",X"35",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"A9",X"00",
		X"00",X"3F",X"AA",X"00",X"00",X"30",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"0E",X"00",X"32",X"00",X"EE",X"EE",X"23",X"22",X"EE",X"E0",X"32",
		X"22",X"EE",X"00",X"20",X"22",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"02",X"00",X"00",
		X"23",X"22",X"00",X"00",X"03",X"22",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"20",X"00",X"00",X"02",X"22",X"00",X"00",X"02",X"02",X"00",X"00",X"02",X"02",X"00",
		X"00",X"02",X"02",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"20",X"00",X"00",X"A6",X"20",X"00",X"00",X"26",X"00",
		X"00",X"00",X"26",X"70",X"00",X"00",X"27",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"7A",X"70",
		X"00",X"00",X"7A",X"00",X"00",X"00",X"AA",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"22",X"00",X"00",X"70",X"00",X"00",X"02",X"03",X"00",X"00",X"02",X"22",X"00",
		X"00",X"02",X"22",X"00",X"00",X"20",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"EE",X"00",X"00",X"2D",X"EB",X"00",X"00",
		X"22",X"DD",X"00",X"00",X"22",X"ED",X"00",X"00",X"72",X"ED",X"00",X"00",X"D7",X"DD",X"00",X"00",
		X"DD",X"EB",X"00",X"00",X"0D",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"02",X"22",X"00",
		X"00",X"02",X"22",X"00",X"00",X"00",X"03",X"00",X"00",X"07",X"70",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FC",X"70",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",
		X"00",X"00",X"C7",X"FF",X"00",X"00",X"FC",X"70",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",
		X"00",X"00",X"C7",X"7F",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"7F",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"7F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"2C",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"FF",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"70",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",
		X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"FF",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"70",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"70",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"F7",X"00",X"00",X"FF",X"77",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"70",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"F7",X"00",X"00",X"FF",X"77",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"77",X"0F",X"00",X"00",X"77",X"FF",X"00",
		X"00",X"00",X"FC",X"F0",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F0",
		X"00",X"00",X"C7",X"F7",X"00",X"00",X"FC",X"F7",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",
		X"CC",X"77",X"FF",X"00",X"77",X"77",X"FC",X"F0",X"00",X"00",X"C7",X"F0",X"00",X"00",X"C7",X"F7",
		X"00",X"00",X"C7",X"F7",X"00",X"00",X"C7",X"F0",X"00",X"00",X"FC",X"00",X"00",X"00",X"7F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"7F",X"00",
		X"00",X"00",X"FC",X"00",X"00",X"00",X"C7",X"00",X"77",X"07",X"7C",X"00",X"CC",X"7F",X"7C",X"70",
		X"CC",X"7F",X"7C",X"70",X"77",X"07",X"7C",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"FC",X"00",
		X"00",X"00",X"7F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"99",X"30",X"33",X"99",X"99",X"93",
		X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"EE",X"44",X"E9",X"99",X"99",X"44",X"9E",X"99",X"99",
		X"C4",X"9E",X"99",X"33",X"44",X"E9",X"9E",X"EE",X"33",X"99",X"9E",X"99",X"00",X"99",X"39",X"33",
		X"00",X"33",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"33",X"00",X"00",
		X"EE",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",
		X"33",X"33",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"33",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"99",X"99",X"EE",X"33",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"99",X"44",X"E9",X"99",X"93",X"44",X"9E",X"99",X"30",
		X"C4",X"9E",X"99",X"30",X"44",X"E9",X"9E",X"93",X"33",X"99",X"9E",X"99",X"00",X"99",X"39",X"99",
		X"00",X"33",X"03",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"03",X"EE",X"00",X"00",
		X"39",X"9E",X"00",X"00",X"3E",X"39",X"00",X"00",X"E9",X"03",X"00",X"00",X"99",X"00",X"00",X"00",
		X"93",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"33",X"00",X"00",
		X"99",X"E9",X"00",X"00",X"33",X"E9",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E9",X"EE",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"4E",X"99",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"4E",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"EE",X"EE",X"00",X"EE",X"CC",X"C9",X"00",
		X"EE",X"EE",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"9E",X"CC",X"11",X"F9",X"9E",X"CC",X"11",X"F9",
		X"9E",X"CC",X"11",X"F9",X"99",X"CC",X"11",X"F9",X"CC",X"CC",X"AC",X"00",X"EE",X"EE",X"CC",X"00",
		X"EE",X"CC",X"C9",X"00",X"99",X"EE",X"EE",X"00",X"99",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"E9",X"00",X"00",X"EE",X"E9",X"00",
		X"00",X"EC",X"E9",X"00",X"00",X"EC",X"E9",X"00",X"00",X"EC",X"E9",X"00",X"00",X"EC",X"E9",X"00",
		X"00",X"EC",X"C0",X"00",X"00",X"EC",X"C0",X"00",X"00",X"EC",X"C0",X"00",X"00",X"EC",X"CF",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"CA",X"CE",X"00",X"00",X"CC",X"9E",X"00",X"00",X"CC",X"90",X"00",X"00",X"C1",X"E0",X"00",
		X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F4",X"00",X"00",X"FF",X"77",X"77",X"00",X"77",X"CC",X"C4",X"00",
		X"77",X"77",X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"F4",X"CC",X"44",X"44",X"F4",X"CC",X"44",X"44",
		X"F4",X"CC",X"44",X"44",X"FF",X"CC",X"44",X"44",X"CC",X"CC",X"CC",X"00",X"77",X"77",X"CC",X"00",
		X"77",X"CC",X"C4",X"00",X"FF",X"77",X"77",X"00",X"FF",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"7F",X"00",X"00",X"77",X"7F",X"00",
		X"00",X"7C",X"7F",X"00",X"00",X"7C",X"7F",X"00",X"00",X"7C",X"7F",X"00",X"00",X"7C",X"7F",X"00",
		X"00",X"7C",X"C0",X"00",X"00",X"7C",X"C0",X"00",X"00",X"7C",X"C0",X"00",X"00",X"7C",X"CF",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"CC",X"C7",X"00",X"00",X"CC",X"C4",X"00",
		X"00",X"CC",X"C7",X"00",X"00",X"CC",X"47",X"00",X"00",X"CC",X"40",X"00",X"00",X"C4",X"70",X"00",
		X"00",X"CC",X"70",X"00",X"00",X"CC",X"70",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"31",X"31",X"31",X"03",X"13",X"13",X"13",X"11",X"31",X"31",X"30",X"11",X"11",X"11",X"10",
		X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"35",X"35",X"35",X"30",
		X"53",X"53",X"53",X"50",X"35",X"35",X"35",X"30",X"53",X"53",X"53",X"50",X"35",X"35",X"35",X"30",
		X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"B0",X"DB",X"DB",X"DB",X"D0",X"BD",X"BD",X"BD",X"B0",
		X"DB",X"DB",X"DB",X"D0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",
		X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"DF",X"DF",X"DF",X"D0",X"0D",X"FD",X"FD",X"FD",X"0F",X"DF",X"DF",X"DF",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"40",
		X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"50",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F5",X"00",X"EA",X"00",X"00",X"00",X"09",X"00",X"FA",X"75",X"A0",
		X"00",X"05",X"07",X"09",X"A0",X"00",X"00",X"97",X"AF",X"00",X"0F",X"00",X"00",X"B0",X"F0",X"00",
		X"40",X"09",X"09",X"00",X"0A",X"A0",X"90",X"00",X"20",X"0B",X"00",X"A5",X"00",X"E0",X"00",X"00",
		X"00",X"02",X"9A",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"0A",X"00",X"90",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"92",X"00",X"00",
		X"09",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"B2",X"00",X"00",X"05",X"0B",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"E3",X"00",X"00",
		X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"04",X"44",X"44",X"00",X"00",
		X"44",X"04",X"00",X"00",X"44",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"07",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"93",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"07",X"77",X"55",X"00",X"05",X"55",
		X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",
		X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",
		X"CC",X"00",X"00",X"C5",X"CC",X"00",X"00",X"C5",X"55",X"05",X"00",X"55",X"00",X"5C",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"CC",X"55",X"CC",X"C5",
		X"CC",X"00",X"5C",X"C5",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"50",
		X"00",X"00",X"50",X"C5",X"00",X"00",X"50",X"C5",X"00",X"00",X"50",X"CC",X"00",X"00",X"50",X"CC",
		X"00",X"00",X"50",X"CC",X"00",X"00",X"50",X"CC",X"00",X"00",X"50",X"C5",X"00",X"00",X"50",X"C5",
		X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",
		X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"66",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"66",X"77",X"66",X"00",X"66",X"77",X"66",X"00",X"22",X"27",X"22",X"00",X"22",X"77",X"22",X"00",
		X"00",X"77",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"77",X"22",X"22",X"00",X"77",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"66",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"66",X"77",X"66",X"00",X"66",X"77",X"66",X"00",X"22",X"27",X"22",X"00",X"22",X"77",X"22",X"00",
		X"00",X"77",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"77",X"22",X"22",X"00",X"77",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"77",X"00",X"00",X"CC",X"77",X"00",X"00",X"CC",
		X"22",X"00",X"00",X"00",X"22",X"CC",X"00",X"00",X"77",X"77",X"CC",X"00",X"77",X"77",X"CC",X"00",
		X"CC",X"22",X"77",X"00",X"CC",X"22",X"77",X"00",X"CC",X"22",X"22",X"00",X"CC",X"22",X"72",X"00",
		X"77",X"77",X"22",X"00",X"77",X"72",X"22",X"00",X"77",X"77",X"22",X"00",X"77",X"77",X"22",X"00",
		X"22",X"77",X"77",X"C0",X"22",X"27",X"77",X"C0",X"22",X"22",X"77",X"00",X"22",X"22",X"77",X"00",
		X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",X"CC",X"22",X"22",X"00",X"CC",X"22",X"22",X"00",
		X"CC",X"77",X"22",X"CC",X"CC",X"77",X"22",X"CC",X"77",X"CC",X"77",X"00",X"77",X"CC",X"77",X"00",
		X"77",X"00",X"CC",X"00",X"77",X"00",X"CC",X"00",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A2",X"00",X"00",X"00",X"32",X"00",X"00",X"10",X"33",X"00",X"10",X"11",X"33",X"00",X"11",
		X"31",X"31",X"01",X"D1",X"33",X"32",X"01",X"D1",X"33",X"31",X"01",X"D1",X"33",X"31",X"11",X"D1",
		X"33",X"31",X"D1",X"D1",X"33",X"32",X"D1",X"D1",X"33",X"31",X"D1",X"D1",X"33",X"31",X"D1",X"D1",
		X"33",X"31",X"D1",X"D1",X"33",X"32",X"D1",X"D1",X"33",X"31",X"D1",X"D1",X"33",X"3A",X"D1",X"D1",
		X"33",X"31",X"21",X"D1",X"33",X"32",X"22",X"D1",X"33",X"22",X"32",X"D1",X"33",X"23",X"33",X"D1",
		X"33",X"23",X"33",X"D1",X"33",X"22",X"32",X"D1",X"33",X"32",X"22",X"D1",X"33",X"31",X"21",X"D1",
		X"33",X"1A",X"D1",X"D1",X"33",X"AD",X"D1",X"D1",X"33",X"11",X"11",X"D1",X"31",X"00",X"01",X"D1",
		X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"00",X"DD",X"DD",X"DD",X"00",X"33",X"33",X"33",X"10",X"11",X"11",X"11",X"11",
		X"2A",X"22",X"22",X"11",X"11",X"11",X"11",X"10",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"11",X"11",X"21",X"00",X"01",X"DD",X"22",X"00",X"01",X"D2",X"D2",X"00",X"01",X"D2",X"D3",X"00",
		X"01",X"D2",X"33",X"00",X"01",X"D2",X"D3",X"00",X"01",X"D2",X"D2",X"00",X"0A",X"DD",X"22",X"00",
		X"11",X"1A",X"21",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"1A",X"1A",X"11",X"00",
		X"01",X"DD",X"DD",X"00",X"01",X"DD",X"DD",X"00",X"01",X"DD",X"DD",X"00",X"11",X"11",X"11",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"11",X"11",X"11",X"10",X"2A",X"22",X"22",X"11",
		X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"10",X"DD",X"DD",X"DD",X"00",X"11",X"11",X"11",X"00",
		X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"50",X"55",X"00",X"00",X"55",X"C5",X"00",X"00",X"2C",
		X"C5",X"00",X"05",X"CC",X"6C",X"00",X"05",X"2C",X"AC",X"20",X"05",X"55",X"6C",X"C5",X"05",X"55",
		X"6C",X"C7",X"05",X"2C",X"6C",X"7C",X"25",X"CC",X"6C",X"C7",X"25",X"2C",X"AC",X"C7",X"25",X"55",
		X"6C",X"7C",X"25",X"55",X"6C",X"77",X"25",X"2C",X"6C",X"55",X"CC",X"CC",X"6C",X"55",X"7C",X"2C",
		X"AC",X"55",X"7C",X"55",X"6C",X"55",X"7C",X"55",X"6C",X"55",X"7C",X"2C",X"6C",X"55",X"7C",X"CC",
		X"6C",X"55",X"7C",X"2C",X"AC",X"55",X"7C",X"55",X"6C",X"55",X"7C",X"55",X"6C",X"55",X"CC",X"2C",
		X"6C",X"77",X"75",X"CC",X"6C",X"CC",X"55",X"2C",X"CC",X"22",X"05",X"55",X"CC",X"22",X"05",X"55",
		X"C5",X"77",X"00",X"50",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"05",
		X"25",X"2C",X"55",X"00",X"25",X"2C",X"55",X"00",X"55",X"CC",X"5C",X"50",X"5A",X"55",X"A5",X"55",
		X"CC",X"C6",X"CC",X"65",X"CC",X"CC",X"CC",X"C5",X"6A",X"66",X"A6",X"55",X"CC",X"CC",X"CC",X"50",
		X"55",X"5C",X"CC",X"00",X"00",X"5C",X"77",X"00",X"00",X"C7",X"77",X"00",X"00",X"77",X"57",X"77",
		X"00",X"77",X"55",X"C0",X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",
		X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",X"00",X"77",X"55",X"C0",
		X"00",X"77",X"57",X"77",X"00",X"C7",X"77",X"00",X"00",X"5C",X"77",X"00",X"55",X"5C",X"CC",X"00",
		X"CC",X"CC",X"CC",X"50",X"6A",X"66",X"A6",X"55",X"CC",X"CC",X"CC",X"C5",X"CC",X"C6",X"CC",X"65",
		X"55",X"55",X"A5",X"55",X"55",X"CC",X"5C",X"50",X"25",X"2C",X"55",X"00",X"C5",X"CC",X"55",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"0F",X"30",X"00",X"00",X"F3",X"30",X"00",
		X"00",X"33",X"3F",X"00",X"55",X"33",X"3F",X"00",X"05",X"35",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"3F",X"00",X"00",X"9A",X"93",X"00",X"0F",X"99",X"59",X"00",
		X"F5",X"55",X"55",X"00",X"0F",X"33",X"93",X"00",X"00",X"39",X"33",X"00",X"00",X"99",X"3F",X"00",
		X"00",X"99",X"55",X"00",X"00",X"55",X"55",X"00",X"09",X"95",X"55",X"00",X"99",X"39",X"95",X"00",
		X"00",X"33",X"FF",X"00",X"00",X"F3",X"00",X"00",X"00",X"0F",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"22",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E2",X"22",X"20",X"22",X"22",X"00",X"00",
		X"22",X"BB",X"00",X"00",X"22",X"EB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"32",X"30",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"32",X"00",X"00",X"20",X"22",X"00",
		X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"02",X"00",X"00",X"20",X"22",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D6",X"EE",X"00",X"00",X"26",X"BE",X"00",X"00",
		X"26",X"BE",X"00",X"00",X"27",X"BE",X"00",X"00",X"77",X"BE",X"00",X"00",X"7D",X"BE",X"00",X"00",
		X"7D",X"BE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"23",X"30",X"00",X"00",X"22",X"22",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"7C",X"00",
		X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",
		X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",
		X"C7",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"00",X"F7",X"F7",X"00",X"00",X"FF",X"CC",X"00",
		X"00",X"FF",X"77",X"00",X"00",X"7F",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"7F",X"00",X"C7",X"00",X"FF",X"00",
		X"C7",X"F7",X"CC",X"00",X"00",X"FF",X"77",X"00",X"00",X"7F",X"CC",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"70",X"FF",X"CC",X"00",X"CC",X"FF",X"77",X"00",
		X"CC",X"FF",X"77",X"00",X"70",X"FF",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"00",X"03",X"99",X"E9",X"00",X"03",X"99",X"E9",X"33",
		X"39",X"9E",X"EE",X"99",X"99",X"99",X"EE",X"EE",X"49",X"99",X"9E",X"99",X"C4",X"99",X"99",X"99",
		X"C4",X"99",X"EE",X"33",X"49",X"9E",X"EE",X"EE",X"33",X"99",X"99",X"99",X"03",X"33",X"99",X"33",
		X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"E9",X"30",X"00",X"00",X"9E",X"93",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",
		X"33",X"9E",X"00",X"00",X"EE",X"39",X"00",X"00",X"99",X"93",X"00",X"00",X"33",X"39",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"39",X"03",X"33",X"33",X"9E",X"03",X"99",X"E9",X"EE",X"03",X"99",X"E9",X"99",
		X"39",X"9E",X"EE",X"99",X"99",X"99",X"EE",X"93",X"49",X"99",X"9E",X"30",X"C4",X"99",X"99",X"00",
		X"C4",X"99",X"EE",X"00",X"49",X"9E",X"EE",X"30",X"33",X"99",X"9E",X"93",X"03",X"33",X"99",X"99",
		X"00",X"00",X"39",X"EE",X"00",X"00",X"03",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"9E",X"30",X"00",X"00",
		X"E9",X"30",X"00",X"00",X"99",X"30",X"00",X"00",X"93",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"99",X"30",X"00",X"00",X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"E0",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"E0",X"00",X"00",X"99",X"E9",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"99",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"99",X"EE",X"00",X"00",X"EE",X"CC",X"9E",X"00",
		X"EE",X"EE",X"CC",X"00",X"CC",X"CC",X"C1",X"00",X"EE",X"CC",X"11",X"99",X"EE",X"CC",X"11",X"99",
		X"EE",X"CC",X"11",X"99",X"EE",X"CC",X"11",X"99",X"CC",X"CC",X"C1",X"00",X"EE",X"EE",X"CC",X"00",
		X"EE",X"CC",X"9E",X"00",X"99",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9E",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"F0",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"47",X"00",X"00",X"FF",X"77",X"00",X"00",X"77",X"CC",X"47",X"00",
		X"77",X"77",X"CC",X"00",X"CC",X"CC",X"C4",X"00",X"4C",X"CC",X"44",X"44",X"4C",X"CC",X"44",X"44",
		X"4C",X"CC",X"44",X"44",X"4C",X"CC",X"44",X"44",X"CC",X"CC",X"C4",X"00",X"77",X"77",X"CC",X"00",
		X"77",X"CC",X"47",X"00",X"FF",X"77",X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"F4",X"F0",X"00",X"00",X"44",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"F0",X"00",
		X"00",X"CC",X"F0",X"00",X"00",X"CC",X"40",X"00",X"00",X"CC",X"40",X"00",X"00",X"CC",X"70",X"00",
		X"00",X"CC",X"70",X"00",X"00",X"CC",X"70",X"00",X"00",X"CC",X"70",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"53",X"53",X"53",X"05",X"35",X"35",X"35",X"03",X"53",X"53",X"53",X"05",X"35",X"35",X"35",
		X"33",X"53",X"53",X"50",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",
		X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",
		X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"35",X"35",X"35",X"00",
		X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",
		X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",
		X"DB",X"DB",X"DB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",
		X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"BD",X"BD",X"BD",X"00",
		X"DB",X"DB",X"DB",X"D0",X"BD",X"BD",X"BD",X"B0",X"DB",X"DB",X"DB",X"D0",X"BD",X"BD",X"BD",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"D0",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"65",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"05",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"06",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"65",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"05",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"0E",X"00",X"05",X"00",X"E0",X"0A",X"00",X"7F",X"09",X"00",X"00",X"F0",X"20",
		X"0A",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"A0",X"AB",X"00",X"0B",X"00",X"F0",X"F0",X"F0",X"00",
		X"0A",X"09",X"09",X"00",X"90",X"20",X"90",X"00",X"0E",X"0B",X"00",X"B0",X"00",X"00",X"00",X"A5",
		X"0E",X"00",X"0B",X"00",X"0A",X"00",X"2E",X"A0",X"00",X"0B",X"00",X"00",X"00",X"09",X"00",X"A7",
		X"00",X"90",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"95",X"00",X"00",X"7E",X"09",X"00",X"00",X"90",X"05",X"00",X"00",
		X"09",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"07",X"00",
		X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"44",X"44",X"00",X"40",X"44",X"40",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"07",X"00",X"00",X"00",
		X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"55",X"00",X"55",X"00",
		X"CC",X"00",X"5C",X"00",X"CC",X"00",X"05",X"00",X"C5",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"55",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"50",X"50",X"00",
		X"50",X"00",X"C5",X"00",X"55",X"50",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"55",X"55",X"00",X"75",X"CC",X"5C",X"00",
		X"75",X"CC",X"5C",X"00",X"75",X"CC",X"5C",X"00",X"75",X"55",X"55",X"00",X"75",X"00",X"00",X"00",
		X"75",X"00",X"00",X"00",X"75",X"00",X"05",X"00",X"75",X"00",X"5C",X"00",X"00",X"00",X"5C",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"75",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5C",X"00",X"75",X"00",X"5C",X"00",X"75",X"00",X"05",X"00",X"75",X"00",X"00",X"00",
		X"75",X"00",X"00",X"00",X"75",X"55",X"55",X"00",X"75",X"CC",X"5C",X"00",X"75",X"CC",X"5C",X"00",
		X"75",X"CC",X"5C",X"00",X"75",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");

begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;