library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity botanic_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of botanic_tile_bit0 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"E6",X"E4",X"00",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"00",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"02",X"02",X"01",X"3F",X"60",X"20",X"3C",X"42",X"A5",X"A5",X"A5",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"0C",X"1A",X"18",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"42",X"A5",X"A5",X"A5",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"03",X"06",X"07",X"17",X"05",X"00",X"00",X"00",X"E0",X"30",X"F8",X"FC",X"B4",
		X"05",X"17",X"07",X"06",X"03",X"00",X"00",X"00",X"B4",X"FC",X"F8",X"30",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"06",X"07",X"17",X"05",X"00",X"00",X"00",X"E0",X"30",X"F8",X"FC",X"B4",
		X"05",X"17",X"07",X"06",X"03",X"00",X"00",X"00",X"B4",X"FC",X"F8",X"30",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"0F",X"1E",X"17",X"00",X"00",X"00",X"40",X"00",X"F0",X"78",X"E8",
		X"17",X"16",X"1F",X"0F",X"06",X"03",X"00",X"00",X"E8",X"68",X"F8",X"F0",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"0F",X"1E",X"17",X"00",X"00",X"00",X"40",X"00",X"F0",X"78",X"E8",
		X"17",X"16",X"1F",X"0F",X"06",X"03",X"00",X"00",X"E8",X"68",X"F8",X"F0",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"19",X"05",X"03",X"13",X"00",X"00",X"00",X"C0",X"1C",X"20",X"F0",X"58",
		X"01",X"13",X"03",X"05",X"19",X"00",X"00",X"00",X"F8",X"58",X"F0",X"20",X"1C",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"05",X"03",X"13",X"00",X"00",X"00",X"98",X"20",X"20",X"F0",X"58",
		X"01",X"13",X"03",X"05",X"09",X"08",X"00",X"00",X"F8",X"58",X"F0",X"20",X"20",X"98",X"00",X"00",
		X"00",X"00",X"00",X"12",X"10",X"08",X"06",X"1F",X"00",X"00",X"00",X"90",X"10",X"20",X"C0",X"F0",
		X"25",X"27",X"0D",X"17",X"13",X"10",X"00",X"00",X"48",X"C8",X"60",X"D0",X"90",X"10",X"00",X"00",
		X"00",X"00",X"00",X"02",X"30",X"08",X"06",X"1F",X"00",X"00",X"00",X"80",X"18",X"20",X"C0",X"F0",
		X"25",X"07",X"1D",X"27",X"23",X"00",X"00",X"00",X"48",X"C0",X"70",X"C8",X"88",X"00",X"00",X"00",
		X"00",X"02",X"1C",X"19",X"10",X"08",X"44",X"69",X"00",X"22",X"C2",X"1C",X"90",X"48",X"3C",X"E6",
		X"7F",X"69",X"44",X"08",X"10",X"19",X"1C",X"02",X"1B",X"E6",X"3C",X"48",X"90",X"1C",X"C2",X"22",
		X"00",X"70",X"B8",X"09",X"05",X"08",X"88",X"D3",X"00",X"01",X"13",X"E4",X"08",X"90",X"78",X"CC",
		X"FE",X"D3",X"88",X"08",X"05",X"09",X"B8",X"70",X"36",X"CC",X"78",X"90",X"08",X"E4",X"13",X"01",
		X"00",X"07",X"03",X"71",X"6B",X"45",X"81",X"23",X"00",X"C0",X"80",X"1C",X"AC",X"44",X"02",X"88",
		X"52",X"4A",X"86",X"35",X"2D",X"26",X"C3",X"01",X"94",X"A4",X"C2",X"58",X"68",X"C8",X"86",X"00",
		X"47",X"83",X"C1",X"C3",X"6D",X"11",X"03",X"32",X"C4",X"82",X"06",X"86",X"6C",X"10",X"80",X"98",
		X"2A",X"26",X"25",X"4D",X"16",X"23",X"41",X"C0",X"A8",X"C8",X"48",X"64",X"D0",X"88",X"04",X"06",
		X"00",X"03",X"02",X"61",X"18",X"06",X"01",X"1A",X"00",X"06",X"0C",X"88",X"8B",X"52",X"24",X"A8",
		X"00",X"1A",X"01",X"06",X"18",X"61",X"02",X"03",X"AC",X"A8",X"24",X"52",X"8B",X"88",X"0C",X"06",
		X"00",X"08",X"04",X"04",X"02",X"02",X"01",X"1A",X"00",X"44",X"89",X"D2",X"52",X"54",X"24",X"A8",
		X"00",X"1A",X"01",X"02",X"02",X"04",X"04",X"08",X"AC",X"A8",X"24",X"54",X"52",X"D2",X"89",X"44",
		X"00",X"20",X"20",X"12",X"12",X"08",X"CA",X"A4",X"00",X"08",X"08",X"90",X"90",X"20",X"A6",X"4A",
		X"33",X"08",X"07",X"08",X"73",X"C5",X"98",X"10",X"98",X"20",X"C0",X"20",X"9C",X"46",X"32",X"10",
		X"00",X"00",X"00",X"02",X"82",X"60",X"1A",X"04",X"00",X"00",X"00",X"80",X"82",X"0C",X"B0",X"40",
		X"63",X"B8",X"07",X"38",X"43",X"8D",X"30",X"40",X"8C",X"3A",X"C0",X"38",X"84",X"62",X"18",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"7F",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"7F",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"1E",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"1E",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"01",X"38",X"CD",X"07",X"00",X"40",X"44",X"24",X"12",X"BC",X"BF",X"BF",
		X"01",X"07",X"CD",X"38",X"01",X"01",X"03",X"00",X"80",X"BF",X"BF",X"BC",X"12",X"24",X"44",X"40",
		X"00",X"00",X"06",X"02",X"01",X"00",X"7D",X"87",X"00",X"04",X"0D",X"11",X"12",X"BC",X"BF",X"BF",
		X"01",X"87",X"7D",X"00",X"01",X"02",X"06",X"00",X"80",X"BF",X"BF",X"BC",X"12",X"11",X"0D",X"04",
		X"04",X"04",X"08",X"08",X"0C",X"06",X"42",X"77",X"40",X"40",X"20",X"20",X"60",X"C0",X"84",X"DC",
		X"0F",X"C0",X"2E",X"1E",X"0E",X"6E",X"16",X"06",X"E0",X"06",X"E8",X"F0",X"E0",X"EC",X"D0",X"C0",
		X"02",X"04",X"04",X"04",X"04",X"46",X"62",X"17",X"80",X"40",X"40",X"40",X"40",X"C4",X"8C",X"D0",
		X"0F",X"00",X"0E",X"3E",X"4E",X"CE",X"16",X"66",X"E0",X"00",X"E0",X"F8",X"E4",X"E6",X"D0",X"CC",
		X"00",X"00",X"00",X"04",X"04",X"07",X"1B",X"0D",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"40",
		X"14",X"0A",X"1A",X"06",X"05",X"01",X"00",X"00",X"CC",X"80",X"88",X"84",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"1F",X"07",X"06",X"05",X"00",X"00",X"00",X"00",X"C0",X"28",X"F4",X"F0",
		X"03",X"07",X"0F",X"1F",X"18",X"00",X"00",X"00",X"FC",X"F0",X"E4",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"07",X"04",X"1B",X"00",X"00",X"00",X"00",X"60",X"70",X"70",X"A0",
		X"3B",X"1B",X"04",X"07",X"06",X"00",X"00",X"00",X"80",X"A0",X"70",X"70",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"40",X"A0",X"40",
		X"02",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"00",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",
		X"00",X"05",X"05",X"05",X"07",X"07",X"00",X"00",X"E0",X"F0",X"10",X"10",X"30",X"20",X"00",X"00",
		X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"03",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",X"10",
		X"02",X"01",X"00",X"07",X"07",X"02",X"00",X"00",X"30",X"F0",X"10",X"F0",X"F0",X"10",X"10",X"00",
		X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"03",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",X"10",
		X"02",X"03",X"07",X"05",X"04",X"04",X"06",X"02",X"30",X"F0",X"90",X"D0",X"D0",X"F0",X"70",X"30",
		X"01",X"03",X"02",X"01",X"03",X"02",X"01",X"03",X"E0",X"10",X"30",X"E0",X"10",X"30",X"E0",X"10",
		X"02",X"05",X"06",X"07",X"05",X"04",X"04",X"00",X"30",X"E0",X"F0",X"90",X"90",X"90",X"30",X"20",
		X"00",X"03",X"0F",X"1F",X"03",X"2F",X"3B",X"1F",X"00",X"F0",X"E0",X"80",X"04",X"84",X"C8",X"A0",
		X"1F",X"1F",X"3B",X"2F",X"03",X"1F",X"0F",X"03",X"D0",X"A0",X"C8",X"84",X"04",X"80",X"E0",X"F0",
		X"00",X"FF",X"0F",X"07",X"03",X"2F",X"3B",X"1F",X"00",X"00",X"C0",X"C0",X"00",X"84",X"CC",X"A0",
		X"1F",X"1F",X"3B",X"2F",X"03",X"07",X"0F",X"FF",X"D0",X"A0",X"CC",X"84",X"00",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"07",X"07",X"71",X"3B",X"17",X"00",X"1E",X"F0",X"C0",X"80",X"86",X"EC",X"F2",
		X"1F",X"17",X"3B",X"71",X"07",X"07",X"00",X"00",X"F8",X"F2",X"EC",X"86",X"80",X"C0",X"F0",X"1E",
		X"00",X"07",X"3F",X"0F",X"07",X"71",X"3B",X"17",X"00",X"F8",X"E0",X"C0",X"86",X"84",X"EC",X"F2",
		X"1F",X"17",X"3B",X"71",X"07",X"0F",X"3F",X"07",X"F8",X"F2",X"EC",X"84",X"86",X"C0",X"E0",X"F8",
		X"00",X"0F",X"10",X"10",X"0F",X"00",X"0F",X"10",X"00",X"F8",X"04",X"04",X"F8",X"00",X"F8",X"04",
		X"10",X"0F",X"00",X"0F",X"10",X"10",X"10",X"0C",X"04",X"F8",X"00",X"04",X"84",X"44",X"24",X"1C",
		X"00",X"0F",X"10",X"10",X"0F",X"00",X"0F",X"10",X"00",X"F8",X"04",X"04",X"F8",X"00",X"F8",X"04",
		X"10",X"0F",X"00",X"00",X"08",X"06",X"01",X"00",X"04",X"F8",X"00",X"10",X"FC",X"10",X"90",X"70",
		X"00",X"0F",X"10",X"10",X"0F",X"00",X"0F",X"10",X"00",X"F8",X"04",X"04",X"F8",X"00",X"F8",X"04",
		X"10",X"0F",X"00",X"0F",X"10",X"10",X"10",X"0F",X"04",X"F8",X"00",X"78",X"84",X"84",X"84",X"78",
		X"1F",X"10",X"1F",X"00",X"1F",X"10",X"1F",X"00",X"FC",X"04",X"FC",X"00",X"FC",X"04",X"FC",X"00",
		X"0C",X"11",X"11",X"0F",X"00",X"00",X"1F",X"10",X"F8",X"04",X"04",X"F8",X"00",X"04",X"FC",X"04",
		X"1F",X"10",X"1F",X"00",X"1F",X"10",X"1F",X"00",X"FC",X"04",X"FC",X"00",X"FC",X"04",X"FC",X"00",
		X"1F",X"10",X"1C",X"00",X"1F",X"10",X"10",X"1C",X"04",X"C4",X"3C",X"00",X"7C",X"84",X"84",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"13",X"3F",X"3F",X"00",X"00",X"00",X"00",X"22",X"77",X"DD",X"DD",
		X"3F",X"3F",X"13",X"03",X"00",X"00",X"00",X"00",X"DD",X"DD",X"77",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"09",X"1F",X"1F",X"00",X"00",X"02",X"17",X"BD",X"ED",X"ED",X"ED",
		X"1F",X"19",X"09",X"07",X"00",X"00",X"00",X"00",X"EF",X"FA",X"90",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"77",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"DD",X"DD",X"77",X"22",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"E8",X"BC",X"B6",X"B7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B7",X"F6",X"5C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"03",X"03",X"0F",X"0F",X"00",X"00",X"C0",X"E0",X"C0",X"C0",X"F0",X"F0",
		X"03",X"07",X"0C",X"07",X"03",X"07",X"0C",X"07",X"C0",X"E0",X"30",X"E0",X"C0",X"E0",X"30",X"E0",
		X"00",X"00",X"00",X"03",X"07",X"09",X"09",X"0F",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"C0",X"F0",
		X"0F",X"03",X"03",X"06",X"03",X"01",X"03",X"01",X"F0",X"E0",X"F0",X"18",X"F0",X"F8",X"0C",X"F8",
		X"03",X"07",X"0C",X"07",X"03",X"07",X"0C",X"07",X"C0",X"E0",X"30",X"E0",X"C0",X"E0",X"30",X"E0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"06",X"03",X"07",X"0C",X"07",X"03",X"01",X"F0",X"18",X"F0",X"E0",X"30",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"0F",X"0F",X"0B",X"03",X"05",X"00",X"01",X"00",X"E0",X"F0",X"E0",X"F8",X"F0",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"07",X"03",X"03",X"07",X"03",X"03",X"07",X"C0",X"C0",X"E0",X"80",X"E0",X"C0",X"E0",X"80",
		X"00",X"02",X"01",X"07",X"03",X"0F",X"0F",X"0F",X"F8",X"F0",X"F8",X"E0",X"F0",X"E0",X"E0",X"C0",
		X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"03",X"01",X"07",X"03",X"03",X"A0",X"80",X"A0",X"C0",X"A0",X"80",X"80",X"C0",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"02",X"06",X"07",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0B",X"03",X"07",X"07",X"07",X"03",X"03",X"05",X"80",X"40",X"C0",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"22",
		X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"02",X"10",X"02",X"12",X"12",X"12",
		X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"10",X"02",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"08",X"40",X"48",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"08",X"40",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",
		X"00",X"00",X"00",X"05",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"F4",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"1F",X"1F",X"1F",X"07",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",
		X"07",X"1F",X"1F",X"1F",X"07",X"00",X"00",X"00",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"1F",X"3F",X"7F",X"7F",X"7F",X"3F",X"0F",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"1F",X"00",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",X"00",
		X"0F",X"1F",X"1F",X"1F",X"0F",X"0E",X"02",X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"D8",X"0C",X"06",
		X"01",X"07",X"1F",X"1F",X"1F",X"0F",X"0F",X"00",X"9A",X"FC",X"F0",X"E0",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"01",X"02",X"04",X"00",X"7F",X"00",X"F5",X"F5",X"77",X"02",X"3E",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7F",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"C0",X"F0",X"3E",X"02",X"77",X"F5",
		X"54",X"50",X"80",X"F0",X"4E",X"1F",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"CE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"1F",X"4E",X"F0",X"80",X"50",X"00",X"00",X"CE",X"FE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"04",X"00",X"03",X"07",X"F5",X"F5",X"77",X"06",X"3E",X"FE",X"FE",X"FE",
		X"1F",X"3F",X"7B",X"00",X"00",X"00",X"00",X"00",X"FE",X"B4",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7B",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"B4",
		X"1F",X"07",X"03",X"00",X"04",X"02",X"01",X"00",X"FE",X"FE",X"FE",X"FE",X"3E",X"06",X"77",X"F5",
		X"54",X"50",X"80",X"F0",X"DE",X"AF",X"DF",X"7D",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",
		X"1B",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"9E",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"9E",
		X"1B",X"7D",X"DF",X"AF",X"DE",X"F0",X"80",X"50",X"F0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"04",X"00",X"03",X"07",X"F5",X"F5",X"77",X"06",X"3E",X"FE",X"FE",X"FE",
		X"0F",X"1F",X"3F",X"7E",X"7F",X"6F",X"7F",X"7C",X"FE",X"FE",X"FE",X"FE",X"DC",X"F8",X"F8",X"00",
		X"00",X"7C",X"7F",X"6F",X"7F",X"7E",X"3F",X"1F",X"00",X"00",X"F8",X"F8",X"DC",X"FE",X"FE",X"FE",
		X"0F",X"07",X"03",X"00",X"04",X"02",X"01",X"00",X"FE",X"FE",X"FE",X"FE",X"3E",X"06",X"77",X"F5",
		X"54",X"50",X"80",X"F8",X"DE",X"EF",X"BF",X"BD",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",
		X"FF",X"77",X"3F",X"3E",X"1C",X"00",X"00",X"00",X"C0",X"E0",X"30",X"1E",X"0E",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"3F",X"77",X"00",X"00",X"00",X"0E",X"0E",X"1E",X"30",X"E0",
		X"FF",X"BD",X"BF",X"EF",X"DE",X"F8",X"80",X"50",X"C0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"62",X"56",X"50",X"33",X"10",X"1B",X"00",
		X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"8C",X"D4",X"14",X"98",X"10",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"18",X"0B",X"08",X"13",X"10",X"40",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",
		X"A0",X"30",X"A0",X"20",X"90",X"10",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"07",X"01",X"05",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"02",X"07",X"00",X"00",X"03",X"01",X"00",X"A2",X"A2",X"B6",X"D0",X"F3",X"9C",X"FF",X"04",
		X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"07",X"00",X"40",X"C0",X"C0",X"00",X"40",X"00",X"C0",
		X"8A",X"8A",X"DB",X"16",X"9E",X"73",X"FF",X"40",X"00",X"80",X"C0",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"7F",X"F8",X"DB",X"F8",X"F3",X"70",X"B0",X"20",
		X"03",X"01",X"01",X"03",X"06",X"02",X"06",X"00",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"3E",X"B6",X"3F",X"9E",X"1C",X"1A",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"C0",X"80",X"C0",X"00",
		X"00",X"F8",X"8C",X"AE",X"8F",X"FF",X"47",X"4F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"7F",X"47",X"57",X"47",X"7F",X"1F",X"0F",X"00",X"E2",X"E2",X"F6",X"F0",X"F3",X"FC",X"FF",X"04",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"00",X"3E",X"62",X"EA",X"E2",X"FE",X"C4",X"E4",
		X"8F",X"8F",X"DF",X"1F",X"9F",X"7F",X"FF",X"40",X"FC",X"C4",X"D4",X"C4",X"FC",X"F0",X"E0",X"00",
		X"01",X"03",X"0F",X"18",X"1A",X"18",X"0E",X"06",X"FF",X"F8",X"FB",X"F8",X"FB",X"30",X"B0",X"20",
		X"03",X"03",X"06",X"0C",X"38",X"28",X"38",X"00",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"BF",X"3E",X"BE",X"18",X"1A",X"08",X"00",X"80",X"E0",X"30",X"B0",X"30",X"E0",X"C0",
		X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"60",X"38",X"28",X"38",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"02",X"03",X"00",X"00",X"00",X"3F",X"3F",X"21",X"21",X"E3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"01",X"01",X"01",X"01",X"00",X"00",X"1B",X"F2",X"FD",X"11",X"11",X"FD",X"01",X"0D",X"CD",X"41",
		X"03",X"03",X"02",X"02",X"03",X"00",X"03",X"00",X"03",X"01",X"01",X"3F",X"FF",X"00",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"05",
		X"FD",X"FF",X"FC",X"FC",X"FC",X"CC",X"84",X"84",X"C0",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",
		X"12",X"1E",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"41",X"CD",X"DD",X"3D",X"FD",X"FD",X"FF",X"FD",
		X"00",X"03",X"00",X"03",X"03",X"00",X"00",X"03",X"00",X"FF",X"C0",X"00",X"FF",X"3F",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"19",X"11",X"31",X"21",X"21",X"40",X"40",
		X"CC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"FD",X"3D",X"1D",X"4D",X"61",X"7F",X"FF",
		X"02",X"82",X"82",X"43",X"40",X"40",X"23",X"22",X"3F",X"03",X"03",X"FF",X"00",X"3F",X"E0",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"4F",X"47",X"47",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"01",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F0",X"F0",X"C0",
		X"22",X"23",X"20",X"23",X"22",X"23",X"22",X"23",X"3F",X"FF",X"00",X"00",X"3F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"23",X"21",X"30",X"10",X"18",X"08",X"0C",
		X"FF",X"FF",X"FF",X"7C",X"7C",X"7C",X"7C",X"3C",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"7F",X"7F",
		X"FF",X"FC",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"0D",X"1D",X"3D",X"FD",X"FD",
		X"20",X"23",X"43",X"42",X"42",X"C3",X"80",X"02",X"00",X"03",X"01",X"01",X"3F",X"FF",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"24",X"24",X"DC",X"FC",X"3C",X"3C",X"1F",X"05",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"0E",X"FD",X"FF",X"FD",X"FD",X"3D",X"7D",X"8D",X"00",
		X"02",X"02",X"02",X"03",X"00",X"00",X"00",X"00",X"21",X"21",X"3F",X"FF",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"02",X"02",X"02",X"02",X"03",X"FF",X"3F",X"00",X"21",X"21",X"21",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"3F",X"3E",X"3C",X"3C",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"7C",X"7C",X"3C",X"3C",X"3C",
		X"3C",X"3C",X"3C",X"3E",X"1F",X"1F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"C3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"3C",X"7C",X"7C",X"7C",X"FC",X"F8",X"F8",X"F0",
		X"07",X"01",X"00",X"00",X"00",X"00",X"38",X"3C",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"1C",X"3C",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"18",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"3C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"0C",
		X"1F",X"18",X"00",X"00",X"00",X"00",X"00",X"31",X"FF",X"0F",X"1F",X"3F",X"7F",X"FF",X"FE",X"FC",
		X"F8",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"0C",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0C",X"FC",X"FC",X"FC",X"FC",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0F",X"1F",X"3F",X"3E",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0C",X"FC",X"FC",X"FC",X"FC",
		X"3C",X"38",X"38",X"38",X"38",X"38",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"F8",X"70",X"70",X"70",X"70",X"70",X"F8",X"FC",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"30",X"38",X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"03",X"3F",X"FF",X"FF",X"E0",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"7C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1E",X"3E",X"3E",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"80",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1C",X"00",X"1C",X"3C",X"FC",X"FC",X"FC",X"FC",X"3C",X"1C",
		X"3E",X"3E",X"3E",X"3E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",
		X"3E",X"3C",X"38",X"38",X"38",X"38",X"38",X"3C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"1C",X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",
		X"3E",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"F8",X"00",X"00",
		X"00",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"1C",X"7C",X"FC",X"FC",X"FC",X"78",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"00",X"00",X"00",X"FC",X"FE",X"FE",X"FE",X"FF",
		X"00",X"00",X"00",X"03",X"1F",X"3F",X"7F",X"F8",X"00",X"00",X"00",X"80",X"F8",X"FC",X"FC",X"7C",
		X"0F",X"1E",X"1C",X"1C",X"1C",X"3C",X"38",X"38",X"1F",X"0F",X"03",X"03",X"01",X"01",X"01",X"03",
		X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"1C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"38",X"3C",X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"07",X"1F",X"FF",X"FF",X"FE",X"C0",X"00",X"00",
		X"E0",X"F8",X"FF",X"FF",X"03",X"00",X"00",X"00",X"1C",X"3C",X"FC",X"FC",X"FC",X"1C",X"00",X"00",
		X"46",X"EB",X"91",X"91",X"81",X"81",X"42",X"00",X"6E",X"91",X"91",X"91",X"91",X"91",X"6E",X"00",
		X"7E",X"91",X"91",X"91",X"91",X"91",X"61",X"00",X"FF",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"C3",X"A5",X"A5",X"A5",X"BD",X"C3",X"7E",X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"00",X"F0",X"F8",X"38",X"18",X"18",
		X"18",X"18",X"38",X"F8",X"F0",X"00",X"00",X"00",X"18",X"18",X"1C",X"1F",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"1C",X"18",X"18",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"02",X"0B",X"1F",X"17",X"37",X"37",X"FB",X"FB",
		X"C0",X"80",X"40",X"40",X"C0",X"EF",X"FE",X"7D",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",
		X"0F",X"1F",X"1B",X"1D",X"1E",X"1F",X"FE",X"3D",X"FA",X"6D",X"73",X"BB",X"BD",X"3D",X"CE",X"F7",
		X"FB",X"F7",X"EF",X"DF",X"DF",X"BC",X"B3",X"CF",X"C0",X"C0",X"E0",X"F8",X"0C",X"F8",X"FF",X"FC",
		X"EF",X"FF",X"1F",X"3E",X"39",X"27",X"3F",X"0F",X"F8",X"E6",X"9F",X"7D",X"FD",X"FA",X"EB",X"D7",
		X"7F",X"7F",X"CF",X"E0",X"F6",X"F3",X"79",X"B8",X"E7",X"FB",X"80",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"75",X"6E",X"2F",X"2F",X"3E",X"12",X"01",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"C0",X"80",X"70",X"3C",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"FF",
		X"E7",X"DB",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"BD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F1",X"E0",X"D8",X"D0",X"A0",X"BB",X"DC",X"C0",X"00",X"00",X"00",X"00",X"00",X"7F",X"FC",
		X"67",X"7F",X"C0",X"E0",X"F0",X"F0",X"78",X"B8",X"E7",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FB",X"3E",X"FA",X"6D",X"73",X"3B",X"3D",X"3D",X"AE",X"7F",
		X"E7",X"FB",X"00",X"00",X"00",X"00",X"03",X"03",X"F8",X"F6",X"1F",X"3D",X"FD",X"FA",X"EB",X"D7",
		X"02",X"03",X"03",X"03",X"03",X"01",X"01",X"03",X"C0",X"80",X"40",X"40",X"C0",X"C0",X"C0",X"80",
		X"03",X"43",X"63",X"BB",X"BD",X"3D",X"CE",X"F7",X"41",X"47",X"E7",X"DF",X"DF",X"BC",X"B3",X"CF",
		X"F8",X"E6",X"9F",X"7D",X"FF",X"C9",X"C2",X"02",X"7F",X"7F",X"CF",X"E0",X"B0",X"B0",X"C0",X"C0",
		X"01",X"03",X"03",X"03",X"01",X"02",X"02",X"01",X"C0",X"40",X"40",X"C0",X"C0",X"C0",X"C0",X"80",
		X"01",X"03",X"07",X"0F",X"0D",X"3D",X"B3",X"7C",X"C0",X"80",X"40",X"00",X"80",X"00",X"00",X"00",
		X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"E7",X"3B",X"0B",X"0F",X"05",X"02",X"02",X"00",X"00",X"00",X"80",X"00",X"80",X"C0",X"C0",
		X"01",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"C0",X"80",X"60",X"70",X"F0",X"BC",X"DB",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1C",
		X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"67",X"5F",X"FC",X"F8",X"A0",X"A0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AD",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"7C",
		X"FF",X"F3",X"05",X"03",X"03",X"01",X"02",X"02",X"E7",X"DF",X"E0",X"40",X"80",X"80",X"C0",X"C0",
		X"01",X"03",X"03",X"03",X"03",X"07",X"AF",X"7E",X"C0",X"80",X"40",X"40",X"C0",X"E0",X"FB",X"7C",
		X"FF",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"03",X"03",X"07",X"AE",X"7E",X"C0",X"80",X"40",X"40",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"F3",X"05",X"03",X"03",X"01",X"02",X"02",X"C0",X"C0",X"C0",X"40",X"80",X"80",X"C0",X"C0",
		X"01",X"03",X"03",X"03",X"03",X"03",X"02",X"02",X"C0",X"80",X"40",X"40",X"C0",X"E0",X"FB",X"FC",
		X"03",X"03",X"03",X"03",X"03",X"01",X"02",X"02",X"E7",X"DF",X"E0",X"40",X"80",X"80",X"C0",X"C0",
		X"01",X"03",X"03",X"03",X"03",X"06",X"AE",X"7D",X"C0",X"80",X"40",X"40",X"C0",X"E0",X"BB",X"FC",
		X"FF",X"F3",X"05",X"03",X"03",X"01",X"02",X"02",X"E7",X"DF",X"E0",X"40",X"80",X"80",X"C0",X"C0",
		X"E0",X"C1",X"83",X"02",X"01",X"0C",X"0D",X"4B",X"00",X"C0",X"70",X"DC",X"B6",X"EF",X"FF",X"FF",
		X"79",X"79",X"4B",X"0B",X"0C",X"00",X"C0",X"E0",X"FF",X"FF",X"FF",X"DE",X"88",X"00",X"00",X"00",
		X"F0",X"90",X"F8",X"58",X"44",X"5C",X"32",X"BE",X"01",X"02",X"04",X"09",X"12",X"24",X"49",X"95",
		X"04",X"09",X"09",X"15",X"15",X"25",X"48",X"93",X"00",X"FF",X"E8",X"CF",X"E8",X"FF",X"00",X"FF",
		X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"49",X"24",X"12",X"09",X"04",X"02",X"01",
		X"93",X"48",X"25",X"15",X"15",X"09",X"09",X"04",X"FF",X"00",X"FF",X"E8",X"CF",X"E8",X"FF",X"00",
		X"03",X"03",X"01",X"FF",X"03",X"03",X"01",X"02",X"40",X"40",X"C0",X"FF",X"40",X"40",X"80",X"C0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"03",X"03",X"01",X"02",
		X"40",X"40",X"C0",X"80",X"40",X"40",X"80",X"C0",X"02",X"01",X"03",X"03",X"03",X"01",X"01",X"02",
		X"C0",X"C0",X"80",X"40",X"40",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"3E",X"3F",X"3E",X"1C",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"3F",X"0F",X"03",
		X"C0",X"F0",X"FC",X"FF",X"FF",X"FC",X"F0",X"C0",X"FF",X"FF",X"7E",X"7E",X"3C",X"3C",X"18",X"18",
		X"18",X"18",X"3C",X"3C",X"7E",X"7E",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"FF",X"FF",X"18",X"18",X"18",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"08",X"08",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"08",X"08",
		X"10",X"10",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"30",X"10",X"10",
		X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
