library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bgchip_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bgchip_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F3",X"F1",X"E1",X"F3",X"F3",X"F1",X"F1",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"EF",X"FF",X"7F",X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"C3",X"E1",X"E1",X"C3",X"C3",X"E1",X"E1",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"68",X"18",X"78",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"78",X"78",X"78",X"69",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"02",X"0A",X"0E",X"00",X"22",X"77",X"FF",X"22",X"27",X"2F",X"2F",
		X"0E",X"08",X"0A",X"0A",X"0E",X"0E",X"00",X"00",X"3C",X"3C",X"3C",X"E1",X"E3",X"26",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"68",X"18",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"18",X"78",X"78",X"78",X"69",X"0F",X"0F",X"0F",X"01",X"07",X"07",X"07",X"03",X"03",X"01",X"00",
		X"00",X"88",X"CC",X"66",X"EE",X"EE",X"EE",X"2A",X"33",X"11",X"C0",X"C0",X"C4",X"7F",X"4F",X"4F",
		X"08",X"08",X"0A",X"0E",X"0E",X"0E",X"0A",X"00",X"69",X"69",X"69",X"4B",X"C3",X"C3",X"0F",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"A0",X"A0",X"0E",X"08",X"00",X"00",X"00",
		X"F0",X"E0",X"E0",X"0F",X"0F",X"0E",X"0E",X"00",X"0F",X"1E",X"1E",X"0F",X"07",X"03",X"00",X"00",
		X"00",X"88",X"CC",X"66",X"33",X"11",X"C0",X"C0",X"00",X"FF",X"77",X"7F",X"2E",X"2E",X"FF",X"1E",
		X"00",X"0C",X"08",X"0F",X"0F",X"78",X"F0",X"0F",X"00",X"07",X"03",X"07",X"07",X"0F",X"3C",X"34",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1E",X"1F",X"17",X"1F",X"1F",X"17",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"3F",X"3F",X"3E",X"3F",X"37",X"3F",X"3F",X"37",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"7F",X"7F",X"7E",X"7F",X"77",X"7F",X"7F",X"77",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"1F",X"1D",X"1F",X"1F",X"1F",X"1F",X"17",X"1F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"3F",X"3D",X"3F",X"3F",X"3F",X"3F",X"37",X"3F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"7F",X"7D",X"7F",X"7F",X"7F",X"7F",X"77",X"7F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1E",X"1F",X"17",X"1F",X"1F",X"17",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"3F",X"3F",X"3E",X"3F",X"37",X"3F",X"3F",X"37",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"7F",X"7F",X"7E",X"7F",X"77",X"7F",X"7F",X"77",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"1F",X"1D",X"1F",X"1F",X"1F",X"1F",X"17",X"1F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"3F",X"3D",X"3F",X"3F",X"3F",X"3F",X"37",X"3F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"7F",X"7D",X"7F",X"7F",X"7F",X"7F",X"77",X"7F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1E",X"1F",X"17",X"1F",X"1F",X"17",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"3F",X"3F",X"3E",X"3F",X"37",X"3F",X"3F",X"37",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"7F",X"7F",X"7E",X"7F",X"77",X"7F",X"7F",X"77",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"1F",X"1D",X"1F",X"1F",X"1F",X"1F",X"17",X"1F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"3F",X"3D",X"3F",X"3F",X"3F",X"3F",X"37",X"3F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"7F",X"7D",X"7F",X"7F",X"7F",X"7F",X"77",X"7F",
		X"FF",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"C3",X"E1",X"E1",X"C3",X"C3",X"E1",X"E1",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"B0",X"F0",X"4F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"90",X"F0",X"CF",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"90",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"10",X"F0",X"CF",X"0F",X"70",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"B0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"B0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"B0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"90",X"F0",X"4F",X"0F",X"F0",X"F0",X"EF",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"10",X"F0",X"EF",X"0F",X"70",X"F0",X"FF",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"10",X"F0",X"FF",X"0F",X"70",X"F0",X"FF",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"30",X"F0",X"EF",X"0F",X"30",X"F0",X"EF",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"CF",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"B0",X"F0",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
