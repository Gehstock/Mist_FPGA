library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sp_graphx is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sp_graphx is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"CC",X"EE",X"FF",X"BB",X"99",X"18",X"19",X"11",X"1D",X"3F",X"BF",X"FF",X"DF",X"CF",X"E7",
		X"00",X"06",X"8E",X"BF",X"FF",X"7F",X"7E",X"FD",X"22",X"66",X"EE",X"EE",X"AA",X"22",X"02",X"02",
		X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"77",X"33",X"33",X"33",X"33",X"11",X"11",X"11",
		X"DD",X"89",X"89",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"33",X"33",X"22",X"02",X"00",X"00",X"00",X"00",X"8B",X"8B",X"EF",X"77",X"E7",X"EB",
		X"00",X"00",X"44",X"CF",X"CF",X"DF",X"FF",X"7F",X"00",X"00",X"00",X"11",X"33",X"EE",X"EE",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"3B",X"33",X"77",X"77",X"22",X"22",X"22",
		X"FE",X"EE",X"AA",X"02",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"44",X"CC",X"CC",X"CD",X"EF",X"77",X"77",X"DF",
		X"00",X"00",X"00",X"2A",X"EE",X"EF",X"CF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"C7",X"77",X"FF",X"FF",X"CC",X"88",X"00",X"00",
		X"FF",X"FF",X"EA",X"04",X"00",X"00",X"00",X"00",X"EE",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"11",X"33",X"77",X"3B",X"33",X"77",X"FB",X"23",
		X"00",X"00",X"00",X"0C",X"9D",X"EE",X"EF",X"FF",X"00",X"00",X"00",X"88",X"00",X"00",X"08",X"08",
		X"00",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"23",X"77",X"EE",X"CC",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"62",X"44",X"09",X"00",X"00",X"00",X"FF",X"EE",X"44",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"13",X"15",X"33",X"77",X"7B",X"77",
		X"CC",X"88",X"88",X"88",X"8E",X"BF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"08",
		X"00",X"00",X"11",X"33",X"66",X"00",X"00",X"00",X"EF",X"EF",X"FF",X"DC",X"01",X"00",X"00",X"00",
		X"EF",X"7F",X"FF",X"99",X"00",X"01",X"00",X"00",X"08",X"00",X"FF",X"EE",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"10",X"7F",X"33",X"77",
		X"11",X"77",X"EE",X"66",X"EF",X"CF",X"FF",X"7F",X"88",X"00",X"00",X"00",X"08",X"08",X"CC",X"88",
		X"11",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"EF",X"FF",X"88",X"13",X"00",X"00",X"00",X"00",
		X"2F",X"FF",X"F7",X"D9",X"00",X"13",X"00",X"00",X"0C",X"0C",X"00",X"CC",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"17",X"00",X"11",X"FF",
		X"00",X"3F",X"00",X"11",X"FB",X"F7",X"FF",X"9F",X"00",X"FF",X"EE",X"CC",X"88",X"8E",X"0E",X"CC",
		X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"11",X"00",X"17",X"00",X"00",X"00",
		X"3F",X"9F",X"FF",X"F7",X"FB",X"11",X"00",X"3F",X"FF",X"CC",X"0E",X"8E",X"88",X"CC",X"EE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"17",X"00",X"11",X"FF",
		X"00",X"3F",X"00",X"11",X"FB",X"F7",X"FF",X"9F",X"00",X"FF",X"EE",X"CC",X"88",X"8E",X"0E",X"CC",
		X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"11",X"00",X"17",X"00",X"00",X"00",
		X"3F",X"9F",X"FF",X"F7",X"FB",X"11",X"00",X"3F",X"FF",X"CC",X"0E",X"8E",X"88",X"CC",X"EE",X"FF",
		X"30",X"70",X"43",X"43",X"52",X"61",X"21",X"30",X"00",X"80",X"80",X"80",X"80",X"81",X"C1",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"04",X"14",X"FE",X"60",X"F0",X"96",X"96",X"D2",X"B4",X"A4",X"E0",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F3",X"73",X"30",X"43",X"C3",X"10",X"10",
		X"FE",X"FE",X"F6",X"E0",X"96",X"96",X"40",X"40",X"F0",X"C0",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"30",X"70",X"30",X"00",X"30",X"70",X"E0",X"80",X"81",X"A3",X"F3",
		X"80",X"A0",X"10",X"10",X"00",X"14",X"04",X"CC",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",
		X"10",X"10",X"00",X"10",X"30",X"00",X"00",X"00",X"F7",X"F7",X"72",X"B4",X"2D",X"61",X"10",X"00",
		X"EE",X"FC",X"FC",X"F0",X"08",X"48",X"20",X"00",X"C0",X"C0",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"10",X"10",X"70",X"30",X"40",X"E0",X"E0",X"2C",X"48",X"48",X"C0",X"C6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"2C",
		X"10",X"00",X"10",X"61",X"01",X"10",X"00",X"00",X"F7",X"FF",X"F7",X"F3",X"A4",X"96",X"90",X"00",
		X"18",X"F8",X"F8",X"F0",X"70",X"00",X"00",X"00",X"A4",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"00",X"10",X"30",X"F0",X"E0",X"D1",X"F3",X"F7",
		X"00",X"E0",X"F0",X"80",X"00",X"0C",X"8A",X"CE",X"00",X"00",X"80",X"40",X"40",X"60",X"60",X"E0",
		X"60",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"F7",X"79",X"79",X"16",X"86",X"10",X"10",X"00",
		X"EE",X"DC",X"F8",X"F0",X"60",X"00",X"00",X"00",X"E0",X"C0",X"80",X"80",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"10",X"21",X"70",X"F0",X"E0",X"E0",X"E7",
		X"00",X"E0",X"68",X"68",X"80",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"12",X"03",X"70",X"21",X"00",X"00",X"00",X"FF",X"FF",X"F7",X"F2",X"58",X"80",X"80",X"00",
		X"00",X"08",X"F8",X"C3",X"F0",X"C0",X"40",X"00",X"00",X"E0",X"78",X"68",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"03",X"00",X"40",X"30",X"70",X"E0",X"F1",X"F7",X"F7",
		X"00",X"00",X"F0",X"F0",X"20",X"00",X"8E",X"88",X"00",X"00",X"00",X"80",X"C0",X"20",X"00",X"30",
		X"43",X"30",X"21",X"01",X"10",X"10",X"00",X"00",X"F3",X"F7",X"7B",X"B0",X"B0",X"00",X"00",X"00",
		X"8E",X"CC",X"80",X"F0",X"F0",X"E0",X"40",X"00",X"60",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"30",X"03",X"C3",X"30",X"10",X"10",X"30",X"30",X"70",X"F7",X"F7",X"F3",
		X"30",X"E1",X"96",X"F0",X"C0",X"88",X"8E",X"88",X"E0",X"3C",X"3C",X"E0",X"00",X"00",X"00",X"00",
		X"C3",X"03",X"30",X"20",X"00",X"00",X"00",X"00",X"F7",X"F7",X"70",X"30",X"30",X"10",X"10",X"00",
		X"8E",X"88",X"C0",X"F0",X"96",X"E1",X"30",X"00",X"00",X"00",X"00",X"E0",X"3C",X"3C",X"E0",X"00",
		X"00",X"00",X"00",X"20",X"30",X"03",X"43",X"30",X"10",X"10",X"30",X"70",X"70",X"F7",X"F7",X"F3",
		X"00",X"80",X"F0",X"F0",X"10",X"88",X"8E",X"88",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"00",
		X"43",X"03",X"30",X"20",X"00",X"00",X"00",X"00",X"F7",X"F7",X"70",X"70",X"30",X"10",X"10",X"00",
		X"8E",X"88",X"10",X"F0",X"F0",X"80",X"00",X"00",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"00",X"00",X"00",X"44",X"DC",X"EF",X"FE",X"FE",
		X"00",X"00",X"00",X"11",X"D1",X"3F",X"F3",X"F3",X"00",X"00",X"00",X"00",X"CC",X"EE",X"CC",X"88",
		X"11",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"EF",X"8B",X"9B",X"98",X"98",X"00",X"00",X"00",
		X"3F",X"0E",X"4E",X"40",X"40",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"EE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"CC",X"CC",X"FE",X"FE",X"47",X"CF",
		X"00",X"00",X"00",X"80",X"D1",X"F3",X"3F",X"7F",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",
		X"11",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"70",X"7C",X"53",X"10",X"00",X"00",X"00",X"00",
		X"C4",X"F3",X"19",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"77",X"77",X"00",X"00",X"11",X"FF",X"FF",X"FF",X"FE",X"67",
		X"00",X"00",X"00",X"20",X"68",X"2C",X"97",X"F3",X"00",X"00",X"00",X"00",X"00",X"88",X"EE",X"CC",
		X"77",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"47",X"51",X"90",X"20",X"00",X"00",X"00",
		X"7F",X"7F",X"19",X"33",X"77",X"55",X"00",X"00",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"11",X"33",X"33",X"99",X"FE",X"12",
		X"00",X"00",X"88",X"88",X"70",X"3C",X"96",X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"47",X"A3",X"41",X"00",X"11",X"00",X"00",
		X"F3",X"5D",X"44",X"66",X"CC",X"88",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"11",X"33",X"00",X"00",X"11",X"11",X"FF",X"FF",X"BB",X"33",X"07",
		X"00",X"44",X"CC",X"EE",X"CC",X"BC",X"96",X"C3",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"03",X"63",X"80",X"11",X"33",X"11",X"00",
		X"7B",X"FF",X"FF",X"77",X"EE",X"CC",X"CC",X"00",X"CC",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"AA",X"31",X"34",
		X"00",X"00",X"00",X"33",X"FF",X"EE",X"BC",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F4",X"34",X"72",X"02",X"11",X"EE",X"00",X"00",
		X"3C",X"3F",X"FF",X"BB",X"88",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"EE",X"FF",X"FF",X"11",X"17",X"C7",X"07",
		X"00",X"22",X"77",X"FF",X"FF",X"EE",X"D2",X"D2",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"C7",X"17",X"11",X"FF",X"FF",X"EE",X"00",X"00",
		X"D2",X"EE",X"FF",X"FF",X"77",X"22",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"17",X"C7",X"07",
		X"00",X"00",X"00",X"77",X"77",X"EE",X"D2",X"D2",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"80",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"C7",X"17",X"11",X"FF",X"00",X"00",X"00",X"00",
		X"D2",X"EE",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"80",X"81",X"D1",X"C1",X"E1",
		X"00",X"00",X"00",X"08",X"0C",X"DC",X"1C",X"3C",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"71",X"33",X"43",X"A3",X"00",X"00",X"00",X"00",
		X"FC",X"EE",X"9E",X"AE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"61",X"61",
		X"00",X"00",X"00",X"04",X"0E",X"EE",X"0E",X"1C",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"33",X"F3",X"57",X"13",X"11",X"00",X"00",X"00",
		X"FC",X"FC",X"0C",X"6C",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"E0",X"D1",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"8E",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"10",X"60",X"00",X"00",X"00",X"00",X"00",X"C3",X"77",X"3F",X"BF",X"47",X"55",X"00",X"00",
		X"1C",X"78",X"F8",X"C8",X"80",X"40",X"40",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"30",X"30",X"31",X"61",X"F7",
		X"00",X"80",X"C0",X"80",X"85",X"CE",X"6F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"3F",X"47",X"9B",X"00",X"10",X"00",X"00",
		X"BE",X"F8",X"C8",X"80",X"80",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"10",X"00",X"30",X"70",X"70",X"70",X"60",X"E1",X"CF",
		X"00",X"80",X"80",X"00",X"00",X"04",X"8E",X"CE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"23",X"01",X"33",X"00",X"00",X"00",X"00",X"00",X"EF",X"EF",X"3E",X"9C",X"20",X"40",X"40",X"00",
		X"4C",X"A0",X"F0",X"F0",X"10",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"B0",X"BF",X"3F",
		X"00",X"00",X"70",X"F0",X"80",X"27",X"2F",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"64",X"20",X"40",X"00",X"00",X"00",
		X"0C",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"80",X"50",X"BE",X"3F",X"FF",
		X"00",X"30",X"70",X"F0",X"E0",X"80",X"2F",X"2F",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"3F",X"BE",X"50",X"80",X"00",X"00",X"00",X"00",
		X"2F",X"80",X"E0",X"F0",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"80",X"50",X"BE",X"3F",X"FF",
		X"00",X"00",X"00",X"70",X"F0",X"80",X"2F",X"2F",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"08",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"3F",X"BE",X"50",X"80",X"00",X"00",X"00",X"00",
		X"2F",X"80",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"46",
		X"00",X"00",X"00",X"00",X"01",X"66",X"22",X"88",X"00",X"33",X"44",X"8A",X"11",X"76",X"80",X"00",
		X"00",X"11",X"11",X"02",X"11",X"00",X"00",X"00",X"8A",X"10",X"08",X"08",X"CC",X"88",X"44",X"88",
		X"CC",X"A8",X"00",X"00",X"00",X"00",X"10",X"F0",X"00",X"00",X"00",X"70",X"00",X"10",X"F0",X"F0",
		X"00",X"00",X"CC",X"02",X"99",X"11",X"00",X"00",X"00",X"00",X"33",X"0C",X"11",X"06",X"10",X"00",
		X"00",X"00",X"00",X"88",X"44",X"02",X"91",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"10",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"E0",X"E0",X"C0",X"F0",
		X"31",X"31",X"01",X"01",X"22",X"44",X"11",X"20",X"08",X"08",X"8C",X"8C",X"88",X"88",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"88",X"04",X"04",X"88",X"A8",X"44",X"54",X"33",
		X"10",X"00",X"00",X"00",X"00",X"CC",X"03",X"91",X"F0",X"10",X"00",X"70",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"44",X"13",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"70",X"F0",X"10",X"00",X"F0",X"00",X"C0",X"E0",X"E0",X"80",X"C0",X"E0",X"F0",X"11",
		X"44",X"44",X"01",X"00",X"20",X"55",X"55",X"2A",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",
		X"00",X"CE",X"02",X"CE",X"02",X"11",X"00",X"00",X"20",X"FF",X"37",X"26",X"04",X"88",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"22",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"89",X"CD",X"03",
		X"00",X"00",X"22",X"33",X"22",X"00",X"11",X"77",X"00",X"00",X"88",X"88",X"04",X"00",X"CC",X"FF",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"44",X"44",X"91",X"11",X"11",X"77",X"FF",X"BB",
		X"66",X"DD",X"FE",X"FD",X"CF",X"46",X"CF",X"CD",X"77",X"BB",X"EE",X"8E",X"0D",X"0D",X"01",X"07",
		X"00",X"00",X"00",X"00",X"00",X"77",X"FF",X"DD",X"00",X"00",X"00",X"80",X"22",X"88",X"AA",X"66",
		X"00",X"00",X"00",X"00",X"00",X"01",X"2A",X"0C",X"00",X"00",X"44",X"44",X"88",X"00",X"00",X"00",
		X"AA",X"EF",X"1E",X"07",X"07",X"02",X"40",X"0E",X"FF",X"19",X"6E",X"1F",X"35",X"1F",X"3F",X"33",
		X"00",X"00",X"EE",X"FF",X"BB",X"66",X"EE",X"CC",X"00",X"88",X"44",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"11",X"11",X"00",X"00",X"00",X"D9",X"BB",X"DD",X"EC",X"CD",X"FF",X"33",X"00",
		X"47",X"8F",X"CE",X"CE",X"CF",X"8B",X"66",X"FF",X"29",X"05",X"08",X"26",X"0E",X"06",X"1D",X"FF",
		X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"00",X"40",X"22",X"DD",X"99",X"00",X"00",X"00",X"00",
		X"66",X"33",X"33",X"11",X"40",X"22",X"22",X"00",X"FF",X"66",X"99",X"FF",X"EE",X"00",X"00",X"00",
		X"84",X"0A",X"01",X"0A",X"0F",X"0D",X"1F",X"C2",X"3F",X"1F",X"35",X"17",X"33",X"3F",X"FF",X"77",
		X"BB",X"FF",X"66",X"BB",X"BB",X"66",X"CC",X"88",X"00",X"44",X"66",X"44",X"66",X"11",X"00",X"00",
		X"FF",X"BB",X"77",X"FF",X"EE",X"00",X"00",X"00",X"AA",X"CC",X"CC",X"88",X"22",X"44",X"00",X"00",
		X"33",X"04",X"A8",X"98",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"00",X"00",
		X"88",X"54",X"22",X"22",X"00",X"33",X"67",X"CF",X"00",X"00",X"91",X"11",X"FF",X"CC",X"0B",X"07",
		X"22",X"FF",X"DD",X"2A",X"0F",X"3F",X"07",X"0F",X"EE",X"FF",X"33",X"1D",X"0E",X"8F",X"0F",X"03",
		X"CE",X"CD",X"EE",X"45",X"EE",X"EF",X"EF",X"FF",X"1E",X"2F",X"4F",X"0F",X"0F",X"07",X"0E",X"6D",
		X"CE",X"87",X"0D",X"0E",X"8F",X"0F",X"01",X"0E",X"0D",X"8F",X"0F",X"06",X"00",X"04",X"0B",X"01",
		X"00",X"11",X"BB",X"CC",X"FF",X"77",X"1E",X"87",X"A2",X"22",X"CC",X"11",X"99",X"BB",X"7F",X"0C",
		X"00",X"01",X"01",X"CC",X"EE",X"BF",X"3F",X"37",X"11",X"22",X"40",X"08",X"40",X"00",X"00",X"00",
		X"0F",X"1F",X"0B",X"03",X"09",X"08",X"83",X"0E",X"0D",X"0F",X"0F",X"09",X"03",X"06",X"05",X"07",
		X"3B",X"2E",X"B7",X"1F",X"0D",X"0F",X"0F",X"0F",X"00",X"00",X"66",X"FF",X"3F",X"3F",X"37",X"6E",
		X"FF",X"11",X"77",X"FF",X"EE",X"66",X"67",X"67",X"3D",X"1F",X"9B",X"17",X"2F",X"0F",X"07",X"5B",
		X"0F",X"0D",X"1A",X"0F",X"0E",X"0D",X"0F",X"8F",X"07",X"01",X"0A",X"04",X"08",X"13",X"07",X"7F",
		X"33",X"11",X"00",X"11",X"11",X"33",X"44",X"00",X"8F",X"8A",X"23",X"23",X"91",X"00",X"00",X"00",
		X"6F",X"0F",X"07",X"0B",X"8C",X"FF",X"77",X"00",X"0F",X"97",X"6F",X"06",X"3F",X"EE",X"88",X"00",
		X"0C",X"08",X"0B",X"84",X"0A",X"03",X"0B",X"0F",X"01",X"07",X"07",X"1A",X"03",X"0B",X"0E",X"4D",
		X"0B",X"85",X"0D",X"1B",X"1F",X"19",X"66",X"FF",X"AA",X"88",X"88",X"CC",X"CC",X"88",X"00",X"00",
		X"1F",X"2F",X"4B",X"8E",X"77",X"FF",X"00",X"00",X"0F",X"0F",X"0B",X"FF",X"BB",X"00",X"00",X"00",
		X"FF",X"CC",X"CC",X"98",X"00",X"40",X"22",X"00",X"00",X"00",X"88",X"88",X"C8",X"62",X"33",X"11",
		X"00",X"00",X"02",X"13",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"09",X"C1",X"03",
		X"00",X"00",X"02",X"03",X"02",X"00",X"11",X"67",X"00",X"00",X"08",X"80",X"40",X"00",X"0C",X"3F",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"04",X"04",X"89",X"01",X"01",X"17",X"3F",X"3B",
		X"06",X"4D",X"0F",X"7C",X"8F",X"06",X"0F",X"0D",X"07",X"0B",X"0E",X"0E",X"0D",X"0D",X"01",X"25",
		X"00",X"00",X"00",X"00",X"00",X"77",X"0F",X"4D",X"00",X"00",X"00",X"80",X"22",X"08",X"AA",X"06",
		X"00",X"00",X"00",X"00",X"00",X"11",X"0A",X"0C",X"00",X"00",X"04",X"04",X"80",X"00",X"00",X"00",
		X"0A",X"0F",X"0F",X"07",X"07",X"02",X"04",X"0E",X"2F",X"09",X"86",X"0F",X"07",X"0F",X"0F",X"03",
		X"00",X"00",X"6E",X"1F",X"0B",X"26",X"2E",X"0C",X"00",X"88",X"44",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"00",X"01",X"01",X"00",X"00",X"00",X"1D",X"1A",X"4D",X"8E",X"8D",X"0F",X"03",X"00",
		X"07",X"0F",X"0E",X"4A",X"0F",X"0B",X"06",X"0F",X"0B",X"05",X"08",X"06",X"0E",X"06",X"0D",X"0F",
		X"00",X"00",X"00",X"00",X"10",X"22",X"22",X"00",X"04",X"02",X"0D",X"09",X"00",X"00",X"00",X"00",
		X"46",X"03",X"03",X"01",X"04",X"22",X"22",X"00",X"0F",X"06",X"09",X"3E",X"CE",X"00",X"00",X"00",
		X"0C",X"28",X"01",X"0A",X"0F",X"0D",X"0F",X"0E",X"1E",X"2F",X"27",X"07",X"03",X"0F",X"0F",X"17",
		X"0B",X"4F",X"66",X"2B",X"2B",X"06",X"CC",X"88",X"00",X"04",X"06",X"04",X"06",X"01",X"00",X"00",
		X"0F",X"0B",X"27",X"87",X"EE",X"00",X"00",X"00",X"2A",X"0C",X"CC",X"08",X"02",X"04",X"00",X"00",
		X"03",X"04",X"0A",X"09",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"30",X"40",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F1",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"70",X"72",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"CC",X"88",X"77",X"00",X"99",X"AA",
		X"00",X"CC",X"22",X"66",X"CC",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"EE",X"00",X"00",X"FF",X"44",X"00",
		X"22",X"22",X"44",X"00",X"22",X"EE",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",
		X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"00",X"0F",X"04",X"02",X"01",
		X"02",X"0C",X"00",X"08",X"0E",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",
		X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"09",X"0A",X"0A",X"0A",X"0E",
		X"02",X"0C",X"00",X"0C",X"02",X"02",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",
		X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",
		X"02",X"0C",X"00",X"0C",X"02",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"80",X"80",X"70",X"00",X"70",X"80",X"80",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"70",X"80",X"80",X"70",X"00",X"F0",
		X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",X"88",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"99",X"AA",X"AA",X"EE",X"00",X"FF",
		X"CC",X"00",X"CC",X"22",X"22",X"44",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",
		X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"08",X"09",X"05",X"03",X"00",X"0F",
		X"0C",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"12",X"1E",X"00",X"00",X"0F",X"00",X"10",X"76",X"1E",X"1E",
		X"00",X"00",X"0F",X"1E",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"1C",X"1C",X"10",X"10",X"DC",X"FE",
		X"3E",X"1E",X"12",X"10",X"00",X"00",X"00",X"00",X"DE",X"1E",X"1E",X"76",X"10",X"00",X"0F",X"00",
		X"1E",X"FE",X"FE",X"FE",X"FE",X"1E",X"0F",X"00",X"1C",X"FE",X"DC",X"10",X"10",X"1C",X"1C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"70",X"80",X"80",X"70",X"00",X"70",
		X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"88",X"88",X"77",X"00",X"77",
		X"CC",X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"70",X"00",X"60",X"90",X"80",X"80",
		X"20",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"77",X"00",X"88",X"DD",X"AA",X"88",
		X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",
		X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",
		X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"27",X"57",X"88",X"22",X"00",X"00",X"00",
		X"4C",X"4C",X"88",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"44",X"11",X"00",X"00",X"02",X"00",X"A2",X"03",X"AB",X"05",
		X"00",X"00",X"10",X"B8",X"44",X"22",X"1B",X"86",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"44",
		X"00",X"11",X"22",X"10",X"10",X"00",X"00",X"00",X"BC",X"21",X"65",X"81",X"44",X"22",X"00",X"00",
		X"BE",X"3C",X"B4",X"54",X"11",X"04",X"00",X"00",X"88",X"80",X"84",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"22",X"01",X"44",X"38",X"20",X"44",X"11",X"88",X"74",X"00",X"8B",X"00",X"44",X"88",
		X"22",X"10",X"22",X"89",X"01",X"22",X"88",X"00",X"20",X"80",X"00",X"08",X"08",X"11",X"C0",X"00",
		X"00",X"DA",X"01",X"03",X"44",X"00",X"11",X"88",X"22",X"C0",X"00",X"22",X"44",X"10",X"02",X"02",
		X"55",X"00",X"15",X"24",X"C0",X"22",X"00",X"44",X"30",X"20",X"E9",X"40",X"65",X"00",X"88",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"04",X"22",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"22",X"11",X"88",X"44",X"00",X"22",
		X"11",X"04",X"00",X"20",X"11",X"00",X"A8",X"20",X"00",X"C0",X"81",X"22",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"04",X"A2",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"11",X"22",X"22",X"00",X"00",X"00",X"00",X"11",X"02",X"00",X"C0",X"00",X"10",X"04",X"44",
		X"00",X"00",X"60",X"00",X"88",X"01",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"80",X"80",X"00",X"11",X"00",X"22",X"00",
		X"22",X"0C",X"00",X"00",X"60",X"20",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"44",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"44",X"00",X"00",X"00",X"10",X"00",X"22",X"04",X"00",X"00",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"22",X"15",X"30",X"00",X"88",X"44",X"01",
		X"88",X"00",X"11",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"11",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"C0",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"80",X"00",X"00",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"11",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",
		X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"10",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"11",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"01",X"03",X"00",X"00",X"01",X"01",X"0F",X"0F",X"0B",X"03",X"77",
		X"00",X"04",X"0C",X"0E",X"0C",X"7C",X"F6",X"F3",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"33",X"53",X"80",X"01",X"03",X"01",X"00",
		X"CB",X"0F",X"0F",X"07",X"0E",X"0C",X"0C",X"00",X"0C",X"08",X"08",X"08",X"00",X"00",X"00",X"00",
		X"0F",X"0C",X"0C",X"0F",X"0F",X"0C",X"0C",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",
		X"0C",X"0C",X"0C",X"0F",X"07",X"00",X"00",X"07",X"03",X"03",X"03",X"0F",X"0E",X"00",X"00",X"0F",
		X"0C",X"0F",X"07",X"00",X"00",X"0C",X"0C",X"0C",X"03",X"0F",X"0E",X"00",X"00",X"03",X"03",X"03",
		X"00",X"00",X"07",X"0F",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"0E",X"0F",X"03",X"03",X"03",X"03",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"11",X"11",X"51",X"D1",X"D5",X"FF",
		X"00",X"00",X"00",X"00",X"40",X"60",X"74",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"31",X"31",X"20",X"20",X"00",X"00",X"00",X"00",X"EF",X"2F",X"07",X"03",X"01",X"00",X"00",X"00",
		X"FF",X"9F",X"0C",X"08",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"20",X"60",X"F3",X"FF",
		X"00",X"00",X"44",X"44",X"CC",X"98",X"BA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"10",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"17",X"03",X"03",X"01",X"00",X"00",X"00",
		X"7F",X"7F",X"1F",X"0C",X"00",X"00",X"00",X"00",X"C0",X"C8",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"00",X"00",X"00",X"10",X"F0",X"F7",X"FF",X"77",
		X"00",X"00",X"11",X"B3",X"22",X"44",X"DD",X"7F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"3F",X"10",X"10",X"20",X"00",X"00",X"80",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"30",X"20",X"00",X"00",X"00",X"00",X"F0",X"F7",X"FF",X"77",X"37",
		X"00",X"00",X"00",X"C0",X"99",X"AA",X"CC",X"7F",X"00",X"00",X"00",X"88",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"27",X"17",X"07",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"32",X"30",X"60",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"20",X"F0",X"F7",X"77",X"37",X"27",
		X"00",X"00",X"00",X"E0",X"CC",X"99",X"EE",X"4C",X"00",X"00",X"00",X"00",X"CC",X"88",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"03",X"00",X"00",X"10",X"00",X"00",
		X"FE",X"FE",X"FE",X"74",X"E0",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F2",X"77",X"37",X"3F",X"0F",
		X"00",X"00",X"00",X"C0",X"E8",X"CC",X"99",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"1F",X"13",X"11",X"30",X"60",X"00",X"00",
		X"CC",X"FC",X"E8",X"C8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"33",X"13",X"17",X"3F",
		X"00",X"00",X"00",X"80",X"C0",X"E8",X"FC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"3F",X"17",X"13",X"33",X"F0",X"00",X"00",
		X"FF",X"88",X"FC",X"E8",X"C0",X"80",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"3F",
		X"00",X"00",X"CC",X"22",X"11",X"88",X"88",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"3B",X"3B",X"19",X"28",X"20",X"00",X"00",X"00",
		X"8B",X"8B",X"03",X"82",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"66",X"99",X"00",X"00",X"11",X"11",X"3F",
		X"00",X"00",X"00",X"88",X"88",X"88",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"05",X"00",X"00",X"00",X"00",X"00",X"3B",X"33",X"22",X"50",X"50",X"00",X"00",X"00",
		X"8E",X"8B",X"03",X"07",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"19",
		X"00",X"00",X"00",X"00",X"33",X"CC",X"EE",X"CC",X"00",X"00",X"00",X"00",X"88",X"44",X"44",X"00",
		X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"3B",X"33",X"62",X"A0",X"20",X"00",X"00",X"00",
		X"8C",X"8A",X"06",X"06",X"0E",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"0E",X"1D",X"3B",
		X"00",X"00",X"EE",X"11",X"11",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"73",X"A0",X"40",X"01",X"00",X"00",X"00",
		X"CC",X"8A",X"06",X"0E",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"0E",X"0D",X"33",
		X"00",X"00",X"00",X"00",X"00",X"77",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"44",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"F7",X"40",X"81",X"03",X"00",X"01",X"00",
		X"CC",X"04",X"04",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"09",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"00",X"00",X"00",X"00",X"88",X"44",X"44",X"88",
		X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"B3",X"77",X"80",X"01",X"07",X"03",X"06",X"00",
		X"EE",X"88",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"0C",X"07",X"0F",X"00",X"B3",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"B3",X"00",X"0F",X"07",X"0C",X"00",X"00",
		X"FF",X"EE",X"08",X"08",X"11",X"00",X"00",X"00",X"88",X"44",X"44",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"02",X"03",X"03",X"01",X"00",X"00",X"01",X"01",X"01",X"03",X"0F",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"09",X"0F",X"87",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"9E",X"CF",X"67",X"01",X"01",X"00",X"00",
		X"0F",X"2E",X"6E",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"08",X"0D",X"0F",X"3C",
		X"00",X"00",X"08",X"08",X"08",X"0C",X"0C",X"87",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"9E",X"CF",X"DF",X"02",X"02",X"00",X"00",
		X"0F",X"0F",X"6E",X"CC",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0C",X"0C",X"0F",X"0F",X"9E",
		X"00",X"00",X"02",X"02",X"04",X"0C",X"0C",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0C",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"AD",X"8F",X"37",X"19",X"00",X"00",X"00",
		X"0F",X"0F",X"4E",X"CC",X"00",X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"04",X"0E",X"0E",X"0F",X"AD",
		X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"00",X"01",X"00",X"00",X"00",X"1E",X"2D",X"8F",X"4F",X"77",X"00",X"00",X"00",
		X"0C",X"87",X"0F",X"8F",X"88",X"00",X"00",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"CF",X"8F",
		X"00",X"04",X"08",X"08",X"00",X"08",X"0F",X"86",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"11",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"9E",X"AD",X"0F",X"77",X"11",X"00",X"00",X"00",
		X"86",X"0E",X"0F",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"47",X"CF",X"8F",
		X"00",X"00",X"0E",X"0C",X"08",X"08",X"0E",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"0F",X"CF",X"FF",X"00",X"00",X"00",X"00",
		X"86",X"84",X"0E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"67",X"CF",X"8F",
		X"00",X"00",X"00",X"07",X"0E",X"0C",X"0C",X"86",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"8F",X"CF",X"67",X"01",X"00",X"00",X"00",
		X"87",X"86",X"0C",X"0C",X"0E",X"07",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"70",X"F0",X"00",X"00",X"00",X"00",X"00",X"1E",X"F0",X"D0",X"10",X"32",X"66",X"00",X"00",
		X"0F",X"F0",X"70",X"00",X"88",X"CC",X"00",X"00",X"0C",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",
		X"00",X"00",X"40",X"40",X"80",X"80",X"80",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"D0",X"10",X"64",X"DD",X"11",X"00",X"00",
		X"0F",X"C3",X"70",X"10",X"00",X"88",X"00",X"00",X"00",X"0C",X"84",X"C0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"00",X"00",X"00",X"10",X"20",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"D2",X"F0",X"30",X"A8",X"EA",X"22",X"22",X"00",
		X"00",X"0E",X"87",X"E1",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"03",X"E1",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"86",
		X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"00",X"00",X"00",X"00",X"D2",X"21",X"50",X"90",X"CC",X"88",X"00",X"00",
		X"00",X"0C",X"0E",X"86",X"C3",X"E1",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"61",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"08",X"0C",X"86",X"86",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"77",X"10",X"11",X"11",X"00",X"00",X"00",X"70",X"E1",X"30",X"B8",X"10",X"10",X"00",X"00",
		X"00",X"08",X"0C",X"0E",X"84",X"86",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"86",X"C2",X"C3",X"43",X"61",X"21",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"33",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"70",X"90",X"B8",X"30",X"30",X"10",X"10",X"10",
		X"80",X"0C",X"0C",X"0C",X"84",X"84",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"33",X"00",X"40",X"61",X"61",X"61",X"61",X"61",X"21",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"33",X"22",X"00",X"00",X"00",X"00",X"00",X"F0",X"21",X"61",X"61",X"61",X"61",X"61",X"40",
		X"F0",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"77",X"44",X"77",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"11",X"99",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"22",
		X"22",X"22",X"22",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"33",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"88",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"1D",X"0F",X"87",X"E1",
		X"44",X"CC",X"CC",X"CC",X"88",X"3B",X"7F",X"7F",X"00",X"00",X"00",X"33",X"FF",X"EE",X"EE",X"88",
		X"11",X"33",X"77",X"44",X"00",X"00",X"00",X"00",X"F8",X"FD",X"BB",X"33",X"77",X"77",X"66",X"44",
		X"4E",X"8E",X"E8",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"A0",X"10",
		X"00",X"00",X"00",X"03",X"21",X"76",X"77",X"11",X"00",X"00",X"00",X"11",X"1F",X"0F",X"C3",X"E9",
		X"44",X"CC",X"CC",X"CC",X"CC",X"0C",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"77",X"77",X"FF",X"EE",X"EE",X"CC",X"88",
		X"F7",X"B7",X"60",X"10",X"00",X"00",X"00",X"00",X"FF",X"EE",X"00",X"00",X"A0",X"40",X"A0",X"10",
		X"00",X"00",X"11",X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"88",X"DD",X"1F",X"87",X"F0",X"70",
		X"22",X"77",X"FF",X"EE",X"CC",X"88",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"33",X"33",X"22",X"00",X"00",X"FD",X"DD",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"A8",X"40",X"A0",X"10",
		X"00",X"00",X"00",X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"1D",X"0F",X"87",X"E1",
		X"44",X"CC",X"CC",X"CC",X"88",X"3B",X"7F",X"7F",X"00",X"00",X"00",X"33",X"FF",X"EE",X"EE",X"88",
		X"11",X"33",X"77",X"44",X"00",X"00",X"00",X"00",X"F8",X"FD",X"BB",X"33",X"77",X"77",X"66",X"44",
		X"4E",X"8E",X"E8",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"A0",X"10",
		X"00",X"00",X"00",X"03",X"21",X"76",X"77",X"11",X"00",X"00",X"00",X"11",X"1F",X"0F",X"C3",X"E9",
		X"44",X"CC",X"CC",X"CC",X"CC",X"0C",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"77",X"77",X"FF",X"EE",X"EE",X"CC",X"88",
		X"F7",X"B7",X"60",X"10",X"00",X"00",X"00",X"00",X"FF",X"EE",X"00",X"00",X"A0",X"40",X"A0",X"10",
		X"00",X"00",X"11",X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"88",X"DD",X"1F",X"87",X"F0",X"70",
		X"22",X"77",X"FF",X"EE",X"CC",X"88",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"33",X"33",X"22",X"00",X"00",X"FD",X"DD",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"A8",X"40",X"A0",X"10",
		X"00",X"00",X"00",X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"1D",X"0F",X"87",X"E1",
		X"44",X"CC",X"CC",X"CC",X"88",X"3B",X"7F",X"7F",X"00",X"00",X"00",X"33",X"FF",X"EE",X"EE",X"88",
		X"11",X"33",X"77",X"44",X"00",X"00",X"00",X"00",X"F8",X"FD",X"BB",X"33",X"77",X"77",X"66",X"44",
		X"4E",X"8E",X"E8",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"A0",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"60",X"71",X"71",X"71",X"60",X"12",X"12",X"74",X"FC",X"FD",X"B9",X"11",X"71",
		X"08",X"08",X"C4",X"E6",X"F7",X"B3",X"11",X"C0",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"60",X"14",X"10",X"10",X"10",X"10",X"00",X"00",X"F0",X"F1",X"F3",X"E7",X"F3",X"E1",X"E1",X"61",
		X"E0",X"F0",X"F8",X"FC",X"F8",X"F0",X"E0",X"C0",X"C0",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"30",X"30",X"30",X"71",X"60",X"24",X"00",X"00",X"32",X"FE",X"FE",X"30",X"11",X"F1",
		X"4A",X"4A",X"C0",X"E2",X"FB",X"FB",X"33",X"91",X"00",X"00",X"00",X"60",X"60",X"60",X"E8",X"C0",
		X"10",X"30",X"30",X"30",X"30",X"30",X"10",X"00",X"F0",X"F3",X"FF",X"DF",X"F7",X"D2",X"B4",X"34",
		X"C0",X"E0",X"E0",X"E8",X"E0",X"E0",X"C0",X"80",X"C0",X"C0",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"30",X"30",X"70",X"04",X"30",X"C0",X"C0",X"F7",X"F7",X"FF",X"10",X"E0",X"F1",
		X"02",X"12",X"E9",X"F0",X"F5",X"FD",X"D9",X"91",X"00",X"08",X"00",X"00",X"00",X"A8",X"F8",X"E8",
		X"30",X"70",X"F1",X"70",X"70",X"70",X"01",X"00",X"F0",X"FE",X"FF",X"BF",X"7D",X"78",X"F0",X"E0",
		X"D1",X"C0",X"D0",X"E0",X"C1",X"C0",X"80",X"00",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"34",X"00",X"30",X"30",X"70",X"E0",X"F3",X"F7",X"44",X"00",X"E0",
		X"00",X"00",X"00",X"CD",X"F8",X"F0",X"F4",X"F9",X"00",X"00",X"48",X"84",X"08",X"00",X"88",X"88",
		X"70",X"F1",X"F1",X"F1",X"F1",X"D2",X"34",X"30",X"F1",X"FA",X"FC",X"7E",X"FE",X"F0",X"F0",X"E0",
		X"11",X"91",X"B3",X"90",X"B0",X"B0",X"02",X"00",X"B8",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"70",X"00",X"10",X"30",X"F0",X"51",X"80",X"F0",X"F0",
		X"40",X"E0",X"C0",X"EE",X"FF",X"30",X"73",X"F6",X"00",X"00",X"00",X"02",X"A4",X"C3",X"C0",X"C4",
		X"71",X"F0",X"F1",X"C3",X"34",X"30",X"30",X"00",X"FC",X"FE",X"7E",X"FE",X"F4",X"F0",X"E0",X"40",
		X"B9",X"D1",X"D1",X"D1",X"B0",X"B0",X"24",X"00",X"CC",X"CC",X"FC",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"00",X"00",X"34",X"30",X"00",X"E0",X"F0",X"F8",
		X"00",X"70",X"F0",X"C4",X"FF",X"77",X"30",X"B3",X"00",X"80",X"80",X"00",X"00",X"8B",X"F0",X"C3",
		X"F1",X"D3",X"3D",X"70",X"70",X"30",X"00",X"00",X"FE",X"7E",X"FC",X"FC",X"F0",X"E0",X"00",X"00",
		X"FC",X"B1",X"91",X"91",X"32",X"F0",X"68",X"00",X"C0",X"CC",X"88",X"88",X"E0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"F1",X"00",X"00",X"12",X"10",X"E0",X"F0",X"F8",X"FC",
		X"00",X"00",X"F0",X"F0",X"77",X"33",X"91",X"B0",X"00",X"00",X"C0",X"C0",X"00",X"88",X"CC",X"C3",
		X"1F",X"F1",X"F0",X"70",X"30",X"00",X"00",X"00",X"7E",X"FC",X"F8",X"F0",X"E0",X"10",X"12",X"00",
		X"FF",X"B0",X"91",X"33",X"77",X"F0",X"F0",X"00",X"F0",X"C3",X"CC",X"88",X"00",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
