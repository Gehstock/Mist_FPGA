library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity survival_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of survival_prog is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"FC",X"4B",X"21",X"07",X"68",X"11",X"0E",X"69",X"01",X"FD",X"7F",X"75",X"78",X"12",
		X"73",X"79",X"12",X"2A",X"4C",X"00",X"EB",X"21",X"00",X"50",X"75",X"EB",X"22",X"FE",X"4B",X"EB",
		X"D1",X"40",X"49",X"36",X"01",X"E5",X"CD",X"4E",X"01",X"E1",X"75",X"F2",X"4E",X"01",X"E1",X"E9",
		X"78",X"B3",X"CA",X"7B",X"03",X"F2",X"AE",X"00",X"B2",X"2E",X"48",X"20",X"E6",X"80",X"07",X"57",
		X"26",X"00",X"31",X"00",X"4C",X"7A",X"00",X"E9",X"CD",X"8C",X"1F",X"01",X"38",X"00",X"C5",X"3A",
		X"F3",X"43",X"B7",X"C2",X"1D",X"08",X"CD",X"08",X"32",X"3A",X"EC",X"43",X"B7",X"CA",X"7B",X"03",
		X"F5",X"AF",X"32",X"00",X"50",X"32",X"9E",X"43",X"CD",X"62",X"1F",X"CD",X"B3",X"20",X"CD",X"94",
		X"17",X"F1",X"B9",X"D2",X"7E",X"00",X"0E",X"02",X"21",X"A2",X"3B",X"C3",X"52",X"3B",X"F5",X"21",
		X"CB",X"1E",X"0E",X"01",X"C5",X"CD",X"5D",X"02",X"C1",X"F1",X"B8",X"06",X"02",X"DA",X"95",X"00",
		X"06",X"06",X"21",X"E8",X"1E",X"C5",X"CD",X"5D",X"02",X"C1",X"3A",X"00",X"70",X"2F",X"A0",X"C8",
		X"F5",X"CD",X"94",X"17",X"F1",X"3D",X"FE",X"01",X"CA",X"AE",X"00",X"48",X"3E",X"02",X"32",X"F3",
		X"43",X"06",X"00",X"21",X"EC",X"43",X"CD",X"FC",X"3B",X"21",X"0E",X"68",X"75",X"24",X"7E",X"F6",
		X"01",X"E6",X"FD",X"77",X"3A",X"BE",X"17",X"32",X"A7",X"43",X"CD",X"BD",X"20",X"CD",X"E9",X"20",
		X"CD",X"FD",X"00",X"3E",X"FD",X"32",X"23",X"43",X"21",X"01",X"50",X"75",X"E5",X"CD",X"82",X"17",
		X"C4",X"EA",X"18",X"3E",X"01",X"32",X"F4",X"43",X"AF",X"32",X"EB",X"43",X"CD",X"FD",X"00",X"3E",
		X"FD",X"32",X"C3",X"40",X"E1",X"2B",X"75",X"3E",X"02",X"32",X"F4",X"43",X"C9",X"21",X"45",X"43",
		X"06",X"5D",X"CD",X"D4",X"3C",X"2E",X"8B",X"36",X"01",X"2E",X"44",X"36",X"01",X"21",X"01",X"00",
		X"22",X"40",X"43",X"CD",X"AB",X"1E",X"CD",X"5D",X"20",X"CD",X"62",X"1F",X"21",X"00",X"00",X"22",
		X"85",X"43",X"3E",X"01",X"32",X"7E",X"43",X"32",X"7D",X"43",X"3E",X"38",X"32",X"9D",X"43",X"21",
		X"01",X"50",X"22",X"9A",X"43",X"CD",X"EB",X"21",X"21",X"81",X"43",X"36",X"00",X"23",X"36",X"00",
		X"23",X"36",X"60",X"2E",X"6C",X"36",X"01",X"2E",X"43",X"36",X"00",X"C3",X"91",X"1D",X"21",X"F0",
		X"4B",X"20",X"3E",X"09",X"CD",X"FE",X"02",X"CD",X"6F",X"01",X"21",X"B8",X"43",X"01",X"09",X"03",
		X"11",X"06",X"00",X"70",X"19",X"0D",X"C8",X"D2",X"63",X"01",X"32",X"8B",X"43",X"76",X"C9",X"01",
		X"00",X"00",X"21",X"00",X"00",X"11",X"00",X"00",X"0A",X"03",X"5F",X"19",X"78",X"E6",X"07",X"C2",
		X"78",X"01",X"79",X"B7",X"C2",X"78",X"01",X"CD",X"AF",X"01",X"78",X"E6",X"40",X"CA",X"72",X"01",
		X"3A",X"EA",X"42",X"B7",X"C8",X"21",X"08",X"07",X"3A",X"00",X"78",X"E6",X"80",X"C2",X"98",X"01",
		X"3A",X"00",X"78",X"E6",X"80",X"CA",X"A0",X"01",X"2B",X"7C",X"B5",X"C2",X"98",X"01",X"C9",X"78",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"3D",X"F5",X"EB",X"07",X"21",X"F9",X"01",X"CD",X"9D",X"02",X"F1",
		X"CC",X"E8",X"01",X"7B",X"BE",X"C2",X"CC",X"01",X"23",X"7A",X"BE",X"C8",X"21",X"09",X"02",X"11",
		X"EA",X"42",X"CD",X"76",X"02",X"78",X"0F",X"0F",X"0F",X"E6",X"0F",X"F6",X"30",X"12",X"06",X"40",
		X"0E",X"03",X"21",X"1F",X"02",X"C3",X"5D",X"02",X"E5",X"7E",X"23",X"86",X"2F",X"6F",X"3E",X"00",
		X"CE",X"00",X"2F",X"67",X"23",X"19",X"EB",X"E1",X"C9",X"2D",X"49",X"E2",X"61",X"C6",X"FC",X"62",
		X"30",X"6F",X"C1",X"47",X"78",X"72",X"0A",X"88",X"E7",X"52",X"45",X"50",X"4C",X"41",X"43",X"45",
		X"20",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"20",X"52",X"4F",X"4D",X"20",X"23",X"00",X"8C",
		X"42",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"5C",X"20",X"31",X"39",X"38",
		X"32",X"00",X"CE",X"42",X"52",X"4F",X"43",X"4B",X"2D",X"4F",X"4C",X"41",X"20",X"4D",X"46",X"47",
		X"2E",X"20",X"43",X"4F",X"52",X"50",X"2E",X"00",X"30",X"42",X"53",X"55",X"52",X"56",X"49",X"56",
		X"41",X"4C",X"00",X"8F",X"49",X"5E",X"00",X"3A",X"F0",X"43",X"E6",X"01",X"C8",X"5E",X"23",X"56",
		X"23",X"CD",X"76",X"02",X"0D",X"C2",X"5D",X"02",X"C9",X"0D",X"FA",X"76",X"02",X"7E",X"23",X"B7",
		X"CA",X"69",X"02",X"C3",X"6D",X"02",X"7E",X"23",X"B7",X"C8",X"FE",X"41",X"DA",X"86",X"02",X"FE",
		X"60",X"D2",X"86",X"02",X"D6",X"40",X"12",X"CD",X"83",X"3C",X"C3",X"76",X"02",X"CD",X"9D",X"02",
		X"7E",X"23",X"66",X"6F",X"C9",X"CD",X"9D",X"02",X"7E",X"BD",X"C3",X"9E",X"02",X"85",X"6F",X"7C",
		X"CE",X"00",X"67",X"C9",X"21",X"00",X"01",X"01",X"00",X"06",X"21",X"A5",X"02",X"3A",X"8B",X"43",
		X"07",X"E6",X"03",X"CD",X"9D",X"02",X"7E",X"21",X"AA",X"02",X"E5",X"15",X"00",X"11",X"37",X"41",
		X"AF",X"21",X"BC",X"02",X"19",X"AE",X"C8",X"11",X"FE",X"FF",X"01",X"A4",X"FF",X"19",X"5E",X"09",
		X"56",X"7B",X"07",X"07",X"07",X"E6",X"03",X"21",X"A5",X"02",X"CD",X"9D",X"02",X"7A",X"BE",X"C8",
		X"E1",X"21",X"96",X"43",X"7E",X"34",X"FE",X"0F",X"D2",X"1E",X"1B",X"C3",X"2E",X"00",X"CD",X"F9",
		X"02",X"21",X"3F",X"43",X"3E",X"3F",X"C3",X"FE",X"02",X"21",X"3F",X"4B",X"3E",X"47",X"36",X"00",
		X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",
		X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",
		X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"36",X"00",X"2B",X"BC",X"C2",
		X"FE",X"02",X"C9",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",
		X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"21",X"A9",X"43",X"7E",X"23",
		X"E5",X"07",X"E6",X"0E",X"21",X"8A",X"03",X"C3",X"42",X"09",X"B2",X"03",X"54",X"04",X"1A",X"3B",
		X"D5",X"37",X"35",X"3A",X"D5",X"37",X"54",X"04",X"1A",X"3B",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"B7",X"C2",X"CA",X"03",X"34",X"CD",X"EE",X"02",X"21",X"85",X"3B",X"0E",X"01",X"CD",
		X"5D",X"02",X"21",X"CD",X"3B",X"0E",X"01",X"C3",X"5D",X"02",X"23",X"34",X"2B",X"C2",X"D1",X"03",
		X"34",X"4E",X"79",X"FE",X"32",X"DA",X"E3",X"03",X"AF",X"23",X"77",X"2B",X"77",X"2B",X"34",X"20",
		X"C3",X"EE",X"02",X"E6",X"01",X"CA",X"FD",X"03",X"79",X"FE",X"01",X"23",X"CA",X"F3",X"03",X"7E",
		X"FE",X"03",X"D8",X"36",X"FF",X"21",X"07",X"04",X"0E",X"02",X"C3",X"5D",X"02",X"23",X"7E",X"FE",
		X"05",X"D8",X"36",X"FF",X"C3",X"83",X"21",X"0A",X"42",X"53",X"55",X"52",X"56",X"49",X"56",X"41",
		X"4C",X"00",X"8C",X"42",X"52",X"4F",X"43",X"4B",X"2D",X"4F",X"4C",X"41",X"20",X"5C",X"20",X"31",
		X"39",X"38",X"32",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B7",X"C2",X"5A",X"04",X"34",X"20",X"23",X"34",X"2B",X"C2",X"61",X"04",
		X"34",X"4E",X"79",X"FE",X"09",X"DA",X"70",X"04",X"AF",X"23",X"77",X"2B",X"77",X"2B",X"34",X"C9",
		X"FE",X"02",X"D2",X"DE",X"04",X"23",X"36",X"FF",X"CD",X"BD",X"20",X"CD",X"FD",X"00",X"3E",X"02",
		X"32",X"9E",X"43",X"21",X"00",X"00",X"22",X"40",X"43",X"3E",X"FD",X"32",X"23",X"43",X"AF",X"32",
		X"6D",X"43",X"32",X"F4",X"43",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"FE",X"03",
		X"D2",X"A1",X"06",X"23",X"36",X"00",X"3E",X"02",X"32",X"9E",X"43",X"CD",X"71",X"22",X"21",X"F5",
		X"43",X"7E",X"FE",X"02",X"D8",X"3E",X"FF",X"32",X"AB",X"43",X"E5",X"CD",X"D3",X"23",X"E1",X"CD",
		X"AB",X"25",X"21",X"15",X"05",X"22",X"75",X"43",X"3A",X"BA",X"43",X"E6",X"10",X"C8",X"21",X"DD",
		X"05",X"22",X"75",X"43",X"C9",X"08",X"08",X"08",X"08",X"08",X"02",X"02",X"02",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"08",X"08",X"03",X"02",X"08",X"08",X"08",X"08",X"08",X"05",X"05",X"05",
		X"05",X"05",X"05",X"06",X"07",X"07",X"07",X"06",X"08",X"08",X"08",X"08",X"00",X"02",X"05",X"00",
		X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"02",X"03",X"03",X"03",
		X"03",X"02",X"01",X"01",X"01",X"01",X"08",X"08",X"08",X"00",X"08",X"08",X"08",X"18",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"07",X"07",X"07",X"07",
		X"07",X"07",X"00",X"02",X"02",X"08",X"08",X"08",X"08",X"04",X"06",X"06",X"06",X"05",X"04",X"02",
		X"01",X"01",X"01",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"D4",X"00",X"D0",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"D4",X"00",X"D0",X"00",X"D4",X"00",X"D0",
		X"00",X"D4",X"00",X"D0",X"00",X"D4",X"00",X"D0",X"00",X"D4",X"00",X"00",X"00",X"08",X"08",X"08",
		X"08",X"08",X"02",X"02",X"08",X"08",X"08",X"01",X"01",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"06",X"06",X"06",X"08",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"02",X"03",X"03",
		X"02",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"18",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"05",X"05",X"05",X"05",X"05",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"06",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"03",X"02",X"02",X"02",X"02",X"02",X"01",X"00",X"00",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"05",X"04",X"02",X"07",X"06",X"05",X"05",X"05",X"06",X"00",
		X"01",X"02",X"03",X"04",X"04",X"02",X"00",X"07",X"07",X"05",X"04",X"02",X"01",X"00",X"00",X"01",
		X"02",X"03",X"04",X"05",X"05",X"05",X"06",X"00",X"01",X"02",X"00",X"00",X"00",X"08",X"02",X"08",
		X"08",X"08",X"04",X"05",X"05",X"05",X"05",X"08",X"01",X"01",X"01",X"01",X"01",X"08",X"08",X"08",
		X"80",X"FE",X"04",X"D2",X"02",X"07",X"23",X"36",X"00",X"CD",X"C0",X"0A",X"2A",X"75",X"43",X"23",
		X"7E",X"FE",X"80",X"C0",X"3E",X"FF",X"32",X"AB",X"43",X"C9",X"00",X"00",X"D4",X"00",X"D4",X"00",
		X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"D4",X"00",X"D0",X"00",X"D4",X"00",X"D0",X"00",X"D4",X"00",
		X"D0",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"D0",X"D5",
		X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",
		X"00",X"00",X"FE",X"05",X"D8",X"FE",X"06",X"D2",X"7C",X"07",X"23",X"36",X"FF",X"CD",X"83",X"21",
		X"CD",X"1C",X"01",X"21",X"01",X"00",X"22",X"40",X"43",X"AF",X"32",X"7F",X"43",X"32",X"9D",X"43",
		X"32",X"9E",X"43",X"CD",X"AB",X"1E",X"21",X"00",X"00",X"22",X"F7",X"43",X"23",X"22",X"F5",X"43",
		X"22",X"6C",X"43",X"C9",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D4",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"00",X"00",X"00",X"D0",X"D5",X"D5",
		X"D5",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",
		X"D5",X"D5",X"D0",X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"D5",
		X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"00",X"FE",X"07",X"D2",X"F7",
		X"07",X"23",X"4E",X"79",X"32",X"9D",X"43",X"D6",X"09",X"D8",X"E6",X"07",X"CC",X"DF",X"07",X"79",
		X"FE",X"38",X"D8",X"C3",X"36",X"09",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"D4",X"00",X"D0",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"C5",
		X"E5",X"11",X"05",X"4B",X"79",X"0F",X"0F",X"0F",X"E6",X"1F",X"83",X"5F",X"21",X"4B",X"23",X"0E",
		X"18",X"CD",X"30",X"3D",X"E1",X"C1",X"C9",X"FE",X"08",X"D0",X"23",X"36",X"00",X"3A",X"F5",X"43",
		X"E6",X"07",X"FE",X"07",X"C2",X"36",X"09",X"36",X"FF",X"21",X"00",X"00",X"22",X"ED",X"43",X"22",
		X"45",X"43",X"22",X"46",X"43",X"22",X"8F",X"43",X"AF",X"32",X"88",X"43",X"D0",X"CD",X"36",X"09",
		X"20",X"C3",X"B3",X"20",X"00",X"00",X"00",X"E7",X"08",X"08",X"08",X"08",X"08",X"18",X"08",X"08",
		X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"08",X"08",X"08",X"02",X"08",X"08",X"08",X"18",X"08",
		X"08",X"18",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"28",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"08",
		X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"08",X"08",X"02",X"08",X"08",X"18",X"08",
		X"18",X"08",X"08",X"08",X"08",X"08",X"18",X"18",X"28",X"08",X"08",X"00",X"00",X"08",X"08",X"02",
		X"08",X"08",X"08",X"18",X"08",X"18",X"08",X"18",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"02",
		X"08",X"18",X"28",X"08",X"18",X"18",X"06",X"18",X"28",X"08",X"18",X"08",X"18",X"00",X"00",X"00",
		X"07",X"06",X"28",X"08",X"18",X"08",X"18",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"07",X"07",X"07",X"11",X"01",X"08",X"06",X"05",X"05",X"05",X"04",X"03",X"04",X"04",X"04",
		X"04",X"05",X"05",X"05",X"00",X"10",X"10",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"12",X"02",X"08",X"06",X"26",X"06",X"02",X"12",X"12",X"02",X"12",X"06",
		X"16",X"06",X"26",X"06",X"15",X"05",X"26",X"06",X"06",X"16",X"15",X"05",X"05",X"05",X"15",X"06",
		X"07",X"10",X"10",X"00",X"07",X"17",X"26",X"02",X"12",X"12",X"22",X"02",X"02",X"04",X"05",X"05",
		X"05",X"08",X"01",X"01",X"01",X"01",X"11",X"18",X"04",X"04",X"04",X"04",X"08",X"01",X"02",X"04",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"06",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"10",X"10",X"01",X"02",X"13",X"13",X"04",X"02",X"11",X"12",X"04",X"05",X"15",
		X"25",X"05",X"03",X"03",X"02",X"80",X"00",X"21",X"F5",X"43",X"7E",X"07",X"E6",X"0E",X"E5",X"21",
		X"98",X"09",X"CD",X"8D",X"02",X"20",X"E3",X"7E",X"C9",X"D0",X"D0",X"D0",X"D5",X"D5",X"D5",X"D5",
		X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",
		X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"22",X"0F",X"11",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"21",X"71",X"22",X"D3",X"23",X"AB",X"25",
		X"00",X"0A",X"AE",X"17",X"62",X"26",X"02",X"2D",X"00",X"0A",X"AE",X"17",X"62",X"26",X"02",X"2D",
		X"00",X"0A",X"AE",X"17",X"62",X"26",X"02",X"2D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",
		X"D0",X"D0",X"00",X"00",X"D0",X"00",X"D0",X"00",X"D0",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",
		X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"F7",X"43",X"7E",X"34",X"07",X"E6",X"1E",X"E5",X"21",X"58",X"0A",X"C3",X"42",X"09",
		X"00",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",
		X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",
		X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"0B",X"85",X"0B",X"8C",X"0B",X"9C",X"0B",
		X"A3",X"0B",X"AD",X"0B",X"B1",X"0B",X"BE",X"0B",X"C5",X"0B",X"CF",X"0B",X"D3",X"0B",X"E3",X"0B",
		X"EA",X"0B",X"F1",X"0B",X"F5",X"0B",X"F9",X"0B",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",
		X"D5",X"D5",X"D0",X"00",X"D4",X"00",X"D0",X"00",X"D4",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"D4",X"00",
		X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"D0",X"D5",X"D5",X"D5",
		X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"D4",X"00",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",
		X"00",X"21",X"F7",X"43",X"7E",X"34",X"07",X"E6",X"1E",X"E5",X"21",X"18",X"0B",X"C3",X"42",X"09",
		X"00",X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",
		X"D0",X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D4",X"00",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",
		X"D4",X"00",X"D0",X"D5",X"D5",X"D5",X"D5",X"D0",X"03",X"0C",X"0A",X"0C",X"11",X"0C",X"1B",X"0C",
		X"22",X"0C",X"29",X"0C",X"30",X"0C",X"37",X"0C",X"3E",X"0C",X"45",X"0C",X"4C",X"0C",X"56",X"0C",
		X"5D",X"0C",X"64",X"0C",X"65",X"0C",X"68",X"0C",X"C9",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",
		X"00",X"D0",X"D0",X"00",X"D0",X"D0",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D0",X"D0",X"D0",X"00",X"00",X"00",
		X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CD",X"8C",X"12",X"C9",X"CD",X"32",X"11",X"CD",X"C9",X"0F",X"C9",X"CD",X"93",X"11",X"CD",
		X"2B",X"19",X"CD",X"7A",X"1C",X"CD",X"5A",X"0D",X"CD",X"CE",X"19",X"C9",X"CD",X"DA",X"12",X"CD",
		X"32",X"11",X"C9",X"CD",X"93",X"11",X"CD",X"90",X"1D",X"CD",X"CA",X"0C",X"C9",X"CD",X"32",X"11",
		X"C9",X"CD",X"93",X"11",X"CD",X"CE",X"19",X"CD",X"7A",X"1C",X"CD",X"5A",X"0D",X"C9",X"CD",X"32",
		X"11",X"CD",X"C9",X"0F",X"C9",X"CD",X"93",X"11",X"CD",X"90",X"1D",X"CD",X"CA",X"0C",X"C9",X"CD",
		X"32",X"11",X"C9",X"CD",X"93",X"11",X"CD",X"2B",X"19",X"CD",X"7A",X"1C",X"CD",X"5A",X"0D",X"CD",
		X"CE",X"19",X"C9",X"CD",X"DA",X"12",X"CD",X"32",X"11",X"C9",X"CD",X"90",X"1D",X"CD",X"E2",X"1D",
		X"C9",X"CD",X"73",X"1E",X"C9",X"CD",X"86",X"1E",X"C9",X"CD",X"93",X"11",X"CD",X"90",X"1D",X"CD",
		X"CA",X"0C",X"C9",X"CD",X"8C",X"12",X"CD",X"CF",X"0D",X"C9",X"CD",X"32",X"11",X"CD",X"C9",X"0F",
		X"C9",X"CD",X"93",X"11",X"CD",X"2B",X"19",X"CD",X"CE",X"19",X"C9",X"CD",X"DA",X"12",X"CD",X"32",
		X"11",X"C9",X"CD",X"93",X"11",X"CD",X"90",X"1D",X"C9",X"CD",X"CF",X"0D",X"CD",X"32",X"11",X"C9",
		X"CD",X"93",X"11",X"CD",X"CE",X"19",X"C9",X"CD",X"32",X"11",X"CD",X"C9",X"0F",X"C9",X"CD",X"93",
		X"11",X"CD",X"90",X"1D",X"C9",X"CD",X"CF",X"0D",X"CD",X"32",X"11",X"C9",X"CD",X"93",X"11",X"CD",
		X"2B",X"19",X"CD",X"CE",X"19",X"C9",X"CD",X"DA",X"12",X"CD",X"32",X"11",X"C9",X"CD",X"93",X"11",
		X"CD",X"90",X"1D",X"C9",X"C9",X"C3",X"38",X"0B",X"CD",X"90",X"1D",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D0",X"D0",X"D0",X"D0",X"00",X"00",X"00",
		X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"17",X"6A",X"11",X"33",X"6C",X"0E",X"10",X"3E",X"20",X"96",X"12",
		X"13",X"2B",X"0D",X"F2",X"BD",X"0C",X"BE",X"CA",X"08",X"32",X"00",X"CD",X"CF",X"0D",X"CD",X"5B",
		X"10",X"21",X"7D",X"43",X"7E",X"B7",X"C0",X"2E",X"6C",X"36",X"01",X"2E",X"4A",X"77",X"2E",X"89",
		X"77",X"2E",X"90",X"36",X"01",X"23",X"36",X"02",X"23",X"77",X"2E",X"87",X"77",X"2E",X"93",X"77",
		X"23",X"77",X"2E",X"4E",X"77",X"23",X"77",X"2E",X"F5",X"34",X"23",X"23",X"3E",X"F8",X"A6",X"77",
		X"2E",X"40",X"7E",X"FE",X"06",X"D8",X"2E",X"43",X"36",X"0F",X"2E",X"48",X"36",X"50",X"C8",X"36",
		X"85",X"C9",X"D0",X"D0",X"D5",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D5",X"D0",X"D0",X"D5",
		X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D5",X"D0",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"D4",X"00",X"00",X"00",X"00",X"D4",X"D4",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"D4",X"D4",X"00",
		X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"40",X"4B",X"3A",X"42",X"43",
		X"4F",X"3A",X"7F",X"43",X"B7",X"C8",X"47",X"E6",X"01",X"C0",X"7E",X"E6",X"10",X"C0",X"7E",X"E6",
		X"E0",X"B8",X"C0",X"7D",X"C6",X"05",X"6F",X"0D",X"C2",X"6A",X"0D",X"78",X"F6",X"01",X"32",X"7F",
		X"43",X"3E",X"0B",X"32",X"92",X"43",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D4",
		X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D4",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"D0",X"D0",X"D4",X"D0",X"00",X"00",X"00",X"00",X"D0",X"D4",X"D0",
		X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",
		X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",
		X"7F",X"43",X"E6",X"01",X"C0",X"21",X"40",X"4B",X"E5",X"7E",X"FE",X"60",X"DA",X"04",X"0E",X"E6",
		X"10",X"C2",X"04",X"0E",X"23",X"56",X"23",X"5E",X"21",X"4F",X"4B",X"7D",X"C6",X"05",X"6F",X"FE",
		X"90",X"D2",X"04",X"0E",X"7E",X"E6",X"E0",X"FE",X"20",X"CC",X"5B",X"0E",X"C2",X"EB",X"0D",X"E1",
		X"E5",X"CD",X"BC",X"0E",X"E1",X"7D",X"C6",X"05",X"6F",X"FE",X"59",X"DA",X"D8",X"0D",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"D0",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"D0",X"00",X"00",X"00",X"00",X"D0",X"D5",
		X"D5",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"B7",X"CA",X"BD",X"0C",X"23",X"7E",X"2B",X"BA",X"CA",
		X"65",X"0E",X"3D",X"BA",X"C0",X"23",X"23",X"7E",X"2B",X"2B",X"BB",X"CA",X"71",X"0E",X"3D",X"BB",
		X"C0",X"36",X"00",X"C9",X"D0",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"D5",X"D0",X"00",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"11",X"51",X"43",X"0E",
		X"05",X"E5",X"1A",X"B7",X"CA",X"D1",X"0E",X"7B",X"C6",X"05",X"5F",X"0D",X"C2",X"C2",X"0E",X"E1",
		X"C9",X"0E",X"03",X"CD",X"3C",X"3C",X"AF",X"12",X"13",X"12",X"D1",X"D5",X"7B",X"D6",X"40",X"21",
		X"C8",X"24",X"CD",X"9D",X"02",X"0E",X"04",X"CD",X"3C",X"3C",X"3E",X"14",X"12",X"21",X"47",X"43",
		X"01",X"00",X"05",X"CD",X"EA",X"3B",X"21",X"01",X"80",X"22",X"90",X"43",X"D1",X"21",X"7F",X"43",
		X"7E",X"B7",X"C2",X"0D",X"0F",X"1A",X"E6",X"E0",X"77",X"C6",X"04",X"4F",X"C9",X"E6",X"E0",X"47",
		X"EB",X"7E",X"E6",X"1F",X"B0",X"77",X"C9",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"D0",
		X"D0",X"D0",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"D0",
		X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"E6",X"E0",X"D6",X"60",X"07",X"07",X"07",X"E6",X"03",
		X"C9",X"D0",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D5",X"D5",
		X"D5",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"D0",X"D4",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"D4",X"21",X"51",X"43",X"01",X"05",X"05",X"7E",
		X"B7",X"CA",X"DB",X"0F",X"E5",X"C5",X"CD",X"2B",X"10",X"C1",X"E1",X"7D",X"81",X"6F",X"05",X"C2",
		X"CF",X"0F",X"C9",X"00",X"00",X"D4",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",
		X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"04",X"00",X"0A",X"03",X"03",X"0B",X"00",X"0A",X"03",X"03",X"04",X"00",X"0A",X"12",X"00",X"16",
		X"09",X"00",X"00",X"00",X"00",X"05",X"00",X"0A",X"09",X"00",X"05",X"00",X"00",X"00",X"00",X"0C",
		X"03",X"0D",X"0E",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"23",X"23",X"23",X"7E",X"34",
		X"2B",X"B7",X"CA",X"44",X"10",X"FE",X"10",X"DA",X"51",X"10",X"2B",X"2B",X"AF",X"77",X"47",X"23",
		X"23",X"CA",X"1F",X"13",X"CD",X"51",X"10",X"21",X"1F",X"F8",X"19",X"EB",X"0E",X"00",X"C3",X"FA",
		X"13",X"07",X"07",X"E6",X"3C",X"C6",X"80",X"47",X"D2",X"1F",X"13",X"21",X"73",X"43",X"56",X"23",
		X"5E",X"21",X"40",X"4B",X"3A",X"42",X"43",X"47",X"7E",X"E6",X"10",X"CC",X"1D",X"11",X"C2",X"B3",
		X"10",X"E5",X"CD",X"9B",X"1E",X"E1",X"3A",X"7D",X"43",X"B7",X"C8",X"20",X"E5",X"21",X"4A",X"43",
		X"36",X"01",X"2E",X"93",X"36",X"B0",X"23",X"36",X"04",X"2E",X"92",X"36",X"00",X"2E",X"72",X"11",
		X"4B",X"43",X"0E",X"03",X"CD",X"3C",X"3C",X"AF",X"EB",X"77",X"23",X"77",X"2E",X"8B",X"77",X"2E",
		X"F7",X"3E",X"F8",X"A6",X"77",X"2E",X"F5",X"34",X"CD",X"58",X"19",X"E1",X"7E",X"CD",X"77",X"0F",
		X"47",X"37",X"C9",X"7D",X"C6",X"05",X"6F",X"05",X"C2",X"68",X"10",X"AF",X"C9",X"00",X"00",X"07",
		X"03",X"03",X"08",X"00",X"0C",X"03",X"03",X"0B",X"00",X"06",X"00",X"00",X"06",X"00",X"06",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"05",X"00",X"00",
		X"05",X"00",X"05",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"1B",
		X"1C",X"00",X"02",X"05",X"00",X"05",X"00",X"00",X"05",X"00",X"05",X"00",X"10",X"0F",X"00",X"1A",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"06",X"00",X"00",
		X"06",X"00",X"06",X"00",X"00",X"06",X"00",X"07",X"03",X"03",X"08",X"00",X"00",X"23",X"7E",X"92",
		X"CD",X"6F",X"3C",X"4F",X"23",X"7E",X"93",X"CD",X"6F",X"3C",X"B1",X"2B",X"2B",X"FE",X"02",X"3F",
		X"9F",X"C9",X"00",X"21",X"40",X"4B",X"3A",X"42",X"43",X"47",X"B7",X"07",X"07",X"80",X"85",X"6F",
		X"3E",X"10",X"90",X"47",X"0E",X"05",X"7E",X"B7",X"CA",X"52",X"11",X"E5",X"C5",X"CD",X"4C",X"1A",
		X"C1",X"E1",X"79",X"85",X"6F",X"05",X"C2",X"46",X"11",X"21",X"90",X"4B",X"3A",X"42",X"43",X"47",
		X"07",X"07",X"80",X"85",X"6F",X"0E",X"05",X"3E",X"10",X"90",X"47",X"7E",X"B7",X"CA",X"77",X"11",
		X"C5",X"E5",X"CD",X"FB",X"11",X"E1",X"C1",X"79",X"85",X"6F",X"05",X"C2",X"6B",X"11",X"11",X"A4",
		X"4B",X"21",X"54",X"4B",X"0E",X"3C",X"C3",X"3C",X"3C",X"3A",X"A5",X"43",X"BA",X"C2",X"52",X"11",
		X"C3",X"77",X"11",X"00",X"AF",X"32",X"98",X"43",X"21",X"40",X"4B",X"3A",X"42",X"43",X"47",X"07",
		X"07",X"80",X"85",X"6F",X"0E",X"05",X"3E",X"10",X"90",X"47",X"7E",X"B7",X"CA",X"B6",X"11",X"E5",
		X"C5",X"CD",X"00",X"12",X"C1",X"E1",X"79",X"85",X"6F",X"05",X"C2",X"AA",X"11",X"21",X"98",X"43",
		X"7E",X"B7",X"C0",X"23",X"23",X"7E",X"23",X"B6",X"C0",X"2E",X"85",X"7E",X"B7",X"CA",X"D4",X"11",
		X"23",X"7E",X"B7",X"C0",X"CD",X"9B",X"1E",X"3A",X"7D",X"43",X"B7",X"C8",X"21",X"4A",X"43",X"7E",
		X"B7",X"C0",X"36",X"03",X"2E",X"89",X"36",X"10",X"AF",X"2E",X"92",X"77",X"2E",X"4E",X"77",X"23",
		X"77",X"2E",X"F5",X"34",X"23",X"23",X"3E",X"F8",X"A6",X"77",X"C9",X"0E",X"00",X"C3",X"01",X"12",
		X"4E",X"C5",X"E5",X"23",X"7E",X"23",X"4E",X"CD",X"92",X"1D",X"21",X"00",X"08",X"19",X"D1",X"C1",
		X"46",X"71",X"79",X"B7",X"C8",X"32",X"98",X"43",X"78",X"FE",X"D0",X"D8",X"32",X"9C",X"43",X"C2",
		X"4A",X"12",X"36",X"D1",X"CD",X"82",X"12",X"3A",X"45",X"43",X"3C",X"32",X"45",X"43",X"E5",X"E5",
		X"E5",X"CD",X"78",X"12",X"E1",X"CD",X"6E",X"12",X"E1",X"CD",X"5C",X"12",X"E1",X"3E",X"D5",X"11",
		X"E0",X"FF",X"19",X"BE",X"C0",X"36",X"D3",X"C3",X"42",X"12",X"FE",X"D4",X"CA",X"64",X"12",X"FE",
		X"D5",X"C0",X"36",X"D3",X"CD",X"82",X"12",X"E5",X"CD",X"3D",X"12",X"E1",X"3E",X"D5",X"11",X"20",
		X"00",X"C3",X"42",X"12",X"36",X"D2",X"CD",X"82",X"12",X"E5",X"CD",X"78",X"12",X"E1",X"3E",X"D4",
		X"23",X"BE",X"C0",X"36",X"D2",X"C3",X"70",X"12",X"3E",X"D4",X"2B",X"BE",X"C0",X"36",X"D2",X"C3",
		X"7A",X"12",X"E5",X"21",X"50",X"00",X"19",X"AF",X"12",X"77",X"E1",X"C9",X"00",X"21",X"40",X"4B",
		X"7E",X"E6",X"10",X"C2",X"9B",X"12",X"E5",X"CD",X"18",X"14",X"E1",X"7D",X"C6",X"05",X"6F",X"FE",
		X"54",X"DA",X"90",X"12",X"7E",X"FE",X"60",X"DA",X"AF",X"12",X"E6",X"10",X"CC",X"18",X"14",X"21",
		X"90",X"4B",X"E5",X"CD",X"C9",X"13",X"E1",X"7D",X"C6",X"05",X"6F",X"FE",X"A4",X"DA",X"B2",X"12",
		X"7E",X"FE",X"60",X"D4",X"C9",X"13",X"CD",X"88",X"13",X"11",X"90",X"4B",X"21",X"40",X"4B",X"3A",
		X"42",X"43",X"4F",X"07",X"07",X"81",X"4F",X"C3",X"3C",X"3C",X"00",X"CD",X"F0",X"18",X"21",X"40",
		X"4B",X"01",X"05",X"05",X"7E",X"E6",X"10",X"CA",X"F1",X"12",X"C5",X"E5",X"CD",X"F9",X"12",X"E1",
		X"C1",X"79",X"85",X"6F",X"05",X"C2",X"E4",X"12",X"C9",X"23",X"23",X"23",X"23",X"7E",X"35",X"B7",
		X"C0",X"77",X"2B",X"7E",X"34",X"2B",X"FE",X"10",X"DA",X"18",X"13",X"2B",X"2B",X"7E",X"E6",X"EF",
		X"77",X"23",X"23",X"06",X"00",X"C3",X"1F",X"13",X"07",X"07",X"E6",X"3C",X"C6",X"40",X"47",X"4E",
		X"2B",X"7E",X"CD",X"92",X"1D",X"21",X"00",X"08",X"19",X"EB",X"48",X"C3",X"FA",X"13",X"3A",X"F0",
		X"43",X"E6",X"03",X"CA",X"8F",X"13",X"FE",X"02",X"C0",X"C3",X"95",X"13",X"3A",X"F0",X"43",X"E6",
		X"03",X"CA",X"BD",X"13",X"FE",X"02",X"C0",X"C3",X"98",X"13",X"00",X"3A",X"F5",X"43",X"E6",X"07",
		X"FE",X"04",X"CA",X"88",X"13",X"FE",X"05",X"CA",X"02",X"18",X"FE",X"07",X"C0",X"3A",X"6C",X"43",
		X"B7",X"C8",X"3A",X"4F",X"43",X"FE",X"04",X"D0",X"B7",X"CA",X"88",X"13",X"3A",X"F0",X"43",X"E6",
		X"03",X"CA",X"8F",X"13",X"FE",X"02",X"CA",X"95",X"13",X"21",X"9F",X"43",X"4E",X"23",X"7E",X"23",
		X"66",X"6F",X"79",X"B7",X"C8",X"C3",X"5D",X"02",X"3A",X"F0",X"43",X"0F",X"DA",X"95",X"13",X"CD",
		X"BD",X"13",X"C3",X"66",X"19",X"CD",X"66",X"19",X"21",X"40",X"4B",X"3A",X"42",X"43",X"47",X"0E",
		X"FB",X"07",X"07",X"80",X"85",X"D6",X"05",X"6F",X"7E",X"E6",X"10",X"C2",X"B5",X"13",X"E5",X"C5",
		X"CD",X"D5",X"13",X"C1",X"E1",X"7D",X"81",X"6F",X"05",X"C2",X"A8",X"13",X"C9",X"21",X"40",X"4B",
		X"3A",X"42",X"43",X"47",X"0E",X"05",X"C3",X"A8",X"13",X"23",X"7E",X"23",X"4E",X"CD",X"92",X"1D",
		X"0E",X"00",X"C3",X"FA",X"13",X"3A",X"F7",X"43",X"3D",X"07",X"E6",X"10",X"4F",X"46",X"78",X"C6",
		X"02",X"07",X"07",X"E6",X"10",X"A9",X"B0",X"E6",X"F0",X"4F",X"78",X"E6",X"03",X"07",X"07",X"B1",
		X"4F",X"C5",X"23",X"7E",X"23",X"4E",X"CD",X"92",X"1D",X"C1",X"79",X"12",X"13",X"B7",X"CA",X"0F",
		X"14",X"0C",X"79",X"12",X"1B",X"CD",X"83",X"3C",X"0C",X"79",X"12",X"13",X"3C",X"12",X"C9",X"12",
		X"CD",X"83",X"3C",X"AF",X"12",X"1B",X"12",X"C9",X"AF",X"32",X"97",X"43",X"7E",X"E6",X"E0",X"47",
		X"7E",X"E6",X"07",X"4F",X"23",X"E5",X"D1",X"23",X"23",X"36",X"00",X"3A",X"44",X"43",X"FE",X"04",
		X"D2",X"BB",X"14",X"3A",X"7E",X"43",X"B7",X"CA",X"BB",X"14",X"21",X"72",X"43",X"7E",X"1F",X"DA",
		X"5E",X"14",X"1F",X"23",X"DA",X"52",X"14",X"23",X"13",X"1A",X"1B",X"BE",X"C2",X"5E",X"14",X"C3",
		X"57",X"14",X"1A",X"BE",X"C2",X"5E",X"14",X"3E",X"01",X"B1",X"4F",X"C3",X"B6",X"14",X"D5",X"E1",
		X"2B",X"3A",X"F0",X"43",X"AE",X"23",X"AE",X"23",X"AE",X"23",X"AE",X"E6",X"57",X"CA",X"51",X"16",
		X"7E",X"B7",X"CA",X"BB",X"14",X"1A",X"FE",X"01",X"CA",X"85",X"14",X"FE",X"0A",X"CA",X"85",X"14",
		X"FE",X"15",X"C2",X"A1",X"14",X"79",X"E6",X"04",X"F6",X"02",X"4F",X"13",X"1A",X"1B",X"FE",X"09",
		X"DA",X"B6",X"14",X"FE",X"0C",X"D2",X"B6",X"14",X"79",X"E6",X"04",X"4F",X"36",X"00",X"C3",X"B6",
		X"14",X"3A",X"F0",X"43",X"E6",X"80",X"CA",X"0B",X"15",X"13",X"1A",X"1B",X"FE",X"0A",X"C2",X"0B",
		X"15",X"79",X"3C",X"E6",X"04",X"4F",X"79",X"B0",X"1B",X"12",X"13",X"7B",X"D6",X"41",X"2E",X"00",
		X"D6",X"05",X"DA",X"C9",X"14",X"2C",X"C3",X"C0",X"14",X"3A",X"F7",X"43",X"07",X"07",X"07",X"67",
		X"E6",X"07",X"BD",X"CA",X"51",X"16",X"3A",X"44",X"43",X"FE",X"06",X"D2",X"51",X"16",X"3A",X"92",
		X"43",X"B7",X"CA",X"F1",X"14",X"E6",X"03",X"BD",X"C2",X"F1",X"14",X"7C",X"E6",X"07",X"CA",X"51",
		X"16",X"3A",X"7E",X"43",X"B7",X"CA",X"0B",X"15",X"7C",X"C6",X"02",X"E6",X"07",X"BD",X"C2",X"0B",
		X"15",X"3A",X"72",X"43",X"E6",X"07",X"4F",X"B0",X"1B",X"12",X"13",X"D5",X"2A",X"73",X"43",X"1A",
		X"95",X"CD",X"6F",X"3C",X"6F",X"13",X"1A",X"1B",X"94",X"CD",X"6F",X"3C",X"B5",X"FE",X"02",X"DA",
		X"6F",X"15",X"FE",X"03",X"D2",X"33",X"15",X"D1",X"3A",X"97",X"43",X"B7",X"CA",X"51",X"16",X"D5",
		X"C3",X"3E",X"15",X"FE",X"04",X"D2",X"3E",X"15",X"E1",X"E5",X"23",X"23",X"36",X"01",X"79",X"07",
		X"21",X"E9",X"16",X"CD",X"9D",X"02",X"1A",X"86",X"FA",X"85",X"15",X"FE",X"17",X"D2",X"9D",X"15",
		X"13",X"23",X"1A",X"86",X"FA",X"A9",X"15",X"FE",X"18",X"D2",X"B6",X"15",X"1B",X"2B",X"CD",X"1C",
		X"1C",X"DA",X"6F",X"15",X"C2",X"D8",X"15",X"1A",X"86",X"12",X"13",X"23",X"1A",X"86",X"12",X"D1",
		X"C9",X"E1",X"3A",X"97",X"43",X"B7",X"C2",X"8F",X"15",X"E5",X"D5",X"E1",X"23",X"23",X"7E",X"B7",
		X"C0",X"F6",X"02",X"77",X"C9",X"D1",X"CD",X"71",X"15",X"79",X"D6",X"04",X"CA",X"C3",X"15",X"32",
		X"97",X"43",X"81",X"E6",X"07",X"4F",X"B0",X"1B",X"12",X"13",X"C3",X"0B",X"15",X"D1",X"CD",X"71",
		X"15",X"79",X"B7",X"CA",X"C3",X"15",X"C3",X"8F",X"15",X"D1",X"CD",X"71",X"15",X"79",X"D6",X"02",
		X"CA",X"C3",X"15",X"C3",X"8F",X"15",X"D1",X"CD",X"71",X"15",X"79",X"D6",X"06",X"CA",X"C3",X"15",
		X"C3",X"8F",X"15",X"D5",X"E1",X"23",X"23",X"7E",X"B7",X"CA",X"51",X"16",X"35",X"3A",X"44",X"43",
		X"FE",X"07",X"D2",X"51",X"16",X"C3",X"24",X"16",X"D1",X"67",X"79",X"07",X"07",X"07",X"07",X"84",
		X"21",X"FD",X"16",X"CD",X"9D",X"02",X"3A",X"97",X"43",X"B7",X"CA",X"F8",X"15",X"3A",X"F0",X"43",
		X"07",X"07",X"E6",X"02",X"3D",X"C3",X"8F",X"15",X"7E",X"32",X"97",X"43",X"B7",X"C8",X"81",X"E6",
		X"07",X"4F",X"B0",X"1B",X"12",X"13",X"13",X"13",X"EB",X"7E",X"F5",X"B7",X"C2",X"11",X"16",X"36",
		X"03",X"35",X"EB",X"1B",X"1B",X"7E",X"E1",X"CD",X"6F",X"3C",X"FE",X"04",X"C2",X"0B",X"15",X"7C",
		X"B7",X"CA",X"0B",X"15",X"2A",X"73",X"43",X"79",X"E6",X"02",X"C2",X"3B",X"16",X"13",X"1A",X"1B",
		X"BC",X"3E",X"02",X"D2",X"44",X"16",X"3E",X"06",X"C3",X"44",X"16",X"1A",X"BD",X"3E",X"00",X"DA",
		X"44",X"16",X"3E",X"04",X"4F",X"B0",X"1B",X"12",X"13",X"3E",X"03",X"32",X"97",X"43",X"C3",X"0B",
		X"15",X"D5",X"C5",X"2A",X"73",X"43",X"EB",X"7B",X"96",X"4F",X"9F",X"E6",X"04",X"5F",X"23",X"7A",
		X"96",X"47",X"9F",X"E6",X"04",X"57",X"78",X"B1",X"C2",X"6E",X"16",X"C1",X"D1",X"C9",X"78",X"CD",
		X"45",X"3C",X"67",X"79",X"CD",X"45",X"3C",X"84",X"67",X"78",X"B7",X"CA",X"96",X"16",X"79",X"B7",
		X"7A",X"C2",X"8A",X"16",X"EE",X"06",X"5F",X"C3",X"96",X"16",X"0F",X"B3",X"0F",X"5F",X"0F",X"DA",
		X"96",X"16",X"3E",X"07",X"AB",X"5F",X"C1",X"7C",X"E1",X"E5",X"23",X"23",X"23",X"BE",X"77",X"E1",
		X"EB",X"DA",X"B8",X"16",X"FE",X"04",X"DA",X"B8",X"16",X"79",X"95",X"E6",X"07",X"D6",X"04",X"3F",
		X"9F",X"E6",X"04",X"D6",X"02",X"C3",X"8F",X"15",X"4D",X"3A",X"44",X"43",X"FE",X"08",X"D2",X"DC",
		X"16",X"3A",X"7E",X"43",X"B7",X"CA",X"DC",X"16",X"2A",X"EF",X"43",X"7C",X"81",X"07",X"CE",X"03",
		X"AD",X"E6",X"16",X"C2",X"DC",X"16",X"79",X"C6",X"04",X"E6",X"07",X"4F",X"79",X"B0",X"1B",X"12",
		X"13",X"3E",X"03",X"32",X"97",X"43",X"C3",X"0B",X"15",X"01",X"00",X"01",X"FF",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"01",X"00",X"01",X"01",X"01",X"11",X"0D",X"17",X"01",X"00",X"00",X"FF",
		X"00",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",
		X"FF",X"01",X"FD",X"01",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",
		X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"FF",X"FD",X"00",X"00",X"01",X"01",X"00",X"00",X"FF",X"FD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"03",X"00",X"3A",X"A1",X"42",
		X"47",X"11",X"11",X"34",X"02",X"21",X"2B",X"1F",X"0E",X"08",X"1A",X"BE",X"13",X"23",X"C0",X"0D",
		X"C8",X"C3",X"8A",X"17",X"3A",X"00",X"78",X"2F",X"E6",X"60",X"0F",X"0F",X"0F",X"0F",X"C6",X"02",
		X"47",X"FE",X"08",X"DA",X"AB",X"17",X"06",X"10",X"0E",X"05",X"C9",X"0F",X"4F",X"C9",X"00",X"34",
		X"3A",X"4A",X"43",X"B7",X"C8",X"35",X"21",X"4F",X"43",X"7E",X"B7",X"C2",X"66",X"18",X"34",X"2E",
		X"90",X"36",X"01",X"23",X"36",X"02",X"2E",X"87",X"36",X"00",X"21",X"85",X"43",X"7E",X"B7",X"CA",
		X"D8",X"17",X"23",X"36",X"00",X"F4",X"A1",X"1C",X"21",X"3F",X"4B",X"11",X"00",X"48",X"01",X"D4",
		X"D0",X"7E",X"B8",X"DA",X"F2",X"17",X"CA",X"F3",X"17",X"B9",X"DA",X"F2",X"17",X"FE",X"D6",X"DA",
		X"F3",X"17",X"73",X"2D",X"C2",X"E1",X"17",X"25",X"7C",X"BA",X"D2",X"E1",X"17",X"C9",X"11",X"C1",
		X"C5",X"21",X"3A",X"4A",X"43",X"B7",X"CA",X"88",X"13",X"3A",X"F0",X"43",X"E6",X"01",X"C2",X"1F",
		X"18",X"3A",X"4A",X"43",X"FE",X"02",X"F5",X"D4",X"2E",X"13",X"F1",X"DC",X"3C",X"13",X"C9",X"3A",
		X"4A",X"43",X"3D",X"4F",X"11",X"A6",X"42",X"21",X"2D",X"18",X"C3",X"69",X"02",X"2A",X"20",X"41",
		X"20",X"56",X"49",X"52",X"55",X"53",X"20",X"47",X"4F",X"54",X"20",X"59",X"4F",X"55",X"21",X"00",
		X"2A",X"20",X"43",X"45",X"4C",X"4C",X"20",X"4C",X"49",X"46",X"45",X"20",X"4F",X"56",X"45",X"52",
		X"21",X"21",X"00",X"2A",X"20",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",X"4D",X"45",X"44",X"49",
		X"43",X"49",X"4E",X"45",X"21",X"00",X"FE",X"02",X"DA",X"92",X"18",X"2B",X"34",X"7E",X"FE",X"40",
		X"D8",X"2E",X"F5",X"34",X"AF",X"32",X"50",X"43",X"32",X"8B",X"43",X"20",X"CD",X"D8",X"17",X"21",
		X"F3",X"43",X"7E",X"B7",X"C8",X"23",X"7E",X"E6",X"01",X"C6",X"ED",X"6F",X"CD",X"19",X"3C",X"C3",
		X"00",X"21",X"2B",X"34",X"7E",X"FE",X"80",X"C2",X"9F",X"18",X"36",X"00",X"23",X"34",X"C9",X"3D",
		X"0F",X"D8",X"E6",X"7F",X"47",X"2F",X"E6",X"02",X"32",X"9E",X"43",X"3A",X"4A",X"43",X"FE",X"02",
		X"CA",X"CA",X"18",X"FE",X"03",X"CA",X"D0",X"18",X"78",X"E6",X"07",X"C0",X"78",X"0F",X"E6",X"3C",
		X"FE",X"20",X"D0",X"C6",X"E0",X"47",X"2B",X"C3",X"1F",X"13",X"11",X"44",X"41",X"C3",X"D3",X"18",
		X"11",X"64",X"41",X"78",X"E6",X"07",X"C0",X"78",X"E6",X"08",X"C2",X"DC",X"21",X"4F",X"12",X"CD",
		X"83",X"3C",X"79",X"12",X"CD",X"83",X"3C",X"79",X"12",X"C9",X"E1",X"26",X"50",X"36",X"01",X"C9",
		X"00",X"2A",X"A2",X"43",X"36",X"01",X"21",X"34",X"02",X"46",X"0E",X"02",X"7E",X"23",X"B7",X"CA",
		X"09",X"19",X"AE",X"86",X"80",X"47",X"C3",X"FC",X"18",X"23",X"23",X"0D",X"C2",X"FC",X"18",X"78",
		X"AE",X"E6",X"09",X"2A",X"A2",X"43",X"AE",X"3D",X"77",X"4F",X"FE",X"07",X"CA",X"22",X"19",X"F0",
		X"C6",X"02",X"B1",X"E6",X"03",X"D6",X"02",X"77",X"C3",X"2E",X"00",X"00",X"CD",X"BA",X"19",X"CD",
		X"D6",X"1A",X"20",X"E6",X"80",X"07",X"32",X"80",X"43",X"CD",X"BC",X"02",X"3A",X"71",X"43",X"E6",
		X"0F",X"FE",X"08",X"D0",X"CD",X"51",X"1B",X"CD",X"58",X"19",X"CD",X"66",X"19",X"21",X"72",X"43",
		X"11",X"77",X"43",X"0E",X"05",X"C3",X"3C",X"3C",X"21",X"78",X"43",X"7E",X"23",X"4E",X"CD",X"92",
		X"1D",X"0E",X"00",X"C3",X"FA",X"13",X"21",X"72",X"43",X"3A",X"F7",X"43",X"E6",X"08",X"07",X"B6",
		X"47",X"E6",X"F0",X"C6",X"08",X"4F",X"E5",X"C5",X"23",X"7E",X"23",X"4E",X"CD",X"92",X"1D",X"C1",
		X"78",X"07",X"E6",X"0E",X"21",X"8A",X"19",X"C3",X"42",X"09",X"9A",X"19",X"9A",X"19",X"A3",X"19",
		X"A3",X"19",X"A3",X"19",X"AB",X"19",X"AB",X"19",X"B4",X"19",X"CD",X"FA",X"13",X"1B",X"78",X"E6",
		X"F7",X"12",X"C9",X"D5",X"CD",X"FA",X"13",X"D1",X"C3",X"9E",X"19",X"D5",X"CD",X"FA",X"13",X"D1",
		X"13",X"C3",X"9E",X"19",X"CD",X"FA",X"13",X"C3",X"9E",X"19",X"00",X"C9",X"3A",X"F7",X"43",X"E6",
		X"03",X"FE",X"01",X"C0",X"3A",X"F2",X"43",X"E6",X"08",X"C0",X"32",X"99",X"43",X"C9",X"21",X"82",
		X"43",X"7E",X"23",X"B6",X"C8",X"3A",X"F3",X"43",X"B7",X"C2",X"F3",X"19",X"06",X"10",X"3A",X"F7",
		X"43",X"E6",X"04",X"CA",X"E8",X"19",X"06",X"20",X"3A",X"71",X"43",X"A0",X"C8",X"21",X"9A",X"43",
		X"C3",X"06",X"1A",X"3A",X"F2",X"43",X"E6",X"08",X"21",X"99",X"43",X"B7",X"C2",X"01",X"1A",X"77",
		X"C9",X"35",X"F0",X"36",X"02",X"23",X"7E",X"23",X"B6",X"C8",X"EB",X"CD",X"BD",X"1A",X"D8",X"E5",
		X"E5",X"EB",X"CD",X"19",X"3C",X"CD",X"EB",X"21",X"E1",X"11",X"72",X"43",X"1A",X"E6",X"07",X"4F",
		X"F6",X"20",X"77",X"13",X"23",X"20",X"1A",X"77",X"13",X"23",X"1A",X"77",X"23",X"79",X"E6",X"01",
		X"3C",X"77",X"3E",X"05",X"32",X"87",X"43",X"E1",X"79",X"D6",X"02",X"FE",X"03",X"D8",X"3C",X"FE",
		X"05",X"D2",X"4C",X"1A",X"B7",X"CA",X"49",X"1A",X"23",X"23",X"34",X"C9",X"AF",X"32",X"97",X"43",
		X"E5",X"7E",X"E6",X"07",X"4F",X"07",X"23",X"EB",X"21",X"E9",X"16",X"CD",X"9D",X"02",X"1A",X"86",
		X"3C",X"FA",X"86",X"1A",X"FE",X"1A",X"D2",X"86",X"1A",X"23",X"13",X"1A",X"86",X"3C",X"FA",X"B0",
		X"1A",X"FE",X"1B",X"D2",X"B0",X"1A",X"3D",X"12",X"2B",X"1B",X"1A",X"86",X"12",X"13",X"13",X"1A",
		X"E1",X"B7",X"F0",X"36",X"00",X"C9",X"E1",X"79",X"B7",X"1F",X"D2",X"B8",X"1A",X"3E",X"02",X"A9",
		X"E6",X"07",X"F6",X"20",X"77",X"3A",X"97",X"43",X"B7",X"C2",X"A9",X"1A",X"7E",X"32",X"97",X"43",
		X"E5",X"23",X"23",X"23",X"35",X"E1",X"C3",X"50",X"1A",X"BE",X"C2",X"50",X"1A",X"36",X"00",X"C9",
		X"E1",X"79",X"1F",X"3E",X"06",X"DA",X"8F",X"1A",X"3E",X"04",X"C3",X"8F",X"1A",X"21",X"54",X"4B",
		X"7E",X"B7",X"C8",X"7D",X"C6",X"05",X"6F",X"FE",X"90",X"DA",X"C0",X"1A",X"37",X"C9",X"2A",X"D7",
		X"1A",X"23",X"22",X"E3",X"47",X"36",X"21",X"6D",X"43",X"34",X"7E",X"23",X"3A",X"F1",X"43",X"77",
		X"23",X"3A",X"AC",X"43",X"77",X"2B",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"E5",X"21",X"26",
		X"1B",X"CD",X"9D",X"02",X"46",X"21",X"7C",X"43",X"4E",X"E1",X"23",X"7E",X"E6",X"01",X"80",X"FE",
		X"08",X"CA",X"05",X"1B",X"81",X"47",X"3A",X"F3",X"43",X"B7",X"C2",X"3E",X"1B",X"2A",X"75",X"43",
		X"46",X"23",X"7E",X"FE",X"80",X"CA",X"3E",X"1B",X"22",X"75",X"43",X"DA",X"3E",X"1B",X"3D",X"CC",
		X"82",X"17",X"C2",X"6A",X"01",X"36",X"08",X"05",X"00",X"06",X"04",X"04",X"08",X"07",X"01",X"08",
		X"00",X"08",X"02",X"08",X"07",X"08",X"ED",X"56",X"FB",X"76",X"CD",X"CE",X"1A",X"C9",X"21",X"71",
		X"43",X"4E",X"70",X"2B",X"79",X"E6",X"0F",X"FE",X"08",X"D8",X"34",X"3E",X"01",X"BE",X"D0",X"77",
		X"C9",X"21",X"82",X"43",X"7E",X"B7",X"C2",X"68",X"1B",X"23",X"B6",X"C8",X"7E",X"FE",X"03",X"D2",
		X"68",X"1B",X"2B",X"2B",X"7E",X"E6",X"02",X"C8",X"21",X"72",X"43",X"7E",X"E6",X"E0",X"47",X"20",
		X"3A",X"71",X"43",X"E6",X"0F",X"FE",X"08",X"D0",X"4F",X"B0",X"77",X"23",X"EB",X"21",X"70",X"43",
		X"7E",X"35",X"B7",X"C0",X"77",X"AF",X"32",X"97",X"43",X"D5",X"79",X"07",X"21",X"E9",X"16",X"CD",
		X"9D",X"02",X"1A",X"86",X"FA",X"BA",X"1B",X"FE",X"17",X"D2",X"CC",X"1B",X"13",X"23",X"1A",X"86",
		X"FA",X"D6",X"1B",X"FE",X"18",X"D2",X"E1",X"1B",X"1B",X"2B",X"CD",X"1C",X"1C",X"C2",X"FC",X"1B",
		X"1A",X"86",X"12",X"13",X"23",X"1A",X"86",X"12",X"D1",X"C9",X"D1",X"CD",X"EC",X"1B",X"79",X"D6",
		X"04",X"C8",X"32",X"97",X"43",X"81",X"E6",X"07",X"4F",X"C3",X"89",X"1B",X"D1",X"CD",X"EC",X"1B",
		X"79",X"B7",X"C8",X"C3",X"C2",X"1B",X"D1",X"CD",X"EC",X"1B",X"79",X"D6",X"02",X"C8",X"C3",X"C2",
		X"1B",X"D1",X"CD",X"EC",X"1B",X"79",X"D6",X"06",X"C8",X"C3",X"C2",X"1B",X"79",X"0F",X"DA",X"F3",
		X"1B",X"E1",X"C9",X"3A",X"97",X"43",X"B7",X"C8",X"E1",X"C3",X"C2",X"1B",X"D1",X"67",X"79",X"07",
		X"07",X"07",X"07",X"84",X"21",X"FD",X"16",X"CD",X"9D",X"02",X"3A",X"97",X"43",X"B7",X"C0",X"7E",
		X"B7",X"C8",X"CD",X"6F",X"3C",X"FE",X"03",X"D0",X"7E",X"C3",X"C2",X"1B",X"E5",X"D5",X"C5",X"CD",
		X"26",X"1C",X"C1",X"D1",X"E1",X"C9",X"13",X"23",X"1A",X"86",X"4F",X"1B",X"2B",X"1A",X"86",X"CD",
		X"92",X"1D",X"21",X"00",X"08",X"19",X"EB",X"1A",X"47",X"13",X"1A",X"4F",X"CD",X"83",X"3C",X"1A",
		X"67",X"1B",X"1A",X"6F",X"B4",X"B0",X"B1",X"C8",X"CD",X"68",X"1C",X"F5",X"11",X"00",X"CF",X"7A",
		X"91",X"7B",X"17",X"5F",X"7A",X"94",X"7B",X"17",X"5F",X"7A",X"95",X"7B",X"17",X"5F",X"7A",X"90",
		X"7B",X"17",X"5F",X"F1",X"7B",X"3D",X"3C",X"C9",X"16",X"20",X"78",X"92",X"BA",X"D8",X"79",X"92",
		X"BA",X"D8",X"7C",X"92",X"BA",X"D8",X"7D",X"92",X"BA",X"C9",X"3A",X"7E",X"43",X"B7",X"C0",X"21",
		X"85",X"43",X"7E",X"B7",X"C2",X"97",X"1C",X"3A",X"F0",X"43",X"07",X"07",X"E6",X"03",X"C6",X"38",
		X"77",X"23",X"36",X"1E",X"C3",X"51",X"1D",X"B7",X"23",X"FA",X"5E",X"1D",X"35",X"2B",X"C2",X"AE",
		X"1C",X"21",X"85",X"43",X"36",X"FF",X"23",X"36",X"00",X"3E",X"00",X"C3",X"51",X"1D",X"3A",X"73",
		X"43",X"B7",X"CA",X"BA",X"1C",X"FE",X"16",X"C2",X"48",X"1D",X"3A",X"74",X"43",X"B7",X"CA",X"C6",
		X"1C",X"FE",X"17",X"C2",X"48",X"1D",X"3E",X"B0",X"32",X"93",X"43",X"7E",X"F6",X"80",X"77",X"23",
		X"36",X"30",X"E6",X"03",X"3C",X"3C",X"07",X"07",X"07",X"07",X"4F",X"06",X"00",X"21",X"9B",X"43",
		X"CD",X"EA",X"3B",X"AF",X"CD",X"51",X"1D",X"2A",X"73",X"43",X"7D",X"4C",X"CD",X"92",X"1D",X"21",
		X"00",X"08",X"19",X"EB",X"3E",X"D1",X"12",X"13",X"12",X"CD",X"83",X"3C",X"3E",X"D1",X"12",X"1B",
		X"12",X"32",X"9C",X"43",X"CD",X"EB",X"21",X"11",X"21",X"42",X"0E",X"04",X"1A",X"B7",X"CA",X"44",
		X"1D",X"CD",X"83",X"3C",X"0D",X"C2",X"0C",X"1D",X"21",X"37",X"1D",X"0E",X"01",X"CD",X"5D",X"02",
		X"21",X"F3",X"43",X"7E",X"B7",X"C8",X"23",X"7E",X"E6",X"01",X"C6",X"ED",X"6F",X"7E",X"C6",X"01",
		X"27",X"77",X"2E",X"88",X"36",X"80",X"C9",X"21",X"42",X"31",X"46",X"52",X"45",X"45",X"20",X"43",
		X"45",X"4C",X"4C",X"00",X"3E",X"4C",X"12",X"C9",X"4E",X"23",X"7E",X"E6",X"02",X"CA",X"51",X"1D",
		X"79",X"32",X"06",X"4B",X"32",X"1E",X"4B",X"32",X"26",X"48",X"32",X"3E",X"48",X"C9",X"7E",X"B7",
		X"C8",X"35",X"01",X"00",X"00",X"CA",X"75",X"1D",X"FE",X"28",X"D0",X"3A",X"85",X"43",X"E6",X"03",
		X"C6",X"32",X"47",X"0E",X"30",X"78",X"32",X"06",X"43",X"32",X"1E",X"43",X"32",X"46",X"40",X"32",
		X"5E",X"40",X"79",X"32",X"E6",X"42",X"32",X"FE",X"42",X"32",X"26",X"40",X"32",X"3E",X"40",X"C9",
		X"C9",X"C9",X"3C",X"07",X"E6",X"3E",X"21",X"A2",X"1D",X"CD",X"9D",X"02",X"7E",X"23",X"56",X"81",
		X"5F",X"C9",X"26",X"43",X"06",X"43",X"E6",X"42",X"C6",X"42",X"A6",X"42",X"86",X"42",X"66",X"42",
		X"46",X"42",X"26",X"42",X"06",X"42",X"E6",X"41",X"C6",X"41",X"A6",X"41",X"86",X"41",X"66",X"41",
		X"46",X"41",X"26",X"41",X"06",X"41",X"E6",X"40",X"C6",X"40",X"A6",X"40",X"86",X"40",X"66",X"40",
		X"46",X"40",X"26",X"40",X"06",X"40",X"26",X"40",X"26",X"40",X"26",X"40",X"26",X"40",X"26",X"40",
		X"26",X"40",X"00",X"21",X"9C",X"43",X"7E",X"B7",X"C8",X"AF",X"32",X"7E",X"43",X"32",X"7D",X"43",
		X"21",X"20",X"4B",X"11",X"00",X"4A",X"01",X"D4",X"D0",X"3A",X"7D",X"43",X"B7",X"CA",X"04",X"1E",
		X"04",X"C3",X"32",X"1E",X"7E",X"B8",X"DA",X"26",X"1E",X"CA",X"1E",X"1E",X"B9",X"DA",X"25",X"1E",
		X"CA",X"18",X"1E",X"FE",X"D5",X"C2",X"26",X"1E",X"32",X"7E",X"43",X"C3",X"26",X"1E",X"32",X"7D",
		X"43",X"04",X"C3",X"51",X"1E",X"73",X"2D",X"C2",X"04",X"1E",X"2B",X"2B",X"7C",X"BA",X"D2",X"04",
		X"1E",X"C9",X"3A",X"7E",X"43",X"B7",X"C2",X"5D",X"1E",X"7E",X"B8",X"DA",X"51",X"1E",X"B9",X"DA",
		X"50",X"1E",X"CA",X"4A",X"1E",X"FE",X"D5",X"C2",X"51",X"1E",X"32",X"7E",X"43",X"C3",X"67",X"1E",
		X"73",X"2D",X"C2",X"39",X"1E",X"2B",X"2B",X"7C",X"BA",X"D2",X"39",X"1E",X"C9",X"7E",X"B8",X"DA",
		X"67",X"1E",X"B9",X"D2",X"67",X"1E",X"73",X"2D",X"C2",X"5D",X"1E",X"2B",X"2B",X"7C",X"BA",X"D2",
		X"5D",X"1E",X"C9",X"00",X"CD",X"31",X"2F",X"21",X"9C",X"43",X"7E",X"B7",X"C8",X"21",X"FF",X"49",
		X"11",X"00",X"49",X"C3",X"F6",X"1D",X"00",X"CD",X"19",X"23",X"21",X"9C",X"43",X"7E",X"B7",X"C8",
		X"36",X"00",X"21",X"FF",X"48",X"11",X"00",X"48",X"C3",X"F6",X"1D",X"AF",X"32",X"7E",X"43",X"32",
		X"7D",X"43",X"21",X"20",X"4B",X"11",X"00",X"48",X"C3",X"F6",X"1D",X"0D",X"7D",X"91",X"47",X"7D",
		X"90",X"A9",X"6F",X"EB",X"2A",X"28",X"3E",X"54",X"19",X"EB",X"21",X"62",X"42",X"19",X"7E",X"23",
		X"22",X"A5",X"43",X"C6",X"04",X"77",X"23",X"36",X"00",X"C9",X"21",X"C9",X"41",X"50",X"55",X"53",
		X"48",X"00",X"CB",X"42",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"CB",X"42",X"31",X"20",X"4F",X"52",X"20",X"32",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"2B",X"42",
		X"47",X"41",X"4D",X"45",X"20",X"20",X"4F",X"56",X"45",X"52",X"00",X"20",X"43",X"48",X"49",X"53",
		X"43",X"4F",X"52",X"45",X"20",X"53",X"55",X"52",X"56",X"49",X"56",X"41",X"4C",X"20",X"EC",X"20",
		X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"00",X"21",X"42",X"20",X"52",X"4F",X"43",X"4B",X"2D",
		X"4F",X"4C",X"41",X"20",X"00",X"42",X"42",X"00",X"23",X"43",X"50",X"31",X"2D",X"20",X"20",X"30",
		X"30",X"20",X"E8",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E9",X"20",X"50",X"32",X"2D",
		X"20",X"20",X"30",X"30",X"00",X"24",X"42",X"E3",X"5A",X"41",X"50",X"53",X"2D",X"30",X"30",X"30",
		X"E1",X"00",X"CD",X"F9",X"02",X"AF",X"CD",X"8C",X"1F",X"CD",X"83",X"21",X"21",X"F5",X"43",X"06",
		X"04",X"CD",X"D4",X"3C",X"2E",X"FE",X"36",X"50",X"20",X"E6",X"80",X"07",X"32",X"80",X"43",X"3A",
		X"00",X"78",X"2F",X"E6",X"0C",X"0F",X"0F",X"C6",X"02",X"2B",X"77",X"AF",X"E6",X"02",X"C2",X"4E",
		X"3D",X"3A",X"00",X"78",X"E6",X"80",X"C2",X"8C",X"1F",X"20",X"F3",X"CD",X"12",X"21",X"CD",X"4A",
		X"13",X"CD",X"BC",X"19",X"3A",X"9E",X"43",X"E6",X"02",X"4F",X"3A",X"F4",X"43",X"E6",X"01",X"B1",
		X"32",X"00",X"50",X"3A",X"9D",X"43",X"32",X"00",X"58",X"3A",X"00",X"78",X"E6",X"80",X"CA",X"B9",
		X"1F",X"21",X"F0",X"43",X"CD",X"7D",X"3C",X"3E",X"0F",X"32",X"00",X"68",X"4A",X"21",X"EB",X"43",
		X"3A",X"00",X"78",X"2F",X"E6",X"10",X"BE",X"CA",X"02",X"20",X"77",X"B7",X"2E",X"A9",X"77",X"23",
		X"77",X"23",X"77",X"2E",X"EC",X"77",X"C2",X"55",X"20",X"2E",X"F5",X"77",X"2E",X"ED",X"77",X"23",
		X"77",X"2E",X"F3",X"77",X"23",X"7E",X"E6",X"01",X"C4",X"B8",X"21",X"FF",X"FF",X"F7",X"EF",X"E7",
		X"DF",X"D7",X"2E",X"EC",X"B7",X"CA",X"09",X"20",X"77",X"2E",X"AC",X"46",X"20",X"E6",X"80",X"07",
		X"4F",X"32",X"95",X"43",X"3A",X"00",X"69",X"77",X"23",X"70",X"3A",X"00",X"70",X"2F",X"2E",X"F1",
		X"46",X"77",X"23",X"70",X"2E",X"AC",X"3A",X"00",X"69",X"BE",X"C2",X"09",X"20",X"3A",X"F1",X"43",
		X"E6",X"01",X"4F",X"78",X"2F",X"A1",X"C8",X"2E",X"EC",X"7E",X"FE",X"99",X"C2",X"49",X"20",X"21",
		X"0E",X"68",X"75",X"24",X"7E",X"E6",X"FE",X"77",X"C9",X"F5",X"01",X"01",X"00",X"CD",X"EA",X"3B",
		X"F1",X"B7",X"C2",X"B3",X"20",X"3A",X"F3",X"43",X"B7",X"C0",X"CD",X"F9",X"02",X"CD",X"F1",X"02",
		X"21",X"0B",X"1F",X"0E",X"05",X"CD",X"5D",X"02",X"11",X"C2",X"42",X"01",X"58",X"50",X"CD",X"9A",
		X"19",X"11",X"62",X"40",X"01",X"58",X"54",X"CD",X"A3",X"19",X"CD",X"DC",X"21",X"11",X"25",X"43",
		X"01",X"18",X"19",X"D5",X"C5",X"C5",X"CD",X"83",X"3C",X"06",X"E0",X"CD",X"26",X"3D",X"EB",X"36",
		X"E5",X"23",X"C1",X"48",X"06",X"E3",X"CD",X"76",X"3C",X"36",X"E7",X"C1",X"E1",X"36",X"E4",X"23",
		X"C5",X"48",X"06",X"E1",X"CD",X"76",X"3C",X"36",X"E6",X"EB",X"CD",X"83",X"3C",X"C1",X"06",X"E2",
		X"C3",X"26",X"3D",X"21",X"EC",X"43",X"11",X"41",X"40",X"20",X"C3",X"A5",X"3C",X"21",X"AE",X"43",
		X"06",X"06",X"CD",X"D4",X"3C",X"3A",X"78",X"00",X"32",X"A4",X"43",X"21",X"45",X"43",X"AF",X"77",
		X"23",X"77",X"23",X"77",X"21",X"B0",X"43",X"11",X"64",X"42",X"CD",X"B4",X"3C",X"21",X"B3",X"43",
		X"11",X"04",X"40",X"CD",X"B4",X"3C",X"C3",X"40",X"31",X"3A",X"00",X"78",X"2F",X"E6",X"03",X"C6",
		X"02",X"21",X"ED",X"43",X"77",X"23",X"77",X"3A",X"F3",X"43",X"D6",X"01",X"C2",X"00",X"21",X"77",
		X"21",X"ED",X"43",X"11",X"63",X"42",X"CD",X"A5",X"3C",X"21",X"EE",X"43",X"11",X"03",X"40",X"C3",
		X"A5",X"3C",X"00",X"3A",X"F3",X"43",X"B7",X"C8",X"CD",X"3E",X"32",X"3A",X"F5",X"43",X"E6",X"07",
		X"FE",X"04",X"D8",X"21",X"47",X"43",X"4E",X"2B",X"46",X"2B",X"7E",X"B0",X"B1",X"C8",X"EB",X"3A",
		X"F4",X"43",X"E6",X"01",X"6F",X"07",X"85",X"21",X"B0",X"43",X"85",X"6F",X"CD",X"EA",X"3B",X"1A",
		X"E6",X"0F",X"47",X"1A",X"E6",X"F0",X"4F",X"AF",X"12",X"13",X"12",X"13",X"12",X"CD",X"EA",X"3B",
		X"E5",X"CD",X"D4",X"20",X"E1",X"11",X"FD",X"43",X"1A",X"FE",X"10",X"D0",X"13",X"13",X"CD",X"DC",
		X"3C",X"D0",X"20",X"21",X"F4",X"43",X"7E",X"E6",X"01",X"C6",X"ED",X"6F",X"7E",X"FE",X"10",X"D2",
		X"7A",X"21",X"C6",X"01",X"27",X"77",X"2E",X"88",X"36",X"80",X"01",X"50",X"03",X"21",X"FE",X"43",
		X"C3",X"EA",X"3B",X"11",X"06",X"43",X"01",X"18",X"19",X"26",X"00",X"C3",X"3B",X"3D",X"00",X"34",
		X"2B",X"7E",X"36",X"00",X"FE",X"02",X"C8",X"77",X"2B",X"7E",X"FE",X"01",X"C8",X"23",X"7E",X"B7",
		X"C2",X"B3",X"21",X"3A",X"EE",X"43",X"B7",X"C8",X"3E",X"01",X"32",X"F4",X"43",X"01",X"01",X"00",
		X"C3",X"BF",X"21",X"3A",X"ED",X"43",X"B7",X"C8",X"AF",X"32",X"F4",X"43",X"01",X"00",X"01",X"21",
		X"00",X"50",X"11",X"A4",X"43",X"70",X"1A",X"71",X"12",X"1C",X"7B",X"FE",X"F7",X"C2",X"C5",X"21",
		X"11",X"E0",X"4B",X"70",X"1A",X"71",X"12",X"20",X"1C",X"C2",X"D3",X"21",X"CD",X"40",X"31",X"CD",
		X"B3",X"20",X"CD",X"D4",X"20",X"CD",X"00",X"21",X"CD",X"91",X"1D",X"11",X"24",X"41",X"21",X"9B",
		X"43",X"C3",X"AA",X"3C",X"3D",X"22",X"8C",X"24",X"14",X"24",X"77",X"25",X"11",X"26",X"F7",X"26",
		X"48",X"24",X"A0",X"26",X"3A",X"F3",X"43",X"B7",X"C8",X"21",X"11",X"22",X"0E",X"01",X"C3",X"5D",
		X"02",X"CB",X"42",X"43",X"41",X"4E",X"20",X"59",X"4F",X"55",X"20",X"44",X"4F",X"20",X"5A",X"41",
		X"50",X"20",X"41",X"4C",X"4C",X"3F",X"00",X"11",X"EB",X"42",X"01",X"16",X"00",X"C3",X"26",X"3D",
		X"3A",X"F3",X"43",X"B7",X"C8",X"CD",X"83",X"21",X"AF",X"32",X"9E",X"43",X"C9",X"E6",X"29",X"4B",
		X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"5E",X"2E",X"5E",
		X"2E",X"5E",X"2E",X"0C",X"2E",X"0C",X"2E",X"0C",X"2E",X"5E",X"2E",X"5E",X"2E",X"5E",X"2E",X"4B",
		X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"E6",X"29",X"4B",
		X"23",X"00",X"CD",X"EE",X"22",X"21",X"6D",X"43",X"7E",X"34",X"F5",X"F5",X"B7",X"CC",X"30",X"22",
		X"F1",X"3C",X"CD",X"A1",X"23",X"F1",X"4F",X"3A",X"6C",X"43",X"B7",X"79",X"CA",X"97",X"22",X"FE",
		X"C9",X"DA",X"63",X"23",X"FE",X"D0",X"D8",X"FE",X"E4",X"D8",X"21",X"7C",X"43",X"22",X"A2",X"43",
		X"2E",X"7D",X"36",X"D0",X"2E",X"6C",X"7E",X"B7",X"CA",X"E1",X"22",X"3A",X"00",X"78",X"2F",X"E6",
		X"10",X"CA",X"E1",X"22",X"3A",X"00",X"70",X"2F",X"E6",X"02",X"CA",X"E1",X"22",X"2E",X"6D",X"35",
		X"2E",X"8B",X"7E",X"B7",X"C0",X"2E",X"97",X"34",X"C0",X"2E",X"6D",X"36",X"00",X"2E",X"41",X"7E",
		X"C6",X"FF",X"9F",X"E6",X"07",X"2B",X"86",X"3C",X"2E",X"8B",X"77",X"CD",X"F9",X"02",X"C3",X"E6",
		X"2E",X"21",X"F5",X"43",X"34",X"2E",X"6D",X"36",X"00",X"2E",X"6C",X"36",X"00",X"C9",X"11",X"21",
		X"42",X"01",X"05",X"00",X"1A",X"FE",X"4C",X"CA",X"02",X"23",X"3A",X"F3",X"43",X"B7",X"C8",X"CD",
		X"26",X"3D",X"21",X"13",X"23",X"0E",X"01",X"CD",X"5D",X"02",X"11",X"01",X"41",X"21",X"44",X"43",
		X"C3",X"A5",X"3C",X"81",X"41",X"20",X"20",X"23",X"00",X"00",X"11",X"4B",X"00",X"3A",X"F5",X"43",
		X"B0",X"47",X"21",X"FA",X"00",X"07",X"81",X"4F",X"E5",X"EB",X"19",X"D1",X"80",X"47",X"4E",X"3E",
		X"3E",X"77",X"50",X"59",X"AE",X"48",X"73",X"5F",X"21",X"EF",X"43",X"7E",X"23",X"AE",X"E6",X"2C",
		X"C0",X"E1",X"7B",X"E6",X"08",X"C8",X"EB",X"D5",X"E5",X"D1",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C6",X"38",X"32",X"9D",X"43",X"F5",X"FE",X"38",X"CC",X"04",X"22",X"F1",X"F5",
		X"FE",X"D4",X"CC",X"27",X"22",X"F1",X"E6",X"07",X"C0",X"3E",X"40",X"32",X"97",X"43",X"3A",X"40",
		X"43",X"07",X"E6",X"0E",X"21",X"F4",X"21",X"CD",X"8D",X"02",X"79",X"0F",X"0F",X"4F",X"E6",X"3E",
		X"CD",X"8D",X"02",X"11",X"06",X"4B",X"79",X"0F",X"E6",X"1F",X"83",X"5F",X"0E",X"18",X"C3",X"30",
		X"3D",X"F5",X"3A",X"F4",X"43",X"B7",X"C2",X"B8",X"23",X"11",X"C2",X"42",X"01",X"58",X"50",X"F1",
		X"E6",X"0F",X"CA",X"9A",X"19",X"C3",X"C4",X"23",X"11",X"62",X"40",X"01",X"58",X"54",X"F1",X"E6",
		X"0F",X"CA",X"A3",X"19",X"FE",X"08",X"C0",X"0E",X"00",X"C3",X"FA",X"13",X"E5",X"21",X"F5",X"43",
		X"B6",X"C0",X"3A",X"00",X"34",X"06",X"20",X"21",X"4A",X"43",X"CD",X"D4",X"3C",X"2E",X"7F",X"7E",
		X"E6",X"E0",X"77",X"CD",X"30",X"22",X"CD",X"7D",X"20",X"3E",X"C0",X"32",X"A8",X"43",X"20",X"3A",
		X"40",X"43",X"07",X"E6",X"0E",X"21",X"7C",X"24",X"CD",X"8D",X"02",X"11",X"40",X"4B",X"3A",X"42",
		X"43",X"4F",X"B7",X"07",X"07",X"81",X"4F",X"CD",X"3C",X"3C",X"AF",X"12",X"13",X"7B",X"FE",X"E0",
		X"DA",X"0A",X"24",X"C9",X"9A",X"03",X"24",X"04",X"4B",X"03",X"63",X"03",X"C5",X"05",X"BA",X"06",
		X"06",X"28",X"1E",X"28",X"D2",X"06",X"E3",X"0F",X"EA",X"06",X"34",X"07",X"34",X"07",X"EA",X"06",
		X"E3",X"0F",X"D2",X"06",X"1E",X"28",X"06",X"28",X"BA",X"06",X"C5",X"05",X"63",X"03",X"4B",X"03",
		X"4B",X"23",X"24",X"04",X"4C",X"07",X"4B",X"23",X"12",X"0D",X"2A",X"0D",X"42",X"0D",X"42",X"0D",
		X"42",X"0D",X"12",X"0D",X"B7",X"0D",X"0F",X"0E",X"87",X"0D",X"9F",X"0D",X"9F",X"0D",X"9F",X"0D",
		X"9F",X"0D",X"87",X"0D",X"0F",X"0E",X"B7",X"0D",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4B",X"23",
		X"12",X"0D",X"42",X"0D",X"42",X"0D",X"2A",X"0D",X"12",X"0D",X"4B",X"23",X"C8",X"24",X"C8",X"24",
		X"E1",X"24",X"FA",X"24",X"2C",X"25",X"13",X"25",X"45",X"25",X"5E",X"25",X"9A",X"03",X"24",X"04",
		X"3C",X"04",X"96",X"04",X"4A",X"26",X"AE",X"04",X"C6",X"04",X"AE",X"04",X"95",X"05",X"47",X"27",
		X"3C",X"04",X"47",X"27",X"5F",X"27",X"AE",X"04",X"C6",X"04",X"AE",X"04",X"95",X"05",X"AE",X"04",
		X"AD",X"05",X"AE",X"04",X"4A",X"26",X"96",X"04",X"33",X"03",X"24",X"04",X"9A",X"03",X"4B",X"23",
		X"21",X"00",X"00",X"39",X"22",X"00",X"44",X"21",X"7B",X"16",X"02",X"00",X"08",X"9D",X"16",X"06",
		X"00",X"1E",X"BD",X"16",X"0A",X"00",X"2D",X"DD",X"16",X"0E",X"00",X"3C",X"7B",X"16",X"15",X"00",
		X"4B",X"7B",X"16",X"02",X"00",X"08",X"9D",X"16",X"06",X"00",X"1E",X"BD",X"16",X"0A",X"00",X"2D",
		X"DD",X"16",X"0E",X"00",X"3C",X"7B",X"16",X"15",X"00",X"4B",X"7B",X"16",X"02",X"00",X"08",X"9D",
		X"16",X"06",X"00",X"1E",X"BD",X"05",X"0D",X"00",X"2D",X"DD",X"16",X"0E",X"00",X"3C",X"7B",X"05",
		X"05",X"00",X"4B",X"7E",X"06",X"00",X"00",X"08",X"9E",X"0A",X"00",X"00",X"1E",X"BE",X"0E",X"00",
		X"00",X"2D",X"DF",X"03",X"0D",X"00",X"3C",X"9D",X"0A",X"0D",X"00",X"4B",X"7B",X"0A",X"05",X"00",
		X"08",X"9D",X"16",X"06",X"00",X"0C",X"BD",X"0A",X"12",X"00",X"10",X"DD",X"16",X"0E",X"00",X"14",
		X"DC",X"07",X"0B",X"00",X"1C",X"7B",X"16",X"02",X"00",X"08",X"9D",X"0B",X"0A",X"00",X"0C",X"BD",
		X"16",X"0A",X"00",X"10",X"DD",X"16",X"0E",X"00",X"14",X"DB",X"02",X"02",X"00",X"1C",X"7B",X"16",
		X"02",X"00",X"08",X"9D",X"16",X"06",X"00",X"0C",X"BD",X"16",X"0A",X"00",X"10",X"DD",X"16",X"0E",
		X"00",X"14",X"9B",X"01",X"14",X"00",X"1C",X"4C",X"07",X"24",X"04",X"4B",X"23",X"4B",X"23",X"64",
		X"07",X"96",X"07",X"AF",X"07",X"C7",X"07",X"64",X"07",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"49",
		X"09",X"96",X"07",X"AF",X"07",X"C7",X"07",X"49",X"09",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"61",
		X"09",X"61",X"09",X"80",X"09",X"B8",X"09",X"4C",X"07",X"4B",X"23",X"00",X"34",X"3A",X"F3",X"43",
		X"B7",X"C2",X"C0",X"25",X"2A",X"26",X"08",X"22",X"EF",X"43",X"2A",X"24",X"08",X"22",X"F7",X"43",
		X"3A",X"AC",X"43",X"32",X"6F",X"43",X"3A",X"F1",X"43",X"32",X"6E",X"43",X"AF",X"32",X"86",X"43",
		X"21",X"9A",X"43",X"7E",X"B7",X"C2",X"E3",X"25",X"23",X"3E",X"50",X"BE",X"DA",X"E3",X"25",X"77",
		X"CD",X"EB",X"21",X"21",X"82",X"43",X"7E",X"B7",X"C2",X"FA",X"25",X"23",X"3E",X"25",X"BE",X"DA",
		X"FA",X"25",X"77",X"2B",X"2B",X"36",X"07",X"CD",X"91",X"1D",X"21",X"45",X"26",X"E5",X"11",X"71",
		X"43",X"0E",X"05",X"3E",X"08",X"12",X"13",X"20",X"CD",X"3C",X"3C",X"E1",X"0E",X"05",X"C3",X"3C",
		X"3C",X"9B",X"28",X"B3",X"28",X"39",X"0B",X"51",X"0B",X"69",X"0B",X"6C",X"0C",X"6C",X"0C",X"69",
		X"0B",X"51",X"0B",X"39",X"0B",X"84",X"0C",X"4B",X"23",X"9C",X"0C",X"4B",X"23",X"84",X"0C",X"39",
		X"0B",X"51",X"0B",X"69",X"0B",X"6C",X"0C",X"6C",X"0C",X"69",X"0B",X"51",X"0B",X"39",X"0B",X"B3",
		X"28",X"9B",X"28",X"4B",X"23",X"42",X"00",X"0A",X"28",X"08",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2E",X"F4",X"7E",X"E6",X"01",X"C6",X"ED",X"6F",X"7E",X"B7",X"C2",X"2E",X"27",
		X"2E",X"F6",X"7E",X"FE",X"FF",X"CA",X"2B",X"27",X"34",X"FE",X"20",X"DA",X"02",X"18",X"C2",X"D4",
		X"26",X"34",X"2E",X"8B",X"36",X"0F",X"CD",X"30",X"22",X"21",X"FE",X"1E",X"0E",X"01",X"CD",X"5D",
		X"02",X"3A",X"F3",X"43",X"B7",X"C8",X"AF",X"21",X"AB",X"43",X"77",X"2B",X"77",X"2B",X"77",X"D0",
		X"9A",X"03",X"A6",X"29",X"BE",X"29",X"E2",X"28",X"FA",X"28",X"12",X"29",X"2A",X"29",X"27",X"0E",
		X"3F",X"0E",X"74",X"0E",X"8C",X"0E",X"A4",X"0E",X"17",X"0F",X"2F",X"0F",X"47",X"0F",X"5F",X"0F",
		X"81",X"0F",X"99",X"0F",X"B1",X"0F",X"8E",X"29",X"4B",X"23",X"4B",X"23",X"4B",X"23",X"4C",X"07",
		X"4C",X"07",X"4B",X"23",X"FE",X"F0",X"D8",X"C2",X"EE",X"26",X"35",X"E5",X"2E",X"50",X"7E",X"34",
		X"F5",X"CD",X"77",X"27",X"F1",X"E1",X"D6",X"C0",X"D8",X"32",X"50",X"43",X"34",X"C9",X"35",X"3A",
		X"8B",X"43",X"B7",X"F8",X"36",X"FF",X"C9",X"D0",X"09",X"E8",X"09",X"10",X"0A",X"4B",X"23",X"44",
		X"28",X"5C",X"28",X"28",X"0A",X"40",X"0A",X"78",X"0A",X"90",X"0A",X"A8",X"0A",X"90",X"0A",X"78",
		X"0A",X"40",X"0A",X"28",X"0A",X"5C",X"28",X"44",X"28",X"4B",X"23",X"D0",X"0A",X"E8",X"0A",X"00",
		X"0B",X"E8",X"0A",X"83",X"28",X"24",X"04",X"4C",X"07",X"4B",X"23",X"CD",X"D8",X"2F",X"21",X"F5",
		X"43",X"34",X"23",X"AF",X"77",X"20",X"21",X"ED",X"43",X"7E",X"23",X"B6",X"C0",X"2E",X"F3",X"77",
		X"23",X"7E",X"B7",X"C2",X"B8",X"21",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"FE",X"80",X"D0",X"1F",X"D8",X"1F",X"D8",X"E6",X"1F",
		X"F5",X"21",X"AE",X"43",X"3A",X"F4",X"43",X"E6",X"01",X"4F",X"07",X"81",X"85",X"6F",X"7E",X"0E",
		X"00",X"E6",X"F0",X"CA",X"9F",X"27",X"0E",X"0A",X"D6",X"10",X"CA",X"9F",X"27",X"0E",X"14",X"7E",
		X"E6",X"0F",X"81",X"D6",X"02",X"D2",X"AA",X"27",X"3E",X"00",X"FE",X"11",X"DA",X"B1",X"27",X"3E",
		X"10",X"C1",X"4F",X"90",X"DA",X"CB",X"28",X"78",X"B7",X"C2",X"F8",X"27",X"C5",X"CD",X"F9",X"02",
		X"CD",X"83",X"21",X"01",X"04",X"13",X"11",X"CB",X"49",X"21",X"42",X"29",X"CD",X"23",X"3C",X"21",
		X"D6",X"29",X"0E",X"02",X"CD",X"5D",X"02",X"3E",X"38",X"32",X"07",X"4B",X"32",X"27",X"48",X"11",
		X"EB",X"4A",X"0E",X"C8",X"CD",X"FA",X"13",X"11",X"CE",X"4A",X"0E",X"C8",X"CD",X"FA",X"13",X"0E",
		X"28",X"11",X"DC",X"48",X"CD",X"FA",X"13",X"C1",X"48",X"21",X"BA",X"49",X"0D",X"FA",X"36",X"28",
		X"36",X"C2",X"2B",X"C3",X"FC",X"27",X"00",X"00",X"D4",X"00",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",
		X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"00",X"D4",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",
		X"D4",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",
		X"D4",X"00",X"D4",X"00",X"00",X"00",X"48",X"21",X"9A",X"49",X"0D",X"FA",X"74",X"28",X"36",X"C3",
		X"2B",X"C3",X"3A",X"28",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"78",X"FE",X"10",X"D8",X"3E",X"C6",X"32",X"AB",X"49",X"3E",X"C7",X"32",
		X"8B",X"49",X"C9",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",X"D5",X"D5",X"D0",
		X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"D5",X"D5",X"D5",
		X"D0",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"D0",X"D5",X"D5",X"D5",X"D0",X"D5",
		X"D5",X"D0",X"00",X"D0",X"00",X"00",X"00",X"00",X"D4",X"00",X"D0",X"D0",X"00",X"00",X"00",X"D0",
		X"D0",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"08",X"D8",X"21",X"FE",
		X"29",X"3A",X"BA",X"43",X"E6",X"10",X"CA",X"DC",X"28",X"21",X"7B",X"2B",X"11",X"C7",X"42",X"C3",
		X"69",X"02",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",
		X"D5",X"D5",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"D0",X"00",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"D0",X"00",X"00",X"00",X"D0",X"D4",X"00",X"00",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D6",X"D7",X"D8",X"DE",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C4",X"3F",X"D9",X"DF",X"C1",X"C1",X"C1",X"C1",X"C1",X"C1",X"C1",
		X"C1",X"C1",X"C1",X"C1",X"C1",X"C1",X"C1",X"C1",X"C5",X"3F",X"DA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"DC",X"DD",X"D0",X"D5",
		X"D5",X"D5",X"D5",X"D5",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D5",X"D5",X"D5",X"D5",
		X"D5",X"D5",X"D0",X"D0",X"D5",X"D0",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D5",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D0",X"00",X"00",X"D0",X"D5",X"D5",X"D5",X"D5",X"D5",
		X"D5",X"D5",X"D0",X"00",X"00",X"00",X"9A",X"42",X"49",X"2E",X"43",X"2E",X"55",X"2E",X"00",X"52",
		X"41",X"33",X"38",X"25",X"43",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"20",X"56",
		X"49",X"54",X"41",X"4C",X"20",X"53",X"49",X"47",X"4E",X"53",X"20",X"47",X"4F",X"4F",X"44",X"21",
		X"21",X"00",X"57",X"45",X"41",X"4B",X"20",X"42",X"55",X"54",X"20",X"49",X"4D",X"50",X"52",X"4F",
		X"56",X"49",X"4E",X"47",X"21",X"21",X"00",X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"20",X"42",X"55",
		X"54",X"20",X"54",X"52",X"59",X"20",X"48",X"41",X"52",X"44",X"45",X"52",X"00",X"4D",X"45",X"44",
		X"49",X"43",X"41",X"54",X"49",X"4F",X"4E",X"20",X"45",X"46",X"46",X"45",X"43",X"54",X"49",X"56",
		X"45",X"21",X"00",X"4F",X"2E",X"4B",X"2E",X"20",X"54",X"4F",X"20",X"50",X"4C",X"41",X"59",X"20",
		X"53",X"50",X"4F",X"52",X"54",X"53",X"21",X"00",X"20",X"44",X"4F",X"49",X"4E",X"47",X"20",X"4D",
		X"55",X"43",X"48",X"20",X"42",X"45",X"54",X"54",X"45",X"52",X"21",X"00",X"4D",X"55",X"43",X"48",
		X"20",X"49",X"4D",X"50",X"52",X"4F",X"56",X"45",X"44",X"20",X"41",X"43",X"54",X"49",X"4F",X"4E",
		X"21",X"00",X"20",X"47",X"4F",X"4F",X"44",X"20",X"43",X"4F",X"4F",X"52",X"44",X"49",X"4E",X"41",
		X"54",X"49",X"4F",X"4E",X"21",X"21",X"00",X"20",X"4E",X"49",X"43",X"45",X"20",X"52",X"45",X"54",
		X"55",X"52",X"4E",X"20",X"50",X"4C",X"41",X"59",X"53",X"21",X"21",X"00",X"46",X"45",X"45",X"4C",
		X"49",X"4E",X"47",X"20",X"50",X"52",X"45",X"54",X"54",X"59",X"20",X"47",X"4F",X"4F",X"44",X"3F",
		X"00",X"59",X"4F",X"55",X"27",X"4C",X"4C",X"20",X"4D",X"41",X"4B",X"45",X"20",X"49",X"54",X"20",
		X"53",X"4F",X"4F",X"4E",X"21",X"00",X"57",X"41",X"54",X"43",X"48",X"20",X"59",X"4F",X"55",X"52",
		X"20",X"42",X"41",X"43",X"4B",X"48",X"41",X"4E",X"44",X"21",X"00",X"20",X"56",X"45",X"52",X"59",
		X"20",X"47",X"4F",X"4F",X"44",X"20",X"48",X"45",X"41",X"4C",X"54",X"48",X"21",X"21",X"00",X"45",
		X"58",X"43",X"45",X"4C",X"4C",X"45",X"4E",X"54",X"20",X"43",X"4F",X"4E",X"44",X"49",X"54",X"49",
		X"4F",X"4E",X"21",X"00",X"53",X"55",X"50",X"45",X"52",X"42",X"20",X"50",X"45",X"52",X"46",X"4F",
		X"52",X"4D",X"41",X"4E",X"43",X"45",X"21",X"21",X"00",X"20",X"55",X"4E",X"42",X"45",X"4C",X"49",
		X"45",X"56",X"41",X"42",X"4C",X"59",X"20",X"47",X"4F",X"4F",X"44",X"21",X"21",X"00",X"20",X"53",
		X"55",X"50",X"45",X"52",X"20",X"48",X"4F",X"54",X"2D",X"53",X"48",X"4F",X"54",X"21",X"21",X"21",
		X"21",X"21",X"00",X"00",X"00",X"05",X"00",X"00",X"06",X"00",X"05",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"05",X"00",X"11",X"13",X"14",X"15",X"05",X"00",X"00",X"43",X"4F",X"4C",X"44",X"20",
		X"42",X"55",X"54",X"20",X"49",X"4D",X"50",X"52",X"4F",X"56",X"49",X"4E",X"47",X"21",X"21",X"00",
		X"55",X"4E",X"55",X"53",X"55",X"41",X"4C",X"20",X"48",X"45",X"41",X"52",X"54",X"20",X"54",X"48",
		X"52",X"4F",X"42",X"3F",X"00",X"47",X"4F",X"4F",X"44",X"20",X"45",X"58",X"45",X"52",X"43",X"49",
		X"53",X"45",X"20",X"54",X"4F",X"44",X"41",X"59",X"21",X"00",X"4D",X"41",X"4B",X"49",X"4E",X"47",
		X"20",X"47",X"4F",X"4F",X"44",X"20",X"50",X"52",X"4F",X"47",X"52",X"45",X"53",X"53",X"21",X"00",
		X"43",X"4F",X"4D",X"49",X"4E",X"47",X"20",X"41",X"4C",X"4F",X"4E",X"47",X"20",X"4E",X"49",X"43",
		X"45",X"4C",X"59",X"21",X"00",X"41",X"42",X"4F",X"55",X"54",X"20",X"4E",X"4F",X"52",X"4D",X"41",
		X"4C",X"20",X"48",X"45",X"41",X"4C",X"54",X"48",X"21",X"00",X"4B",X"45",X"45",X"50",X"20",X"55",
		X"50",X"20",X"54",X"48",X"45",X"20",X"47",X"4F",X"4F",X"44",X"20",X"57",X"4F",X"52",X"4B",X"00",
		X"53",X"48",X"4F",X"57",X"49",X"4E",X"47",X"20",X"4D",X"55",X"43",X"48",X"20",X"54",X"41",X"4C",
		X"45",X"4E",X"54",X"21",X"21",X"00",X"44",X"4F",X"4E",X"27",X"54",X"20",X"43",X"41",X"54",X"43",
		X"48",X"20",X"43",X"4F",X"4C",X"44",X"20",X"4E",X"4F",X"57",X"21",X"00",X"48",X"49",X"47",X"48",
		X"20",X"54",X"45",X"43",X"48",X"4E",X"49",X"51",X"55",X"45",X"20",X"53",X"48",X"4F",X"57",X"4E",
		X"21",X"00",X"57",X"41",X"54",X"43",X"48",X"20",X"59",X"4F",X"55",X"52",X"20",X"52",X"49",X"47",
		X"48",X"54",X"20",X"53",X"49",X"44",X"45",X"00",X"20",X"55",X"53",X"45",X"20",X"4C",X"45",X"53",
		X"53",X"20",X"4D",X"45",X"44",X"49",X"43",X"49",X"4E",X"45",X"21",X"00",X"47",X"4C",X"4F",X"52",
		X"49",X"4F",X"55",X"53",X"20",X"50",X"4C",X"41",X"59",X"2F",X"41",X"43",X"54",X"49",X"4F",X"4E",
		X"21",X"00",X"56",X"45",X"52",X"59",X"20",X"53",X"50",X"49",X"52",X"49",X"54",X"45",X"44",X"20",
		X"41",X"43",X"54",X"49",X"4F",X"4E",X"21",X"00",X"46",X"49",X"4E",X"45",X"20",X"52",X"45",X"43",
		X"4F",X"52",X"44",X"20",X"42",X"52",X"45",X"41",X"4B",X"45",X"52",X"21",X"21",X"00",X"54",X"4F",
		X"50",X"20",X"41",X"43",X"54",X"49",X"4F",X"4E",X"2F",X"42",X"45",X"53",X"54",X"20",X"50",X"4C",
		X"41",X"59",X"21",X"00",X"4F",X"56",X"45",X"52",X"20",X"54",X"48",X"45",X"20",X"54",X"4F",X"50",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"0B",X"00",X"00",X"05",X"00",X"00",X"06",X"00",X"05",X"17",X"18",X"19",X"05",
		X"00",X"00",X"00",X"34",X"AF",X"32",X"6D",X"43",X"3A",X"6C",X"43",X"B7",X"C8",X"35",X"21",X"4F",
		X"43",X"7E",X"B7",X"C2",X"3A",X"2D",X"2B",X"34",X"7E",X"FE",X"30",X"D8",X"CD",X"D8",X"17",X"C3",
		X"42",X"2D",X"00",X"00",X"05",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"05",X"00",
		X"10",X"0F",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"FE",X"02",X"D2",X"7A",X"2D",X"C3",
		X"42",X"2D",X"21",X"4F",X"43",X"34",X"2B",X"36",X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"2E",X"00",X"00",X"1A",X"00",X"00",X"00",X"1A",X"00",X"01",X"03",X"03",X"04",X"00",X"0A",
		X"03",X"03",X"04",X"00",X"01",X"03",X"03",X"04",X"2D",X"2F",X"FE",X"03",X"D2",X"DF",X"2D",X"2B",
		X"34",X"7E",X"FE",X"30",X"D8",X"35",X"21",X"86",X"2E",X"22",X"A0",X"43",X"3E",X"01",X"32",X"9F",
		X"43",X"21",X"9A",X"43",X"7E",X"23",X"B6",X"CA",X"42",X"2D",X"3A",X"84",X"43",X"B7",X"C0",X"CD",
		X"19",X"3C",X"20",X"CD",X"EB",X"21",X"2E",X"84",X"36",X"08",X"2E",X"45",X"36",X"30",X"C9",X"00",
		X"00",X"05",X"00",X"1F",X"00",X"05",X"00",X"05",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"06",
		X"00",X"07",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"1D",X"1E",X"04",X"05",X"00",X"0C",
		X"03",X"03",X"05",X"00",X"0C",X"03",X"0D",X"0E",X"00",X"00",X"02",X"03",X"04",X"00",X"00",X"FE",
		X"04",X"D2",X"CB",X"2E",X"3A",X"43",X"43",X"FE",X"0F",X"CA",X"F0",X"2D",X"2B",X"36",X"FF",X"23",
		X"2B",X"34",X"7E",X"B7",X"C2",X"24",X"2E",X"2E",X"41",X"7E",X"C6",X"FF",X"9F",X"E6",X"07",X"2B",
		X"86",X"3C",X"2E",X"8B",X"77",X"20",X"CD",X"38",X"22",X"C3",X"42",X"2D",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F5",X"3E",X"02",X"32",X"9E",X"43",X"21",X"96",X"2E",X"22",X"A0",X"43",
		X"3E",X"06",X"32",X"9F",X"43",X"21",X"49",X"43",X"11",X"6D",X"41",X"CD",X"AF",X"3C",X"F1",X"FE",
		X"80",X"D8",X"21",X"48",X"43",X"7E",X"B7",X"C8",X"3E",X"80",X"32",X"4E",X"43",X"3A",X"84",X"43",
		X"B7",X"C0",X"CD",X"19",X"3C",X"2B",X"2B",X"34",X"3E",X"08",X"32",X"84",X"43",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3E",X"3E",X"3E",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"42",X"35",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",
		X"53",X"2F",X"53",X"45",X"43",X"00",X"46",X"42",X"33",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",
		X"53",X"2F",X"5A",X"41",X"50",X"00",X"86",X"42",X"49",X"4E",X"53",X"55",X"52",X"41",X"4E",X"43",
		X"45",X"20",X"52",X"45",X"42",X"41",X"54",X"45",X"00",X"E9",X"41",X"42",X"4F",X"4E",X"55",X"53",
		X"00",X"EC",X"41",X"E4",X"E0",X"E0",X"E0",X"E0",X"E5",X"00",X"ED",X"41",X"E1",X"00",X"4D",X"41",
		X"E3",X"00",X"EE",X"41",X"E6",X"E2",X"E2",X"E2",X"E2",X"E7",X"00",X"4F",X"3E",X"02",X"32",X"9E",
		X"43",X"79",X"FE",X"05",X"DA",X"59",X"2F",X"CD",X"38",X"22",X"21",X"F5",X"43",X"34",X"34",X"CD",
		X"1C",X"01",X"AF",X"32",X"9F",X"43",X"21",X"44",X"43",X"01",X"01",X"00",X"CD",X"EA",X"3B",X"2E",
		X"40",X"34",X"7E",X"FE",X"08",X"DA",X"17",X"2F",X"36",X"01",X"23",X"34",X"7E",X"FE",X"02",X"DA",
		X"07",X"2F",X"36",X"01",X"2B",X"36",X"05",X"2E",X"F4",X"7E",X"E6",X"01",X"21",X"22",X"43",X"CA",
		X"15",X"2F",X"21",X"C2",X"40",X"36",X"1E",X"CD",X"82",X"17",X"F5",X"CD",X"AB",X"1E",X"CD",X"38",
		X"22",X"F1",X"CA",X"31",X"2F",X"21",X"96",X"43",X"7E",X"34",X"FE",X"17",X"D8",X"77",X"CA",X"A4",
		X"43",X"00",X"21",X"6F",X"43",X"7E",X"E6",X"01",X"2B",X"7E",X"CA",X"4D",X"2F",X"E6",X"F0",X"CA",
		X"25",X"2F",X"FE",X"20",X"CA",X"25",X"2F",X"FE",X"40",X"CA",X"25",X"2F",X"C9",X"E6",X"F0",X"C8",
		X"FE",X"20",X"C8",X"FE",X"40",X"C2",X"25",X"2F",X"C9",X"2B",X"7E",X"34",X"FE",X"80",X"CA",X"42",
		X"2D",X"0F",X"E6",X"3F",X"4F",X"CD",X"C5",X"2F",X"21",X"B2",X"41",X"79",X"FE",X"0C",X"DA",X"7F",
		X"2F",X"CA",X"AD",X"2F",X"06",X"00",X"D6",X"33",X"4F",X"D8",X"FE",X"0C",X"CA",X"B2",X"2F",X"79",
		X"FE",X"0C",X"D0",X"0F",X"0F",X"0F",X"5F",X"E6",X"1F",X"57",X"7B",X"E6",X"E0",X"5F",X"19",X"7D",
		X"91",X"6F",X"0C",X"79",X"07",X"5F",X"51",X"70",X"2C",X"70",X"2C",X"15",X"C2",X"97",X"2F",X"EB",
		X"7B",X"91",X"91",X"5F",X"CD",X"83",X"3C",X"EB",X"1D",X"C2",X"96",X"2F",X"C9",X"C5",X"CD",X"F9",
		X"02",X"C1",X"11",X"06",X"43",X"0E",X"18",X"C3",X"26",X"3D",X"CD",X"F9",X"02",X"21",X"1F",X"02",
		X"0E",X"02",X"C3",X"5D",X"02",X"3A",X"40",X"43",X"E6",X"03",X"06",X"FE",X"C8",X"06",X"FD",X"3D",
		X"C8",X"06",X"FF",X"3D",X"C8",X"06",X"4C",X"C9",X"3A",X"B4",X"43",X"B7",X"C2",X"44",X"30",X"3A",
		X"F4",X"43",X"E6",X"01",X"4F",X"07",X"81",X"11",X"B0",X"43",X"83",X"5F",X"21",X"BA",X"43",X"01",
		X"01",X"06",X"CD",X"DC",X"3C",X"D2",X"03",X"30",X"78",X"85",X"6F",X"0C",X"79",X"FE",X"0A",X"C2",
		X"F2",X"2F",X"C9",X"D5",X"E5",X"79",X"32",X"B4",X"43",X"21",X"E4",X"43",X"11",X"EA",X"43",X"3E",
		X"09",X"91",X"CA",X"22",X"30",X"07",X"4F",X"07",X"81",X"4F",X"7E",X"12",X"2B",X"1B",X"0D",X"C2",
		X"1A",X"30",X"E1",X"D1",X"1A",X"77",X"2B",X"1B",X"1A",X"77",X"2B",X"1B",X"1A",X"77",X"21",X"5F",
		X"31",X"0E",X"08",X"CD",X"5D",X"02",X"CD",X"F9",X"02",X"AF",X"32",X"EF",X"43",X"3D",X"32",X"6D",
		X"43",X"3A",X"B4",X"43",X"00",X"47",X"B7",X"FA",X"F4",X"30",X"E6",X"0F",X"07",X"4F",X"07",X"81",
		X"21",X"AF",X"43",X"85",X"6F",X"11",X"D2",X"41",X"C5",X"E5",X"D5",X"0E",X"03",X"CD",X"30",X"3D",
		X"D1",X"D5",X"13",X"01",X"03",X"E2",X"CD",X"26",X"3D",X"D1",X"E1",X"C1",X"78",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"03",X"4F",X"85",X"6F",X"0D",X"FA",X"80",X"30",X"CD",X"83",X"3C",X"C3",X"76",X"30",
		X"13",X"3E",X"1E",X"12",X"11",X"F0",X"43",X"1A",X"E6",X"0F",X"C2",X"EE",X"30",X"1B",X"1A",X"FE",
		X"0A",X"D2",X"A5",X"30",X"3A",X"00",X"70",X"2F",X"4F",X"E6",X"08",X"CA",X"B3",X"30",X"3A",X"6D",
		X"43",X"3C",X"CA",X"EE",X"30",X"E1",X"21",X"6D",X"43",X"3E",X"80",X"77",X"2E",X"B4",X"B6",X"77",
		X"C3",X"83",X"21",X"3E",X"F0",X"32",X"6D",X"43",X"79",X"E6",X"40",X"CA",X"C5",X"30",X"78",X"D6",
		X"10",X"DA",X"EE",X"30",X"47",X"79",X"E6",X"20",X"CA",X"D4",X"30",X"78",X"C6",X"10",X"FE",X"30",
		X"D2",X"EE",X"30",X"47",X"79",X"E6",X"80",X"CA",X"E0",X"30",X"7E",X"3D",X"FA",X"EE",X"30",X"77",
		X"79",X"E6",X"10",X"CA",X"EE",X"30",X"7E",X"3C",X"FE",X"1B",X"D2",X"EE",X"30",X"77",X"78",X"32",
		X"B4",X"43",X"E1",X"C9",X"21",X"6D",X"43",X"7E",X"34",X"FE",X"F7",X"DA",X"04",X"31",X"AF",X"77",
		X"32",X"B4",X"43",X"C9",X"E6",X"08",X"C2",X"30",X"31",X"11",X"89",X"42",X"D5",X"21",X"F3",X"3A",
		X"CD",X"76",X"02",X"D1",X"13",X"D5",X"23",X"23",X"CD",X"76",X"02",X"D1",X"1B",X"0E",X"01",X"C5",
		X"D5",X"79",X"CD",X"8A",X"3A",X"D1",X"C1",X"0C",X"79",X"FE",X"0A",X"DA",X"1F",X"31",X"E1",X"C9",
		X"11",X"E9",X"42",X"E1",X"78",X"17",X"E6",X"1E",X"83",X"5F",X"01",X"14",X"00",X"C3",X"26",X"3D",
		X"21",X"BA",X"43",X"11",X"B0",X"43",X"CD",X"DC",X"3C",X"DA",X"4D",X"31",X"EB",X"11",X"B3",X"43",
		X"CD",X"DC",X"3C",X"DA",X"57",X"31",X"EB",X"11",X"61",X"42",X"C3",X"B4",X"3C",X"E5",X"21",X"E7",
		X"42",X"54",X"48",X"41",X"54",X"27",X"53",X"20",X"41",X"20",X"48",X"45",X"41",X"4C",X"54",X"48",
		X"59",X"20",X"53",X"43",X"4F",X"52",X"45",X"21",X"00",X"0F",X"43",X"55",X"50",X"2F",X"44",X"4F",
		X"57",X"4E",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",X"53",X"20",X"4C",X"45",X"54",X"54",X"45",
		X"52",X"2E",X"2E",X"00",X"11",X"42",X"E4",X"E0",X"E0",X"E0",X"E0",X"E0",X"E5",X"00",X"F2",X"42",
		X"59",X"4F",X"55",X"52",X"20",X"3E",X"20",X"E1",X"20",X"44",X"57",X"46",X"20",X"E3",X"20",X"3C",
		X"20",X"43",X"4F",X"44",X"45",X"00",X"13",X"42",X"E6",X"E2",X"E2",X"E2",X"E2",X"E2",X"E7",X"00",
		X"15",X"43",X"4C",X"45",X"46",X"54",X"2F",X"52",X"49",X"47",X"48",X"54",X"20",X"4D",X"4F",X"56",
		X"45",X"53",X"20",X"41",X"52",X"52",X"4F",X"57",X"2E",X"2E",X"00",X"DA",X"42",X"22",X"5A",X"41",
		X"50",X"22",X"20",X"57",X"48",X"45",X"4E",X"20",X"41",X"4C",X"4C",X"20",X"53",X"45",X"54",X"2E",
		X"00",X"DB",X"42",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"00",X"00",X"01",X"30",X"32",X"16",X"69",X"21",X"00",X"68",
		X"7D",X"23",X"77",X"FE",X"07",X"C2",X"25",X"32",X"EB",X"3E",X"C0",X"A6",X"77",X"0A",X"03",X"B6",
		X"77",X"EB",X"C3",X"28",X"32",X"0A",X"12",X"03",X"3E",X"0D",X"BD",X"C2",X"10",X"32",X"75",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"00",X"00",X"00",X"0E",X"0E",X"00",X"CD",X"98",
		X"34",X"CD",X"64",X"32",X"CD",X"D2",X"33",X"CD",X"85",X"33",X"CD",X"FB",X"32",X"3A",X"92",X"43",
		X"FE",X"09",X"DC",X"18",X"33",X"CD",X"F9",X"33",X"3A",X"8B",X"43",X"B7",X"F8",X"CD",X"AF",X"33",
		X"CD",X"35",X"33",X"C9",X"21",X"93",X"43",X"7E",X"B7",X"C8",X"34",X"FE",X"D0",X"D8",X"FE",X"FF",
		X"CA",X"BE",X"33",X"FE",X"E0",X"C2",X"90",X"32",X"21",X"94",X"43",X"34",X"35",X"CA",X"90",X"32",
		X"35",X"C2",X"8B",X"32",X"AF",X"32",X"93",X"43",X"C3",X"BE",X"33",X"3E",X"D0",X"32",X"93",X"43",
		X"D6",X"10",X"07",X"E6",X"7E",X"21",X"9B",X"32",X"C3",X"6D",X"34",X"42",X"00",X"3E",X"00",X"3A",
		X"00",X"37",X"00",X"34",X"00",X"31",X"00",X"2E",X"00",X"2C",X"00",X"29",X"00",X"27",X"00",X"25",
		X"00",X"23",X"00",X"21",X"00",X"23",X"00",X"25",X"00",X"27",X"00",X"29",X"00",X"2C",X"00",X"2E",
		X"00",X"31",X"00",X"34",X"00",X"37",X"00",X"3A",X"00",X"3E",X"00",X"42",X"00",X"46",X"00",X"4A",
		X"00",X"4E",X"00",X"53",X"00",X"58",X"00",X"5D",X"00",X"62",X"00",X"68",X"00",X"6E",X"00",X"75",
		X"00",X"7C",X"00",X"83",X"00",X"8B",X"00",X"93",X"00",X"9C",X"00",X"A5",X"00",X"AF",X"00",X"BA",
		X"00",X"C5",X"00",X"D0",X"00",X"DD",X"00",X"EA",X"00",X"00",X"00",X"21",X"90",X"43",X"7E",X"B7",
		X"C8",X"23",X"35",X"35",X"7E",X"FE",X"20",X"D2",X"0F",X"33",X"2B",X"35",X"C3",X"BE",X"33",X"3E",
		X"D0",X"96",X"4F",X"06",X"00",X"C3",X"73",X"34",X"21",X"87",X"43",X"7E",X"B7",X"C8",X"35",X"CA",
		X"BE",X"33",X"D6",X"02",X"07",X"E6",X"06",X"21",X"2D",X"33",X"C3",X"6D",X"34",X"7C",X"00",X"62",
		X"00",X"53",X"00",X"3E",X"00",X"21",X"8F",X"43",X"34",X"7E",X"FE",X"0C",X"D8",X"36",X"00",X"3A",
		X"F5",X"43",X"E6",X"07",X"FE",X"04",X"C0",X"3A",X"71",X"43",X"E6",X"0F",X"FE",X"08",X"D0",X"07",
		X"C6",X"20",X"4F",X"06",X"00",X"E1",X"11",X"00",X"69",X"21",X"04",X"68",X"75",X"79",X"12",X"23",
		X"75",X"78",X"12",X"23",X"23",X"75",X"1A",X"F6",X"3F",X"E6",X"FB",X"12",X"23",X"75",X"AF",X"12",
		X"23",X"75",X"12",X"23",X"75",X"3E",X"10",X"12",X"23",X"75",X"3E",X"0E",X"12",X"23",X"75",X"12",
		X"23",X"75",X"AF",X"12",X"C9",X"21",X"89",X"43",X"7E",X"B7",X"C8",X"23",X"7E",X"35",X"FE",X"0A",
		X"D2",X"AD",X"33",X"B7",X"C0",X"36",X"0C",X"2B",X"35",X"7E",X"E6",X"03",X"FE",X"02",X"D8",X"01",
		X"BA",X"00",X"E6",X"01",X"CA",X"55",X"33",X"01",X"8B",X"00",X"C3",X"55",X"33",X"E1",X"C9",X"21",
		X"84",X"43",X"7E",X"B7",X"C8",X"35",X"3D",X"C0",X"01",X"6E",X"00",X"C3",X"55",X"33",X"3E",X"02",
		X"21",X"07",X"68",X"75",X"24",X"B6",X"77",X"C9",X"3E",X"01",X"C3",X"C0",X"33",X"3E",X"04",X"C3",
		X"C0",X"33",X"21",X"88",X"43",X"7E",X"B7",X"C8",X"35",X"C2",X"E2",X"33",X"CD",X"BE",X"33",X"C3",
		X"00",X"21",X"E1",X"0F",X"0F",X"E6",X"02",X"21",X"ED",X"33",X"C3",X"6D",X"34",X"9C",X"00",X"5D",
		X"00",X"3E",X"00",X"6E",X"00",X"C5",X"00",X"5E",X"01",X"21",X"92",X"43",X"7E",X"B7",X"C8",X"2B",
		X"FE",X"0A",X"DA",X"10",X"34",X"CD",X"61",X"34",X"E6",X"06",X"21",X"F1",X"33",X"C3",X"6D",X"34",
		X"00",X"FE",X"06",X"DA",X"2B",X"34",X"CD",X"61",X"34",X"E6",X"1F",X"01",X"6E",X"00",X"B7",X"CA",
		X"73",X"34",X"FE",X"04",X"C0",X"01",X"3E",X"00",X"C3",X"73",X"34",X"FE",X"02",X"DA",X"45",X"34",
		X"CD",X"61",X"34",X"E6",X"0F",X"01",X"6E",X"00",X"B7",X"CA",X"73",X"34",X"FE",X"04",X"C0",X"01",
		X"3E",X"00",X"C3",X"73",X"34",X"7E",X"FE",X"40",X"DA",X"4D",X"34",X"36",X"40",X"35",X"7E",X"E6",
		X"07",X"01",X"6E",X"00",X"B7",X"CA",X"73",X"34",X"FE",X"04",X"C0",X"01",X"3E",X"00",X"C3",X"73",
		X"34",X"35",X"7E",X"FE",X"40",X"D8",X"36",X"3F",X"23",X"35",X"2B",X"7E",X"C9",X"CD",X"9D",X"02",
		X"4E",X"23",X"46",X"E1",X"21",X"07",X"69",X"11",X"09",X"68",X"7D",X"12",X"7E",X"F6",X"3F",X"E6",
		X"FD",X"77",X"00",X"7B",X"12",X"36",X"0F",X"3D",X"12",X"36",X"00",X"3C",X"3C",X"12",X"36",X"00",
		X"3E",X"02",X"12",X"71",X"3C",X"12",X"70",X"C9",X"3A",X"F5",X"43",X"E6",X"07",X"FE",X"07",X"C2",
		X"AD",X"34",X"3A",X"4F",X"43",X"FE",X"04",X"D8",X"3A",X"88",X"43",X"B7",X"C0",X"21",X"8B",X"43",
		X"7E",X"B7",X"C8",X"FA",X"C2",X"34",X"F6",X"80",X"77",X"21",X"FF",X"00",X"22",X"8C",X"43",X"22",
		X"8D",X"43",X"E1",X"3A",X"8B",X"43",X"E6",X"0F",X"3D",X"07",X"21",X"68",X"36",X"CD",X"9D",X"02",
		X"5E",X"23",X"56",X"1A",X"13",X"4F",X"21",X"8C",X"43",X"34",X"7E",X"D6",X"03",X"C0",X"77",X"23",
		X"34",X"7E",X"FE",X"04",X"DA",X"EE",X"34",X"D6",X"10",X"D8",X"77",X"23",X"34",X"2B",X"E5",X"23",
		X"6E",X"26",X"00",X"19",X"46",X"78",X"E1",X"FE",X"FF",X"C2",X"01",X"35",X"AF",X"32",X"8B",X"43",
		X"C9",X"FE",X"80",X"C2",X"0D",X"35",X"7E",X"FE",X"01",X"C0",X"36",X"0E",X"C9",X"07",X"07",X"07",
		X"E6",X"06",X"EB",X"21",X"23",X"35",X"CD",X"9D",X"02",X"7E",X"EB",X"BE",X"D2",X"2B",X"35",X"13",
		X"1A",X"77",X"C9",X"00",X"0F",X"01",X"0E",X"01",X"0A",X"01",X"06",X"78",X"E6",X"3F",X"81",X"B7",
		X"17",X"5F",X"3E",X"00",X"17",X"57",X"21",X"9E",X"35",X"19",X"C5",X"E5",X"01",X"00",X"68",X"11",
		X"00",X"69",X"3E",X"06",X"CD",X"9D",X"02",X"CD",X"8C",X"35",X"3E",X"0A",X"CD",X"9D",X"02",X"CD",
		X"8C",X"35",X"E1",X"7E",X"23",X"66",X"6F",X"D5",X"E5",X"D1",X"29",X"19",X"11",X"B8",X"0B",X"19",
		X"D1",X"EB",X"E3",X"EB",X"53",X"19",X"D1",X"3E",X"0B",X"02",X"7D",X"12",X"3E",X"0C",X"02",X"7C",
		X"12",X"21",X"0A",X"68",X"AF",X"75",X"2B",X"12",X"3E",X"10",X"75",X"2B",X"12",X"75",X"2B",X"12",
		X"75",X"1A",X"F6",X"3F",X"E6",X"FC",X"12",X"36",X"0D",X"AF",X"12",X"C9",X"79",X"03",X"02",X"7E",
		X"23",X"12",X"79",X"03",X"02",X"7E",X"23",X"12",X"C9",X"D5",X"E5",X"0E",X"4C",X"21",X"E6",X"06",
		X"83",X"06",X"26",X"06",X"CD",X"05",X"7A",X"05",X"2B",X"05",X"E1",X"04",X"9B",X"04",X"59",X"04",
		X"1A",X"04",X"DF",X"03",X"A8",X"03",X"73",X"03",X"42",X"03",X"13",X"03",X"E7",X"02",X"BD",X"02",
		X"96",X"02",X"71",X"02",X"4D",X"02",X"2D",X"02",X"0D",X"02",X"F0",X"01",X"D4",X"01",X"B9",X"01",
		X"A1",X"01",X"89",X"01",X"73",X"01",X"5E",X"01",X"4B",X"01",X"38",X"01",X"27",X"01",X"16",X"01",
		X"08",X"01",X"F8",X"00",X"EA",X"00",X"DD",X"00",X"D0",X"00",X"C5",X"00",X"BA",X"00",X"AF",X"00",
		X"A5",X"00",X"9C",X"00",X"93",X"00",X"8B",X"00",X"83",X"00",X"7C",X"00",X"75",X"00",X"6E",X"00",
		X"68",X"00",X"62",X"00",X"5D",X"00",X"58",X"00",X"53",X"00",X"4E",X"00",X"4A",X"00",X"46",X"00",
		X"42",X"00",X"3E",X"00",X"3A",X"00",X"37",X"00",X"34",X"00",X"31",X"00",X"2E",X"00",X"2C",X"00",
		X"29",X"00",X"27",X"00",X"25",X"00",X"23",X"00",X"21",X"00",X"1F",X"00",X"1D",X"00",X"1C",X"00",
		X"1A",X"00",X"19",X"00",X"17",X"00",X"16",X"00",X"15",X"00",X"13",X"00",X"12",X"00",X"11",X"00",
		X"10",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",
		X"0A",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"07",X"00",
		X"3A",X"8B",X"43",X"B7",X"C2",X"68",X"36",X"11",X"88",X"36",X"A7",X"36",X"C5",X"36",X"E0",X"36",
		X"00",X"37",X"40",X"37",X"24",X"37",X"77",X"37",X"A7",X"36",X"C5",X"36",X"E0",X"36",X"00",X"37",
		X"40",X"37",X"24",X"37",X"9C",X"37",X"9C",X"37",X"24",X"80",X"80",X"80",X"80",X"64",X"60",X"61",
		X"5C",X"5E",X"5B",X"5D",X"58",X"80",X"96",X"95",X"94",X"93",X"92",X"91",X"90",X"52",X"55",X"53",
		X"99",X"55",X"50",X"92",X"54",X"D8",X"FF",X"18",X"80",X"80",X"80",X"80",X"D9",X"80",X"99",X"60",
		X"A0",X"80",X"60",X"9B",X"80",X"5C",X"9B",X"D9",X"80",X"80",X"80",X"A0",X"A3",X"E5",X"80",X"A3",
		X"A0",X"A2",X"9E",X"E0",X"FF",X"18",X"80",X"80",X"80",X"80",X"9C",X"9E",X"5C",X"99",X"99",X"59",
		X"99",X"57",X"99",X"5A",X"D9",X"80",X"9A",X"97",X"5C",X"D9",X"80",X"95",X"92",X"57",X"D0",X"FF",
		X"18",X"80",X"80",X"80",X"80",X"55",X"99",X"9C",X"59",X"9C",X"9E",X"DC",X"99",X"9C",X"DE",X"80",
		X"9C",X"80",X"99",X"9C",X"DC",X"59",X"9A",X"99",X"D7",X"95",X"97",X"D9",X"97",X"D5",X"80",X"FF",
		X"18",X"80",X"80",X"80",X"5C",X"1C",X"9C",X"97",X"60",X"20",X"A0",X"9C",X"5C",X"60",X"E3",X"23",
		X"61",X"60",X"DE",X"80",X"5E",X"60",X"A1",X"A1",X"60",X"1E",X"A0",X"9C",X"5C",X"60",X"9E",X"97",
		X"5B",X"1E",X"DC",X"FF",X"17",X"80",X"80",X"80",X"80",X"99",X"DC",X"9E",X"A0",X"80",X"62",X"A0",
		X"DE",X"80",X"9B",X"D7",X"59",X"9B",X"DC",X"99",X"99",X"80",X"57",X"99",X"DB",X"97",X"D4",X"FF",
		X"18",X"80",X"80",X"80",X"9C",X"5C",X"1C",X"5C",X"1A",X"59",X"1C",X"61",X"23",X"65",X"25",X"65",
		X"23",X"A1",X"61",X"20",X"5E",X"1E",X"5E",X"20",X"61",X"20",X"61",X"1E",X"5C",X"1E",X"5C",X"19",
		X"9C",X"9C",X"5C",X"1C",X"5C",X"1A",X"59",X"1C",X"61",X"23",X"65",X"25",X"65",X"23",X"E1",X"80",
		X"61",X"A3",X"A3",X"A1",X"A0",X"E1",X"FF",X"18",X"80",X"80",X"80",X"DC",X"5A",X"59",X"1C",X"61",
		X"23",X"E5",X"A1",X"80",X"DE",X"60",X"61",X"20",X"61",X"1E",X"DC",X"D9",X"80",X"DC",X"5A",X"59",
		X"1C",X"61",X"23",X"E5",X"A1",X"A1",X"A3",X"A3",X"A1",X"A0",X"E1",X"FF",X"18",X"80",X"80",X"80",
		X"80",X"AB",X"A5",X"A7",X"A2",X"E0",X"80",X"80",X"80",X"80",X"AB",X"A5",X"A7",X"A2",X"E0",X"80",
		X"80",X"80",X"80",X"80",X"80",X"6A",X"68",X"67",X"69",X"66",X"65",X"67",X"68",X"66",X"64",X"5F",
		X"62",X"60",X"5D",X"DC",X"80",X"80",X"80",X"80",X"AB",X"A5",X"A7",X"A2",X"E0",X"80",X"80",X"80",
		X"80",X"FF",X"3A",X"8B",X"43",X"00",X"B7",X"C2",X"E0",X"37",X"34",X"E5",X"CD",X"EE",X"02",X"E1",
		X"23",X"34",X"2B",X"C2",X"E7",X"37",X"34",X"4E",X"79",X"FE",X"0E",X"DA",X"1B",X"38",X"23",X"AF",
		X"77",X"2B",X"77",X"2B",X"34",X"E5",X"11",X"A9",X"31",X"21",X"13",X"38",X"0E",X"06",X"1A",X"2F",
		X"AE",X"C2",X"0C",X"38",X"13",X"23",X"0D",X"C2",X"FE",X"37",X"E1",X"C9",X"E1",X"35",X"35",X"C9",
		X"B7",X"C0",X"01",X"BB",X"A8",X"B9",X"DF",X"1C",X"DF",X"00",X"C9",X"FE",X"0C",X"D2",X"AA",X"38",
		X"23",X"FE",X"01",X"C2",X"6C",X"38",X"3E",X"FE",X"32",X"9D",X"43",X"32",X"00",X"58",X"21",X"BB",
		X"38",X"0E",X"03",X"CD",X"5D",X"02",X"11",X"21",X"43",X"01",X"18",X"08",X"CD",X"83",X"20",X"11",
		X"A5",X"42",X"01",X"58",X"50",X"CD",X"9A",X"19",X"11",X"45",X"41",X"0E",X"70",X"CD",X"FA",X"13",
		X"3E",X"D1",X"32",X"85",X"48",X"3E",X"D0",X"32",X"66",X"48",X"32",X"A4",X"48",X"3E",X"20",X"32",
		X"E5",X"49",X"32",X"65",X"49",X"32",X"65",X"4A",X"32",X"C5",X"48",X"C9",X"7E",X"FE",X"30",X"D8",
		X"36",X"FF",X"2B",X"7E",X"3D",X"4F",X"FE",X"08",X"DA",X"A4",X"38",X"0C",X"FE",X"08",X"C2",X"93",
		X"38",X"3E",X"38",X"32",X"98",X"4A",X"3E",X"3A",X"32",X"38",X"4A",X"3E",X"4C",X"32",X"58",X"40",
		X"C3",X"A4",X"38",X"FE",X"0A",X"D2",X"A4",X"38",X"0C",X"C5",X"11",X"DB",X"42",X"01",X"05",X"4C",
		X"CD",X"26",X"3D",X"C1",X"21",X"09",X"39",X"C3",X"5D",X"02",X"FE",X"0D",X"D0",X"23",X"7E",X"FE",
		X"50",X"C0",X"21",X"EC",X"39",X"0E",X"03",X"C3",X"5D",X"02",X"21",X"00",X"43",X"3D",X"3D",X"3D",
		X"3D",X"3D",X"20",X"48",X"4F",X"57",X"20",X"54",X"4F",X"20",X"50",X"4C",X"41",X"59",X"20",X"20",
		X"3D",X"3D",X"3D",X"3D",X"3D",X"00",X"02",X"43",X"2A",X"20",X"5A",X"41",X"50",X"20",X"56",X"45",
		X"49",X"4E",X"53",X"20",X"41",X"4E",X"44",X"20",X"47",X"45",X"52",X"4D",X"53",X"20",X"20",X"2A",
		X"00",X"C8",X"42",X"43",X"45",X"4C",X"4C",X"20",X"20",X"20",X"20",X"20",X"20",X"47",X"45",X"52",
		X"4D",X"53",X"20",X"56",X"45",X"49",X"4E",X"53",X"00",X"2A",X"42",X"20",X"53",X"43",X"4F",X"52",
		X"49",X"4E",X"47",X"20",X"00",X"0C",X"43",X"2A",X"20",X"41",X"4E",X"59",X"20",X"47",X"45",X"52",
		X"4D",X"20",X"20",X"35",X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"CD",X"42",
		X"41",X"4C",X"4C",X"20",X"31",X"43",X"4F",X"4C",X"4F",X"52",X"2D",X"2D",X"2D",X"20",X"4E",X"4F",
		X"20",X"4B",X"49",X"4C",X"4C",X"21",X"00",X"0F",X"43",X"2A",X"20",X"41",X"4E",X"59",X"20",X"56",
		X"45",X"49",X"4E",X"20",X"20",X"31",X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",
		X"11",X"43",X"2A",X"20",X"5A",X"41",X"50",X"53",X"20",X"4C",X"45",X"46",X"54",X"20",X"20",X"33",
		X"30",X"2F",X"5A",X"41",X"50",X"00",X"13",X"43",X"00",X"35",X"43",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"24",X"24",X"24",X"20",X"53",X"50",X"45",X"43",X"49",X"41",X"4C",X"53",X"20",X"24",X"24",X"24",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"00",X"17",X"43",X"2A",X"20",X"47",X"4F",X"20",X"54",X"4F",X"20",
		X"46",X"4C",X"41",X"53",X"48",X"49",X"4E",X"47",X"20",X"43",X"4F",X"52",X"4E",X"45",X"52",X"53",
		X"00",X"F8",X"41",X"47",X"45",X"54",X"20",X"5A",X"41",X"50",X"53",X"2B",X"54",X"49",X"4E",X"59",
		X"00",X"1A",X"43",X"2A",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"43",X"45",X"4C",X"4C",X"53",
		X"20",X"41",X"54",X"20",X"53",X"43",X"4F",X"52",X"45",X"53",X"00",X"3B",X"42",X"20",X"3D",X"20",
		X"31",X"46",X"52",X"45",X"45",X"20",X"43",X"45",X"4C",X"4C",X"00",X"00",X"9D",X"42",X"53",X"55",
		X"52",X"56",X"49",X"56",X"41",X"4C",X"20",X"20",X"5C",X"20",X"31",X"39",X"38",X"32",X"00",X"BE",
		X"42",X"52",X"4F",X"43",X"4B",X"2D",X"4F",X"4C",X"41",X"20",X"4D",X"46",X"47",X"2E",X"20",X"43",
		X"4F",X"52",X"50",X"2E",X"00",X"3F",X"43",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"00",X"3A",X"8B",X"43",X"B7",X"C2",X"3D",X"3A",X"34",X"C3",X"EE",X"02",X"23",X"34",X"2B",
		X"C2",X"44",X"3A",X"34",X"4E",X"79",X"FE",X"10",X"DA",X"53",X"3A",X"AF",X"23",X"77",X"2B",X"77",
		X"2B",X"34",X"C9",X"FE",X"05",X"D2",X"65",X"3A",X"23",X"7E",X"FE",X"10",X"D8",X"36",X"FF",X"21",
		X"B9",X"3A",X"C3",X"5D",X"02",X"FE",X"06",X"D2",X"79",X"3A",X"23",X"7E",X"FE",X"15",X"D8",X"36",
		X"FF",X"21",X"EC",X"39",X"0E",X"03",X"C3",X"5D",X"02",X"FE",X"0F",X"D0",X"23",X"7E",X"FE",X"30",
		X"D8",X"36",X"FF",X"11",X"84",X"42",X"79",X"D6",X"05",X"4F",X"13",X"13",X"3D",X"C2",X"8A",X"3A",
		X"3E",X"2A",X"12",X"CD",X"83",X"3C",X"3E",X"30",X"B1",X"12",X"CD",X"83",X"3C",X"CD",X"83",X"3C",
		X"79",X"07",X"4F",X"07",X"81",X"21",X"AF",X"43",X"85",X"6F",X"0E",X"03",X"CD",X"30",X"3D",X"23",
		X"23",X"15",X"CD",X"83",X"3C",X"C3",X"B4",X"3C",X"21",X"00",X"43",X"2A",X"20",X"54",X"4F",X"44",
		X"41",X"59",X"27",X"53",X"20",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"53",
		X"20",X"20",X"2A",X"00",X"21",X"43",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"00",X"83",X"42",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"20",X"20",X"20",X"53",X"43",X"4F",
		X"52",X"45",X"00",X"84",X"42",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"20",X"20",X"20",X"20",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"00",X"00",X"3A",X"8B",X"43",X"B7",X"C2",X"22",X"3B",X"34",X"C3",
		X"EE",X"02",X"23",X"34",X"2B",X"C2",X"29",X"3B",X"34",X"4E",X"79",X"FE",X"32",X"DA",X"3B",X"3B",
		X"AF",X"23",X"77",X"2B",X"77",X"2B",X"34",X"20",X"C3",X"EE",X"02",X"E6",X"01",X"CA",X"7B",X"3B",
		X"79",X"FE",X"01",X"23",X"CA",X"4B",X"3B",X"7E",X"FE",X"03",X"D8",X"36",X"FF",X"21",X"85",X"3B",
		X"0E",X"04",X"CD",X"5D",X"02",X"CD",X"94",X"17",X"78",X"E6",X"0F",X"F6",X"30",X"32",X"ED",X"42",
		X"78",X"E6",X"F0",X"CA",X"6B",X"3B",X"3E",X"31",X"32",X"0D",X"43",X"79",X"F6",X"30",X"32",X"EA",
		X"42",X"FE",X"31",X"C8",X"20",X"3E",X"13",X"32",X"2A",X"42",X"C9",X"23",X"7E",X"FE",X"05",X"D8",
		X"36",X"FF",X"C3",X"83",X"21",X"21",X"43",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",
		X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",
		X"3D",X"00",X"AA",X"42",X"43",X"4F",X"49",X"4E",X"20",X"20",X"46",X"4F",X"52",X"20",X"31",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"AD",X"42",X"43",X"4F",X"49",X"4E",X"53",X"20",X"46",
		X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"3F",X"43",X"3D",
		X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",
		X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"00",X"7E",X"81",X"27",X"77",X"2B",X"7E",
		X"88",X"27",X"77",X"2B",X"7E",X"CE",X"00",X"27",X"77",X"23",X"23",X"C9",X"37",X"3E",X"99",X"CE",
		X"00",X"91",X"86",X"27",X"77",X"2B",X"3E",X"99",X"CE",X"00",X"90",X"86",X"27",X"77",X"2B",X"3E",
		X"99",X"CE",X"00",X"86",X"27",X"77",X"23",X"23",X"C9",X"C5",X"01",X"01",X"00",X"CD",X"FC",X"3B",
		X"C1",X"7E",X"C9",X"D5",X"C5",X"7E",X"12",X"23",X"13",X"05",X"C2",X"25",X"3C",X"C1",X"D1",X"0D",
		X"C8",X"7B",X"F5",X"CD",X"83",X"3C",X"F1",X"BB",X"C8",X"C3",X"23",X"3C",X"7E",X"12",X"23",X"13",
		X"0D",X"C2",X"3C",X"3C",X"C9",X"E5",X"D5",X"C5",X"CD",X"6F",X"3C",X"5F",X"16",X"00",X"21",X"00",
		X"00",X"0E",X"08",X"0D",X"CA",X"60",X"3C",X"29",X"17",X"D2",X"53",X"3C",X"19",X"C3",X"53",X"3C",
		X"7C",X"1F",X"7D",X"1F",X"FE",X"80",X"DA",X"6B",X"3C",X"3E",X"7F",X"C1",X"D1",X"E1",X"C9",X"B7",
		X"F0",X"2F",X"3C",X"C9",X"06",X"00",X"70",X"23",X"0D",X"C2",X"76",X"3C",X"C9",X"34",X"C0",X"2B",
		X"34",X"23",X"C9",X"7B",X"D6",X"20",X"5F",X"7A",X"DE",X"00",X"57",X"E6",X"07",X"FE",X"07",X"C0",
		X"20",X"7B",X"C6",X"20",X"5F",X"7A",X"CE",X"00",X"57",X"E6",X"03",X"FE",X"03",X"C0",X"7B",X"FE",
		X"40",X"D2",X"83",X"3C",X"C9",X"06",X"02",X"C3",X"B6",X"3C",X"06",X"03",X"C3",X"B6",X"3C",X"06",
		X"04",X"C3",X"B6",X"3C",X"06",X"06",X"7E",X"E6",X"0F",X"F6",X"30",X"12",X"CD",X"91",X"3C",X"05",
		X"C8",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"F6",X"30",X"12",X"CD",X"91",X"3C",X"2B",X"05",
		X"C2",X"B6",X"3C",X"C9",X"AF",X"77",X"23",X"05",X"C2",X"D5",X"3C",X"C9",X"1A",X"96",X"1B",X"2B",
		X"1A",X"9E",X"1B",X"2B",X"1A",X"9E",X"13",X"23",X"13",X"23",X"D8",X"C0",X"1A",X"AE",X"C0",X"1B",
		X"2B",X"1A",X"AE",X"13",X"23",X"C0",X"37",X"C9",X"11",X"3F",X"43",X"21",X"3E",X"43",X"01",X"1F",
		X"19",X"C5",X"D5",X"E5",X"7E",X"12",X"1B",X"2B",X"0D",X"C2",X"04",X"3D",X"E1",X"D1",X"CD",X"83",
		X"3C",X"EB",X"CD",X"83",X"3C",X"EB",X"C1",X"05",X"C2",X"01",X"3D",X"11",X"20",X"43",X"7C",X"E6",
		X"08",X"B2",X"57",X"01",X"19",X"00",X"78",X"12",X"CD",X"83",X"3C",X"0D",X"C2",X"26",X"3D",X"C9",
		X"7E",X"12",X"23",X"CD",X"83",X"3C",X"0D",X"C2",X"30",X"3D",X"C9",X"C5",X"D5",X"7C",X"12",X"13",
		X"05",X"C2",X"3D",X"3D",X"D1",X"CD",X"83",X"3C",X"C1",X"0D",X"C2",X"3B",X"3D",X"C9",X"21",X"00",
		X"44",X"22",X"00",X"00",X"2A",X"06",X"00",X"C1",X"E5",X"11",X"5C",X"00",X"0E",X"13",X"C9",X"41",
		X"4C",X"4C",X"20",X"47",X"41",X"4D",X"45",X"20",X"46",X"45",X"41",X"54",X"55",X"52",X"45",X"53",
		X"20",X"49",X"4E",X"43",X"4C",X"55",X"44",X"49",X"4E",X"47",X"20",X"4E",X"41",X"4D",X"45",X"2C",
		X"20",X"47",X"41",X"4D",X"45",X"20",X"49",X"44",X"45",X"41",X"2C",X"20",X"44",X"45",X"53",X"49",
		X"47",X"4E",X"2C",X"20",X"53",X"48",X"41",X"50",X"45",X"53",X"2C",X"20",X"43",X"4F",X"4C",X"4F",
		X"52",X"53",X"2C",X"20",X"53",X"4F",X"55",X"4E",X"44",X"53",X"2C",X"20",X"4D",X"55",X"53",X"49",
		X"43",X"20",X"41",X"4E",X"44",X"20",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"20",X"43",X"4F",
		X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"42",X"59",X"20",
		X"4D",X"49",X"43",X"52",X"4F",X"54",X"52",X"41",X"49",X"4E",X"20",X"4C",X"54",X"44",X"2E",X"20",
		X"41",X"4E",X"44",X"20",X"41",X"53",X"53",X"49",X"47",X"4E",X"45",X"44",X"20",X"54",X"4F",X"20",
		X"52",X"4F",X"43",X"4B",X"2D",X"4F",X"4C",X"41",X"20",X"4D",X"46",X"47",X"2E",X"20",X"43",X"4F",
		X"52",X"50",X"2E",X"20",X"50",X"4C",X"41",X"47",X"49",X"41",X"52",X"49",X"53",X"54",X"53",X"20",
		X"57",X"49",X"4C",X"4C",X"20",X"42",X"45",X"20",X"50",X"52",X"4F",X"53",X"45",X"43",X"55",X"54",
		X"45",X"44",X"2E",X"00",X"2B",X"3E",X"00",X"00",X"DF",X"00",X"DF",X"0F",X"E6",X"04",X"3E",X"5C",
		X"CD",X"FF",X"40",X"C9",X"7E",X"B7",X"C8",X"CD",X"25",X"42",X"FE",X"20",X"D2",X"56",X"3E",X"FE",
		X"0A",X"CA",X"56",X"3E",X"FE",X"07",X"CA",X"56",X"3E",X"FE",X"09",X"CA",X"56",X"3E",X"3E",X"07",
		X"CD",X"FF",X"40",X"C3",X"37",X"3E",X"77",X"CD",X"D9",X"42",X"23",X"04",X"15",X"C2",X"34",X"3E",
		X"C9",X"36",X"00",X"48",X"16",X"FF",X"CD",X"D3",X"3D",X"CD",X"25",X"42",X"FE",X"7F",X"CA",X"9C",
		X"3E",X"FE",X"08",X"CA",X"9E",X"3E",X"FE",X"0D",X"CA",X"02",X"3F",X"FE",X"1B",X"C8",X"FE",X"08",
		X"CA",X"9E",X"3E",X"FE",X"0A",X"CA",X"BC",X"3E",X"FE",X"07",X"CA",X"BC",X"3E",X"FE",X"09",X"CA",
		X"BC",X"3E",X"FE",X"20",X"DA",X"69",X"3E",X"FE",X"5F",X"C2",X"BC",X"3E",X"3E",X"5F",X"05",X"04",
		X"CA",X"C4",X"3E",X"CD",X"D9",X"42",X"2B",X"05",X"11",X"69",X"3E",X"D5",X"E5",X"0D",X"7E",X"B7",
		X"37",X"CA",X"5C",X"27",X"23",X"7E",X"2B",X"77",X"23",X"C3",X"AE",X"3E",X"F5",X"79",X"FE",X"FF",
		X"DA",X"CC",X"3E",X"F1",X"3E",X"07",X"CD",X"FF",X"40",X"C3",X"69",X"3E",X"90",X"0C",X"04",X"C5",
		X"EB",X"6F",X"26",X"00",X"19",X"44",X"4D",X"23",X"CD",X"ED",X"42",X"C1",X"F1",X"77",X"CD",X"D9",
		X"42",X"23",X"C3",X"C9",X"3E",X"78",X"B7",X"C8",X"2B",X"3E",X"08",X"CD",X"D9",X"42",X"05",X"15",
		X"C2",X"F4",X"3E",X"C9",X"78",X"B7",X"C8",X"05",X"2B",X"7E",X"CD",X"D9",X"42",X"15",X"C2",X"F4",
		X"3E",X"C9",X"CD",X"F6",X"20",X"CD",X"51",X"42",X"C1",X"D1",X"7A",X"A3",X"3C",X"21",X"84",X"09",
		X"C8",X"37",X"F5",X"23",X"C3",X"37",X"0E",X"C1",X"D1",X"7A",X"A3",X"3C",X"CA",X"4C",X"42",X"C3",
		X"AA",X"0D",X"CD",X"1E",X"1A",X"CD",X"3A",X"2A",X"CD",X"07",X"44",X"3B",X"EB",X"2A",X"27",X"0C",
		X"C3",X"3C",X"3F",X"3A",X"C9",X"0A",X"B7",X"CA",X"46",X"3F",X"D1",X"EB",X"E5",X"AF",X"32",X"C9",
		X"0A",X"BA",X"F5",X"D5",X"46",X"B0",X"CA",X"4A",X"14",X"23",X"4E",X"23",X"66",X"69",X"C3",X"70",
		X"3F",X"58",X"E5",X"0E",X"02",X"7E",X"23",X"FE",X"5C",X"CA",X"BC",X"40",X"FE",X"20",X"C2",X"66",
		X"3F",X"0C",X"05",X"C2",X"55",X"3F",X"E1",X"43",X"3E",X"5C",X"CD",X"F5",X"40",X"CD",X"FF",X"40",
		X"AF",X"5F",X"57",X"CD",X"F5",X"40",X"57",X"7E",X"23",X"FE",X"21",X"CA",X"B9",X"40",X"FE",X"23",
		X"CA",X"CC",X"3F",X"FE",X"26",X"CA",X"B4",X"40",X"05",X"CA",X"92",X"40",X"FE",X"2B",X"3E",X"08",
		X"CA",X"73",X"3F",X"2B",X"7E",X"23",X"FE",X"2E",X"CA",X"EB",X"3F",X"FE",X"5F",X"CA",X"A8",X"40",
		X"FE",X"5C",X"CA",X"51",X"3F",X"BE",X"C2",X"6A",X"3F",X"FE",X"24",X"CA",X"C5",X"3F",X"FE",X"2A",
		X"C2",X"6A",X"3F",X"78",X"23",X"FE",X"02",X"DA",X"BD",X"3F",X"7E",X"FE",X"24",X"3E",X"20",X"C2",
		X"C9",X"3F",X"05",X"1C",X"FE",X"AF",X"C6",X"10",X"23",X"1C",X"82",X"57",X"1C",X"0E",X"00",X"05",
		X"CA",X"21",X"40",X"7E",X"23",X"FE",X"2E",X"CA",X"F6",X"3F",X"FE",X"23",X"CA",X"CC",X"3F",X"FE",
		X"2C",X"C2",X"02",X"40",X"7A",X"F6",X"40",X"57",X"C3",X"CC",X"3F",X"7E",X"FE",X"23",X"3E",X"2E",
		X"C2",X"6A",X"3F",X"0E",X"01",X"23",X"0C",X"05",X"CA",X"21",X"40",X"7E",X"23",X"FE",X"23",X"C9");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
