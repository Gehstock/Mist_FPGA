-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity INVADERS_ROM_F is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of INVADERS_ROM_F is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"CD",x"74",x"14",x"00",x"C5",x"E5",x"1A", -- 0x0400
    x"D3",x"04",x"DB",x"03",x"B6",x"77",x"23",x"13", -- 0x0408
    x"AF",x"D3",x"04",x"DB",x"03",x"B6",x"77",x"E1", -- 0x0410
    x"01",x"20",x"00",x"09",x"C1",x"05",x"C2",x"05", -- 0x0418
    x"14",x"C9",x"00",x"00",x"CD",x"74",x"14",x"C5", -- 0x0420
    x"E5",x"AF",x"77",x"23",x"77",x"23",x"E1",x"01", -- 0x0428
    x"20",x"00",x"09",x"C1",x"05",x"C2",x"27",x"14", -- 0x0430
    x"C9",x"C5",x"1A",x"77",x"13",x"01",x"20",x"00", -- 0x0438
    x"09",x"C1",x"05",x"C2",x"39",x"14",x"C9",x"00", -- 0x0440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"CD",x"74",x"14",x"C5",x"E5",x"1A", -- 0x0450
    x"D3",x"04",x"DB",x"03",x"2F",x"A6",x"77",x"23", -- 0x0458
    x"13",x"AF",x"D3",x"04",x"DB",x"03",x"2F",x"A6", -- 0x0460
    x"77",x"E1",x"01",x"20",x"00",x"09",x"C1",x"05", -- 0x0468
    x"C2",x"55",x"14",x"C9",x"7D",x"E6",x"07",x"D3", -- 0x0470
    x"02",x"C3",x"47",x"1A",x"C5",x"E5",x"7E",x"12", -- 0x0478
    x"13",x"23",x"0D",x"C2",x"7E",x"14",x"E1",x"01", -- 0x0480
    x"20",x"00",x"09",x"C1",x"05",x"C2",x"7C",x"14", -- 0x0488
    x"C9",x"CD",x"74",x"14",x"AF",x"32",x"61",x"20", -- 0x0490
    x"C5",x"E5",x"1A",x"D3",x"04",x"DB",x"03",x"F5", -- 0x0498
    x"A6",x"CA",x"A9",x"14",x"3E",x"01",x"32",x"61", -- 0x04A0
    x"20",x"F1",x"B6",x"77",x"23",x"13",x"AF",x"D3", -- 0x04A8
    x"04",x"DB",x"03",x"F5",x"A6",x"CA",x"BD",x"14", -- 0x04B0
    x"3E",x"01",x"32",x"61",x"20",x"F1",x"B6",x"77", -- 0x04B8
    x"E1",x"01",x"20",x"00",x"09",x"C1",x"05",x"C2", -- 0x04C0
    x"98",x"14",x"C9",x"AF",x"C5",x"77",x"01",x"20", -- 0x04C8
    x"00",x"09",x"C1",x"05",x"C2",x"CC",x"14",x"C9", -- 0x04D0
    x"3A",x"25",x"20",x"FE",x"05",x"C8",x"FE",x"02", -- 0x04D8
    x"C0",x"3A",x"29",x"20",x"FE",x"D8",x"47",x"D2", -- 0x04E0
    x"30",x"15",x"3A",x"02",x"20",x"A7",x"C8",x"78", -- 0x04E8
    x"FE",x"CE",x"D2",x"79",x"15",x"C6",x"06",x"47", -- 0x04F0
    x"3A",x"09",x"20",x"FE",x"90",x"D2",x"04",x"15", -- 0x04F8
    x"B8",x"D2",x"30",x"15",x"68",x"CD",x"62",x"15", -- 0x0500
    x"3A",x"2A",x"20",x"67",x"CD",x"6F",x"15",x"22", -- 0x0508
    x"64",x"20",x"3E",x"05",x"32",x"25",x"20",x"CD", -- 0x0510
    x"81",x"15",x"7E",x"A7",x"CA",x"30",x"15",x"36", -- 0x0518
    x"00",x"CD",x"5F",x"0A",x"CD",x"3B",x"1A",x"CD", -- 0x0520
    x"D3",x"15",x"3E",x"10",x"32",x"03",x"20",x"C9", -- 0x0528
    x"3E",x"03",x"32",x"25",x"20",x"C3",x"4A",x"15", -- 0x0530
    x"21",x"03",x"20",x"35",x"C0",x"2A",x"64",x"20", -- 0x0538
    x"06",x"10",x"CD",x"24",x"14",x"3E",x"04",x"32", -- 0x0540
    x"25",x"20",x"AF",x"32",x"02",x"20",x"06",x"F7", -- 0x0548
    x"C3",x"DC",x"19",x"00",x"0E",x"00",x"BC",x"D4", -- 0x0550
    x"90",x"15",x"BC",x"D0",x"C6",x"10",x"0C",x"C3", -- 0x0558
    x"5A",x"15",x"3A",x"09",x"20",x"65",x"CD",x"54", -- 0x0560
    x"15",x"41",x"05",x"DE",x"10",x"6F",x"C9",x"3A", -- 0x0568
    x"0A",x"20",x"CD",x"54",x"15",x"DE",x"10",x"67", -- 0x0570
    x"C9",x"3E",x"01",x"32",x"85",x"20",x"C3",x"45", -- 0x0578
    x"15",x"78",x"07",x"07",x"07",x"80",x"80",x"80", -- 0x0580
    x"81",x"3D",x"6F",x"3A",x"67",x"20",x"67",x"C9", -- 0x0588
    x"0C",x"C6",x"10",x"FA",x"90",x"15",x"C9",x"3A", -- 0x0590
    x"0D",x"20",x"A7",x"C2",x"B7",x"15",x"21",x"A4", -- 0x0598
    x"3E",x"CD",x"C5",x"15",x"D0",x"06",x"FE",x"3E", -- 0x05A0
    x"01",x"32",x"0D",x"20",x"78",x"32",x"08",x"20", -- 0x05A8
    x"3A",x"0E",x"20",x"32",x"07",x"20",x"C9",x"21", -- 0x05B0
    x"24",x"25",x"CD",x"C5",x"15",x"D0",x"CD",x"F1", -- 0x05B8
    x"18",x"AF",x"C3",x"A9",x"15",x"06",x"17",x"7E", -- 0x05C0
    x"A7",x"C2",x"6B",x"16",x"23",x"05",x"C2",x"C7", -- 0x05C8
    x"15",x"C9",x"00",x"CD",x"74",x"14",x"E5",x"C5", -- 0x05D0
    x"E5",x"1A",x"D3",x"04",x"DB",x"03",x"77",x"23", -- 0x05D8
    x"13",x"AF",x"D3",x"04",x"DB",x"03",x"77",x"E1", -- 0x05E0
    x"01",x"20",x"00",x"09",x"C1",x"05",x"C2",x"D7", -- 0x05E8
    x"15",x"E1",x"C9",x"CD",x"11",x"16",x"01",x"00", -- 0x05F0
    x"37",x"7E",x"A7",x"CA",x"FF",x"15",x"0C",x"23", -- 0x05F8
    x"05",x"C2",x"F9",x"15",x"79",x"32",x"82",x"20", -- 0x0600
    x"FE",x"01",x"C0",x"21",x"6B",x"20",x"36",x"01", -- 0x0608
    x"C9",x"2E",x"00",x"3A",x"67",x"20",x"67",x"C9", -- 0x0610
    x"3A",x"15",x"20",x"FE",x"FF",x"C0",x"21",x"10", -- 0x0618
    x"20",x"7E",x"23",x"46",x"B0",x"C0",x"3A",x"25", -- 0x0620
    x"20",x"A7",x"C0",x"3A",x"EF",x"20",x"A7",x"CA", -- 0x0628
    x"52",x"16",x"3A",x"2D",x"20",x"A7",x"C2",x"48", -- 0x0630
    x"16",x"CD",x"C0",x"17",x"E6",x"10",x"C8",x"3E", -- 0x0638
    x"01",x"32",x"25",x"20",x"32",x"2D",x"20",x"C9", -- 0x0640
    x"CD",x"C0",x"17",x"E6",x"10",x"C0",x"32",x"2D", -- 0x0648
    x"20",x"C9",x"21",x"25",x"20",x"36",x"01",x"2A", -- 0x0650
    x"ED",x"20",x"23",x"7D",x"FE",x"7E",x"DA",x"63", -- 0x0658
    x"16",x"2E",x"74",x"22",x"ED",x"20",x"7E",x"32", -- 0x0660
    x"1D",x"20",x"C9",x"37",x"C9",x"AF",x"CD",x"8B", -- 0x0668
    x"1A",x"CD",x"10",x"19",x"36",x"00",x"CD",x"CA", -- 0x0670
    x"09",x"23",x"11",x"F5",x"20",x"1A",x"BE",x"1B", -- 0x0678
    x"2B",x"1A",x"CA",x"8B",x"16",x"D2",x"98",x"16", -- 0x0680
    x"C3",x"8F",x"16",x"BE",x"D2",x"98",x"16",x"7E", -- 0x0688
    x"12",x"13",x"23",x"7E",x"12",x"CD",x"50",x"19", -- 0x0690
    x"3A",x"CE",x"20",x"A7",x"CA",x"C9",x"16",x"21", -- 0x0698
    x"03",x"28",x"11",x"A6",x"1A",x"0E",x"14",x"CD", -- 0x06A0
    x"93",x"0A",x"25",x"25",x"06",x"1B",x"3A",x"67", -- 0x06A8
    x"20",x"0F",x"DA",x"B7",x"16",x"06",x"1C",x"78", -- 0x06B0
    x"CD",x"FF",x"08",x"CD",x"B1",x"0A",x"CD",x"E7", -- 0x06B8
    x"18",x"7E",x"A7",x"CA",x"C9",x"16",x"C3",x"ED", -- 0x06C0
    x"02",x"21",x"18",x"2D",x"11",x"A6",x"1A",x"0E", -- 0x06C8
    x"0A",x"CD",x"93",x"0A",x"CD",x"B6",x"0A",x"CD", -- 0x06D0
    x"D6",x"09",x"AF",x"32",x"EF",x"20",x"D3",x"05", -- 0x06D8
    x"CD",x"D1",x"19",x"C3",x"89",x"0B",x"31",x"00", -- 0x06E0
    x"24",x"FB",x"AF",x"32",x"15",x"20",x"CD",x"D8", -- 0x06E8
    x"14",x"06",x"04",x"CD",x"FA",x"18",x"CD",x"59", -- 0x06F0
    x"0A",x"C2",x"EE",x"16",x"CD",x"D7",x"19",x"21", -- 0x06F8
    x"01",x"27",x"CD",x"FA",x"19",x"AF",x"CD",x"8B", -- 0x0700
    x"1A",x"06",x"FB",x"C3",x"6B",x"19",x"CD",x"CA", -- 0x0708
    x"09",x"23",x"7E",x"11",x"B8",x"1C",x"21",x"A1", -- 0x0710
    x"1A",x"0E",x"04",x"47",x"1A",x"B8",x"D2",x"27", -- 0x0718
    x"17",x"23",x"13",x"0D",x"C2",x"1C",x"17",x"7E", -- 0x0720
    x"32",x"CF",x"20",x"C9",x"3A",x"25",x"20",x"FE", -- 0x0728
    x"00",x"C2",x"39",x"17",x"06",x"FD",x"C3",x"DC", -- 0x0730
    x"19",x"06",x"02",x"C3",x"FA",x"18",x"00",x"00", -- 0x0738
    x"21",x"9B",x"20",x"35",x"CC",x"6D",x"17",x"3A", -- 0x0740
    x"68",x"20",x"A7",x"CA",x"6D",x"17",x"21",x"96", -- 0x0748
    x"20",x"35",x"C0",x"21",x"98",x"20",x"7E",x"D3", -- 0x0750
    x"05",x"3A",x"82",x"20",x"A7",x"CA",x"6D",x"17", -- 0x0758
    x"2B",x"7E",x"2B",x"77",x"2B",x"36",x"01",x"3E", -- 0x0760
    x"04",x"32",x"9B",x"20",x"C9",x"3A",x"98",x"20", -- 0x0768
    x"E6",x"30",x"D3",x"05",x"C9",x"3A",x"95",x"20", -- 0x0770
    x"A7",x"CA",x"AA",x"17",x"21",x"11",x"1A",x"11", -- 0x0778
    x"21",x"1A",x"3A",x"82",x"20",x"BE",x"D2",x"8E", -- 0x0780
    x"17",x"23",x"13",x"C3",x"85",x"17",x"1A",x"32", -- 0x0788
    x"97",x"20",x"21",x"98",x"20",x"7E",x"E6",x"30", -- 0x0790
    x"47",x"7E",x"E6",x"0F",x"07",x"FE",x"10",x"C2", -- 0x0798
    x"A4",x"17",x"3E",x"01",x"B0",x"77",x"AF",x"32", -- 0x07A0
    x"95",x"20",x"21",x"99",x"20",x"35",x"C0",x"06", -- 0x07A8
    x"EF",x"C3",x"DC",x"19",x"06",x"EF",x"21",x"98", -- 0x07B0
    x"20",x"7E",x"A0",x"77",x"D3",x"05",x"C9",x"00", -- 0x07B8
    x"3A",x"67",x"20",x"0F",x"D2",x"CA",x"17",x"DB", -- 0x07C0
    x"01",x"C9",x"DB",x"02",x"C9",x"DB",x"02",x"E6", -- 0x07C8
    x"04",x"C8",x"3A",x"9A",x"20",x"A7",x"C0",x"31", -- 0x07D0
    x"00",x"24",x"06",x"04",x"CD",x"D6",x"09",x"05", -- 0x07D8
    x"C2",x"DC",x"17",x"3E",x"01",x"32",x"9A",x"20", -- 0x07E0
    x"CD",x"D7",x"19",x"FB",x"11",x"BC",x"1C",x"21", -- 0x07E8
    x"16",x"30",x"0E",x"04",x"CD",x"93",x"0A",x"CD", -- 0x07F0
    x"B1",x"0A",x"AF",x"32",x"9A",x"20",x"32",x"93"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
