library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj3 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"04",X"1C",X"65",X"E1",X"F9",X"E9",X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"05",X"1D",X"65",X"E1",X"F9",X"D9",X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",
		X"00",X"03",X"07",X"07",X"1F",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"3F",X"3F",X"1C",X"00",X"00",
		X"00",X"07",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"3F",X"1F",X"03",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"03",
		X"00",X"00",X"01",X"03",X"1B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"1B",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E3",X"1F",X"1F",X"1F",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E1",X"F9",X"E9",X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E7",X"1F",X"1F",X"1F",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"64",X"E1",X"F9",X"E9",X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"71",X"1F",X"1F",X"1F",X"2A",X"26",X"22",X"02",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",
		X"01",X"03",X"07",X"1F",X"65",X"E1",X"F9",X"E9",X"C1",X"55",X"4D",X"45",X"05",X"01",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"6C",X"6F",X"7F",X"FF",X"DF",X"DF",X"DF",X"9F",X"1F",X"0F",X"0F",X"07",X"06",X"04",
		X"01",X"01",X"3B",X"7F",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"DF",X"67",X"31",X"10",X"10",X"00",
		X"10",X"10",X"3F",X"77",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"5F",X"77",X"3F",X"10",X"10",
		X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"06",X"06",X"03",X"01",
		X"00",X"00",X"03",X"07",X"0F",X"0D",X"1E",X"1F",X"1F",X"19",X"09",X"0F",X"07",X"03",X"00",X"00",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",
		X"00",X"00",X"00",X"1F",X"3F",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"3F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"0C",X"1B",X"1A",X"19",X"18",X"0C",X"0F",X"07",X"03",X"00",X"00",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1E",X"3F",X"3F",X"3F",X"7D",X"7F",X"3E",X"1E",X"3F",X"7D",X"3F",X"1F",X"0C",X"00",X"0F",
		X"00",X"1E",X"3F",X"3F",X"3F",X"6F",X"7F",X"3E",X"1E",X"3F",X"7F",X"3F",X"1B",X"0C",X"00",X"0F",
		X"00",X"1E",X"3B",X"3F",X"3F",X"7F",X"7F",X"3E",X"1E",X"3F",X"77",X"3F",X"1F",X"0C",X"00",X"0F",
		X"0F",X"01",X"09",X"1F",X"3F",X"3F",X"1A",X"0E",X"1A",X"3F",X"3F",X"1F",X"09",X"01",X"01",X"0F",
		X"0F",X"01",X"09",X"1F",X"3F",X"3F",X"1A",X"0E",X"1A",X"3F",X"3F",X"1F",X"09",X"01",X"01",X"0F",
		X"38",X"FC",X"FF",X"EF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"EF",X"FF",X"FC",X"38",
		X"00",X"00",X"09",X"00",X"00",X"08",X"08",X"08",X"08",X"04",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"08",X"00",X"00",X"48",X"B4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"3C",X"7C",X"7F",X"FF",X"FC",X"FC",X"FC",X"78",X"20",X"00",X"00",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"60",X"00",X"10",X"08",X"08",X"04",X"02",X"02",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"04",X"04",X"01",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"C0",X"78",X"00",X"00",X"00",X"00",X"00",X"17",X"E7",X"87",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"40",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"87",X"C7",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"08",X"09",X"09",X"08",X"10",X"10",X"10",
		X"03",X"07",X"07",X"03",X"08",X"1C",X"1E",X"3F",X"3F",X"3B",X"1F",X"03",X"03",X"03",X"01",X"00",
		X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"80",X"C0",X"40",X"61",X"3A",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"32",X"41",X"40",X"80",X"00",X"00",
		X"60",X"F0",X"A0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"0E",X"08",X"00",X"00",
		X"0C",X"0C",X"06",X"06",X"06",X"04",X"08",X"10",X"20",X"00",X"80",X"60",X"18",X"0C",X"00",X"00",
		X"00",X"18",X"20",X"40",X"80",X"00",X"00",X"21",X"11",X"09",X"04",X"04",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"15",X"15",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"02",X"01",X"05",X"43",X"0F",X"16",X"03",X"0E",X"5B",X"21",X"00",X"00",X"00",X"00",
		X"00",X"00",X"28",X"87",X"33",X"1E",X"0C",X"44",X"32",X"1E",X"0D",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"12",X"01",X"00",X"22",X"00",X"02",X"40",X"10",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"20",X"00",X"43",X"10",X"00",X"00",X"40",X"21",X"02",X"00",X"00",X"00",X"00",
		X"80",X"0A",X"75",X"1A",X"09",X"04",X"2F",X"50",X"9C",X"0E",X"06",X"35",X"4A",X"07",X"00",X"20",
		X"08",X"80",X"00",X"00",X"09",X"86",X"40",X"01",X"02",X"14",X"09",X"00",X"01",X"A6",X"43",X"00",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"0D",X"2D",X"0D",X"2F",X"07",X"03",X"31",X"79",X"79",X"31",X"03",X"07",X"2F",X"0D",X"2D",X"0D",
		X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"7F",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"01",X"06",X"0D",X"05",X"07",X"02",X"07",X"02",X"02",X"01",X"01",X"00",X"00",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7E",X"F9",X"F8",X"70",X"30",X"10",
		X"02",X"00",X"05",X"02",X"01",X"03",X"06",X"04",X"09",X"09",X"09",X"09",X"0C",X"06",X"03",X"00",
		X"00",X"00",X"01",X"00",X"01",X"03",X"06",X"04",X"09",X"09",X"09",X"09",X"0D",X"06",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0C",X"18",X"30",X"30",X"30",X"30",X"30",X"30",X"18",X"0C",X"07",X"03",X"00",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"0C",X"0C",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"38",X"00",X"00",X"04",X"08",X"10",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"1E",X"3F",X"3F",X"7F",X"7E",X"7E",X"7F",X"7E",X"7F",X"3F",X"3F",X"1E",X"0F",X"07",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1D",X"08",X"02",X"17",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",
		X"00",X"01",X"0D",X"1C",X"61",X"C9",X"ED",X"C7",X"C7",X"ED",X"C9",X"61",X"9C",X"0D",X"01",X"00",
		X"03",X"07",X"05",X"08",X"1B",X"19",X"05",X"3F",X"3F",X"0F",X"05",X"37",X"3F",X"3F",X"3E",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"0C",X"0E",X"0F",X"0F",X"07",X"03",X"00",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"09",X"0A",X"0A",X"0A",X"0E",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
