library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_cpu is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"C3",X"40",X"00",X"00",X"00",X"C3",X"C6",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"08",X"3A",X"7C",X"E0",X"A7",X"C0",X"08",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"C9",
		X"08",X"3A",X"7C",X"E0",X"A7",X"C0",X"3A",X"AE",X"E2",X"47",X"08",X"B8",X"C8",X"32",X"AE",X"E2",
		X"18",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"CD",X"4B",X"2F",X"FB",X"ED",X"4D",X"00",
		X"31",X"00",X"E8",X"3E",X"55",X"06",X"03",X"D9",X"21",X"00",X"E0",X"11",X"01",X"E0",X"01",X"FF",
		X"07",X"77",X"BE",X"C2",X"F6",X"1E",X"ED",X"A0",X"EA",X"52",X"00",X"D9",X"87",X"30",X"01",X"AF",
		X"10",X"E5",X"CD",X"9A",X"09",X"D7",X"CD",X"8C",X"01",X"21",X"34",X"12",X"22",X"68",X"E0",X"CD",
		X"BA",X"04",X"CD",X"30",X"0B",X"FB",X"3E",X"01",X"32",X"7C",X"E0",X"3A",X"00",X"E0",X"A7",X"20",
		X"02",X"18",X"F8",X"AF",X"32",X"7C",X"E0",X"CD",X"B1",X"2C",X"21",X"50",X"E0",X"06",X"B0",X"CD",
		X"E9",X"1E",X"06",X"06",X"CD",X"EE",X"1E",X"CD",X"E0",X"05",X"CD",X"EF",X"0A",X"CD",X"B3",X"09",
		X"3A",X"00",X"D0",X"2F",X"E6",X"03",X"4F",X"3A",X"00",X"E0",X"CB",X"3F",X"28",X"04",X"CB",X"49",
		X"20",X"06",X"CB",X"41",X"20",X"02",X"18",X"E2",X"79",X"CB",X"3F",X"4F",X"3A",X"0B",X"E0",X"E6",
		X"01",X"CB",X"27",X"81",X"21",X"00",X"E0",X"5F",X"0F",X"30",X"0D",X"35",X"CB",X"EB",X"3E",X"64",
		X"32",X"F9",X"E0",X"3E",X"01",X"32",X"F8",X"E0",X"35",X"CB",X"E3",X"3E",X"64",X"32",X"F0",X"E0",
		X"3E",X"01",X"32",X"EF",X"E0",X"CB",X"BB",X"7B",X"32",X"6A",X"E0",X"AF",X"32",X"6D",X"E0",X"CD",
		X"4A",X"02",X"3E",X"1C",X"D7",X"06",X"0C",X"3E",X"FF",X"CD",X"DE",X"1E",X"10",X"F9",X"3E",X"01",
		X"32",X"6D",X"E0",X"3A",X"C8",X"E4",X"A7",X"20",X"FA",X"3E",X"01",X"32",X"63",X"E0",X"3A",X"A8",
		X"E2",X"47",X"3A",X"6B",X"E0",X"80",X"28",X"F6",X"21",X"63",X"E0",X"4E",X"AF",X"77",X"79",X"FE",
		X"03",X"20",X"05",X"3E",X"01",X"32",X"C8",X"E4",X"CD",X"1F",X"10",X"21",X"6A",X"E0",X"28",X"1F",
		X"CB",X"BE",X"79",X"FE",X"03",X"C4",X"F5",X"1D",X"CD",X"97",X"05",X"3A",X"6B",X"E0",X"A7",X"C2",
		X"EB",X"00",X"CD",X"E0",X"05",X"CD",X"6D",X"05",X"21",X"6A",X"E0",X"CB",X"AE",X"18",X"1D",X"CB",
		X"FE",X"79",X"FE",X"03",X"C4",X"D6",X"1D",X"CD",X"7E",X"05",X"3A",X"6B",X"E0",X"A7",X"C2",X"EB",
		X"00",X"CD",X"E0",X"05",X"CD",X"36",X"05",X"21",X"6A",X"E0",X"CB",X"A6",X"7E",X"E6",X"30",X"C2",
		X"EB",X"00",X"CD",X"A0",X"05",X"C3",X"76",X"00",X"8F",X"C0",X"14",X"40",X"8F",X"C0",X"15",X"30",
		X"8F",X"C0",X"00",X"40",X"8F",X"C0",X"00",X"30",X"8F",X"C0",X"00",X"40",X"AF",X"21",X"A0",X"C9",
		X"06",X"60",X"CD",X"E9",X"1E",X"C9",X"3A",X"83",X"E2",X"0F",X"D0",X"3A",X"6D",X"E0",X"A7",X"C8",
		X"FE",X"01",X"CC",X"04",X"02",X"CD",X"CB",X"01",X"CD",X"08",X"02",X"21",X"6D",X"E0",X"34",X"7E",
		X"FE",X"C0",X"D8",X"AF",X"32",X"C8",X"E4",X"32",X"6D",X"E0",X"21",X"E0",X"E1",X"06",X"0C",X"CD",
		X"E9",X"1E",X"21",X"B8",X"E1",X"06",X"08",X"CD",X"E9",X"1E",X"C9",X"DD",X"21",X"E0",X"E1",X"3A",
		X"6D",X"E0",X"FE",X"35",X"D8",X"FE",X"6A",X"38",X"1E",X"FE",X"9F",X"38",X"0D",X"DD",X"36",X"01",
		X"03",X"DD",X"36",X"05",X"02",X"DD",X"36",X"09",X"01",X"C9",X"DD",X"36",X"01",X"03",X"DD",X"36",
		X"05",X"03",X"DD",X"36",X"09",X"03",X"C9",X"DD",X"36",X"01",X"02",X"DD",X"36",X"05",X"02",X"DD",
		X"36",X"09",X"03",X"C9",X"3E",X"11",X"D7",X"C9",X"DD",X"21",X"B8",X"E1",X"3A",X"6D",X"E0",X"4F",
		X"21",X"43",X"02",X"06",X"07",X"7E",X"B9",X"28",X"04",X"23",X"10",X"F9",X"C9",X"78",X"ED",X"44",
		X"C6",X"07",X"CB",X"27",X"4F",X"06",X"00",X"21",X"35",X"02",X"09",X"7E",X"DD",X"77",X"02",X"23",
		X"7E",X"DD",X"77",X"06",X"C9",X"AB",X"AC",X"AD",X"AC",X"AE",X"AF",X"B0",X"AF",X"B1",X"B2",X"B3",
		X"B4",X"B5",X"B6",X"78",X"85",X"92",X"A0",X"A4",X"A6",X"A8",X"CD",X"E0",X"05",X"AF",X"32",X"6B",
		X"E0",X"21",X"6A",X"E0",X"CB",X"46",X"28",X"32",X"CB",X"7E",X"28",X"1F",X"CB",X"6E",X"28",X"1B",
		X"CB",X"FE",X"CB",X"4E",X"28",X"05",X"21",X"01",X"D0",X"CB",X"C6",X"21",X"F7",X"E0",X"11",X"C7",
		X"E4",X"01",X"09",X"00",X"ED",X"B0",X"CD",X"F3",X"04",X"18",X"1D",X"CB",X"66",X"28",X"DD",X"CB",
		X"BE",X"CB",X"4E",X"28",X"05",X"21",X"01",X"D0",X"CB",X"86",X"21",X"EE",X"E0",X"11",X"C7",X"E4",
		X"01",X"09",X"00",X"ED",X"B0",X"CD",X"F9",X"04",X"3E",X"FF",X"32",X"C0",X"E4",X"3A",X"7C",X"E0",
		X"A7",X"20",X"07",X"F3",X"CD",X"C8",X"2B",X"FB",X"18",X"03",X"CD",X"C8",X"2B",X"CD",X"F3",X"05",
		X"CD",X"72",X"1A",X"CD",X"05",X"17",X"CD",X"6F",X"17",X"CD",X"15",X"06",X"3A",X"6A",X"E0",X"0F",
		X"DC",X"59",X"06",X"CD",X"F6",X"02",X"3A",X"C8",X"E4",X"0F",X"DC",X"CE",X"02",X"C9",X"21",X"E2",
		X"02",X"11",X"E0",X"E1",X"01",X"0C",X"00",X"ED",X"B0",X"11",X"B8",X"E1",X"01",X"08",X"00",X"ED",
		X"B0",X"C9",X"88",X"03",X"FF",X"D8",X"98",X"02",X"FE",X"D8",X"A8",X"03",X"FF",X"D8",X"50",X"45",
		X"A9",X"60",X"50",X"45",X"AA",X"50",X"06",X"03",X"11",X"60",X"E1",X"C5",X"21",X"78",X"01",X"01",
		X"14",X"00",X"ED",X"B0",X"E5",X"21",X"4C",X"00",X"19",X"EB",X"E1",X"C1",X"10",X"ED",X"DD",X"21",
		X"C0",X"E1",X"3A",X"CB",X"E4",X"FE",X"A0",X"3E",X"18",X"30",X"02",X"ED",X"44",X"4F",X"DD",X"E5",
		X"DD",X"21",X"C4",X"E1",X"CD",X"7B",X"1F",X"DD",X"E1",X"D0",X"DD",X"E5",X"11",X"04",X"00",X"DD",
		X"7E",X"00",X"81",X"06",X"04",X"CD",X"9E",X"1E",X"DD",X"19",X"10",X"F9",X"DD",X"E1",X"18",X"DD",
		X"AF",X"DD",X"21",X"C0",X"E1",X"DD",X"E5",X"D9",X"5F",X"06",X"02",X"FD",X"7E",X"00",X"A7",X"28",
		X"2F",X"FD",X"7E",X"02",X"A7",X"28",X"29",X"DD",X"7E",X"00",X"A7",X"28",X"23",X"DD",X"7E",X"02",
		X"A7",X"28",X"1D",X"DD",X"7E",X"00",X"C6",X"04",X"FD",X"56",X"00",X"CD",X"A6",X"03",X"A7",X"CA",
		X"80",X"03",X"DD",X"7E",X"03",X"C6",X"04",X"FD",X"56",X"03",X"CD",X"8E",X"03",X"A7",X"20",X"0A",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"C1",X"D9",X"DD",X"E1",X"C9",X"67",X"2E",
		X"30",X"CB",X"43",X"20",X"0D",X"CD",X"B3",X"03",X"A7",X"C0",X"7C",X"C6",X"08",X"67",X"CD",X"B3",
		X"03",X"C9",X"2E",X"20",X"18",X"EF",X"67",X"2E",X"20",X"CB",X"43",X"CA",X"95",X"03",X"2E",X"10",
		X"C3",X"95",X"03",X"7C",X"BA",X"38",X"08",X"7A",X"85",X"BC",X"38",X"03",X"3E",X"01",X"C9",X"AF",
		X"C9",X"3A",X"7B",X"E0",X"F5",X"A7",X"20",X"12",X"CD",X"E0",X"05",X"CD",X"FE",X"2C",X"CD",X"C0",
		X"2C",X"CD",X"98",X"0A",X"CD",X"D2",X"09",X"CD",X"B3",X"09",X"F1",X"C6",X"01",X"38",X"04",X"32",
		X"7B",X"E0",X"C9",X"AF",X"32",X"7B",X"E0",X"21",X"7C",X"E0",X"34",X"28",X"FD",X"CD",X"B1",X"2C",
		X"C9",X"3A",X"7B",X"E0",X"F5",X"A7",X"20",X"E2",X"CD",X"E0",X"05",X"CD",X"FE",X"2C",X"CD",X"09",
		X"04",X"CD",X"63",X"04",X"CD",X"B3",X"09",X"18",X"D1",X"21",X"43",X"04",X"11",X"2D",X"8B",X"01",
		X"0E",X"00",X"CF",X"21",X"35",X"04",X"11",X"2C",X"8B",X"01",X"0E",X"00",X"CF",X"11",X"27",X"8C",
		X"06",X"05",X"C5",X"D5",X"21",X"51",X"04",X"01",X"12",X"00",X"CF",X"D1",X"21",X"FC",X"FF",X"19",
		X"EB",X"C1",X"10",X"EE",X"C9",X"42",X"45",X"53",X"54",X"20",X"35",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"53",X"09",X"09",X"09",X"09",X"09",X"05",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"09",X"06",X"06",X"06",X"05",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"05",X"05",X"05",X"11",X"26",X"8C",X"21",X"13",X"E0",X"06",X"05",X"E5",X"DD",X"E1",X"E5",X"D5",
		X"C5",X"21",X"98",X"04",X"01",X"04",X"00",X"CF",X"1B",X"E3",X"7C",X"E3",X"ED",X"44",X"C6",X"36",
		X"12",X"CD",X"9C",X"04",X"CD",X"A9",X"04",X"C1",X"D1",X"21",X"FC",X"FF",X"19",X"EB",X"E1",X"D5",
		X"11",X"09",X"00",X"19",X"D1",X"10",X"D4",X"C9",X"4E",X"4F",X"2E",X"20",X"21",X"80",X"FE",X"19",
		X"EB",X"DD",X"E5",X"E1",X"EB",X"CD",X"99",X"06",X"C9",X"11",X"80",X"FE",X"19",X"EB",X"DD",X"E5",
		X"E1",X"01",X"06",X"00",X"09",X"01",X"03",X"00",X"CF",X"C9",X"21",X"C6",X"04",X"11",X"13",X"E0",
		X"01",X"2D",X"00",X"ED",X"B0",X"C9",X"00",X"00",X"00",X"02",X"00",X"00",X"48",X"45",X"42",X"00",
		X"00",X"00",X"02",X"00",X"00",X"54",X"41",X"4B",X"00",X"00",X"00",X"02",X"00",X"00",X"41",X"4E",
		X"4A",X"00",X"00",X"00",X"02",X"00",X"00",X"53",X"41",X"4F",X"00",X"00",X"00",X"02",X"00",X"00",
		X"43",X"4F",X"4D",X"21",X"21",X"05",X"C3",X"FC",X"04",X"21",X"29",X"05",X"3A",X"7C",X"E0",X"A7",
		X"C0",X"3A",X"C8",X"E4",X"A7",X"C8",X"11",X"26",X"8A",X"01",X"08",X"00",X"CF",X"21",X"31",X"05",
		X"11",X"A2",X"89",X"01",X"05",X"00",X"CF",X"06",X"06",X"3E",X"FF",X"CD",X"DE",X"1E",X"10",X"F9",
		X"C9",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",
		X"31",X"52",X"45",X"41",X"44",X"59",X"CD",X"6D",X"07",X"3A",X"6A",X"E0",X"0F",X"D0",X"21",X"5B",
		X"05",X"E5",X"CD",X"E0",X"05",X"E1",X"11",X"26",X"8A",X"01",X"08",X"00",X"CF",X"21",X"63",X"05",
		X"11",X"A2",X"8A",X"01",X"0A",X"00",X"CF",X"CD",X"CC",X"05",X"C9",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"20",X"31",X"47",X"41",X"4D",X"45",X"20",X"20",X"4F",X"56",X"45",X"52",X"CD",X"7A",X"07",
		X"21",X"76",X"05",X"C3",X"41",X"05",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"21",X"C7",
		X"E4",X"11",X"EE",X"E0",X"01",X"09",X"00",X"ED",X"B0",X"AF",X"32",X"A6",X"E2",X"21",X"00",X"E1",
		X"06",X"06",X"CD",X"EE",X"1E",X"D7",X"C9",X"21",X"C7",X"E4",X"11",X"F7",X"E0",X"C3",X"84",X"05",
		X"AF",X"21",X"63",X"E0",X"06",X"9D",X"CD",X"E9",X"1E",X"06",X"06",X"CD",X"EE",X"1E",X"32",X"01",
		X"D0",X"D7",X"CD",X"E0",X"05",X"3E",X"1B",X"D7",X"21",X"D6",X"05",X"11",X"22",X"8A",X"01",X"0A",
		X"00",X"CF",X"11",X"23",X"8A",X"06",X"0A",X"3E",X"05",X"CD",X"D3",X"1E",X"06",X"0B",X"3E",X"FF",
		X"CD",X"DE",X"1E",X"10",X"F9",X"C9",X"47",X"41",X"4D",X"45",X"20",X"20",X"4F",X"56",X"45",X"52",
		X"AF",X"21",X"00",X"80",X"06",X"10",X"CD",X"EE",X"1E",X"32",X"00",X"90",X"32",X"00",X"A0",X"CD",
		X"8C",X"01",X"C9",X"21",X"C3",X"06",X"11",X"BC",X"8F",X"01",X"08",X"00",X"CF",X"11",X"BD",X"8F",
		X"01",X"08",X"00",X"CF",X"11",X"BB",X"8F",X"01",X"08",X"00",X"CF",X"CD",X"28",X"07",X"21",X"3A",
		X"8F",X"CD",X"99",X"06",X"C9",X"3A",X"63",X"E0",X"A7",X"CA",X"37",X"06",X"CD",X"1F",X"10",X"C2",
		X"37",X"06",X"3A",X"83",X"E2",X"CB",X"5F",X"CA",X"37",X"06",X"21",X"E9",X"06",X"11",X"38",X"8F",
		X"01",X"03",X"00",X"CF",X"C3",X"4F",X"06",X"21",X"DB",X"06",X"11",X"38",X"8F",X"01",X"03",X"00",
		X"CF",X"11",X"39",X"8F",X"01",X"03",X"00",X"CF",X"11",X"B7",X"8F",X"01",X"08",X"00",X"CF",X"11",
		X"50",X"E0",X"21",X"36",X"8F",X"CD",X"99",X"06",X"C9",X"3A",X"63",X"E0",X"A7",X"CA",X"7B",X"06",
		X"CD",X"1F",X"10",X"CA",X"7B",X"06",X"3A",X"83",X"E2",X"CB",X"5F",X"CA",X"7B",X"06",X"21",X"E9",
		X"06",X"11",X"34",X"8F",X"01",X"03",X"00",X"CF",X"C3",X"93",X"06",X"21",X"EC",X"06",X"11",X"34",
		X"8F",X"01",X"03",X"00",X"CF",X"11",X"35",X"8F",X"01",X"03",X"00",X"CF",X"11",X"B3",X"8F",X"01",
		X"08",X"00",X"CF",X"11",X"59",X"E0",X"21",X"32",X"8F",X"06",X"06",X"1A",X"F5",X"13",X"10",X"FB",
		X"06",X"06",X"11",X"80",X"FF",X"F1",X"A7",X"C2",X"B9",X"06",X"AF",X"77",X"19",X"10",X"F6",X"A7",
		X"ED",X"52",X"3E",X"30",X"77",X"19",X"77",X"C9",X"F1",X"C6",X"30",X"77",X"19",X"10",X"F9",X"3E",
		X"30",X"77",X"C9",X"48",X"49",X"2D",X"53",X"43",X"4F",X"52",X"45",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"55",X"50",X"0D",X"0D",
		X"0D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"32",X"55",X"50",X"0D",
		X"0D",X"0D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"CD",X"1F",X"10",X"C2",X"0C",X"07",
		X"3A",X"7C",X"E0",X"A7",X"C0",X"21",X"50",X"E0",X"CD",X"0F",X"07",X"C9",X"21",X"59",X"E0",X"78",
		X"A7",X"C8",X"0E",X"06",X"5D",X"54",X"34",X"7E",X"FE",X"0A",X"38",X"07",X"36",X"00",X"23",X"0D",
		X"20",X"F4",X"C9",X"6B",X"62",X"10",X"EB",X"C9",X"11",X"5E",X"E0",X"21",X"55",X"E0",X"CD",X"56",
		X"07",X"A7",X"CA",X"3B",X"07",X"11",X"5E",X"E0",X"C3",X"3E",X"07",X"11",X"55",X"E0",X"21",X"18",
		X"E0",X"CD",X"56",X"07",X"A7",X"C2",X"4C",X"07",X"11",X"13",X"E0",X"C9",X"EB",X"05",X"48",X"06",
		X"00",X"A7",X"ED",X"42",X"EB",X"C9",X"06",X"06",X"4E",X"1A",X"B9",X"DA",X"68",X"07",X"CA",X"64",
		X"07",X"C3",X"6A",X"07",X"2B",X"1B",X"10",X"F0",X"AF",X"C9",X"3E",X"01",X"C9",X"11",X"55",X"E0",
		X"CD",X"87",X"07",X"3A",X"8D",X"E2",X"CD",X"E0",X"07",X"C9",X"11",X"5E",X"E0",X"CD",X"87",X"07",
		X"3A",X"8D",X"E2",X"CD",X"E0",X"07",X"C9",X"21",X"18",X"E0",X"06",X"05",X"E5",X"D5",X"C5",X"CD",
		X"56",X"07",X"A7",X"C2",X"A7",X"07",X"C1",X"D1",X"E1",X"D5",X"11",X"09",X"00",X"19",X"D1",X"10",
		X"EB",X"3E",X"0F",X"32",X"8D",X"E2",X"C9",X"C1",X"78",X"ED",X"44",X"C6",X"05",X"32",X"8D",X"E2",
		X"78",X"01",X"FB",X"FF",X"E1",X"09",X"D1",X"EB",X"09",X"EB",X"3D",X"47",X"A7",X"C4",X"C6",X"07",
		X"01",X"09",X"00",X"ED",X"B0",X"C9",X"E5",X"D5",X"C5",X"EB",X"3E",X"09",X"CD",X"0E",X"20",X"3A",
		X"87",X"E2",X"3D",X"06",X"00",X"4F",X"09",X"11",X"3F",X"E0",X"ED",X"B8",X"C1",X"D1",X"E1",X"C9",
		X"FE",X"05",X"D0",X"F5",X"3E",X"21",X"D7",X"CD",X"F2",X"07",X"CD",X"28",X"08",X"F1",X"CD",X"55",
		X"08",X"C9",X"21",X"04",X"08",X"11",X"2E",X"8B",X"01",X"10",X"00",X"CF",X"11",X"2A",X"8C",X"01",
		X"14",X"00",X"CF",X"C9",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",
		X"4F",X"4E",X"53",X"21",X"59",X"4F",X"55",X"20",X"41",X"52",X"45",X"20",X"47",X"52",X"45",X"41",
		X"54",X"20",X"52",X"49",X"44",X"45",X"52",X"2E",X"CD",X"40",X"08",X"21",X"F7",X"31",X"11",X"A6",
		X"8B",X"06",X"0A",X"C5",X"D5",X"01",X"10",X"00",X"CF",X"D1",X"1B",X"1B",X"C1",X"10",X"F4",X"C9",
		X"11",X"95",X"8B",X"06",X"0A",X"C5",X"D5",X"06",X"10",X"3E",X"A7",X"CD",X"D3",X"1E",X"D1",X"13",
		X"13",X"C1",X"10",X"F1",X"C9",X"AF",X"32",X"BD",X"E2",X"21",X"9C",X"88",X"E5",X"EB",X"13",X"3E",
		X"08",X"06",X"03",X"CD",X"D3",X"1E",X"E1",X"AF",X"32",X"BB",X"E2",X"3E",X"41",X"77",X"32",X"BE",
		X"E2",X"E5",X"06",X"03",X"3E",X"70",X"CD",X"DE",X"1E",X"CD",X"C3",X"08",X"FE",X"03",X"CA",X"96",
		X"08",X"FE",X"02",X"F5",X"CC",X"42",X"09",X"F1",X"FE",X"01",X"CC",X"53",X"09",X"CD",X"35",X"09",
		X"DA",X"9E",X"08",X"C3",X"74",X"08",X"A7",X"11",X"80",X"00",X"ED",X"52",X"10",X"D6",X"11",X"13",
		X"E0",X"3A",X"8D",X"E2",X"06",X"09",X"CD",X"0E",X"20",X"2A",X"87",X"E2",X"19",X"11",X"06",X"00",
		X"19",X"EB",X"E1",X"06",X"03",X"C5",X"7E",X"12",X"01",X"80",X"00",X"A7",X"ED",X"42",X"13",X"C1",
		X"10",X"F3",X"C9",X"0E",X"03",X"3A",X"6A",X"E0",X"CB",X"47",X"28",X"34",X"CB",X"7F",X"20",X"30",
		X"3A",X"01",X"D0",X"2F",X"E6",X"04",X"CB",X"57",X"20",X"18",X"3A",X"11",X"E0",X"CB",X"97",X"32",
		X"11",X"E0",X"3A",X"02",X"D0",X"2F",X"E6",X"0C",X"CB",X"57",X"20",X"46",X"CB",X"5F",X"20",X"41",
		X"18",X"3E",X"3A",X"11",X"E0",X"CB",X"57",X"20",X"E9",X"CB",X"D7",X"32",X"11",X"E0",X"18",X"33",
		X"3A",X"01",X"D0",X"2F",X"E6",X"80",X"CB",X"7F",X"20",X"18",X"3A",X"11",X"E0",X"CB",X"BF",X"32",
		X"11",X"E0",X"3A",X"01",X"D0",X"2F",X"E6",X"03",X"CB",X"4F",X"20",X"16",X"CB",X"47",X"20",X"11",
		X"18",X"0E",X"3A",X"11",X"E0",X"CB",X"7F",X"20",X"E9",X"CB",X"FF",X"32",X"11",X"E0",X"18",X"03",
		X"0D",X"0D",X"0D",X"79",X"C9",X"3A",X"BE",X"E2",X"77",X"3A",X"BB",X"E2",X"C6",X"01",X"32",X"BB",
		X"E2",X"C9",X"AF",X"32",X"BB",X"E2",X"3A",X"BD",X"E2",X"D6",X"01",X"D2",X"61",X"09",X"3E",X"24",
		X"C3",X"61",X"09",X"AF",X"32",X"BB",X"E2",X"3A",X"BD",X"E2",X"3C",X"FE",X"25",X"DA",X"61",X"09",
		X"AF",X"C5",X"32",X"BD",X"E2",X"E5",X"21",X"75",X"09",X"4F",X"06",X"00",X"09",X"7E",X"E1",X"77",
		X"32",X"BE",X"E2",X"C1",X"C9",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",
		X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"2E",
		X"2C",X"21",X"22",X"23",X"26",X"3D",X"2D",X"3A",X"3F",X"20",X"21",X"AC",X"09",X"11",X"B8",X"83",
		X"01",X"07",X"00",X"CF",X"F5",X"3E",X"FF",X"CD",X"DE",X"1E",X"F1",X"C9",X"52",X"41",X"4D",X"20",
		X"20",X"4F",X"4B",X"21",X"CB",X"09",X"11",X"02",X"85",X"01",X"07",X"00",X"D5",X"CF",X"D1",X"13",
		X"06",X"07",X"3E",X"01",X"CD",X"D3",X"1E",X"CD",X"B8",X"0A",X"C9",X"43",X"52",X"45",X"44",X"49",
		X"54",X"20",X"0E",X"00",X"3A",X"03",X"E0",X"57",X"CB",X"3F",X"CA",X"DF",X"09",X"CB",X"C1",X"3A",
		X"05",X"E0",X"5F",X"CB",X"3F",X"CA",X"EA",X"09",X"CB",X"C9",X"21",X"48",X"0A",X"D5",X"E5",X"79",
		X"06",X"14",X"CD",X"0E",X"20",X"2A",X"87",X"E2",X"EB",X"E1",X"19",X"11",X"9C",X"8C",X"01",X"14",
		X"00",X"CF",X"D1",X"7A",X"C6",X"30",X"32",X"9C",X"8C",X"7B",X"C6",X"30",X"32",X"9C",X"87",X"D5",
		X"21",X"84",X"0A",X"11",X"98",X"8C",X"01",X"14",X"00",X"CF",X"D1",X"7A",X"CB",X"27",X"FE",X"0A",
		X"DA",X"2C",X"0A",X"D6",X"0A",X"47",X"3E",X"31",X"32",X"18",X"8D",X"78",X"C6",X"30",X"32",X"98",
		X"8C",X"7B",X"CB",X"27",X"FE",X"0A",X"DA",X"42",X"0A",X"D6",X"0A",X"47",X"3E",X"31",X"32",X"18",
		X"88",X"78",X"C6",X"30",X"32",X"98",X"87",X"C9",X"20",X"20",X"20",X"43",X"4F",X"49",X"4E",X"20",
		X"20",X"20",X"20",X"20",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"20",X"20",X"20",X"43",
		X"4F",X"49",X"4E",X"53",X"20",X"20",X"20",X"20",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"20",
		X"20",X"20",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"20",X"20",X"20",X"20",X"43",X"52",X"45",
		X"44",X"49",X"54",X"53",X"20",X"20",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"20",X"20",X"20",
		X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"21",X"AD",X"0A",X"11",X"94",X"8A",X"01",X"0B",
		X"00",X"CF",X"11",X"95",X"8A",X"06",X"0B",X"3E",X"07",X"CD",X"D3",X"1E",X"C9",X"49",X"4E",X"53",
		X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"06",X"00",X"3A",X"00",X"E0",X"FD",X"21",X"82",
		X"81",X"FE",X"0A",X"38",X"05",X"04",X"D6",X"0A",X"18",X"F7",X"4F",X"78",X"CB",X"27",X"CB",X"27",
		X"CB",X"27",X"CB",X"27",X"81",X"FE",X"63",X"38",X"04",X"0E",X"09",X"06",X"09",X"78",X"C6",X"30",
		X"FD",X"77",X"00",X"79",X"C6",X"30",X"01",X"80",X"FF",X"FD",X"09",X"FD",X"77",X"00",X"C9",X"21",
		X"10",X"0B",X"3A",X"00",X"E0",X"CB",X"3F",X"CA",X"FE",X"0A",X"11",X"10",X"00",X"19",X"11",X"A6",
		X"8B",X"01",X"10",X"00",X"CF",X"11",X"A7",X"8B",X"06",X"10",X"3E",X"08",X"CD",X"D3",X"1E",X"C9",
		X"50",X"55",X"53",X"48",X"20",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",
		X"50",X"55",X"53",X"48",X"20",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",
		X"3A",X"03",X"D0",X"2F",X"E6",X"07",X"21",X"91",X"0B",X"A7",X"CA",X"43",X"0B",X"23",X"23",X"3D",
		X"C3",X"39",X"0B",X"7E",X"32",X"03",X"E0",X"23",X"7E",X"32",X"05",X"E0",X"3A",X"03",X"D0",X"2F",
		X"E6",X"18",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"A1",X"0B",X"A7",X"CA",X"65",X"0B",X"23",
		X"23",X"3D",X"C3",X"5B",X"0B",X"7E",X"32",X"04",X"E0",X"23",X"7E",X"32",X"06",X"E0",X"3A",X"04",
		X"D0",X"2F",X"4F",X"CB",X"3F",X"E6",X"01",X"32",X"07",X"E0",X"79",X"CB",X"3F",X"CB",X"3F",X"E6",
		X"01",X"32",X"0A",X"E0",X"79",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"01",X"32",X"0B",X"E0",
		X"C9",X"01",X"01",X"02",X"01",X"01",X"03",X"04",X"01",X"01",X"02",X"03",X"01",X"01",X"05",X"05",
		X"01",X"01",X"01",X"02",X"01",X"01",X"02",X"03",X"01",X"3A",X"BE",X"E5",X"A7",X"C8",X"4F",X"06",
		X"0A",X"C5",X"41",X"CD",X"FA",X"06",X"C1",X"10",X"F8",X"AF",X"32",X"BE",X"E5",X"3A",X"A7",X"E2",
		X"A7",X"C2",X"D6",X"0B",X"3A",X"C9",X"E4",X"C6",X"06",X"FE",X"65",X"DA",X"D0",X"0B",X"3E",X"64",
		X"32",X"C9",X"E4",X"CD",X"6F",X"17",X"21",X"CA",X"E4",X"34",X"C9",X"CD",X"EB",X"0B",X"79",X"47",
		X"CB",X"20",X"CB",X"27",X"CB",X"27",X"80",X"32",X"98",X"E2",X"C9",X"0E",X"05",X"3A",X"CC",X"E4",
		X"A7",X"C2",X"00",X"0C",X"3A",X"C5",X"E2",X"A7",X"C2",X"FE",X"0B",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"C9",X"3A",X"A6",X"E2",X"A7",X"C0",X"CD",X"E8",X"10",X"3A",X"82",X"E2",X"CB",X"5F",X"CA",X"1B",
		X"0C",X"3E",X"08",X"CD",X"1B",X"0C",X"3A",X"82",X"E2",X"D6",X"08",X"16",X"00",X"5F",X"2A",X"80",
		X"E2",X"19",X"22",X"80",X"E2",X"CD",X"34",X"0C",X"2A",X"80",X"E2",X"7C",X"32",X"00",X"A0",X"7D",
		X"32",X"00",X"90",X"C9",X"CB",X"3D",X"CB",X"3D",X"CB",X"85",X"4D",X"06",X"00",X"A7",X"CB",X"0C",
		X"38",X"08",X"21",X"BE",X"8B",X"09",X"CB",X"FD",X"18",X"0B",X"21",X"FE",X"8B",X"3E",X"80",X"91",
		X"CB",X"BF",X"4F",X"ED",X"42",X"CD",X"6B",X"0D",X"EB",X"A7",X"2A",X"94",X"E2",X"3A",X"80",X"E2",
		X"D6",X"08",X"E6",X"F8",X"CB",X"BF",X"06",X"00",X"4F",X"09",X"09",X"09",X"D5",X"D9",X"CD",X"34",
		X"0D",X"D9",X"CD",X"83",X"0C",X"01",X"18",X"00",X"CF",X"D1",X"13",X"21",X"E8",X"E4",X"01",X"18",
		X"00",X"CF",X"C9",X"D5",X"C5",X"3A",X"B8",X"E2",X"A7",X"CA",X"94",X"0C",X"11",X"D0",X"E4",X"01",
		X"18",X"00",X"ED",X"B0",X"21",X"D0",X"E4",X"C1",X"D1",X"FD",X"21",X"C3",X"E4",X"FD",X"7E",X"00",
		X"A7",X"C8",X"FD",X"7E",X"01",X"A7",X"CC",X"AF",X"0C",X"E5",X"CD",X"BE",X"0C",X"E1",X"C9",X"79",
		X"FD",X"BE",X"02",X"CA",X"B8",X"0C",X"F1",X"C9",X"3E",X"01",X"FD",X"77",X"01",X"C9",X"D5",X"E5",
		X"21",X"24",X"0D",X"C5",X"FD",X"4E",X"00",X"0D",X"CB",X"21",X"06",X"00",X"09",X"5E",X"23",X"56",
		X"FD",X"6E",X"01",X"FD",X"34",X"01",X"C1",X"3A",X"B8",X"E2",X"A7",X"C2",X"E5",X"0C",X"FD",X"35",
		X"01",X"2D",X"CA",X"EC",X"0C",X"2D",X"CB",X"25",X"CB",X"25",X"CB",X"25",X"26",X"00",X"19",X"EB",
		X"E1",X"FD",X"7E",X"03",X"C5",X"4F",X"06",X"00",X"09",X"C5",X"EB",X"01",X"04",X"00",X"ED",X"B0",
		X"C1",X"EB",X"21",X"E8",X"E4",X"09",X"EB",X"01",X"04",X"00",X"ED",X"B0",X"FD",X"7E",X"01",X"FE",
		X"05",X"DA",X"21",X"0D",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",
		X"03",X"C1",X"D1",X"C9",X"B7",X"30",X"D7",X"30",X"F7",X"30",X"17",X"31",X"37",X"31",X"57",X"31",
		X"4D",X"4D",X"4D",X"4C",X"3A",X"B8",X"E2",X"A7",X"C8",X"2A",X"A4",X"E2",X"11",X"E8",X"E4",X"3A",
		X"CC",X"E4",X"4F",X"3A",X"CF",X"E4",X"81",X"4F",X"CA",X"59",X"0D",X"06",X"18",X"C5",X"7E",X"E6",
		X"F0",X"81",X"12",X"23",X"13",X"C1",X"10",X"F5",X"C9",X"01",X"18",X"00",X"ED",X"B0",X"3A",X"C7",
		X"E4",X"A7",X"C8",X"FE",X"07",X"D0",X"1B",X"1B",X"1B",X"12",X"C9",X"AF",X"32",X"B8",X"E2",X"3A",
		X"74",X"E0",X"47",X"7D",X"B8",X"C8",X"3E",X"01",X"32",X"B8",X"E2",X"7D",X"32",X"74",X"E0",X"E6",
		X"1F",X"C0",X"CD",X"1F",X"10",X"CA",X"AD",X"0D",X"E5",X"2A",X"66",X"E0",X"23",X"22",X"66",X"E0",
		X"CD",X"F1",X"0D",X"CD",X"54",X"0E",X"CD",X"D2",X"0D",X"CD",X"E7",X"0E",X"CD",X"DC",X"24",X"CD",
		X"31",X"10",X"CD",X"86",X"24",X"CD",X"07",X"2B",X"CD",X"D6",X"0E",X"E1",X"C9",X"E5",X"2A",X"64",
		X"E0",X"23",X"22",X"64",X"E0",X"CD",X"F1",X"0D",X"CD",X"5A",X"0E",X"CD",X"D8",X"0D",X"CD",X"E7",
		X"0E",X"CD",X"DC",X"24",X"CD",X"31",X"10",X"CD",X"8E",X"24",X"CD",X"FA",X"2A",X"CD",X"D0",X"0E",
		X"E1",X"C9",X"3A",X"66",X"E0",X"C3",X"DB",X"0D",X"3A",X"64",X"E0",X"47",X"3A",X"8E",X"E2",X"4F",
		X"A7",X"CA",X"EA",X"0D",X"CB",X"27",X"CB",X"27",X"3D",X"4F",X"78",X"A1",X"B9",X"CC",X"3C",X"17",
		X"C9",X"E5",X"EB",X"21",X"A8",X"0E",X"06",X"12",X"7E",X"23",X"BB",X"C2",X"03",X"0E",X"7E",X"BA",
		X"CA",X"0D",X"0E",X"23",X"10",X"F2",X"AF",X"32",X"C7",X"E4",X"C3",X"1E",X"0E",X"78",X"ED",X"44",
		X"C6",X"13",X"FE",X"07",X"DA",X"1B",X"0E",X"D6",X"06",X"18",X"F7",X"32",X"C7",X"E4",X"21",X"CC",
		X"0E",X"06",X"02",X"7E",X"23",X"BB",X"C2",X"2E",X"0E",X"7E",X"BA",X"CA",X"34",X"0E",X"23",X"10",
		X"F2",X"C3",X"52",X"0E",X"CD",X"1F",X"10",X"CA",X"40",X"0E",X"21",X"85",X"E0",X"C3",X"43",X"0E",
		X"21",X"84",X"E0",X"78",X"ED",X"44",X"C6",X"03",X"BE",X"CA",X"52",X"0E",X"77",X"3E",X"02",X"32",
		X"63",X"E0",X"E1",X"C9",X"ED",X"5B",X"66",X"E0",X"18",X"04",X"ED",X"5B",X"64",X"E0",X"21",X"A2",
		X"0E",X"06",X"03",X"C5",X"D5",X"4E",X"23",X"46",X"E5",X"EB",X"A7",X"ED",X"42",X"38",X"09",X"7C",
		X"A7",X"20",X"05",X"7D",X"FE",X"11",X"38",X"0B",X"E1",X"D1",X"C1",X"23",X"10",X"E5",X"AF",X"32",
		X"CF",X"E2",X"C9",X"E1",X"D1",X"C1",X"78",X"ED",X"44",X"C6",X"04",X"47",X"CD",X"1F",X"10",X"28",
		X"05",X"3A",X"83",X"E0",X"18",X"03",X"3A",X"82",X"E0",X"B8",X"3E",X"01",X"20",X"E1",X"3C",X"C3",
		X"7F",X"0E",X"B5",X"01",X"29",X"04",X"1F",X"06",X"BF",X"01",X"C0",X"01",X"C1",X"01",X"C2",X"01",
		X"C3",X"01",X"C4",X"01",X"33",X"04",X"34",X"04",X"35",X"04",X"36",X"04",X"37",X"04",X"38",X"04",
		X"29",X"06",X"2A",X"06",X"2B",X"06",X"2C",X"06",X"2D",X"06",X"2E",X"06",X"16",X"04",X"14",X"06",
		X"3A",X"64",X"E0",X"C3",X"D9",X"0E",X"3A",X"66",X"E0",X"E6",X"03",X"C0",X"06",X"02",X"CD",X"FA",
		X"06",X"3E",X"01",X"32",X"C1",X"E5",X"C9",X"FD",X"21",X"C3",X"E4",X"3A",X"CE",X"E2",X"47",X"3A",
		X"B9",X"E2",X"80",X"20",X"2F",X"3A",X"CD",X"E4",X"A7",X"20",X"41",X"3A",X"BA",X"E2",X"A7",X"20",
		X"42",X"3A",X"CF",X"E2",X"A7",X"20",X"0A",X"AF",X"21",X"C3",X"E4",X"06",X"04",X"CD",X"E9",X"1E",
		X"C9",X"FD",X"21",X"C3",X"E4",X"06",X"06",X"80",X"FD",X"77",X"00",X"FD",X"36",X"02",X"20",X"FD",
		X"36",X"03",X"0B",X"C9",X"0E",X"02",X"CD",X"EB",X"1F",X"E6",X"07",X"CA",X"37",X"0F",X"E6",X"01",
		X"81",X"FD",X"77",X"00",X"C3",X"53",X"0F",X"3E",X"05",X"C3",X"31",X"0F",X"FD",X"36",X"00",X"01",
		X"C3",X"47",X"0F",X"FD",X"36",X"00",X"04",X"CD",X"EB",X"1F",X"E6",X"07",X"C2",X"53",X"0F",X"FD",
		X"36",X"00",X"06",X"FD",X"21",X"C3",X"E4",X"CD",X"5B",X"0F",X"C9",X"CD",X"1F",X"10",X"CA",X"67",
		X"0F",X"3A",X"8A",X"E2",X"C3",X"6A",X"0F",X"3A",X"89",X"E2",X"FE",X"05",X"38",X"02",X"18",X"07",
		X"A7",X"28",X"0C",X"FE",X"02",X"38",X"04",X"0E",X"07",X"18",X"06",X"0E",X"06",X"18",X"02",X"0E",
		X"03",X"CD",X"EB",X"1F",X"E6",X"07",X"B9",X"D2",X"81",X"0F",X"4F",X"FD",X"7E",X"00",X"C3",X"A5",
		X"0F",X"79",X"21",X"B7",X"0F",X"CB",X"27",X"4F",X"06",X"00",X"09",X"7E",X"FD",X"77",X"03",X"23",
		X"7E",X"FD",X"77",X"02",X"C9",X"3A",X"B9",X"E2",X"A7",X"CA",X"91",X"0F",X"79",X"FE",X"06",X"D2",
		X"91",X"0F",X"AF",X"FD",X"77",X"00",X"C9",X"14",X"08",X"00",X"60",X"02",X"38",X"11",X"40",X"04",
		X"10",X"0E",X"00",X"0B",X"58",X"08",X"20",X"4F",X"A7",X"C2",X"D2",X"0F",X"21",X"2D",X"4E",X"3E",
		X"32",X"C9",X"E6",X"F0",X"FE",X"10",X"C2",X"EB",X"0F",X"79",X"E6",X"0F",X"C2",X"E5",X"0F",X"21",
		X"76",X"4E",X"3E",X"72",X"C9",X"21",X"1F",X"4F",X"3E",X"7E",X"C9",X"FE",X"20",X"C2",X"19",X"10",
		X"79",X"E6",X"0F",X"A7",X"C2",X"FD",X"0F",X"21",X"DA",X"4F",X"3E",X"C2",X"C9",X"FE",X"01",X"C2",
		X"08",X"10",X"21",X"FB",X"50",X"3E",X"A4",X"C9",X"FE",X"02",X"C2",X"13",X"10",X"21",X"DA",X"4F",
		X"3E",X"C2",X"C9",X"21",X"EF",X"51",X"3E",X"86",X"C9",X"21",X"B6",X"52",X"3E",X"98",X"C9",X"3A",
		X"6A",X"E0",X"CB",X"47",X"CA",X"2F",X"10",X"CB",X"7F",X"CA",X"2F",X"10",X"3E",X"01",X"C9",X"AF",
		X"C9",X"CD",X"1F",X"10",X"28",X"11",X"ED",X"5B",X"77",X"E0",X"ED",X"4B",X"66",X"E0",X"C5",X"3A",
		X"6F",X"E0",X"CD",X"C7",X"0F",X"18",X"0F",X"ED",X"5B",X"75",X"E0",X"ED",X"4B",X"64",X"E0",X"C5",
		X"3A",X"6E",X"E0",X"CD",X"C7",X"0F",X"08",X"C1",X"79",X"A7",X"C2",X"69",X"10",X"CB",X"40",X"C2",
		X"69",X"10",X"16",X"00",X"1E",X"00",X"C3",X"7E",X"10",X"CD",X"1F",X"10",X"CA",X"75",X"10",X"3A",
		X"7A",X"E0",X"C3",X"78",X"10",X"3A",X"79",X"E0",X"A7",X"C2",X"84",X"10",X"13",X"13",X"CD",X"A6",
		X"10",X"C3",X"BE",X"10",X"19",X"5E",X"23",X"56",X"EB",X"22",X"94",X"E2",X"11",X"18",X"00",X"A7",
		X"ED",X"52",X"22",X"A4",X"E2",X"CD",X"1F",X"10",X"CA",X"A1",X"10",X"21",X"7A",X"E0",X"C3",X"A4",
		X"10",X"21",X"79",X"E0",X"35",X"C9",X"CD",X"1F",X"10",X"CA",X"B5",X"10",X"ED",X"53",X"77",X"E0",
		X"AF",X"32",X"81",X"E0",X"C9",X"ED",X"53",X"75",X"E0",X"AF",X"32",X"80",X"E0",X"C9",X"E5",X"C5",
		X"D5",X"08",X"4F",X"06",X"00",X"09",X"CB",X"3B",X"CB",X"3A",X"D2",X"CF",X"10",X"CB",X"FB",X"19",
		X"CD",X"1F",X"10",X"CA",X"DD",X"10",X"7E",X"32",X"7A",X"E0",X"C3",X"E1",X"10",X"7E",X"32",X"79",
		X"E0",X"D1",X"C1",X"E1",X"19",X"C3",X"85",X"10",X"3A",X"BF",X"E2",X"FE",X"02",X"D2",X"04",X"12",
		X"A7",X"C2",X"FB",X"10",X"3A",X"B0",X"E2",X"A7",X"CA",X"FF",X"10",X"AF",X"C3",X"92",X"11",X"3A",
		X"CC",X"E4",X"47",X"3A",X"CD",X"E4",X"B0",X"CA",X"1A",X"11",X"3A",X"96",X"E2",X"A7",X"C2",X"1A",
		X"11",X"3A",X"83",X"E2",X"E6",X"3F",X"C0",X"C3",X"20",X"11",X"3A",X"83",X"E2",X"E6",X"0F",X"C0",
		X"3A",X"96",X"E2",X"A7",X"C2",X"F8",X"11",X"3A",X"C9",X"E4",X"A7",X"CA",X"F8",X"11",X"3A",X"82",
		X"E2",X"A7",X"C2",X"36",X"11",X"3C",X"47",X"3A",X"AC",X"E2",X"FE",X"03",X"D2",X"D3",X"11",X"CD",
		X"1F",X"10",X"CA",X"6E",X"11",X"3A",X"87",X"E0",X"2F",X"E6",X"0C",X"CB",X"5F",X"C2",X"BA",X"11",
		X"CB",X"57",X"C2",X"D3",X"11",X"3A",X"8C",X"E2",X"A7",X"CA",X"6A",X"11",X"78",X"D6",X"02",X"DA",
		X"67",X"11",X"FE",X"02",X"D2",X"69",X"11",X"3E",X"02",X"47",X"78",X"C3",X"92",X"11",X"3A",X"87",
		X"E0",X"2F",X"E6",X"A0",X"CB",X"6F",X"20",X"42",X"CB",X"7F",X"20",X"57",X"3A",X"8C",X"E2",X"A7",
		X"CA",X"91",X"11",X"78",X"D6",X"02",X"DA",X"8E",X"11",X"FE",X"02",X"D2",X"90",X"11",X"3E",X"02",
		X"47",X"78",X"32",X"82",X"E2",X"F5",X"CB",X"3F",X"CB",X"3F",X"E6",X"03",X"32",X"8E",X"E2",X"3A",
		X"07",X"E0",X"A7",X"C2",X"AB",X"11",X"06",X"13",X"C3",X"AD",X"11",X"06",X"0C",X"F1",X"CD",X"0E",
		X"20",X"3A",X"87",X"E2",X"CB",X"87",X"32",X"93",X"E2",X"C9",X"78",X"3C",X"CD",X"2A",X"12",X"D2",
		X"CF",X"11",X"F5",X"3A",X"83",X"E2",X"E6",X"3F",X"CC",X"3C",X"17",X"F1",X"C3",X"92",X"11",X"79",
		X"C3",X"92",X"11",X"78",X"CB",X"87",X"A7",X"CA",X"F3",X"11",X"FE",X"02",X"DA",X"F3",X"11",X"D6",
		X"02",X"FE",X"02",X"DA",X"F3",X"11",X"FE",X"0D",X"D2",X"F3",X"11",X"F5",X"3E",X"17",X"D7",X"F1",
		X"C3",X"92",X"11",X"3E",X"02",X"C3",X"92",X"11",X"3A",X"82",X"E2",X"D6",X"01",X"D2",X"92",X"11",
		X"AF",X"32",X"8C",X"E2",X"3A",X"C9",X"E4",X"A7",X"CA",X"1D",X"12",X"3A",X"CA",X"E2",X"FE",X"30",
		X"DA",X"16",X"12",X"32",X"6B",X"E0",X"CD",X"6F",X"17",X"AF",X"C3",X"92",X"11",X"21",X"A6",X"E2",
		X"7E",X"A7",X"C2",X"16",X"12",X"34",X"AF",X"C3",X"92",X"11",X"F5",X"0E",X"0C",X"3A",X"97",X"E2",
		X"A7",X"C2",X"3E",X"12",X"3A",X"C5",X"E2",X"A7",X"C2",X"42",X"12",X"C3",X"44",X"12",X"0D",X"0D",
		X"0D",X"0D",X"0D",X"0D",X"F1",X"B9",X"C9",X"DD",X"21",X"C0",X"E1",X"26",X"04",X"3A",X"96",X"E2",
		X"A7",X"C2",X"F6",X"12",X"3A",X"83",X"E2",X"0F",X"D8",X"CD",X"15",X"13",X"3A",X"AC",X"E2",X"FE",
		X"03",X"DA",X"6B",X"12",X"3A",X"AD",X"E2",X"0F",X"DA",X"C5",X"12",X"CD",X"1F",X"10",X"CA",X"98",
		X"12",X"3A",X"87",X"E0",X"2F",X"E6",X"0C",X"CB",X"5F",X"C2",X"D2",X"12",X"CB",X"57",X"C2",X"F4",
		X"12",X"3A",X"8C",X"E2",X"21",X"11",X"E0",X"CB",X"5E",X"CA",X"BF",X"12",X"3A",X"82",X"E2",X"CB",
		X"3F",X"3C",X"32",X"8C",X"E2",X"CB",X"9E",X"C9",X"3A",X"87",X"E0",X"2F",X"E6",X"A0",X"CB",X"6F",
		X"C2",X"CA",X"12",X"CB",X"7F",X"C2",X"F4",X"12",X"3A",X"8C",X"E2",X"21",X"11",X"E0",X"CB",X"6E",
		X"CA",X"BF",X"12",X"3A",X"82",X"E2",X"CB",X"3F",X"3C",X"32",X"8C",X"E2",X"CB",X"AE",X"C9",X"A7",
		X"C8",X"21",X"8C",X"E2",X"35",X"26",X"01",X"C3",X"F6",X"12",X"21",X"11",X"E0",X"CB",X"EE",X"C3",
		X"D7",X"12",X"21",X"11",X"E0",X"CB",X"DE",X"06",X"04",X"11",X"04",X"00",X"DD",X"7E",X"03",X"3C",
		X"4F",X"78",X"FE",X"04",X"C2",X"EB",X"12",X"79",X"FE",X"60",X"D0",X"79",X"CD",X"BC",X"1E",X"DD",
		X"19",X"10",X"E9",X"C9",X"26",X"02",X"06",X"04",X"11",X"04",X"00",X"DD",X"7E",X"03",X"CB",X"87",
		X"94",X"4F",X"78",X"FE",X"04",X"C2",X"0C",X"13",X"79",X"FE",X"30",X"D8",X"79",X"CD",X"BC",X"1E",
		X"DD",X"19",X"10",X"E7",X"C9",X"DD",X"E5",X"3A",X"B0",X"E2",X"A7",X"C2",X"45",X"13",X"3A",X"83",
		X"E2",X"CB",X"3F",X"E6",X"01",X"4F",X"3A",X"8E",X"E2",X"A7",X"CA",X"3E",X"13",X"FE",X"01",X"CA",
		X"4A",X"13",X"3E",X"01",X"CB",X"41",X"CA",X"53",X"13",X"3E",X"20",X"C3",X"53",X"13",X"3E",X"0C",
		X"CB",X"41",X"CA",X"53",X"13",X"3E",X"0E",X"C3",X"53",X"13",X"3E",X"10",X"CB",X"41",X"CA",X"53",
		X"13",X"3E",X"12",X"CD",X"B2",X"1E",X"11",X"04",X"00",X"DD",X"19",X"3C",X"CD",X"B2",X"1E",X"DD",
		X"19",X"AF",X"CD",X"B2",X"1E",X"DD",X"19",X"CD",X"B2",X"1E",X"DD",X"E1",X"C9",X"3A",X"82",X"E2",
		X"A7",X"C8",X"DD",X"21",X"C0",X"E1",X"3A",X"99",X"E2",X"D6",X"01",X"32",X"99",X"E2",X"D2",X"23",
		X"14",X"AF",X"32",X"99",X"E2",X"3A",X"9A",X"E2",X"D6",X"01",X"32",X"9A",X"E2",X"D2",X"70",X"14",
		X"AF",X"32",X"9A",X"E2",X"CD",X"1F",X"10",X"CA",X"AD",X"13",X"3A",X"88",X"E0",X"2F",X"E6",X"0C",
		X"CB",X"5F",X"C2",X"DA",X"13",X"CB",X"57",X"C2",X"04",X"14",X"C3",X"BD",X"13",X"3A",X"87",X"E0",
		X"2F",X"E6",X"03",X"CB",X"47",X"C2",X"C5",X"13",X"CB",X"4F",X"C2",X"EF",X"13",X"AF",X"32",X"91",
		X"E2",X"32",X"92",X"E2",X"C9",X"3A",X"11",X"E0",X"CB",X"47",X"C2",X"1E",X"14",X"CD",X"DB",X"0B",
		X"32",X"99",X"E2",X"AF",X"32",X"9A",X"E2",X"C3",X"23",X"14",X"3A",X"12",X"E0",X"CB",X"5F",X"C2",
		X"1E",X"14",X"CD",X"DB",X"0B",X"32",X"99",X"E2",X"AF",X"32",X"9A",X"E2",X"C3",X"23",X"14",X"3A",
		X"11",X"E0",X"CB",X"4F",X"C2",X"19",X"14",X"CD",X"DB",X"0B",X"32",X"9A",X"E2",X"AF",X"32",X"99",
		X"E2",X"C3",X"70",X"14",X"3A",X"12",X"E0",X"CB",X"57",X"C2",X"19",X"14",X"CD",X"DB",X"0B",X"32",
		X"9A",X"E2",X"AF",X"32",X"99",X"E2",X"C3",X"70",X"14",X"AF",X"32",X"9A",X"E2",X"C9",X"AF",X"32",
		X"99",X"E2",X"C9",X"DD",X"7E",X"00",X"FE",X"F8",X"D2",X"BF",X"14",X"06",X"04",X"11",X"04",X"00",
		X"3A",X"82",X"E2",X"ED",X"44",X"E6",X"0F",X"CB",X"3F",X"CB",X"3F",X"FE",X"03",X"DA",X"42",X"14",
		X"3E",X"02",X"DD",X"86",X"00",X"CD",X"9E",X"1E",X"DD",X"19",X"10",X"E4",X"3A",X"AC",X"E2",X"A7",
		X"C0",X"D5",X"11",X"F4",X"FF",X"DD",X"19",X"DD",X"7E",X"00",X"C6",X"10",X"D1",X"DD",X"19",X"CD",
		X"9E",X"1E",X"DD",X"19",X"CD",X"9E",X"1E",X"21",X"91",X"E2",X"34",X"AF",X"32",X"92",X"E2",X"C9",
		X"DD",X"7E",X"00",X"FE",X"39",X"DA",X"BF",X"14",X"06",X"04",X"11",X"04",X"00",X"3A",X"82",X"E2",
		X"ED",X"44",X"E6",X"0F",X"CB",X"3F",X"CB",X"3F",X"FE",X"03",X"DA",X"8F",X"14",X"3E",X"02",X"ED",
		X"44",X"DD",X"86",X"00",X"CD",X"9E",X"1E",X"DD",X"19",X"10",X"E2",X"3A",X"AC",X"E2",X"A7",X"C0",
		X"D5",X"11",X"F4",X"FF",X"DD",X"19",X"DD",X"7E",X"00",X"D6",X"10",X"D1",X"DD",X"19",X"CD",X"9E",
		X"1E",X"DD",X"19",X"CD",X"9E",X"1E",X"21",X"92",X"E2",X"34",X"AF",X"32",X"91",X"E2",X"C9",X"AF",
		X"32",X"A7",X"E5",X"3C",X"32",X"96",X"E2",X"C9",X"3A",X"83",X"E2",X"0F",X"D8",X"DD",X"21",X"C0",
		X"E1",X"3A",X"AC",X"E2",X"A7",X"C8",X"0F",X"38",X"05",X"CD",X"70",X"14",X"18",X"03",X"CD",X"23",
		X"14",X"3A",X"AD",X"E2",X"D6",X"01",X"38",X"04",X"32",X"AD",X"E2",X"C9",X"AF",X"32",X"AC",X"E2",
		X"32",X"AD",X"E2",X"C9",X"3A",X"83",X"E2",X"0F",X"D8",X"3A",X"AC",X"E2",X"A7",X"C0",X"CD",X"1F",
		X"10",X"CA",X"0B",X"15",X"CD",X"12",X"15",X"CD",X"64",X"15",X"C9",X"CD",X"B6",X"15",X"CD",X"08",
		X"16",X"C9",X"3A",X"92",X"E2",X"57",X"3A",X"99",X"E2",X"A7",X"20",X"0A",X"3A",X"88",X"E0",X"2F",
		X"E6",X"0C",X"CB",X"5F",X"28",X"1B",X"3A",X"91",X"E2",X"FE",X"02",X"D8",X"7A",X"A7",X"C0",X"21",
		X"8F",X"E2",X"34",X"7E",X"FE",X"06",X"38",X"03",X"3E",X"06",X"77",X"0E",X"00",X"CD",X"5A",X"16",
		X"C9",X"21",X"8F",X"E2",X"7E",X"A7",X"28",X"0C",X"0E",X"00",X"CD",X"5A",X"16",X"35",X"21",X"12",
		X"E0",X"CB",X"D6",X"C9",X"21",X"12",X"E0",X"CB",X"96",X"AF",X"32",X"8F",X"E2",X"32",X"91",X"E2",
		X"32",X"99",X"E2",X"C9",X"3A",X"91",X"E2",X"57",X"3A",X"9A",X"E2",X"A7",X"20",X"0A",X"3A",X"88",
		X"E0",X"2F",X"E6",X"0C",X"CB",X"57",X"28",X"1B",X"3A",X"92",X"E2",X"FE",X"02",X"D8",X"7A",X"A7",
		X"C0",X"21",X"90",X"E2",X"34",X"7E",X"FE",X"06",X"38",X"03",X"3E",X"06",X"77",X"0E",X"01",X"CD",
		X"5A",X"16",X"C9",X"21",X"90",X"E2",X"7E",X"A7",X"28",X"0C",X"0E",X"01",X"CD",X"5A",X"16",X"35",
		X"21",X"12",X"E0",X"CB",X"DE",X"C9",X"21",X"12",X"E0",X"CB",X"9E",X"AF",X"32",X"90",X"E2",X"32",
		X"92",X"E2",X"32",X"9A",X"E2",X"C9",X"3A",X"92",X"E2",X"57",X"3A",X"99",X"E2",X"A7",X"20",X"0A",
		X"3A",X"87",X"E0",X"2F",X"E6",X"03",X"CB",X"47",X"28",X"1B",X"3A",X"91",X"E2",X"FE",X"02",X"D8",
		X"7A",X"A7",X"C0",X"21",X"8F",X"E2",X"34",X"7E",X"FE",X"06",X"38",X"03",X"3E",X"06",X"77",X"0E",
		X"00",X"CD",X"5A",X"16",X"C9",X"21",X"8F",X"E2",X"7E",X"A7",X"28",X"0C",X"0E",X"00",X"CD",X"5A",
		X"16",X"35",X"21",X"11",X"E0",X"CB",X"CE",X"C9",X"21",X"11",X"E0",X"CB",X"8E",X"AF",X"32",X"8F",
		X"E2",X"32",X"91",X"E2",X"32",X"99",X"E2",X"C9",X"3A",X"91",X"E2",X"57",X"3A",X"9A",X"E2",X"A7",
		X"20",X"0A",X"3A",X"87",X"E0",X"2F",X"E6",X"03",X"CB",X"4F",X"28",X"1B",X"3A",X"92",X"E2",X"FE",
		X"02",X"D8",X"7A",X"A7",X"C0",X"21",X"90",X"E2",X"34",X"7E",X"FE",X"06",X"38",X"03",X"3E",X"06",
		X"77",X"0E",X"01",X"CD",X"5A",X"16",X"C9",X"21",X"90",X"E2",X"7E",X"A7",X"28",X"0C",X"0E",X"01",
		X"CD",X"5A",X"16",X"35",X"21",X"11",X"E0",X"CB",X"C6",X"C9",X"21",X"11",X"E0",X"CB",X"86",X"AF",
		X"32",X"90",X"E2",X"32",X"92",X"E2",X"32",X"9A",X"E2",X"C9",X"DD",X"21",X"C0",X"E1",X"E5",X"C5",
		X"3D",X"CB",X"27",X"CB",X"27",X"4F",X"06",X"00",X"3A",X"8E",X"E2",X"A7",X"CA",X"80",X"16",X"FE",
		X"01",X"CA",X"7A",X"16",X"21",X"DA",X"16",X"C3",X"83",X"16",X"21",X"C2",X"16",X"C3",X"83",X"16",
		X"21",X"AA",X"16",X"09",X"C1",X"06",X"04",X"11",X"04",X"00",X"7E",X"CD",X"B2",X"1E",X"79",X"A7",
		X"CA",X"98",X"16",X"3E",X"40",X"C3",X"9A",X"16",X"3E",X"C0",X"CD",X"A8",X"1E",X"23",X"DD",X"19",
		X"10",X"E8",X"E1",X"7E",X"FE",X"06",X"D8",X"35",X"35",X"C9",X"16",X"17",X"00",X"00",X"16",X"17",
		X"00",X"00",X"18",X"19",X"1A",X"1B",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"1C",X"1D",
		X"0B",X"1F",X"5A",X"5B",X"00",X"00",X"5A",X"5B",X"00",X"00",X"5C",X"5D",X"00",X"00",X"5C",X"5D",
		X"00",X"00",X"5E",X"5F",X"60",X"61",X"62",X"5F",X"63",X"61",X"03",X"04",X"00",X"00",X"03",X"04",
		X"00",X"00",X"05",X"06",X"00",X"00",X"05",X"06",X"00",X"00",X"07",X"08",X"00",X"00",X"09",X"0A",
		X"00",X"00",X"06",X"03",X"D9",X"06",X"00",X"D9",X"D9",X"CD",X"B6",X"1A",X"11",X"80",X"00",X"FD",
		X"19",X"D9",X"10",X"F4",X"C9",X"21",X"38",X"17",X"11",X"06",X"8F",X"01",X"04",X"00",X"CF",X"11",
		X"07",X"8F",X"06",X"04",X"3E",X"07",X"CD",X"D3",X"1E",X"11",X"05",X"8E",X"06",X"03",X"3E",X"01",
		X"CD",X"D3",X"1E",X"3A",X"CA",X"E4",X"A7",X"CA",X"32",X"17",X"FD",X"21",X"04",X"8D",X"CD",X"F2",
		X"16",X"C9",X"3E",X"09",X"32",X"04",X"8D",X"C9",X"42",X"55",X"4D",X"50",X"3A",X"A7",X"E2",X"A7",
		X"C0",X"21",X"87",X"17",X"11",X"12",X"8F",X"01",X"04",X"00",X"CF",X"11",X"13",X"8F",X"06",X"04",
		X"3E",X"07",X"CD",X"D3",X"1E",X"3E",X"25",X"32",X"10",X"8C",X"3A",X"63",X"E0",X"A7",X"CA",X"6F",
		X"17",X"3A",X"C9",X"E4",X"A7",X"CA",X"7D",X"17",X"3D",X"CA",X"7D",X"17",X"32",X"C9",X"E4",X"CD",
		X"8B",X"17",X"3A",X"C9",X"E4",X"FD",X"21",X"10",X"8D",X"CD",X"F2",X"16",X"C9",X"3E",X"09",X"32",
		X"10",X"8D",X"AF",X"32",X"C9",X"E4",X"C9",X"46",X"55",X"45",X"4C",X"3A",X"C9",X"E4",X"FE",X"14",
		X"DA",X"9E",X"17",X"FE",X"64",X"D2",X"A5",X"17",X"06",X"01",X"AF",X"C3",X"A8",X"17",X"06",X"08",
		X"3E",X"01",X"C3",X"A8",X"17",X"06",X"07",X"AF",X"32",X"C4",X"E2",X"78",X"11",X"11",X"8E",X"06",
		X"03",X"CD",X"D3",X"1E",X"C9",X"3A",X"A6",X"E2",X"A7",X"C0",X"3A",X"C4",X"E2",X"47",X"3A",X"CB",
		X"E2",X"80",X"C8",X"3A",X"83",X"E2",X"E6",X"3F",X"C0",X"3E",X"14",X"D7",X"C9",X"DD",X"21",X"C4",
		X"E1",X"3A",X"A7",X"E5",X"A7",X"C8",X"FE",X"01",X"C2",X"FF",X"17",X"3A",X"AA",X"E2",X"C6",X"08",
		X"47",X"DD",X"7E",X"00",X"C6",X"08",X"B8",X"38",X"04",X"06",X"01",X"18",X"02",X"06",X"02",X"3A",
		X"AB",X"E2",X"D6",X"10",X"4F",X"DD",X"7E",X"03",X"B9",X"30",X"02",X"CB",X"D0",X"78",X"C9",X"AF",
		X"32",X"AC",X"E2",X"C9",X"F5",X"3A",X"AC",X"E2",X"47",X"F1",X"B8",X"CA",X"3D",X"18",X"32",X"AC",
		X"E2",X"3E",X"19",X"D7",X"CD",X"1F",X"10",X"A7",X"CA",X"21",X"18",X"3A",X"8B",X"E0",X"C3",X"24",
		X"18",X"3A",X"8A",X"E0",X"06",X"0D",X"A7",X"20",X"02",X"06",X"08",X"3A",X"82",X"E2",X"80",X"47",
		X"3A",X"A7",X"E2",X"A7",X"CA",X"39",X"18",X"CB",X"38",X"78",X"32",X"AD",X"E2",X"AF",X"32",X"96",
		X"E2",X"32",X"A7",X"E5",X"C9",X"3A",X"96",X"E2",X"FE",X"20",X"D0",X"FE",X"15",X"D2",X"BC",X"18",
		X"FE",X"02",X"D2",X"76",X"18",X"CD",X"CD",X"17",X"A7",X"C2",X"04",X"18",X"3E",X"01",X"32",X"C6",
		X"E2",X"3E",X"1F",X"D7",X"3A",X"C0",X"E1",X"32",X"D0",X"E1",X"3A",X"C3",X"E1",X"32",X"D3",X"E1",
		X"CD",X"D8",X"18",X"C3",X"B7",X"18",X"3A",X"83",X"E2",X"0F",X"D8",X"3A",X"96",X"E2",X"DD",X"21",
		X"D0",X"E1",X"21",X"8F",X"30",X"3D",X"CB",X"27",X"4F",X"06",X"00",X"09",X"46",X"3A",X"C0",X"E1",
		X"FE",X"A0",X"DA",X"99",X"18",X"78",X"ED",X"44",X"47",X"78",X"DD",X"86",X"00",X"FE",X"F0",X"D2",
		X"BC",X"18",X"FE",X"40",X"DA",X"BC",X"18",X"CD",X"9E",X"1E",X"3E",X"22",X"CD",X"B2",X"1E",X"23",
		X"7E",X"DD",X"86",X"03",X"CD",X"BC",X"1E",X"21",X"96",X"E2",X"34",X"C9",X"21",X"96",X"E2",X"34",
		X"7E",X"FE",X"20",X"D8",X"3A",X"7C",X"E0",X"A7",X"CA",X"D1",X"18",X"21",X"7B",X"E0",X"CB",X"FE",
		X"C9",X"3A",X"C0",X"E1",X"32",X"CB",X"E4",X"C9",X"3A",X"BF",X"E2",X"A7",X"C2",X"20",X"19",X"3A",
		X"82",X"E2",X"47",X"CB",X"27",X"CB",X"27",X"80",X"3C",X"32",X"9B",X"E2",X"AF",X"32",X"9C",X"E2",
		X"DD",X"21",X"C0",X"E1",X"DD",X"56",X"00",X"DD",X"5E",X"03",X"06",X"04",X"21",X"FF",X"2F",X"7E",
		X"82",X"CD",X"9E",X"1E",X"23",X"3E",X"41",X"CD",X"A8",X"1E",X"7E",X"CD",X"B2",X"1E",X"23",X"7E",
		X"83",X"CD",X"BC",X"1E",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"23",X"10",X"E0",X"C9",
		X"AF",X"06",X"04",X"11",X"04",X"00",X"DD",X"21",X"C0",X"E1",X"CD",X"B2",X"1E",X"DD",X"19",X"10",
		X"F9",X"C9",X"3A",X"82",X"E2",X"0E",X"02",X"FE",X"05",X"DA",X"44",X"19",X"FE",X"09",X"DA",X"45",
		X"19",X"C3",X"46",X"19",X"0D",X"0D",X"79",X"C9",X"3A",X"BF",X"E2",X"A7",X"C2",X"19",X"1A",X"3A",
		X"9B",X"E2",X"A7",X"C8",X"DD",X"21",X"C0",X"E1",X"3A",X"83",X"E2",X"47",X"CD",X"32",X"19",X"A7",
		X"CA",X"6B",X"19",X"FE",X"01",X"CA",X"74",X"19",X"C3",X"77",X"19",X"CB",X"40",X"C8",X"CB",X"48",
		X"C8",X"C3",X"77",X"19",X"CB",X"40",X"C8",X"21",X"FF",X"2F",X"11",X"0C",X"00",X"3A",X"9C",X"E2",
		X"A7",X"CA",X"88",X"19",X"47",X"19",X"10",X"FD",X"DD",X"7E",X"00",X"FE",X"E8",X"DA",X"98",X"19",
		X"D6",X"05",X"CD",X"9E",X"1E",X"C3",X"A2",X"19",X"FE",X"48",X"D2",X"A2",X"19",X"C6",X"05",X"CD",
		X"9E",X"1E",X"32",X"9E",X"E2",X"DD",X"7E",X"03",X"32",X"9F",X"E2",X"11",X"04",X"00",X"06",X"04",
		X"C5",X"3A",X"9C",X"E2",X"FE",X"06",X"D2",X"DC",X"19",X"7E",X"ED",X"44",X"47",X"3A",X"9E",X"E2",
		X"80",X"CD",X"9E",X"1E",X"3E",X"C0",X"CD",X"A8",X"1E",X"23",X"7E",X"CD",X"B2",X"1E",X"23",X"7E",
		X"47",X"3A",X"9F",X"E2",X"80",X"CD",X"BC",X"1E",X"23",X"C3",X"FB",X"19",X"7E",X"47",X"3A",X"9E",
		X"E2",X"80",X"CD",X"9E",X"1E",X"AF",X"CD",X"A8",X"1E",X"23",X"7E",X"CD",X"B2",X"1E",X"23",X"7E",
		X"ED",X"44",X"47",X"3A",X"9F",X"E2",X"80",X"CD",X"BC",X"1E",X"23",X"DD",X"19",X"C1",X"10",X"B0",
		X"21",X"9C",X"E2",X"34",X"7E",X"FE",X"0C",X"DA",X"0C",X"1A",X"AF",X"77",X"3A",X"9B",X"E2",X"D6",
		X"01",X"D2",X"15",X"1A",X"AF",X"32",X"9B",X"E2",X"C9",X"3A",X"96",X"E2",X"FE",X"08",X"D2",X"69",
		X"1A",X"3D",X"3D",X"4F",X"CB",X"27",X"81",X"4F",X"06",X"00",X"21",X"2F",X"1A",X"09",X"E9",X"C3",
		X"42",X"1A",X"C3",X"48",X"1A",X"C3",X"4E",X"1A",X"C3",X"48",X"1A",X"C3",X"4E",X"1A",X"C3",X"54",
		X"1A",X"C9",X"21",X"77",X"31",X"C3",X"57",X"1A",X"21",X"97",X"31",X"C3",X"57",X"1A",X"21",X"B7",
		X"31",X"C3",X"57",X"1A",X"21",X"D7",X"31",X"ED",X"5B",X"C0",X"E2",X"06",X"08",X"C5",X"D5",X"01",
		X"04",X"00",X"CF",X"D1",X"13",X"C1",X"10",X"F5",X"C9",X"FE",X"20",X"D8",X"3E",X"02",X"32",X"BF",
		X"E2",X"C9",X"21",X"E2",X"1A",X"11",X"0C",X"8F",X"01",X"05",X"00",X"CF",X"3E",X"07",X"11",X"0D",
		X"8F",X"06",X"05",X"CD",X"D3",X"1E",X"3E",X"01",X"11",X"0B",X"8E",X"06",X"03",X"CD",X"D3",X"1E",
		X"CD",X"EF",X"1A",X"3A",X"93",X"E2",X"A7",X"CA",X"DC",X"1A",X"47",X"3A",X"8B",X"E2",X"B8",X"CA",
		X"AB",X"1A",X"DA",X"AA",X"1A",X"3D",X"3D",X"C3",X"AB",X"1A",X"3C",X"32",X"8B",X"E2",X"FD",X"21",
		X"0A",X"8D",X"CD",X"F2",X"16",X"C9",X"FE",X"0A",X"DA",X"C1",X"1A",X"D6",X"0A",X"04",X"C3",X"B6",
		X"1A",X"4F",X"A7",X"C2",X"D2",X"1A",X"78",X"A7",X"C2",X"D0",X"1A",X"0E",X"F7",X"C3",X"D2",X"1A",
		X"0E",X"00",X"79",X"C6",X"09",X"FD",X"77",X"00",X"78",X"06",X"00",X"C9",X"3E",X"09",X"32",X"0A",
		X"8D",X"C9",X"53",X"50",X"45",X"45",X"44",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"21",
		X"0A",X"8C",X"11",X"8A",X"8C",X"3A",X"07",X"E0",X"A7",X"C2",X"02",X"1B",X"3E",X"02",X"77",X"3D",
		X"12",X"C9",X"3E",X"04",X"C3",X"FE",X"1A",X"DD",X"21",X"C0",X"E1",X"3A",X"96",X"E2",X"A7",X"C0",
		X"CD",X"7B",X"1F",X"D2",X"3B",X"1B",X"AF",X"32",X"A7",X"E5",X"3C",X"32",X"96",X"E2",X"3A",X"BA",
		X"E2",X"A7",X"C8",X"FD",X"7E",X"00",X"FE",X"D0",X"D8",X"FE",X"D4",X"D0",X"3E",X"01",X"32",X"BF",
		X"E2",X"11",X"FC",X"00",X"FD",X"19",X"FD",X"22",X"C0",X"E2",X"C9",X"CD",X"ED",X"1B",X"3A",X"CE",
		X"E4",X"A7",X"CA",X"7E",X"1B",X"4F",X"CD",X"1F",X"10",X"28",X"05",X"3A",X"83",X"E0",X"18",X"03",
		X"3A",X"82",X"E0",X"B9",X"28",X"28",X"3A",X"B0",X"E2",X"A7",X"20",X"22",X"FD",X"7E",X"00",X"FE",
		X"59",X"38",X"04",X"FE",X"5C",X"38",X"08",X"FE",X"6A",X"38",X"13",X"FE",X"6D",X"30",X"0F",X"FD",
		X"E5",X"E1",X"24",X"22",X"B6",X"E2",X"CD",X"09",X"1C",X"21",X"B0",X"E2",X"34",X"C9",X"FD",X"7E",
		X"01",X"FE",X"28",X"C0",X"FD",X"7E",X"00",X"FE",X"14",X"D8",X"FE",X"18",X"D0",X"06",X"64",X"CD",
		X"FA",X"06",X"3E",X"12",X"D7",X"3A",X"A7",X"E2",X"A7",X"C2",X"AB",X"1B",X"3A",X"C9",X"E4",X"C6",
		X"0A",X"FE",X"65",X"DA",X"A8",X"1B",X"3E",X"64",X"32",X"C9",X"E4",X"CD",X"B2",X"1B",X"CD",X"6F",
		X"17",X"C9",X"3A",X"CE",X"E2",X"A7",X"C2",X"C7",X"1B",X"3A",X"B9",X"E2",X"A7",X"C2",X"C7",X"1B",
		X"3E",X"04",X"0E",X"84",X"C3",X"CB",X"1B",X"3E",X"63",X"0E",X"01",X"FD",X"E5",X"E1",X"11",X"7E",
		X"00",X"19",X"EB",X"06",X"03",X"C5",X"F5",X"D5",X"06",X"03",X"CD",X"D3",X"1E",X"79",X"D1",X"13",
		X"D5",X"06",X"03",X"CD",X"D3",X"1E",X"D1",X"F1",X"13",X"C1",X"10",X"E9",X"C9",X"06",X"00",X"3A",
		X"C5",X"E2",X"A7",X"CA",X"04",X"1C",X"FD",X"7E",X"00",X"FE",X"60",X"DA",X"04",X"1C",X"FE",X"69",
		X"D2",X"04",X"1C",X"04",X"78",X"32",X"97",X"E2",X"C9",X"11",X"80",X"FF",X"FD",X"19",X"FD",X"7E",
		X"00",X"A7",X"C2",X"09",X"1C",X"FD",X"7E",X"01",X"32",X"B4",X"E2",X"C9",X"3A",X"B0",X"E2",X"A7",
		X"C8",X"21",X"33",X"1C",X"3A",X"B0",X"E2",X"3D",X"CB",X"27",X"4F",X"06",X"00",X"09",X"5E",X"23",
		X"56",X"EB",X"E9",X"54",X"1C",X"92",X"1C",X"AB",X"1C",X"AB",X"1C",X"AB",X"1C",X"AB",X"1C",X"AB",
		X"1C",X"AB",X"1C",X"AB",X"1C",X"AB",X"1C",X"AB",X"1C",X"AB",X"1C",X"C2",X"1C",X"F1",X"1C",X"21",
		X"B0",X"E2",X"34",X"C9",X"DD",X"21",X"C0",X"E1",X"3E",X"0E",X"CD",X"B2",X"1E",X"DD",X"21",X"C4",
		X"E1",X"3C",X"CD",X"B2",X"1E",X"AF",X"DD",X"21",X"C8",X"E1",X"CD",X"B2",X"1E",X"DD",X"21",X"CC",
		X"E1",X"CD",X"B2",X"1E",X"AF",X"32",X"82",X"E2",X"32",X"93",X"E2",X"21",X"CA",X"1D",X"3A",X"B4",
		X"E2",X"3D",X"CB",X"27",X"4F",X"06",X"00",X"09",X"5E",X"23",X"56",X"EB",X"22",X"B1",X"E2",X"C3",
		X"4F",X"1C",X"2A",X"B6",X"E2",X"E5",X"23",X"3E",X"E0",X"77",X"E1",X"3E",X"2B",X"77",X"11",X"80",
		X"00",X"19",X"06",X"08",X"AF",X"CD",X"E9",X"1E",X"C3",X"4F",X"1C",X"2A",X"B6",X"E2",X"11",X"80",
		X"00",X"3A",X"B0",X"E2",X"3D",X"47",X"19",X"10",X"FD",X"AF",X"06",X"08",X"CD",X"E9",X"1E",X"C3",
		X"4F",X"1C",X"CD",X"23",X"1D",X"2A",X"B1",X"E2",X"7D",X"A7",X"C2",X"D2",X"1C",X"7C",X"A7",X"CA",
		X"E8",X"1C",X"E5",X"06",X"0A",X"CD",X"FA",X"06",X"CD",X"80",X"1D",X"E1",X"2B",X"22",X"B1",X"E2",
		X"7D",X"E6",X"1F",X"C0",X"3E",X"15",X"D7",X"C9",X"21",X"00",X"00",X"22",X"B1",X"E2",X"C3",X"4F",
		X"1C",X"CD",X"1F",X"10",X"CA",X"FD",X"1C",X"21",X"83",X"E0",X"C3",X"00",X"1D",X"21",X"82",X"E0",
		X"3A",X"CE",X"E4",X"77",X"AF",X"32",X"CE",X"E4",X"32",X"B0",X"E2",X"32",X"B4",X"E2",X"32",X"93",
		X"E2",X"32",X"8B",X"E2",X"32",X"C7",X"E4",X"21",X"00",X"00",X"22",X"B1",X"E2",X"3E",X"01",X"32",
		X"82",X"E2",X"C9",X"2A",X"B6",X"E2",X"11",X"04",X"05",X"19",X"EB",X"21",X"5B",X"1D",X"01",X"07",
		X"00",X"CF",X"01",X"7F",X"FF",X"EB",X"09",X"3A",X"B4",X"E2",X"C6",X"30",X"77",X"3A",X"B4",X"E2",
		X"3D",X"4F",X"CB",X"27",X"CB",X"27",X"81",X"4F",X"06",X"00",X"2A",X"B6",X"E2",X"11",X"02",X"03",
		X"19",X"EB",X"21",X"62",X"1D",X"09",X"01",X"05",X"00",X"CF",X"C9",X"42",X"4F",X"4E",X"55",X"53",
		X"20",X"23",X"32",X"30",X"30",X"30",X"30",X"31",X"35",X"30",X"30",X"30",X"31",X"30",X"30",X"30",
		X"30",X"20",X"38",X"30",X"30",X"30",X"20",X"35",X"30",X"30",X"30",X"20",X"33",X"30",X"30",X"30",
		X"3A",X"B1",X"E2",X"0F",X"D0",X"21",X"C9",X"E4",X"34",X"7E",X"FE",X"65",X"38",X"06",X"CD",X"98",
		X"1D",X"3E",X"64",X"77",X"CD",X"6F",X"17",X"C9",X"E5",X"2A",X"B6",X"E2",X"11",X"8E",X"05",X"19",
		X"EB",X"D5",X"21",X"B9",X"1D",X"01",X"11",X"00",X"CF",X"D1",X"13",X"3E",X"08",X"06",X"11",X"CD",
		X"D3",X"1E",X"3E",X"01",X"32",X"A7",X"E2",X"E1",X"C9",X"46",X"55",X"45",X"4C",X"20",X"4F",X"56",
		X"45",X"52",X"20",X"43",X"48",X"41",X"52",X"47",X"45",X"21",X"C8",X"00",X"96",X"00",X"64",X"00",
		X"50",X"00",X"32",X"00",X"1E",X"00",X"2A",X"75",X"E0",X"ED",X"5B",X"64",X"E0",X"3A",X"79",X"E0",
		X"3C",X"47",X"3A",X"6E",X"E0",X"4F",X"CD",X"14",X"1E",X"22",X"75",X"E0",X"ED",X"53",X"64",X"E0",
		X"78",X"32",X"79",X"E0",X"C9",X"2A",X"77",X"E0",X"ED",X"5B",X"66",X"E0",X"3A",X"7A",X"E0",X"3C",
		X"47",X"3A",X"6F",X"E0",X"4F",X"CD",X"14",X"1E",X"22",X"77",X"E0",X"ED",X"53",X"66",X"E0",X"78",
		X"32",X"7A",X"E0",X"C9",X"78",X"C6",X"10",X"E5",X"F5",X"D5",X"EB",X"79",X"CD",X"C7",X"0F",X"C5",
		X"06",X"00",X"4F",X"09",X"C1",X"CB",X"3B",X"CB",X"3A",X"30",X"02",X"CB",X"FB",X"19",X"D1",X"7E",
		X"67",X"F1",X"BC",X"28",X"10",X"38",X"0E",X"94",X"E1",X"C5",X"01",X"02",X"00",X"A7",X"ED",X"42",
		X"C1",X"38",X"1D",X"18",X"D2",X"E1",X"47",X"CD",X"70",X"1E",X"C5",X"EB",X"01",X"F0",X"FF",X"09",
		X"C1",X"EB",X"7B",X"A7",X"20",X"04",X"CB",X"42",X"28",X"06",X"3E",X"04",X"32",X"7E",X"E0",X"C9",
		X"79",X"E6",X"F0",X"0F",X"0F",X"0F",X"57",X"1E",X"00",X"21",X"00",X"00",X"06",X"00",X"18",X"EA",
		X"7A",X"FE",X"04",X"28",X"16",X"FE",X"06",X"C0",X"7B",X"FE",X"14",X"D8",X"FE",X"25",X"D0",X"11",
		X"15",X"06",X"21",X"00",X"00",X"06",X"03",X"F1",X"C3",X"5A",X"1E",X"7B",X"FE",X"16",X"D8",X"FE",
		X"27",X"D0",X"11",X"17",X"04",X"21",X"0A",X"00",X"06",X"0B",X"F1",X"C3",X"5A",X"1E",X"DD",X"77",
		X"A0",X"DD",X"77",X"00",X"DD",X"77",X"60",X"C9",X"DD",X"77",X"A1",X"DD",X"77",X"01",X"DD",X"77",
		X"61",X"C9",X"DD",X"77",X"A2",X"DD",X"77",X"02",X"DD",X"77",X"62",X"C9",X"DD",X"77",X"A3",X"DD",
		X"77",X"03",X"DD",X"77",X"63",X"C9",X"ED",X"A0",X"E0",X"E5",X"21",X"7F",X"FF",X"EB",X"19",X"EB",
		X"E1",X"18",X"F3",X"E5",X"EB",X"11",X"80",X"FF",X"77",X"19",X"10",X"FC",X"E1",X"C9",X"C5",X"06",
		X"00",X"4F",X"10",X"FE",X"0D",X"20",X"FB",X"C1",X"C9",X"77",X"23",X"10",X"FC",X"C9",X"77",X"2C",
		X"20",X"FC",X"24",X"10",X"F9",X"C9",X"F3",X"76",X"3A",X"00",X"D0",X"2F",X"CB",X"5F",X"20",X"09",
		X"3A",X"10",X"E0",X"CB",X"9F",X"32",X"10",X"E0",X"C9",X"3A",X"10",X"E0",X"CB",X"5F",X"C0",X"CB",
		X"DF",X"32",X"10",X"E0",X"3A",X"03",X"E0",X"47",X"3A",X"01",X"E0",X"3C",X"32",X"01",X"E0",X"B8",
		X"C0",X"AF",X"32",X"01",X"E0",X"3A",X"05",X"E0",X"47",X"3A",X"00",X"E0",X"80",X"FE",X"99",X"38",
		X"02",X"3E",X"99",X"32",X"00",X"E0",X"3E",X"01",X"D7",X"3A",X"00",X"D0",X"2F",X"CB",X"7F",X"20",
		X"09",X"3A",X"10",X"E0",X"CB",X"BF",X"32",X"10",X"E0",X"C9",X"3A",X"10",X"E0",X"CB",X"7F",X"C0",
		X"CB",X"FF",X"32",X"10",X"E0",X"3A",X"04",X"E0",X"47",X"3A",X"02",X"E0",X"3C",X"32",X"02",X"E0",
		X"B8",X"C0",X"AF",X"32",X"02",X"E0",X"3A",X"06",X"E0",X"47",X"3A",X"00",X"E0",X"80",X"FE",X"99",
		X"38",X"02",X"3E",X"99",X"32",X"00",X"E0",X"3E",X"01",X"D7",X"C9",X"E5",X"C5",X"2A",X"80",X"E2",
		X"DD",X"7E",X"03",X"E6",X"F8",X"CB",X"3F",X"CB",X"3F",X"47",X"7D",X"E6",X"F8",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"0C",X"38",X"03",X"80",X"18",X"16",X"C6",X"40",X"CB",X"7F",X"28",X"07",X"80",X"CB",
		X"7F",X"28",X"09",X"18",X"09",X"80",X"CB",X"7F",X"20",X"02",X"18",X"02",X"D6",X"80",X"CB",X"87",
		X"6F",X"DD",X"7E",X"00",X"C6",X"08",X"4F",X"E6",X"F0",X"2F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"C6",X"80",X"67",X"CB",X"59",X"20",X"04",X"3E",X"80",X"85",X"6F",X"E5",X"FD",X"E1",
		X"21",X"E7",X"1F",X"FD",X"7E",X"01",X"E6",X"F0",X"07",X"07",X"E6",X"0F",X"4F",X"06",X"00",X"09",
		X"7E",X"FD",X"BE",X"00",X"C1",X"E1",X"C9",X"9A",X"74",X"B8",X"C8",X"C5",X"E5",X"2A",X"68",X"E0",
		X"44",X"4D",X"29",X"09",X"79",X"84",X"67",X"22",X"68",X"E0",X"B5",X"CA",X"02",X"20",X"7C",X"C3",
		X"09",X"20",X"21",X"5A",X"36",X"22",X"68",X"E0",X"7C",X"E6",X"0F",X"E1",X"C1",X"C9",X"D5",X"E5",
		X"16",X"00",X"5F",X"2E",X"00",X"60",X"06",X"08",X"29",X"30",X"01",X"19",X"10",X"FA",X"22",X"87",
		X"E2",X"E1",X"D1",X"C9",X"3A",X"83",X"E2",X"E6",X"0F",X"C0",X"21",X"3B",X"20",X"3A",X"A9",X"E2",
		X"CB",X"27",X"4F",X"06",X"00",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"9C",X"21",X"5B",X"20",X"0E",
		X"22",X"0E",X"22",X"0E",X"22",X"FF",X"21",X"1A",X"22",X"DD",X"20",X"0A",X"21",X"50",X"23",X"0E",
		X"22",X"0E",X"22",X"7A",X"22",X"0E",X"22",X"0E",X"22",X"C9",X"22",X"3A",X"63",X"E0",X"FE",X"03",
		X"C2",X"FB",X"22",X"3E",X"20",X"E7",X"CD",X"EB",X"1F",X"E6",X"03",X"CA",X"63",X"20",X"3D",X"32",
		X"C7",X"E2",X"3C",X"FE",X"03",X"DA",X"79",X"20",X"AF",X"32",X"C8",X"E2",X"3C",X"FE",X"03",X"DA",
		X"83",X"20",X"AF",X"32",X"C9",X"E2",X"3A",X"C7",X"E2",X"DD",X"21",X"B0",X"E1",X"16",X"58",X"CD",
		X"AD",X"20",X"3A",X"C8",X"E2",X"DD",X"21",X"10",X"E2",X"16",X"90",X"CD",X"AD",X"20",X"3A",X"C9",
		X"E2",X"DD",X"21",X"70",X"E2",X"16",X"C8",X"CD",X"AD",X"20",X"C3",X"FB",X"22",X"21",X"BB",X"23",
		X"CB",X"27",X"CB",X"27",X"4F",X"06",X"00",X"09",X"7E",X"DD",X"77",X"01",X"23",X"7E",X"DD",X"77",
		X"02",X"23",X"7E",X"DD",X"77",X"05",X"23",X"7E",X"DD",X"77",X"06",X"DD",X"72",X"00",X"7A",X"C6",
		X"10",X"DD",X"77",X"04",X"DD",X"36",X"03",X"99",X"DD",X"36",X"07",X"99",X"C9",X"3A",X"63",X"E0",
		X"FE",X"03",X"C2",X"FB",X"22",X"3A",X"C0",X"E1",X"FE",X"84",X"D2",X"F3",X"20",X"3A",X"C7",X"E2",
		X"C3",X"01",X"21",X"FE",X"BC",X"D2",X"FE",X"20",X"3A",X"C8",X"E2",X"C3",X"01",X"21",X"3A",X"C9",
		X"E2",X"32",X"CD",X"E2",X"CD",X"57",X"21",X"C3",X"FB",X"22",X"3A",X"63",X"E0",X"FE",X"03",X"C2",
		X"FB",X"22",X"3A",X"CD",X"E2",X"21",X"A8",X"23",X"CB",X"27",X"4F",X"06",X"00",X"09",X"5E",X"23",
		X"56",X"EB",X"06",X"0A",X"E5",X"CD",X"FA",X"06",X"CD",X"1F",X"10",X"CA",X"34",X"21",X"CD",X"59",
		X"06",X"C3",X"3F",X"21",X"CD",X"15",X"06",X"3E",X"03",X"CD",X"DE",X"1E",X"CD",X"F8",X"1E",X"E1",
		X"11",X"01",X"00",X"A7",X"ED",X"52",X"F5",X"7D",X"E6",X"0F",X"C2",X"50",X"21",X"3E",X"13",X"D7",
		X"F1",X"D2",X"22",X"21",X"C3",X"FB",X"22",X"F5",X"CD",X"B1",X"2C",X"F1",X"21",X"AE",X"23",X"11",
		X"A0",X"88",X"01",X"0D",X"00",X"CF",X"DD",X"21",X"C0",X"E1",X"21",X"BB",X"23",X"CB",X"27",X"CB",
		X"27",X"4F",X"06",X"00",X"09",X"7E",X"DD",X"77",X"01",X"23",X"7E",X"DD",X"77",X"02",X"23",X"7E",
		X"DD",X"77",X"05",X"23",X"7E",X"DD",X"77",X"06",X"DD",X"36",X"00",X"90",X"DD",X"36",X"04",X"A0",
		X"3E",X"70",X"DD",X"77",X"03",X"DD",X"77",X"07",X"CD",X"F3",X"21",X"C9",X"3A",X"63",X"E0",X"FE",
		X"03",X"CA",X"BD",X"21",X"CD",X"B1",X"2C",X"21",X"C7",X"23",X"11",X"BC",X"E1",X"01",X"14",X"00",
		X"ED",X"B0",X"11",X"20",X"E2",X"01",X"04",X"00",X"ED",X"B0",X"C3",X"FB",X"22",X"3A",X"80",X"E2",
		X"E6",X"80",X"32",X"00",X"90",X"21",X"C0",X"E1",X"11",X"C0",X"8F",X"01",X"14",X"00",X"ED",X"B0",
		X"CD",X"B1",X"2C",X"21",X"C0",X"8F",X"11",X"60",X"E1",X"06",X"03",X"C5",X"E5",X"D5",X"01",X"14",
		X"00",X"ED",X"B0",X"D1",X"21",X"60",X"00",X"19",X"EB",X"E1",X"C1",X"10",X"EE",X"CD",X"F3",X"21",
		X"C3",X"FB",X"22",X"21",X"DF",X"23",X"11",X"D4",X"E1",X"01",X"10",X"00",X"ED",X"B0",X"C9",X"AF",
		X"21",X"00",X"80",X"06",X"0C",X"CD",X"EE",X"1E",X"32",X"00",X"90",X"32",X"00",X"A0",X"06",X"04",
		X"3E",X"FF",X"CD",X"DE",X"1E",X"10",X"F9",X"C3",X"FB",X"22",X"3A",X"63",X"E0",X"FE",X"03",X"CA",
		X"FB",X"22",X"CD",X"1F",X"10",X"CA",X"2E",X"22",X"3A",X"85",X"E0",X"C3",X"31",X"22",X"3A",X"84",
		X"E0",X"FE",X"01",X"C2",X"3C",X"22",X"21",X"EF",X"23",X"C3",X"3F",X"22",X"21",X"01",X"24",X"11",
		X"2D",X"8A",X"01",X"12",X"00",X"CF",X"21",X"13",X"24",X"11",X"2C",X"8A",X"01",X"12",X"00",X"CF",
		X"3E",X"20",X"11",X"2B",X"8A",X"06",X"12",X"CD",X"D3",X"1E",X"3E",X"28",X"32",X"2A",X"8A",X"3E",
		X"05",X"32",X"AA",X"87",X"3E",X"07",X"32",X"2A",X"87",X"3E",X"05",X"32",X"AA",X"84",X"3C",X"32",
		X"2A",X"84",X"3E",X"29",X"32",X"AA",X"81",X"C3",X"FB",X"22",X"21",X"9B",X"23",X"11",X"98",X"88",
		X"01",X"0D",X"00",X"CF",X"3A",X"CA",X"E4",X"F5",X"A7",X"C2",X"94",X"22",X"3E",X"09",X"32",X"14",
		X"87",X"C3",X"9B",X"22",X"FD",X"21",X"14",X"87",X"CD",X"F2",X"16",X"3E",X"13",X"D7",X"21",X"95",
		X"23",X"11",X"14",X"86",X"01",X"06",X"00",X"CF",X"F1",X"4F",X"06",X"0A",X"C5",X"41",X"CD",X"FA",
		X"06",X"C1",X"10",X"F8",X"3E",X"05",X"D7",X"CD",X"1F",X"10",X"CA",X"C3",X"22",X"CD",X"59",X"06",
		X"C3",X"0E",X"22",X"CD",X"15",X"06",X"C3",X"0E",X"22",X"CD",X"B1",X"2C",X"3A",X"63",X"E0",X"FE",
		X"03",X"D2",X"00",X"23",X"CD",X"6F",X"17",X"CD",X"C8",X"2B",X"CD",X"F6",X"02",X"3E",X"01",X"32",
		X"63",X"E0",X"AF",X"32",X"BA",X"E5",X"32",X"82",X"E2",X"32",X"93",X"E2",X"32",X"8B",X"E2",X"32",
		X"A9",X"E2",X"21",X"00",X"E5",X"06",X"A0",X"CD",X"E9",X"1E",X"C9",X"21",X"A9",X"E2",X"34",X"C9",
		X"CD",X"1F",X"10",X"CA",X"26",X"23",X"21",X"00",X"00",X"22",X"66",X"E0",X"22",X"77",X"E0",X"AF",
		X"32",X"7A",X"E0",X"32",X"6F",X"E0",X"32",X"83",X"E0",X"32",X"85",X"E0",X"32",X"CA",X"E4",X"21",
		X"8B",X"E0",X"34",X"C3",X"43",X"23",X"21",X"00",X"00",X"22",X"64",X"E0",X"22",X"75",X"E0",X"AF",
		X"32",X"79",X"E0",X"32",X"6E",X"E0",X"32",X"82",X"E0",X"32",X"84",X"E0",X"32",X"CA",X"E4",X"21",
		X"8A",X"E0",X"34",X"3E",X"64",X"32",X"C9",X"E4",X"3E",X"01",X"32",X"6B",X"E0",X"AF",X"D7",X"C9",
		X"3A",X"C9",X"E4",X"A7",X"CA",X"FB",X"22",X"F5",X"47",X"C5",X"CD",X"3C",X"17",X"06",X"0A",X"CD",
		X"1F",X"10",X"CA",X"6E",X"23",X"CD",X"0C",X"07",X"CD",X"59",X"06",X"C3",X"74",X"23",X"CD",X"00",
		X"07",X"CD",X"15",X"06",X"CD",X"F3",X"05",X"CD",X"F8",X"1E",X"C1",X"78",X"E6",X"0F",X"C2",X"84",
		X"23",X"3E",X"13",X"D7",X"3E",X"10",X"CD",X"DE",X"1E",X"10",X"CE",X"CD",X"3C",X"17",X"F1",X"32",
		X"C9",X"E4",X"C3",X"FB",X"22",X"40",X"31",X"30",X"30",X"3C",X"3E",X"42",X"4F",X"4E",X"55",X"53",
		X"20",X"4F",X"46",X"20",X"42",X"55",X"4D",X"50",X"C8",X"00",X"F4",X"01",X"E8",X"03",X"53",X"50",
		X"45",X"43",X"49",X"41",X"4C",X"20",X"42",X"4F",X"4E",X"55",X"53",X"42",X"27",X"42",X"24",X"40",
		X"26",X"40",X"24",X"43",X"25",X"43",X"24",X"70",X"40",X"A8",X"80",X"80",X"40",X"A7",X"80",X"90",
		X"40",X"A5",X"80",X"A0",X"40",X"A3",X"80",X"B0",X"40",X"A1",X"80",X"C0",X"40",X"9F",X"80",X"80",
		X"40",X"A6",X"D8",X"90",X"40",X"A4",X"D8",X"A0",X"40",X"A2",X"D8",X"B0",X"40",X"A0",X"D8",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"27",X"27",X"27",X"27",X"27",
		X"37",X"20",X"20",X"20",X"20",X"20",X"20",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"37",X"5C",X"5D",X"5D",X"5D",X"5D",X"5D",X"5C",X"5D",X"5D",X"5D",X"5D",X"5D",X"5C",
		X"5D",X"5D",X"5D",X"5D",X"5C",X"3A",X"96",X"E2",X"FE",X"02",X"DA",X"5B",X"24",X"3A",X"CA",X"E2",
		X"FE",X"30",X"D0",X"3A",X"83",X"E2",X"E6",X"03",X"C0",X"CD",X"60",X"24",X"C5",X"CD",X"3C",X"17",
		X"C1",X"21",X"CA",X"E2",X"34",X"3A",X"0A",X"E0",X"A7",X"20",X"05",X"7E",X"B8",X"D8",X"18",X"07",
		X"78",X"C6",X"05",X"47",X"7E",X"B8",X"D8",X"3E",X"30",X"77",X"C9",X"AF",X"32",X"CA",X"E2",X"C9",
		X"CD",X"1F",X"10",X"28",X"05",X"3A",X"8B",X"E0",X"18",X"03",X"3A",X"8A",X"E0",X"FE",X"02",X"3E",
		X"0F",X"30",X"02",X"D6",X"05",X"47",X"3A",X"C9",X"E4",X"A7",X"C0",X"3A",X"A6",X"E2",X"A7",X"C0",
		X"3E",X"01",X"32",X"A6",X"E2",X"C9",X"2A",X"66",X"E0",X"11",X"6F",X"E0",X"18",X"06",X"2A",X"64",
		X"E0",X"11",X"6E",X"E0",X"CD",X"A8",X"24",X"23",X"1A",X"E6",X"0F",X"47",X"7C",X"CB",X"27",X"CB",
		X"27",X"CB",X"27",X"E6",X"F0",X"80",X"12",X"C9",X"7D",X"FE",X"FF",X"C0",X"7C",X"FE",X"01",X"28",
		X"1B",X"FE",X"03",X"28",X"07",X"FE",X"05",X"C0",X"3E",X"30",X"12",X"C9",X"EB",X"3A",X"C0",X"E1",
		X"FE",X"A0",X"38",X"04",X"CB",X"C6",X"EB",X"C9",X"CB",X"86",X"18",X"FA",X"EB",X"3A",X"C0",X"E1",
		X"FE",X"A0",X"38",X"04",X"CB",X"CE",X"18",X"EE",X"CB",X"8E",X"18",X"EA",X"CD",X"1F",X"10",X"28",
		X"0A",X"ED",X"5B",X"66",X"E0",X"3A",X"6F",X"E0",X"4F",X"18",X"08",X"ED",X"5B",X"64",X"E0",X"3A",
		X"6E",X"E0",X"4F",X"D5",X"16",X"00",X"21",X"54",X"25",X"06",X"09",X"7E",X"B9",X"CA",X"05",X"25",
		X"14",X"23",X"10",X"F7",X"76",X"21",X"44",X"25",X"7A",X"CB",X"27",X"4F",X"06",X"00",X"09",X"5E",
		X"23",X"56",X"EB",X"D1",X"2B",X"46",X"23",X"C5",X"4E",X"23",X"46",X"2B",X"78",X"BA",X"CA",X"27",
		X"25",X"DA",X"2C",X"25",X"C3",X"2F",X"25",X"7B",X"B9",X"DA",X"2F",X"25",X"CD",X"37",X"25",X"01",
		X"05",X"00",X"09",X"C1",X"10",X"E1",X"C9",X"E5",X"D5",X"23",X"23",X"5E",X"23",X"56",X"23",X"7E",
		X"12",X"D1",X"E1",X"C9",X"5D",X"25",X"8B",X"25",X"54",X"26",X"F5",X"26",X"D2",X"27",X"F5",X"26",
		X"9B",X"28",X"91",X"29",X"00",X"10",X"12",X"20",X"21",X"22",X"23",X"30",X"09",X"00",X"00",X"7E",
		X"E0",X"00",X"00",X"00",X"CE",X"E4",X"00",X"BF",X"01",X"CE",X"E4",X"01",X"C7",X"01",X"CE",X"E4",
		X"00",X"C8",X"00",X"7E",X"E0",X"02",X"2F",X"01",X"7E",X"E0",X"04",X"44",X"01",X"7E",X"E0",X"01",
		X"E4",X"01",X"7E",X"E0",X"03",X"FC",X"01",X"7E",X"E0",X"04",X"28",X"00",X"02",X"CE",X"E2",X"00",
		X"00",X"02",X"B9",X"E2",X"00",X"00",X"02",X"CF",X"E4",X"00",X"00",X"02",X"AF",X"E2",X"00",X"1E",
		X"02",X"AF",X"E2",X"1A",X"BB",X"02",X"AF",X"E2",X"00",X"21",X"02",X"CE",X"E2",X"01",X"5F",X"02",
		X"CE",X"E2",X"00",X"65",X"02",X"B9",X"E2",X"01",X"87",X"02",X"B9",X"E2",X"00",X"8D",X"02",X"CE",
		X"E2",X"01",X"A6",X"02",X"CE",X"E2",X"00",X"AD",X"02",X"CE",X"E2",X"01",X"BB",X"02",X"CE",X"E2",
		X"00",X"31",X"03",X"CF",X"E4",X"0E",X"BF",X"03",X"CF",X"E4",X"00",X"00",X"02",X"7E",X"E0",X"04",
		X"0D",X"02",X"7E",X"E0",X"01",X"23",X"02",X"7E",X"E0",X"04",X"8F",X"02",X"7E",X"E0",X"00",X"A7",
		X"02",X"7E",X"E0",X"04",X"AF",X"02",X"7E",X"E0",X"00",X"BC",X"02",X"7E",X"E0",X"02",X"DA",X"02",
		X"7E",X"E0",X"04",X"E0",X"02",X"7E",X"E0",X"01",X"EB",X"02",X"7E",X"E0",X"03",X"12",X"03",X"7E",
		X"E0",X"02",X"1B",X"03",X"7E",X"E0",X"04",X"21",X"03",X"7E",X"E0",X"01",X"4B",X"03",X"7E",X"E0",
		X"04",X"54",X"03",X"7E",X"E0",X"02",X"69",X"03",X"7E",X"E0",X"00",X"A2",X"03",X"7E",X"E0",X"02",
		X"AC",X"03",X"7E",X"E0",X"04",X"B6",X"03",X"7E",X"E0",X"01",X"C4",X"03",X"7E",X"E0",X"04",X"CF",
		X"03",X"7E",X"E0",X"02",X"D4",X"03",X"7E",X"E0",X"04",X"DA",X"03",X"7E",X"E0",X"01",X"E8",X"03",
		X"7E",X"E0",X"03",X"20",X"00",X"02",X"CD",X"E4",X"00",X"00",X"02",X"CF",X"E4",X"00",X"00",X"02",
		X"C5",X"E2",X"00",X"00",X"02",X"AF",X"E2",X"00",X"2F",X"02",X"AF",X"E2",X"1A",X"C3",X"02",X"AF",
		X"E2",X"00",X"32",X"02",X"CD",X"E4",X"01",X"68",X"02",X"CD",X"E4",X"00",X"71",X"02",X"C5",X"E2",
		X"01",X"C3",X"02",X"C5",X"E2",X"00",X"69",X"03",X"CF",X"E4",X"0E",X"B7",X"03",X"CF",X"E4",X"00",
		X"00",X"02",X"7E",X"E0",X"04",X"04",X"02",X"7E",X"E0",X"02",X"08",X"02",X"7E",X"E0",X"04",X"0E",
		X"02",X"7E",X"E0",X"01",X"21",X"02",X"7E",X"E0",X"03",X"BF",X"02",X"7E",X"E0",X"04",X"C8",X"02",
		X"7E",X"E0",X"01",X"E5",X"02",X"7E",X"E0",X"03",X"03",X"03",X"7E",X"E0",X"00",X"3E",X"03",X"7E",
		X"E0",X"03",X"4C",X"03",X"7E",X"E0",X"02",X"54",X"03",X"7E",X"E0",X"04",X"5B",X"03",X"7E",X"E0",
		X"01",X"84",X"03",X"7E",X"E0",X"04",X"AF",X"03",X"7E",X"E0",X"01",X"C7",X"03",X"7E",X"E0",X"04",
		X"CF",X"03",X"7E",X"E0",X"02",X"D4",X"03",X"7E",X"E0",X"04",X"DB",X"03",X"7E",X"E0",X"01",X"E8",
		X"03",X"7E",X"E0",X"03",X"2C",X"00",X"04",X"CE",X"E4",X"00",X"00",X"04",X"CF",X"E4",X"00",X"34",
		X"04",X"CE",X"E4",X"02",X"3D",X"04",X"CE",X"E4",X"00",X"6E",X"04",X"CF",X"E4",X"0E",X"72",X"04",
		X"CF",X"E4",X"00",X"DF",X"04",X"CF",X"E4",X"0E",X"19",X"05",X"CF",X"E4",X"00",X"1B",X"05",X"CF",
		X"E4",X"0E",X"1F",X"05",X"CF",X"E4",X"00",X"97",X"05",X"CF",X"E4",X"0E",X"D3",X"05",X"CF",X"E4",
		X"00",X"00",X"04",X"7E",X"E0",X"04",X"19",X"04",X"7E",X"E0",X"00",X"20",X"04",X"7E",X"E0",X"04",
		X"29",X"04",X"7E",X"E0",X"01",X"4F",X"04",X"7E",X"E0",X"04",X"56",X"04",X"7E",X"E0",X"02",X"65",
		X"04",X"7E",X"E0",X"04",X"6C",X"04",X"7E",X"E0",X"01",X"7F",X"04",X"7E",X"E0",X"03",X"82",X"04",
		X"7E",X"E0",X"02",X"9E",X"04",X"7E",X"E0",X"04",X"A6",X"04",X"7E",X"E0",X"01",X"AE",X"04",X"7E",
		X"E0",X"03",X"D4",X"04",X"7E",X"E0",X"04",X"DD",X"04",X"7E",X"E0",X"01",X"E8",X"04",X"7E",X"E0",
		X"00",X"06",X"05",X"7E",X"E0",X"04",X"14",X"05",X"7E",X"E0",X"01",X"19",X"05",X"7E",X"E0",X"04",
		X"2D",X"05",X"7E",X"E0",X"01",X"2C",X"05",X"7E",X"E0",X"03",X"43",X"05",X"7E",X"E0",X"00",X"72",
		X"05",X"7E",X"E0",X"03",X"8A",X"05",X"7E",X"E0",X"02",X"92",X"05",X"7E",X"E0",X"04",X"9A",X"05",
		X"7E",X"E0",X"01",X"A0",X"05",X"7E",X"E0",X"04",X"A8",X"05",X"7E",X"E0",X"00",X"C1",X"05",X"7E",
		X"E0",X"04",X"CD",X"05",X"7E",X"E0",X"01",X"D7",X"05",X"7E",X"E0",X"02",X"EA",X"05",X"7E",X"E0",
		X"00",X"29",X"00",X"04",X"CE",X"E4",X"00",X"00",X"04",X"BA",X"E2",X"00",X"00",X"04",X"CC",X"E4",
		X"00",X"00",X"04",X"CF",X"E4",X"00",X"00",X"04",X"AF",X"E2",X"00",X"60",X"04",X"AF",X"E2",X"1A",
		X"E5",X"04",X"AF",X"E2",X"00",X"34",X"04",X"CE",X"E4",X"02",X"3D",X"04",X"CE",X"E4",X"00",X"63",
		X"04",X"BA",X"E2",X"01",X"85",X"04",X"BA",X"E2",X"00",X"8E",X"04",X"CC",X"E4",X"05",X"E5",X"04",
		X"CC",X"E4",X"00",X"2E",X"05",X"CF",X"E4",X"0E",X"84",X"05",X"CF",X"E4",X"00",X"00",X"04",X"7E",
		X"E0",X"04",X"19",X"04",X"7E",X"E0",X"00",X"20",X"04",X"7E",X"E0",X"04",X"29",X"04",X"7E",X"E0",
		X"01",X"53",X"04",X"7E",X"E0",X"03",X"BB",X"04",X"7E",X"E0",X"00",X"C9",X"04",X"7E",X"E0",X"02",
		X"DE",X"04",X"7E",X"E0",X"04",X"E5",X"04",X"7E",X"E0",X"01",X"EE",X"04",X"7E",X"E0",X"03",X"15",
		X"05",X"7E",X"E0",X"02",X"1F",X"05",X"7E",X"E0",X"04",X"26",X"05",X"7E",X"E0",X"01",X"3F",X"05",
		X"7E",X"E0",X"04",X"47",X"05",X"7E",X"E0",X"02",X"5A",X"05",X"7E",X"E0",X"00",X"73",X"05",X"7E",
		X"E0",X"04",X"7A",X"05",X"7E",X"E0",X"01",X"8B",X"05",X"7E",X"E0",X"04",X"92",X"05",X"7E",X"E0",
		X"02",X"A3",X"05",X"7E",X"E0",X"00",X"CB",X"05",X"7E",X"E0",X"02",X"D5",X"05",X"7E",X"E0",X"04",
		X"EB",X"05",X"7E",X"E0",X"02",X"EA",X"05",X"7E",X"E0",X"00",X"32",X"00",X"04",X"CE",X"E4",X"00",
		X"00",X"04",X"CE",X"E2",X"00",X"00",X"04",X"CF",X"E4",X"00",X"00",X"04",X"B9",X"E2",X"00",X"00",
		X"04",X"AF",X"E2",X"00",X"60",X"04",X"AF",X"E2",X"1A",X"F2",X"04",X"AF",X"E2",X"00",X"34",X"04",
		X"CE",X"E4",X"02",X"3D",X"04",X"CE",X"E4",X"00",X"63",X"04",X"CE",X"E2",X"01",X"88",X"04",X"CE",
		X"E2",X"00",X"8F",X"04",X"B9",X"E2",X"01",X"A8",X"04",X"B9",X"E2",X"00",X"AD",X"04",X"CE",X"E2",
		X"01",X"C6",X"04",X"CE",X"E2",X"00",X"CC",X"04",X"B9",X"E2",X"01",X"DB",X"04",X"B9",X"E2",X"00",
		X"E1",X"04",X"CE",X"E2",X"01",X"E6",X"04",X"CE",X"E2",X"00",X"65",X"05",X"CF",X"E4",X"0E",X"D9",
		X"05",X"CF",X"E4",X"00",X"00",X"04",X"7E",X"E0",X"04",X"19",X"04",X"7E",X"E0",X"00",X"20",X"04",
		X"7E",X"E0",X"04",X"29",X"04",X"7E",X"E0",X"01",X"4F",X"04",X"7E",X"E0",X"04",X"57",X"04",X"7E",
		X"E0",X"02",X"66",X"04",X"7E",X"E0",X"00",X"89",X"04",X"7E",X"E0",X"01",X"AE",X"04",X"7E",X"E0",
		X"00",X"C7",X"04",X"7E",X"E0",X"01",X"E2",X"04",X"7E",X"E0",X"00",X"E6",X"04",X"7E",X"E0",X"04",
		X"EE",X"04",X"7E",X"E0",X"00",X"F2",X"04",X"7E",X"E0",X"02",X"10",X"05",X"7E",X"E0",X"04",X"17",
		X"05",X"7E",X"E0",X"01",X"20",X"05",X"7E",X"E0",X"03",X"49",X"05",X"7E",X"E0",X"02",X"51",X"05",
		X"7E",X"E0",X"04",X"59",X"05",X"7E",X"E0",X"01",X"81",X"05",X"7E",X"E0",X"04",X"89",X"05",X"7E",
		X"E0",X"02",X"9C",X"05",X"7E",X"E0",X"00",X"C0",X"05",X"7E",X"E0",X"02",X"C9",X"05",X"7E",X"E0",
		X"04",X"D8",X"05",X"7E",X"E0",X"01",X"E1",X"05",X"7E",X"E0",X"04",X"EA",X"05",X"7E",X"E0",X"00",
		X"1A",X"00",X"06",X"CE",X"E4",X"00",X"00",X"06",X"CF",X"E4",X"00",X"FF",X"07",X"63",X"E0",X"03",
		X"00",X"06",X"AF",X"E2",X"00",X"EC",X"07",X"AF",X"E2",X"1E",X"29",X"06",X"CE",X"E4",X"03",X"31",
		X"06",X"CE",X"E4",X"00",X"FE",X"06",X"CF",X"E4",X"0E",X"38",X"07",X"CF",X"E4",X"00",X"00",X"06",
		X"7E",X"E0",X"00",X"16",X"06",X"7E",X"E0",X"04",X"1F",X"06",X"7E",X"E0",X"01",X"67",X"06",X"7E",
		X"E0",X"04",X"6F",X"06",X"7E",X"E0",X"02",X"7D",X"06",X"7E",X"E0",X"04",X"89",X"06",X"7E",X"E0",
		X"00",X"AB",X"06",X"7E",X"E0",X"02",X"C2",X"06",X"7E",X"E0",X"04",X"CB",X"06",X"7E",X"E0",X"03",
		X"F8",X"06",X"7E",X"E0",X"04",X"01",X"07",X"7E",X"E0",X"01",X"0F",X"07",X"7E",X"E0",X"04",X"1A",
		X"07",X"7E",X"E0",X"00",X"29",X"07",X"7E",X"E0",X"04",X"40",X"07",X"7E",X"E0",X"00",X"C5",X"07",
		X"7E",X"E0",X"04",X"CD",X"A4",X"2B",X"21",X"50",X"2A",X"11",X"30",X"8F",X"01",X"06",X"00",X"CF",
		X"11",X"31",X"8F",X"01",X"06",X"00",X"CF",X"11",X"16",X"8F",X"01",X"06",X"00",X"CF",X"11",X"17",
		X"8F",X"01",X"06",X"00",X"CF",X"21",X"18",X"8F",X"11",X"98",X"8C",X"06",X"0C",X"C5",X"3E",X"A3",
		X"77",X"12",X"23",X"13",X"3E",X"70",X"77",X"3E",X"60",X"12",X"23",X"13",X"C1",X"10",X"EE",X"C9",
		X"A4",X"70",X"70",X"70",X"70",X"A4",X"50",X"40",X"40",X"40",X"40",X"40",X"A4",X"6F",X"A6",X"6E",
		X"A5",X"A4",X"70",X"60",X"60",X"60",X"60",X"60",X"3A",X"A7",X"E2",X"A7",X"C8",X"3A",X"CC",X"E2",
		X"A7",X"C2",X"93",X"2A",X"06",X"20",X"21",X"BA",X"2A",X"5E",X"23",X"56",X"1A",X"E6",X"F0",X"C6",
		X"0C",X"12",X"23",X"10",X"F4",X"21",X"CC",X"E2",X"34",X"7E",X"FE",X"11",X"D8",X"AF",X"77",X"32",
		X"A7",X"E2",X"C9",X"3A",X"83",X"E2",X"E6",X"3F",X"C0",X"21",X"BA",X"2A",X"3A",X"CC",X"E2",X"3D",
		X"CB",X"27",X"CB",X"27",X"4F",X"06",X"00",X"09",X"5E",X"23",X"56",X"1A",X"E6",X"F0",X"12",X"23",
		X"5E",X"23",X"56",X"1A",X"E6",X"F0",X"12",X"C3",X"85",X"2A",X"31",X"8E",X"B1",X"8D",X"B1",X"8E",
		X"31",X"8D",X"31",X"8F",X"B1",X"8C",X"2F",X"8F",X"AF",X"8C",X"2D",X"8F",X"AD",X"8C",X"2B",X"8F",
		X"AB",X"8C",X"29",X"8F",X"A9",X"8C",X"27",X"8F",X"A7",X"8C",X"25",X"8F",X"A5",X"8C",X"23",X"8F",
		X"A3",X"8C",X"21",X"8F",X"A1",X"8C",X"1F",X"8F",X"9F",X"8C",X"1D",X"8F",X"9D",X"8C",X"1B",X"8F",
		X"9B",X"8C",X"19",X"8F",X"99",X"8C",X"17",X"8F",X"97",X"8C",X"2A",X"64",X"E0",X"ED",X"5B",X"75",
		X"E0",X"3A",X"6E",X"E0",X"C3",X"11",X"2B",X"2A",X"66",X"E0",X"ED",X"5B",X"77",X"E0",X"3A",X"6F",
		X"E0",X"2C",X"20",X"03",X"CB",X"0C",X"D8",X"CD",X"C7",X"0F",X"19",X"06",X"03",X"0E",X"00",X"E5",
		X"5E",X"23",X"56",X"EB",X"11",X"19",X"00",X"A7",X"ED",X"52",X"7E",X"E1",X"B9",X"20",X"06",X"4F",
		X"23",X"23",X"C3",X"1F",X"2B",X"4F",X"CD",X"3E",X"2B",X"23",X"23",X"10",X"E2",X"C9",X"78",X"FE",
		X"02",X"20",X"0D",X"79",X"FE",X"06",X"28",X"05",X"FE",X"09",X"28",X"01",X"AF",X"32",X"CB",X"E2",
		X"3A",X"BA",X"E2",X"A7",X"28",X"07",X"79",X"FE",X"15",X"20",X"02",X"0E",X"13",X"E5",X"C5",X"11",
		X"98",X"8E",X"21",X"C0",X"E4",X"78",X"ED",X"44",X"C6",X"03",X"47",X"85",X"6F",X"78",X"CB",X"27",
		X"CB",X"27",X"CB",X"27",X"83",X"5F",X"CB",X"B9",X"CB",X"B1",X"7E",X"B9",X"CA",X"84",X"2B",X"71",
		X"41",X"CD",X"87",X"2B",X"C1",X"E1",X"C9",X"D5",X"21",X"ED",X"4A",X"11",X"20",X"00",X"05",X"CA",
		X"95",X"2B",X"19",X"10",X"FD",X"D1",X"06",X"08",X"C5",X"D5",X"01",X"04",X"00",X"CF",X"D1",X"13",
		X"C1",X"10",X"F5",X"C9",X"21",X"B0",X"2B",X"11",X"18",X"8C",X"01",X"04",X"00",X"ED",X"B0",X"C9",
		X"11",X"A8",X"10",X"A8",X"3A",X"A7",X"E2",X"A7",X"20",X"0A",X"3A",X"AF",X"E2",X"A7",X"20",X"02",
		X"3E",X"23",X"E7",X"C9",X"3E",X"22",X"18",X"FA",X"CD",X"31",X"10",X"CD",X"DC",X"24",X"CD",X"13",
		X"2A",X"CD",X"1F",X"10",X"28",X"05",X"2A",X"66",X"E0",X"18",X"03",X"2A",X"64",X"E0",X"EB",X"D5",
		X"3E",X"01",X"32",X"82",X"E2",X"CD",X"09",X"0C",X"CD",X"F8",X"1E",X"CD",X"39",X"1F",X"CD",X"1F",
		X"10",X"CA",X"FA",X"2B",X"2A",X"66",X"E0",X"C3",X"FD",X"2B",X"2A",X"64",X"E0",X"D1",X"A7",X"ED",
		X"52",X"7D",X"FE",X"03",X"D0",X"C3",X"DF",X"2B",X"3A",X"83",X"E2",X"A7",X"C0",X"3A",X"84",X"E2",
		X"E6",X"03",X"C0",X"CD",X"1F",X"10",X"C2",X"29",X"2C",X"3A",X"52",X"E0",X"47",X"3A",X"51",X"E0",
		X"21",X"BC",X"E0",X"11",X"89",X"E2",X"C3",X"36",X"2C",X"3A",X"5B",X"E0",X"47",X"3A",X"5A",X"E0",
		X"21",X"BD",X"E0",X"11",X"8A",X"E2",X"CB",X"20",X"CB",X"20",X"CB",X"20",X"CB",X"20",X"80",X"46",
		X"77",X"90",X"27",X"12",X"C9",X"3A",X"85",X"E0",X"47",X"3A",X"8A",X"E2",X"CD",X"1F",X"10",X"20",
		X"07",X"3A",X"84",X"E0",X"47",X"3A",X"89",X"E2",X"4F",X"3A",X"00",X"E3",X"B9",X"C8",X"79",X"32",
		X"00",X"E3",X"80",X"FE",X"05",X"D8",X"E6",X"01",X"47",X"3A",X"7E",X"E0",X"B0",X"20",X"0B",X"00",
		X"3A",X"BF",X"E5",X"A7",X"C0",X"3C",X"32",X"AF",X"E5",X"C9",X"3A",X"AF",X"E5",X"A7",X"C0",X"3E",
		X"01",X"32",X"BF",X"E5",X"C9",X"3A",X"A6",X"E2",X"A7",X"C8",X"CD",X"6F",X"17",X"AF",X"32",X"6B",
		X"E0",X"3A",X"C9",X"E4",X"A7",X"C2",X"AC",X"2C",X"3A",X"83",X"E2",X"E6",X"03",X"C0",X"21",X"A6",
		X"E2",X"34",X"7E",X"FE",X"40",X"D8",X"3E",X"01",X"32",X"A8",X"E2",X"C9",X"AF",X"32",X"A6",X"E2",
		X"C9",X"AF",X"21",X"00",X"E1",X"06",X"01",X"CD",X"EE",X"1E",X"06",X"80",X"CD",X"E9",X"1E",X"C9",
		X"06",X"05",X"21",X"A0",X"8D",X"16",X"B8",X"1E",X"AA",X"C5",X"06",X"0C",X"72",X"23",X"73",X"23",
		X"14",X"10",X"F9",X"D5",X"11",X"68",X"FF",X"19",X"D1",X"C1",X"10",X"ED",X"21",X"36",X"7F",X"11",
		X"60",X"E1",X"01",X"58",X"00",X"ED",X"B0",X"21",X"8E",X"7F",X"11",X"C0",X"E1",X"01",X"40",X"00",
		X"ED",X"B0",X"21",X"CE",X"7F",X"11",X"20",X"E2",X"01",X"20",X"00",X"ED",X"B0",X"C9",X"3E",X"5B",
		X"32",X"06",X"8E",X"3E",X"13",X"32",X"86",X"8D",X"3E",X"08",X"32",X"08",X"8E",X"21",X"45",X"2D",
		X"11",X"10",X"8C",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"71",X"2D",X"11",X"0C",X"89",X"01",X"05",X"00",X"CF",X"11",X"0A",X"89",X"01",
		X"05",X"00",X"CF",X"11",X"06",X"8D",X"01",X"04",X"00",X"CF",X"21",X"5E",X"2D",X"11",X"86",X"8A",
		X"01",X"13",X"00",X"CF",X"C9",X"54",X"41",X"49",X"54",X"4F",X"20",X"43",X"4F",X"52",X"50",X"4F",
		X"52",X"41",X"54",X"49",X"4F",X"4E",X"4E",X"4E",X"53",X"45",X"44",X"20",X"42",X"59",X"53",X"45",
		X"49",X"42",X"55",X"20",X"4B",X"41",X"49",X"48",X"41",X"54",X"53",X"55",X"20",X"49",X"4E",X"43",
		X"2E",X"1B",X"19",X"1F",X"1D",X"5F",X"1A",X"18",X"1E",X"1C",X"5E",X"31",X"39",X"38",X"35",X"3A",
		X"7C",X"E0",X"0F",X"D2",X"93",X"2D",X"CB",X"47",X"CA",X"8F",X"2D",X"CD",X"F1",X"03",X"C9",X"CD",
		X"C1",X"03",X"C9",X"21",X"7B",X"E0",X"CB",X"7E",X"C2",X"AC",X"2D",X"CB",X"46",X"C2",X"A8",X"2D",
		X"E5",X"CD",X"D3",X"2D",X"E1",X"CB",X"C6",X"C9",X"F1",X"C3",X"A0",X"2F",X"21",X"00",X"00",X"22",
		X"64",X"E0",X"22",X"75",X"E0",X"AF",X"32",X"7B",X"E0",X"32",X"6A",X"E0",X"32",X"6E",X"E0",X"32",
		X"CE",X"E2",X"21",X"00",X"E1",X"06",X"06",X"CD",X"EE",X"1E",X"21",X"7C",X"E0",X"34",X"21",X"89",
		X"E0",X"34",X"C9",X"21",X"6A",X"E0",X"CB",X"E6",X"AF",X"32",X"A6",X"E2",X"32",X"C8",X"E4",X"3E",
		X"64",X"32",X"F0",X"E0",X"CD",X"EB",X"2D",X"CD",X"4A",X"02",X"C9",X"3A",X"89",X"E0",X"E6",X"01",
		X"21",X"14",X"2E",X"4F",X"CB",X"27",X"CB",X"27",X"81",X"4F",X"06",X"00",X"09",X"5E",X"23",X"56",
		X"ED",X"53",X"64",X"E0",X"23",X"7E",X"32",X"75",X"E0",X"23",X"7E",X"32",X"79",X"E0",X"23",X"7E",
		X"32",X"6E",X"E0",X"C9",X"00",X"00",X"00",X"8C",X"00",X"21",X"02",X"0A",X"41",X"10",X"3A",X"83",
		X"E2",X"E6",X"1F",X"C0",X"DD",X"21",X"C0",X"E1",X"3A",X"C2",X"E2",X"2F",X"47",X"CD",X"EB",X"1F",
		X"FE",X"08",X"D2",X"56",X"2E",X"0F",X"D2",X"3E",X"2E",X"0E",X"80",X"C3",X"40",X"2E",X"0E",X"C0",
		X"DD",X"7E",X"00",X"B9",X"DA",X"50",X"2E",X"CA",X"56",X"2E",X"CD",X"AB",X"2E",X"C3",X"59",X"2E",
		X"CD",X"B0",X"2E",X"C3",X"59",X"2E",X"CD",X"C4",X"2E",X"DD",X"21",X"D4",X"E1",X"3A",X"C0",X"E1",
		X"DD",X"77",X"00",X"3A",X"C3",X"E1",X"C6",X"40",X"DD",X"77",X"03",X"CD",X"7B",X"1F",X"D2",X"9C",
		X"2E",X"DD",X"7E",X"00",X"C6",X"10",X"DD",X"77",X"00",X"CD",X"7B",X"1F",X"D2",X"93",X"2E",X"DD",
		X"7E",X"00",X"D6",X"20",X"DD",X"77",X"00",X"CD",X"7B",X"1F",X"D2",X"A2",X"2E",X"CD",X"BA",X"2E",
		X"C3",X"C9",X"2E",X"CD",X"B0",X"2E",X"CD",X"BA",X"2E",X"C3",X"C9",X"2E",X"CD",X"B5",X"2E",X"C3",
		X"C9",X"2E",X"CD",X"AB",X"2E",X"CD",X"BA",X"2E",X"C3",X"C9",X"2E",X"CB",X"80",X"CB",X"C8",X"C9",
		X"CB",X"88",X"CB",X"C0",X"C9",X"CB",X"B8",X"CB",X"E8",X"C9",X"CB",X"A8",X"CB",X"F8",X"C9",X"CB",
		X"A8",X"CB",X"B8",X"C9",X"CB",X"80",X"CB",X"88",X"C9",X"78",X"2F",X"32",X"C2",X"E2",X"C9",X"3A",
		X"A7",X"E2",X"0F",X"D0",X"DD",X"21",X"C0",X"E1",X"11",X"04",X"00",X"DD",X"7E",X"01",X"E6",X"F0",
		X"C6",X"03",X"06",X"04",X"CD",X"A8",X"1E",X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"7C",X"E0",X"A7",
		X"CA",X"FF",X"2E",X"21",X"C2",X"E2",X"11",X"87",X"E0",X"01",X"02",X"00",X"ED",X"B0",X"C9",X"21",
		X"01",X"D0",X"11",X"87",X"E0",X"01",X"02",X"00",X"ED",X"B0",X"C9",X"3A",X"A6",X"E2",X"A7",X"C0",
		X"3A",X"B0",X"E2",X"A7",X"C0",X"CD",X"47",X"12",X"CD",X"07",X"1B",X"3A",X"AC",X"E2",X"A7",X"CA",
		X"2B",X"2F",X"CD",X"C8",X"14",X"3A",X"83",X"E2",X"E6",X"03",X"C0",X"3A",X"7C",X"E0",X"A7",X"C4",
		X"1E",X"2E",X"CD",X"6D",X"13",X"CD",X"F4",X"14",X"C9",X"3A",X"A6",X"E2",X"A7",X"C0",X"CD",X"47",
		X"12",X"CD",X"45",X"18",X"CD",X"48",X"19",X"CD",X"25",X"24",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",
		X"E5",X"FD",X"E5",X"21",X"7F",X"E2",X"11",X"7F",X"C8",X"01",X"40",X"00",X"ED",X"B8",X"0E",X"20",
		X"1E",X"3F",X"ED",X"B8",X"11",X"7F",X"C9",X"0E",X"40",X"ED",X"B8",X"0E",X"20",X"1E",X"3F",X"ED",
		X"B8",X"11",X"FF",X"C8",X"0E",X"40",X"ED",X"B8",X"0E",X"20",X"1E",X"BF",X"ED",X"B8",X"3A",X"7C",
		X"E0",X"A7",X"28",X"05",X"CD",X"7F",X"2D",X"18",X"60",X"3A",X"C8",X"E4",X"A7",X"C4",X"96",X"01",
		X"3A",X"63",X"E0",X"A7",X"28",X"53",X"FE",X"01",X"28",X"06",X"CD",X"24",X"20",X"C3",X"E9",X"2F",
		X"3A",X"96",X"E2",X"A7",X"20",X"09",X"AF",X"32",X"96",X"E2",X"CD",X"0B",X"2F",X"18",X"03",X"CD",
		X"39",X"2F",X"CD",X"45",X"2C",X"CD",X"F0",X"32",X"CD",X"85",X"2C",X"CD",X"EC",X"2E",X"CD",X"B5",
		X"17",X"CD",X"B4",X"2B",X"CD",X"72",X"1A",X"CD",X"05",X"17",X"CD",X"01",X"0C",X"CD",X"1C",X"1C",
		X"CD",X"68",X"2A",X"CD",X"08",X"2C",X"CD",X"A9",X"0B",X"CD",X"CF",X"2E",X"CD",X"F3",X"05",X"CD",
		X"15",X"06",X"3A",X"6A",X"E0",X"0F",X"DC",X"59",X"06",X"CD",X"F8",X"1E",X"CD",X"39",X"1F",X"2A",
		X"83",X"E2",X"23",X"22",X"83",X"E2",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"00",
		X"65",X"00",X"F0",X"67",X"09",X"00",X"64",X"10",X"00",X"66",X"F0",X"00",X"6D",X"00",X"F0",X"6F",
		X"00",X"00",X"6C",X"10",X"08",X"6E",X"F6",X"00",X"71",X"00",X"FB",X"73",X"0A",X"FB",X"72",X"FA",
		X"08",X"70",X"FA",X"00",X"6A",X"00",X"F0",X"69",X"00",X"10",X"6B",X"00",X"F6",X"68",X"F0",X"00",
		X"74",X"00",X"F0",X"76",X"00",X"00",X"75",X"F0",X"0C",X"77",X"06",X"00",X"79",X"00",X"F0",X"7B",
		X"F3",X"00",X"7A",X"F0",X"06",X"78",X"0B",X"00",X"65",X"00",X"F0",X"67",X"09",X"00",X"64",X"10",
		X"00",X"66",X"F0",X"00",X"6D",X"00",X"F0",X"6F",X"00",X"00",X"6C",X"10",X"08",X"6E",X"F6",X"00",
		X"71",X"00",X"FB",X"73",X"0A",X"FB",X"72",X"FA",X"08",X"70",X"FA",X"00",X"6A",X"00",X"F0",X"69",
		X"00",X"10",X"6B",X"00",X"F6",X"68",X"F0",X"00",X"74",X"00",X"F0",X"76",X"00",X"00",X"75",X"F0",
		X"0C",X"77",X"06",X"00",X"79",X"00",X"F0",X"7B",X"F3",X"00",X"7A",X"F0",X"06",X"78",X"0B",X"0E",
		X"14",X"0C",X"0F",X"0B",X"0A",X"0B",X"09",X"09",X"06",X"08",X"05",X"08",X"04",X"07",X"02",X"06",
		X"01",X"05",X"00",X"06",X"00",X"05",X"FF",X"07",X"FE",X"0A",X"FC",X"0A",X"FB",X"08",X"FA",X"0B",
		X"F7",X"0A",X"F6",X"0C",X"F1",X"0D",X"E6",X"B3",X"B1",X"AF",X"AD",X"A9",X"A9",X"A9",X"A9",X"B2",
		X"B0",X"AE",X"AC",X"A9",X"A9",X"A9",X"A9",X"EF",X"ED",X"E7",X"E5",X"E9",X"E9",X"E9",X"E9",X"EE",
		X"EC",X"E6",X"E4",X"E9",X"E9",X"E9",X"E9",X"BD",X"BE",X"BF",X"C0",X"E1",X"E1",X"E1",X"E1",X"C4",
		X"D5",X"CF",X"C2",X"E1",X"E1",X"E1",X"E1",X"BE",X"D4",X"CE",X"BD",X"E1",X"E1",X"E1",X"E1",X"BD",
		X"BF",X"BE",X"BF",X"E1",X"E1",X"E1",X"E1",X"BE",X"BF",X"BC",X"BE",X"E1",X"E1",X"E1",X"E1",X"CB",
		X"C9",X"D6",X"C3",X"E1",X"E1",X"E1",X"E1",X"CA",X"C8",X"CD",X"CC",X"E1",X"E1",X"E1",X"E1",X"C0",
		X"C1",X"C3",X"BD",X"E1",X"E1",X"E1",X"E1",X"08",X"09",X"0A",X"0B",X"84",X"84",X"84",X"84",X"0A",
		X"D3",X"D1",X"08",X"94",X"EB",X"EB",X"94",X"08",X"D2",X"D0",X"08",X"84",X"EB",X"EB",X"94",X"0B",
		X"08",X"0A",X"09",X"94",X"84",X"94",X"94",X"63",X"63",X"99",X"63",X"01",X"01",X"01",X"01",X"99",
		X"17",X"15",X"74",X"01",X"28",X"28",X"01",X"63",X"16",X"14",X"99",X"01",X"28",X"28",X"01",X"99",
		X"74",X"63",X"74",X"01",X"01",X"01",X"01",X"08",X"09",X"0A",X"0B",X"84",X"84",X"84",X"84",X"0A",
		X"17",X"15",X"0B",X"84",X"28",X"28",X"84",X"09",X"16",X"14",X"0A",X"84",X"28",X"28",X"84",X"0B",
		X"09",X"08",X"0A",X"84",X"84",X"84",X"84",X"2D",X"2D",X"2D",X"2D",X"94",X"94",X"94",X"94",X"2D",
		X"2F",X"2F",X"2D",X"94",X"D6",X"C6",X"94",X"2D",X"2F",X"2F",X"2D",X"94",X"F6",X"E6",X"94",X"2D",
		X"2D",X"2D",X"2D",X"94",X"94",X"94",X"94",X"D8",X"DA",X"DA",X"D8",X"D7",X"D7",X"C7",X"C7",X"D9",
		X"DB",X"DB",X"D9",X"D7",X"D7",X"C7",X"C7",X"D9",X"DB",X"DB",X"D9",X"F7",X"F7",X"E7",X"E7",X"D8",
		X"DA",X"DA",X"D8",X"F7",X"F7",X"E7",X"E7",X"DC",X"DE",X"DE",X"DC",X"D7",X"D7",X"C7",X"C7",X"DD",
		X"DF",X"DF",X"DD",X"D7",X"D7",X"C7",X"C7",X"DD",X"DF",X"DF",X"DD",X"F7",X"F7",X"E7",X"E7",X"DC",
		X"DE",X"DE",X"DC",X"F7",X"F7",X"E7",X"E7",X"EA",X"E8",X"E2",X"E0",X"C9",X"C9",X"C9",X"C9",X"EB",
		X"E9",X"E3",X"E1",X"C9",X"C9",X"C9",X"C9",X"EB",X"E9",X"E3",X"E1",X"E9",X"E9",X"E9",X"E9",X"EA",
		X"E8",X"E2",X"E0",X"E9",X"E9",X"E9",X"E9",X"22",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"48",
		X"48",X"48",X"48",X"48",X"48",X"48",X"20",X"48",X"4E",X"4C",X"46",X"44",X"4F",X"4D",X"47",X"45",
		X"4A",X"48",X"92",X"90",X"8A",X"88",X"48",X"48",X"B7",X"B5",X"3F",X"A1",X"50",X"52",X"3F",X"3E",
		X"3E",X"48",X"93",X"91",X"8B",X"89",X"48",X"48",X"42",X"40",X"3F",X"3F",X"43",X"41",X"48",X"48",
		X"48",X"48",X"96",X"94",X"8E",X"8C",X"48",X"48",X"9A",X"98",X"56",X"54",X"48",X"48",X"48",X"48",
		X"48",X"48",X"97",X"95",X"8F",X"8D",X"48",X"48",X"9B",X"99",X"57",X"55",X"00",X"00",X"00",X"00",
		X"00",X"48",X"3F",X"3F",X"3F",X"3F",X"48",X"48",X"9E",X"9C",X"5A",X"58",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"48",X"3C",X"3D",X"3D",X"3C",X"48",X"48",X"9F",X"9D",X"5B",X"59",X"53",X"51",X"4B",X"49",
		X"48",X"48",X"3C",X"3D",X"3D",X"3C",X"48",X"48",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"AA",X"A8",X"A6",X"A4",X"A2",X"48",X"23",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"48",
		X"48",X"AB",X"A9",X"A7",X"A5",X"A3",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"63",X"E0",X"FE",X"02",X"D0",X"CD",X"5C",X"33",X"CD",X"6F",X"39",X"CD",X"9B",X"43",X"CD",
		X"5D",X"48",X"CD",X"06",X"33",X"C9",X"3A",X"B6",X"E5",X"A7",X"C0",X"DD",X"21",X"A8",X"E1",X"CD",
		X"46",X"33",X"DD",X"21",X"08",X"E2",X"CD",X"46",X"33",X"DD",X"21",X"68",X"E2",X"CD",X"46",X"33",
		X"DD",X"21",X"D8",X"E1",X"CD",X"46",X"33",X"DD",X"21",X"F0",X"E1",X"01",X"04",X"02",X"CD",X"48",
		X"33",X"DD",X"21",X"F8",X"E1",X"01",X"04",X"02",X"CD",X"48",X"33",X"DD",X"21",X"00",X"E2",X"01",
		X"04",X"02",X"CD",X"48",X"33",X"C9",X"0E",X"0C",X"CD",X"8C",X"35",X"C0",X"41",X"CD",X"51",X"33",
		X"C9",X"DD",X"36",X"00",X"00",X"DD",X"23",X"DD",X"23",X"10",X"F6",X"C9",X"3A",X"83",X"E2",X"E6",
		X"03",X"C0",X"3A",X"B6",X"E5",X"A7",X"C0",X"DD",X"21",X"A8",X"E1",X"FD",X"21",X"00",X"E5",X"CD",
		X"8D",X"33",X"DD",X"21",X"08",X"E2",X"FD",X"21",X"10",X"E5",X"CD",X"8D",X"33",X"DD",X"21",X"68",
		X"E2",X"FD",X"21",X"20",X"E5",X"CD",X"8D",X"33",X"AF",X"32",X"A0",X"E5",X"C9",X"3A",X"C6",X"E2",
		X"A7",X"C2",X"F0",X"33",X"3A",X"B0",X"E2",X"A7",X"C2",X"F0",X"33",X"3A",X"A6",X"E2",X"A7",X"C2",
		X"F0",X"33",X"FD",X"7E",X"01",X"A7",X"CA",X"DB",X"33",X"CD",X"8C",X"35",X"CC",X"9D",X"35",X"DD",
		X"E5",X"FD",X"E5",X"CD",X"A5",X"38",X"FD",X"E1",X"DD",X"E1",X"CD",X"F8",X"38",X"CD",X"3F",X"39",
		X"AF",X"32",X"BD",X"E5",X"CD",X"18",X"34",X"CD",X"FD",X"34",X"CD",X"1D",X"37",X"CD",X"5B",X"37",
		X"CD",X"64",X"38",X"3A",X"A0",X"E5",X"3C",X"32",X"A0",X"E5",X"C9",X"CD",X"8C",X"35",X"CA",X"AC",
		X"33",X"CD",X"EB",X"34",X"CD",X"1D",X"37",X"CD",X"19",X"38",X"CD",X"64",X"38",X"C3",X"D3",X"33",
		X"FD",X"7E",X"01",X"A7",X"C2",X"03",X"34",X"CD",X"1D",X"37",X"CD",X"19",X"38",X"CD",X"64",X"38",
		X"C3",X"D3",X"33",X"FD",X"36",X"01",X"0B",X"06",X"00",X"CD",X"18",X"34",X"CD",X"1D",X"37",X"CD",
		X"5B",X"37",X"CD",X"64",X"38",X"C3",X"D3",X"33",X"CD",X"EB",X"1F",X"FD",X"86",X"00",X"FD",X"77",
		X"00",X"FD",X"7E",X"01",X"FE",X"F0",X"DA",X"2D",X"34",X"FD",X"36",X"01",X"02",X"A7",X"CA",X"EB",
		X"34",X"3A",X"82",X"E2",X"47",X"FD",X"7E",X"01",X"B8",X"C2",X"8A",X"34",X"3A",X"BD",X"E5",X"A7",
		X"CA",X"54",X"34",X"FE",X"01",X"C2",X"4E",X"34",X"FD",X"35",X"01",X"C3",X"C9",X"34",X"FD",X"34",
		X"01",X"C3",X"C9",X"34",X"CD",X"1F",X"10",X"3A",X"8A",X"E0",X"CA",X"60",X"34",X"3A",X"8B",X"E0",
		X"FE",X"04",X"D2",X"66",X"34",X"3C",X"FD",X"86",X"01",X"FE",X"0F",X"D2",X"71",X"34",X"FD",X"77",
		X"01",X"3A",X"82",X"E2",X"FE",X"09",X"DA",X"C9",X"34",X"FD",X"7E",X"00",X"CD",X"EB",X"1F",X"FE",
		X"0C",X"D2",X"C9",X"34",X"FD",X"35",X"01",X"C3",X"C9",X"34",X"3A",X"BD",X"E5",X"A7",X"C2",X"C9",
		X"34",X"FD",X"7E",X"04",X"FE",X"01",X"C2",X"C9",X"34",X"DD",X"7E",X"03",X"FE",X"1E",X"DA",X"C9",
		X"34",X"3A",X"82",X"E2",X"FE",X"05",X"D2",X"B5",X"34",X"FD",X"7E",X"01",X"3C",X"FE",X"0F",X"D2",
		X"C9",X"34",X"FD",X"77",X"01",X"3A",X"82",X"E2",X"FE",X"09",X"D2",X"C9",X"34",X"FD",X"7E",X"01",
		X"3C",X"FE",X"0F",X"D2",X"C9",X"34",X"FD",X"77",X"01",X"FD",X"7E",X"01",X"90",X"FD",X"66",X"04",
		X"FD",X"6E",X"05",X"D2",X"E0",X"34",X"ED",X"44",X"06",X"00",X"4F",X"ED",X"42",X"C3",X"E4",X"34",
		X"06",X"00",X"4F",X"09",X"FD",X"74",X"04",X"FD",X"75",X"05",X"C9",X"01",X"0D",X"00",X"FD",X"66",
		X"04",X"FD",X"6E",X"05",X"ED",X"42",X"FD",X"74",X"04",X"FD",X"75",X"05",X"C9",X"DD",X"7E",X"00",
		X"FE",X"40",X"D8",X"FE",X"FA",X"D0",X"CD",X"1F",X"10",X"3A",X"82",X"E0",X"47",X"3A",X"89",X"E2",
		X"CA",X"1A",X"35",X"3A",X"83",X"E0",X"47",X"3A",X"8A",X"E2",X"80",X"FE",X"03",X"D8",X"FD",X"7E",
		X"02",X"A7",X"C2",X"44",X"35",X"3A",X"C0",X"E1",X"DD",X"46",X"00",X"B8",X"D2",X"3A",X"35",X"CD",
		X"EB",X"1F",X"E6",X"07",X"FD",X"77",X"02",X"C3",X"44",X"35",X"CD",X"EB",X"1F",X"E6",X"07",X"C6",
		X"F0",X"FD",X"77",X"02",X"FD",X"7E",X"02",X"FE",X"10",X"D2",X"55",X"35",X"DD",X"35",X"00",X"FD",
		X"35",X"02",X"C3",X"5E",X"35",X"FE",X"F0",X"D8",X"DD",X"34",X"00",X"FD",X"34",X"02",X"3A",X"A0",
		X"E5",X"FE",X"01",X"DA",X"77",X"35",X"CA",X"70",X"35",X"06",X"C4",X"0E",X"D8",X"C3",X"7B",X"35",
		X"06",X"84",X"0E",X"9C",X"C3",X"7B",X"35",X"06",X"48",X"0E",X"5C",X"DD",X"7E",X"00",X"B8",X"D2",
		X"86",X"35",X"DD",X"34",X"00",X"C9",X"B9",X"D8",X"DD",X"35",X"00",X"C9",X"06",X"06",X"AF",X"DD",
		X"E5",X"E1",X"23",X"23",X"11",X"04",X"00",X"B6",X"19",X"10",X"FC",X"A7",X"C9",X"3A",X"A7",X"E2",
		X"A7",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"C7",X"E5",X"FE",X"FF",X"28",X"22",X"3C",
		X"32",X"C7",X"E5",X"CD",X"1F",X"10",X"21",X"55",X"E0",X"28",X"02",X"2E",X"5E",X"06",X"F0",X"37",
		X"7E",X"2B",X"CB",X"18",X"A7",X"28",X"F9",X"80",X"47",X"CD",X"EB",X"1F",X"3A",X"69",X"E0",X"B8",
		X"D0",X"3A",X"7E",X"E0",X"06",X"02",X"3D",X"28",X"19",X"06",X"00",X"3D",X"28",X"14",X"3D",X"C8",
		X"3D",X"28",X"07",X"3A",X"AF",X"E5",X"A7",X"C0",X"18",X"0D",X"3A",X"A0",X"E5",X"FE",X"01",X"C0",
		X"18",X"05",X"3A",X"A0",X"E5",X"B8",X"C8",X"FD",X"36",X"0A",X"0F",X"FD",X"36",X"02",X"00",X"FD",
		X"36",X"0C",X"00",X"3A",X"C0",X"E5",X"A7",X"C0",X"18",X"11",X"3A",X"B9",X"E5",X"3C",X"FE",X"05",
		X"38",X"01",X"AF",X"32",X"B9",X"E5",X"87",X"FD",X"77",X"03",X"C9",X"3A",X"A0",X"E5",X"47",X"04",
		X"3E",X"20",X"0E",X"38",X"81",X"10",X"FD",X"DD",X"77",X"00",X"3A",X"96",X"E2",X"A7",X"3E",X"08",
		X"20",X"05",X"CD",X"E1",X"36",X"A7",X"C8",X"FD",X"77",X"01",X"47",X"3A",X"82",X"E2",X"90",X"38",
		X"25",X"3A",X"C7",X"E5",X"FE",X"0F",X"D8",X"11",X"D0",X"01",X"CD",X"8B",X"36",X"C0",X"CD",X"C5",
		X"36",X"C8",X"CD",X"0A",X"36",X"FD",X"36",X"04",X"01",X"FD",X"36",X"05",X"F8",X"FD",X"36",X"0C",
		X"01",X"AF",X"32",X"C7",X"E5",X"C9",X"3A",X"C7",X"E5",X"FE",X"40",X"D8",X"11",X"D0",X"00",X"CD",
		X"8B",X"36",X"C0",X"CD",X"C5",X"36",X"C8",X"CD",X"0A",X"36",X"FD",X"36",X"04",X"00",X"FD",X"36",
		X"05",X"D8",X"FD",X"36",X"0C",X"01",X"AF",X"32",X"C7",X"E5",X"C9",X"AF",X"32",X"AA",X"E5",X"FD",
		X"E5",X"FD",X"21",X"30",X"E5",X"CD",X"AD",X"36",X"FD",X"21",X"40",X"E5",X"CD",X"AD",X"36",X"FD",
		X"21",X"50",X"E5",X"CD",X"AD",X"36",X"FD",X"E1",X"3A",X"AA",X"E5",X"A7",X"C9",X"FD",X"66",X"04",
		X"FD",X"6E",X"05",X"ED",X"52",X"D8",X"7C",X"A7",X"C0",X"7D",X"FE",X"60",X"D0",X"3A",X"AA",X"E5",
		X"3C",X"32",X"AA",X"E5",X"C9",X"3A",X"68",X"E5",X"FE",X"01",X"C0",X"DD",X"36",X"00",X"00",X"A7",
		X"C9",X"3A",X"82",X"E2",X"47",X"CD",X"EB",X"1F",X"E6",X"03",X"D6",X"02",X"38",X"01",X"3C",X"80",
		X"C9",X"3A",X"82",X"E2",X"4F",X"FE",X"0A",X"30",X"1C",X"3A",X"C1",X"E5",X"A7",X"C8",X"CD",X"1F",
		X"10",X"3A",X"8A",X"E0",X"28",X"03",X"3A",X"8B",X"E0",X"FE",X"04",X"38",X"02",X"3E",X"03",X"47",
		X"79",X"C6",X"02",X"80",X"C9",X"3A",X"C6",X"E5",X"3C",X"E6",X"03",X"32",X"C6",X"E5",X"21",X"19",
		X"37",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",X"C9",X"03",X"06",X"04",X"05",X"DD",X"7E",X"00",
		X"DD",X"77",X"08",X"DD",X"77",X"10",X"C6",X"10",X"DD",X"77",X"04",X"DD",X"77",X"0C",X"DD",X"77",
		X"14",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"01",X"10",X"00",X"DD",X"75",X"03",X"DD",X"75",X"07",
		X"09",X"FD",X"74",X"06",X"FD",X"75",X"07",X"DD",X"75",X"0B",X"DD",X"75",X"0F",X"09",X"FD",X"74",
		X"08",X"FD",X"75",X"09",X"DD",X"75",X"13",X"DD",X"75",X"17",X"C9",X"21",X"8D",X"37",X"FD",X"7E",
		X"03",X"3C",X"CB",X"47",X"20",X"02",X"D6",X"02",X"FD",X"77",X"03",X"CB",X"27",X"06",X"00",X"4F",
		X"09",X"5E",X"23",X"56",X"EB",X"DD",X"E5",X"06",X"06",X"11",X"04",X"00",X"7E",X"DD",X"77",X"01",
		X"23",X"7E",X"DD",X"77",X"02",X"23",X"DD",X"19",X"10",X"F2",X"DD",X"E1",X"C9",X"A1",X"37",X"AD",
		X"37",X"B9",X"37",X"C5",X"37",X"D1",X"37",X"DD",X"37",X"E9",X"37",X"F5",X"37",X"01",X"38",X"0D",
		X"38",X"C0",X"2A",X"40",X"2A",X"C0",X"29",X"40",X"29",X"C0",X"28",X"40",X"28",X"C0",X"3C",X"40",
		X"3C",X"C0",X"3B",X"40",X"3B",X"C0",X"3A",X"40",X"3A",X"C0",X"33",X"40",X"33",X"C0",X"32",X"40",
		X"32",X"C0",X"31",X"40",X"31",X"C0",X"45",X"40",X"45",X"C0",X"44",X"40",X"44",X"C0",X"43",X"40",
		X"43",X"C4",X"39",X"44",X"39",X"C4",X"38",X"44",X"38",X"C4",X"37",X"44",X"37",X"C4",X"4B",X"44",
		X"4B",X"C4",X"4A",X"44",X"4A",X"C4",X"49",X"44",X"49",X"C6",X"36",X"46",X"36",X"C6",X"35",X"46",
		X"35",X"C6",X"34",X"46",X"34",X"C6",X"48",X"46",X"48",X"C6",X"47",X"46",X"47",X"C6",X"46",X"46",
		X"46",X"40",X"2F",X"40",X"2D",X"40",X"40",X"40",X"2C",X"40",X"30",X"40",X"2B",X"40",X"41",X"40",
		X"3F",X"40",X"40",X"40",X"2C",X"40",X"42",X"40",X"3D",X"FD",X"34",X"0D",X"FD",X"7E",X"0D",X"CB",
		X"47",X"C2",X"3E",X"38",X"21",X"58",X"38",X"11",X"04",X"00",X"DD",X"E5",X"06",X"06",X"7E",X"DD",
		X"36",X"01",X"40",X"DD",X"77",X"02",X"23",X"DD",X"19",X"10",X"F3",X"DD",X"E1",X"C9",X"21",X"5E",
		X"38",X"11",X"04",X"00",X"DD",X"E5",X"06",X"06",X"7E",X"DD",X"36",X"01",X"40",X"DD",X"77",X"02",
		X"23",X"DD",X"19",X"10",X"F3",X"DD",X"E1",X"C9",X"00",X"00",X"88",X"86",X"87",X"85",X"00",X"00",
		X"8C",X"8A",X"8B",X"89",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"01",X"08",X"00",X"09",X"7C",X"FE",
		X"01",X"CA",X"7C",X"38",X"DD",X"36",X"02",X"00",X"DD",X"36",X"06",X"00",X"FD",X"66",X"06",X"FD",
		X"6E",X"07",X"09",X"7C",X"FE",X"01",X"CA",X"91",X"38",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0E",
		X"00",X"FD",X"66",X"08",X"FD",X"6E",X"09",X"09",X"7C",X"FE",X"01",X"C8",X"DD",X"36",X"12",X"00",
		X"DD",X"36",X"16",X"00",X"C9",X"3A",X"96",X"E2",X"A7",X"C0",X"FD",X"21",X"A8",X"E1",X"CD",X"BC",
		X"38",X"FD",X"21",X"08",X"E2",X"CD",X"BC",X"38",X"FD",X"21",X"68",X"E2",X"CD",X"40",X"03",X"4F",
		X"A7",X"C8",X"3A",X"96",X"E2",X"81",X"32",X"96",X"E2",X"3E",X"02",X"32",X"A7",X"E5",X"FD",X"7E",
		X"00",X"32",X"AA",X"E2",X"FD",X"7E",X"03",X"32",X"AB",X"E2",X"C9",X"FD",X"36",X"01",X"00",X"3E",
		X"18",X"D7",X"FD",X"7E",X"0E",X"A7",X"C8",X"FD",X"7E",X"0F",X"FE",X"02",X"D0",X"FD",X"7E",X"03",
		X"3C",X"32",X"BE",X"E5",X"FD",X"34",X"0F",X"C9",X"AF",X"32",X"A8",X"E5",X"FD",X"7E",X"0A",X"A7",
		X"C8",X"FD",X"E5",X"FD",X"21",X"C0",X"E1",X"CD",X"1C",X"39",X"FD",X"E1",X"3A",X"A8",X"E5",X"A7",
		X"C8",X"FD",X"35",X"01",X"FD",X"35",X"01",X"FD",X"36",X"0A",X"00",X"C9",X"0E",X"00",X"DD",X"7E",
		X"00",X"D6",X"08",X"47",X"FD",X"7E",X"00",X"90",X"D8",X"FE",X"20",X"D0",X"FD",X"7E",X"03",X"DD",
		X"96",X"03",X"D8",X"FE",X"48",X"D0",X"3A",X"A8",X"E5",X"C6",X"02",X"32",X"A8",X"E5",X"C9",X"DD",
		X"46",X"03",X"DD",X"36",X"03",X"E0",X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"70",X"03",
		X"30",X"04",X"FD",X"36",X"01",X"01",X"DD",X"7E",X"03",X"47",X"C6",X"30",X"DD",X"77",X"03",X"FD",
		X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"70",X"03",X"D0",X"FD",X"36",X"01",X"00",X"C9",X"3A",
		X"83",X"E2",X"E6",X"03",X"FE",X"01",X"C0",X"DD",X"21",X"F0",X"E1",X"FD",X"21",X"30",X"E5",X"CD",
		X"99",X"39",X"DD",X"21",X"F8",X"E1",X"FD",X"21",X"40",X"E5",X"CD",X"99",X"39",X"DD",X"21",X"00",
		X"E2",X"FD",X"21",X"50",X"E5",X"CD",X"99",X"39",X"C9",X"3A",X"C6",X"E2",X"A7",X"C2",X"1D",X"3A",
		X"3A",X"B0",X"E2",X"A7",X"C2",X"1D",X"3A",X"3A",X"A6",X"E2",X"A7",X"C2",X"1D",X"3A",X"FD",X"7E",
		X"01",X"A7",X"CA",X"03",X"3A",X"06",X"02",X"FD",X"34",X"0A",X"FD",X"7E",X"0A",X"FE",X"10",X"DA",
		X"C6",X"39",X"FD",X"36",X"0E",X"00",X"CD",X"8E",X"35",X"CC",X"4A",X"3A",X"CD",X"81",X"3B",X"CD",
		X"23",X"43",X"CD",X"F7",X"39",X"DD",X"E5",X"FD",X"E5",X"CD",X"58",X"40",X"FD",X"E1",X"DD",X"E1",
		X"3E",X"01",X"32",X"BD",X"E5",X"06",X"01",X"CD",X"18",X"34",X"CD",X"4E",X"3D",X"CD",X"18",X"3E",
		X"CD",X"F7",X"39",X"CD",X"6E",X"3F",X"C9",X"CD",X"FB",X"3D",X"CD",X"4B",X"3F",X"06",X"02",X"CD",
		X"27",X"3F",X"C9",X"06",X"02",X"CD",X"8E",X"35",X"CA",X"C9",X"39",X"CD",X"EB",X"34",X"CD",X"FB",
		X"3D",X"CD",X"C1",X"3E",X"CD",X"4B",X"3F",X"06",X"02",X"CD",X"27",X"3F",X"C9",X"FD",X"7E",X"01",
		X"A7",X"20",X"0F",X"CD",X"FB",X"3D",X"CD",X"C1",X"3E",X"CD",X"4B",X"3F",X"06",X"02",X"CD",X"27",
		X"3F",X"C9",X"FD",X"36",X"01",X"0B",X"06",X"00",X"CD",X"18",X"34",X"CD",X"18",X"3E",X"CD",X"FB",
		X"3D",X"CD",X"4B",X"3F",X"06",X"02",X"CD",X"27",X"3F",X"C9",X"AF",X"FD",X"77",X"08",X"FD",X"77",
		X"09",X"FD",X"77",X"0B",X"FD",X"77",X"0C",X"FD",X"77",X"0D",X"FD",X"77",X"0E",X"FD",X"77",X"0F",
		X"FD",X"7E",X"00",X"FE",X"B0",X"D8",X"3A",X"CA",X"E4",X"FE",X"FA",X"D0",X"CD",X"EB",X"1F",X"E6",
		X"07",X"FE",X"05",X"30",X"F7",X"FD",X"77",X"03",X"3A",X"7E",X"E0",X"CB",X"27",X"21",X"22",X"3B",
		X"06",X"00",X"4F",X"09",X"5E",X"23",X"56",X"EB",X"CD",X"EB",X"1F",X"E6",X"03",X"4F",X"06",X"00",
		X"09",X"7E",X"4F",X"3A",X"A3",X"E5",X"B9",X"C8",X"79",X"32",X"A3",X"E5",X"DD",X"77",X"00",X"3A",
		X"96",X"E2",X"A7",X"3E",X"09",X"C2",X"E8",X"3A",X"3A",X"C1",X"E5",X"A7",X"C8",X"3A",X"82",X"E2",
		X"FE",X"05",X"D2",X"BA",X"3A",X"C6",X"06",X"C3",X"E8",X"3A",X"FD",X"7E",X"03",X"FE",X"01",X"CA",
		X"DC",X"3A",X"FE",X"04",X"CA",X"DC",X"3A",X"FE",X"02",X"CA",X"E3",X"3A",X"CD",X"D1",X"36",X"47",
		X"3A",X"82",X"E2",X"B8",X"30",X"03",X"3D",X"18",X"0F",X"3C",X"18",X"0C",X"3A",X"82",X"E2",X"C6",
		X"02",X"18",X"05",X"3A",X"82",X"E2",X"D6",X"02",X"FD",X"77",X"01",X"47",X"3A",X"82",X"E2",X"90",
		X"38",X"18",X"11",X"D0",X"01",X"CD",X"40",X"3B",X"C0",X"DD",X"36",X"02",X"8E",X"DD",X"36",X"06",
		X"8D",X"FD",X"36",X"04",X"01",X"FD",X"36",X"05",X"F8",X"C9",X"11",X"D0",X"00",X"CD",X"40",X"3B",
		X"C0",X"DD",X"36",X"02",X"8E",X"DD",X"36",X"06",X"8D",X"FD",X"36",X"04",X"00",X"FD",X"36",X"05",
		X"E8",X"C9",X"2C",X"3B",X"30",X"3B",X"34",X"3B",X"38",X"3B",X"3C",X"3B",X"58",X"80",X"B0",X"D0",
		X"50",X"78",X"A0",X"78",X"90",X"B8",X"D0",X"B8",X"58",X"D0",X"D0",X"58",X"88",X"88",X"A8",X"A8",
		X"AF",X"32",X"A6",X"E5",X"FD",X"E5",X"FD",X"21",X"00",X"E5",X"CD",X"69",X"3B",X"FD",X"21",X"10",
		X"E5",X"CD",X"69",X"3B",X"FD",X"21",X"20",X"E5",X"CD",X"69",X"3B",X"FD",X"21",X"60",X"E5",X"CD",
		X"69",X"3B",X"FD",X"E1",X"3A",X"A6",X"E5",X"A7",X"C9",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"ED",
		X"52",X"D8",X"7C",X"A7",X"C0",X"7D",X"FE",X"60",X"D0",X"3A",X"A6",X"E5",X"3C",X"32",X"A6",X"E5",
		X"C9",X"FD",X"E5",X"AF",X"32",X"A2",X"E5",X"DD",X"7E",X"00",X"D6",X"10",X"DD",X"77",X"00",X"DD",
		X"7E",X"03",X"C6",X"20",X"DD",X"77",X"03",X"CD",X"FF",X"3B",X"79",X"A7",X"28",X"08",X"3A",X"A2",
		X"E5",X"CB",X"C7",X"32",X"A2",X"E5",X"DD",X"7E",X"03",X"D6",X"40",X"DD",X"77",X"03",X"CD",X"FF",
		X"3B",X"79",X"A7",X"28",X"08",X"3A",X"A2",X"E5",X"CB",X"CF",X"32",X"A2",X"E5",X"DD",X"7E",X"00",
		X"C6",X"20",X"DD",X"77",X"00",X"CD",X"FF",X"3B",X"79",X"A7",X"28",X"08",X"3A",X"A2",X"E5",X"CB",
		X"D7",X"32",X"A2",X"E5",X"DD",X"7E",X"03",X"C6",X"40",X"DD",X"77",X"03",X"CD",X"FF",X"3B",X"79",
		X"A7",X"28",X"08",X"3A",X"A2",X"E5",X"CB",X"DF",X"32",X"A2",X"E5",X"DD",X"7E",X"00",X"D6",X"10",
		X"DD",X"77",X"00",X"DD",X"7E",X"03",X"D6",X"20",X"DD",X"77",X"03",X"FD",X"E1",X"18",X"27",X"FD",
		X"21",X"A8",X"E1",X"06",X"03",X"0E",X"00",X"AF",X"DD",X"E5",X"CD",X"45",X"03",X"DD",X"E1",X"A7",
		X"28",X"01",X"0C",X"11",X"60",X"00",X"FD",X"19",X"10",X"ED",X"FD",X"21",X"D8",X"E1",X"AF",X"CD",
		X"45",X"03",X"A7",X"C8",X"0C",X"C9",X"DD",X"7E",X"00",X"FE",X"FA",X"D0",X"FE",X"38",X"D8",X"FD",
		X"36",X"02",X"00",X"3A",X"A2",X"E5",X"A7",X"28",X"15",X"CB",X"47",X"C2",X"C6",X"3C",X"CB",X"4F",
		X"C2",X"DD",X"3C",X"CB",X"57",X"C2",X"F4",X"3C",X"CB",X"5F",X"C2",X"0B",X"3D",X"C9",X"3A",X"B0",
		X"E2",X"A7",X"C0",X"3A",X"B8",X"E5",X"A7",X"C0",X"CD",X"1F",X"10",X"28",X"06",X"3A",X"8A",X"E2",
		X"C3",X"66",X"3C",X"3A",X"89",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",X"47",
		X"FD",X"7E",X"0B",X"B8",X"D0",X"FD",X"7E",X"03",X"FE",X"01",X"C8",X"FE",X"04",X"C8",X"3A",X"C4",
		X"E1",X"DD",X"4E",X"00",X"91",X"38",X"08",X"FE",X"08",X"D2",X"AC",X"3C",X"C3",X"C1",X"3C",X"FE",
		X"F8",X"DA",X"97",X"3C",X"C3",X"C1",X"3C",X"FD",X"7E",X"03",X"FE",X"03",X"CA",X"A4",X"3C",X"FD",
		X"36",X"02",X"10",X"C9",X"DD",X"35",X"00",X"FD",X"36",X"02",X"10",X"C9",X"FD",X"7E",X"03",X"FE",
		X"03",X"CA",X"B9",X"3C",X"FD",X"36",X"02",X"F0",X"C9",X"DD",X"34",X"00",X"FD",X"36",X"02",X"F0",
		X"C9",X"FD",X"36",X"02",X"00",X"C9",X"CB",X"57",X"C2",X"22",X"3D",X"CB",X"5F",X"C2",X"42",X"3D",
		X"DD",X"7E",X"00",X"C6",X"02",X"FE",X"D8",X"DA",X"39",X"3D",X"C3",X"42",X"3D",X"CB",X"5F",X"C2",
		X"22",X"3D",X"CB",X"57",X"C2",X"3E",X"3D",X"DD",X"7E",X"00",X"C6",X"02",X"FE",X"D8",X"DA",X"39",
		X"3D",X"C3",X"3E",X"3D",X"CB",X"47",X"C2",X"22",X"3D",X"CB",X"4F",X"C2",X"3E",X"3D",X"DD",X"7E",
		X"00",X"D6",X"02",X"FE",X"58",X"D2",X"34",X"3D",X"C3",X"3E",X"3D",X"CB",X"4F",X"C2",X"22",X"3D",
		X"CB",X"47",X"C2",X"42",X"3D",X"DD",X"7E",X"00",X"D6",X"02",X"FE",X"58",X"D2",X"34",X"3D",X"C3",
		X"42",X"3D",X"FD",X"36",X"02",X"00",X"CD",X"EB",X"1F",X"FE",X"0E",X"D2",X"3E",X"3D",X"FE",X"02",
		X"DA",X"42",X"3D",X"C9",X"FD",X"36",X"02",X"10",X"C9",X"FD",X"36",X"02",X"F0",X"C9",X"FD",X"34",
		X"01",X"C9",X"FD",X"35",X"01",X"FD",X"7E",X"01",X"A7",X"C0",X"FD",X"34",X"01",X"C9",X"DD",X"7E",
		X"00",X"FE",X"38",X"D8",X"FE",X"FA",X"D0",X"FD",X"7E",X"0D",X"A7",X"C2",X"C6",X"3D",X"FD",X"7E",
		X"02",X"A7",X"C8",X"FE",X"10",X"C2",X"96",X"3D",X"DD",X"7E",X"00",X"D6",X"03",X"FE",X"50",X"D8",
		X"FD",X"7E",X"03",X"FE",X"01",X"CA",X"85",X"3D",X"FE",X"03",X"D2",X"8D",X"3D",X"DD",X"7E",X"00",
		X"D6",X"02",X"C3",X"92",X"3D",X"DD",X"7E",X"00",X"D6",X"01",X"C3",X"92",X"3D",X"DD",X"7E",X"00",
		X"D6",X"03",X"DD",X"77",X"00",X"C9",X"FE",X"F0",X"C0",X"DD",X"7E",X"00",X"C6",X"03",X"FE",X"E0",
		X"D0",X"FD",X"7E",X"03",X"FE",X"01",X"CA",X"B6",X"3D",X"FE",X"03",X"D2",X"BD",X"3D",X"DD",X"7E",
		X"00",X"C6",X"02",X"C3",X"C2",X"3D",X"DD",X"7E",X"00",X"3C",X"C3",X"C2",X"3D",X"DD",X"7E",X"00",
		X"C6",X"03",X"DD",X"77",X"00",X"C9",X"FD",X"7E",X"0D",X"FE",X"10",X"DA",X"E2",X"3D",X"FE",X"F0",
		X"D8",X"DD",X"7E",X"00",X"C6",X"03",X"FE",X"F0",X"D2",X"F3",X"3D",X"DD",X"77",X"00",X"FD",X"34",
		X"0D",X"C9",X"DD",X"7E",X"00",X"D6",X"03",X"FE",X"40",X"DA",X"F3",X"3D",X"DD",X"77",X"00",X"FD",
		X"35",X"0D",X"C9",X"AF",X"FD",X"77",X"0D",X"CD",X"DB",X"38",X"C9",X"DD",X"7E",X"00",X"DD",X"77",
		X"04",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"01",X"10",X"00",X"DD",X"75",X"03",X"09",X"FD",X"74",
		X"06",X"FD",X"75",X"07",X"DD",X"75",X"07",X"C9",X"21",X"B9",X"3E",X"FD",X"7E",X"02",X"A7",X"CA",
		X"60",X"3E",X"FD",X"7E",X"0C",X"3C",X"FE",X"04",X"D2",X"40",X"3E",X"FD",X"77",X"0C",X"CB",X"27",
		X"06",X"00",X"4F",X"09",X"7E",X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"06",X"C3",X"89",X"3E",
		X"DD",X"7E",X"02",X"3C",X"3C",X"FE",X"98",X"C2",X"55",X"3E",X"DD",X"36",X"02",X"94",X"DD",X"36",
		X"06",X"93",X"C3",X"89",X"3E",X"DD",X"36",X"02",X"96",X"DD",X"36",X"06",X"95",X"C3",X"89",X"3E",
		X"FD",X"7E",X"0C",X"A7",X"CA",X"6E",X"3E",X"3D",X"FD",X"77",X"0C",X"C3",X"2E",X"3E",X"DD",X"7E",
		X"02",X"FE",X"8E",X"CA",X"81",X"3E",X"DD",X"36",X"02",X"8E",X"DD",X"36",X"06",X"8D",X"C3",X"89",
		X"3E",X"DD",X"36",X"02",X"98",X"DD",X"36",X"06",X"97",X"FD",X"7E",X"02",X"FE",X"10",X"CA",X"A5",
		X"3E",X"3E",X"C0",X"47",X"FD",X"7E",X"03",X"A7",X"C2",X"9D",X"3E",X"3E",X"08",X"80",X"DD",X"77",
		X"01",X"DD",X"77",X"05",X"C9",X"3E",X"40",X"47",X"FD",X"7E",X"03",X"A7",X"C2",X"B1",X"3E",X"3E",
		X"08",X"80",X"DD",X"77",X"01",X"DD",X"77",X"05",X"C9",X"8E",X"8D",X"90",X"8F",X"92",X"91",X"94",
		X"93",X"DD",X"36",X"01",X"40",X"DD",X"36",X"05",X"40",X"FD",X"34",X"08",X"FD",X"7E",X"08",X"FE",
		X"03",X"D2",X"EE",X"3E",X"FD",X"7E",X"08",X"CB",X"4F",X"CA",X"E5",X"3E",X"DD",X"36",X"02",X"82",
		X"DD",X"36",X"06",X"81",X"C9",X"DD",X"36",X"02",X"84",X"DD",X"36",X"06",X"83",X"C9",X"FE",X"10",
		X"D2",X"15",X"3F",X"FD",X"7E",X"0F",X"A7",X"CA",X"D4",X"3E",X"FD",X"7E",X"03",X"21",X"22",X"3F",
		X"06",X"00",X"4F",X"09",X"7E",X"DD",X"36",X"02",X"00",X"DD",X"77",X"06",X"FD",X"36",X"04",X"01",
		X"FD",X"36",X"05",X"40",X"C9",X"DD",X"36",X"02",X"00",X"DD",X"36",X"06",X"00",X"FD",X"36",X"04",
		X"00",X"C9",X"99",X"9E",X"FD",X"7D",X"7E",X"DD",X"E5",X"DD",X"7E",X"00",X"CD",X"9E",X"1E",X"DD",
		X"7E",X"01",X"CD",X"A8",X"1E",X"DD",X"7E",X"02",X"CD",X"B2",X"1E",X"DD",X"7E",X"03",X"CD",X"BC",
		X"1E",X"11",X"04",X"00",X"DD",X"19",X"10",X"E1",X"DD",X"E1",X"C9",X"FD",X"66",X"04",X"FD",X"6E",
		X"05",X"01",X"08",X"00",X"09",X"7C",X"FE",X"01",X"28",X"04",X"DD",X"36",X"02",X"00",X"FD",X"66",
		X"06",X"FD",X"6E",X"07",X"09",X"7C",X"FE",X"01",X"C8",X"DD",X"36",X"06",X"00",X"C9",X"DD",X"7E",
		X"00",X"FE",X"40",X"D8",X"FE",X"FA",X"D0",X"DD",X"7E",X"02",X"DD",X"86",X"06",X"A7",X"C8",X"AF",
		X"32",X"A9",X"E5",X"FD",X"E5",X"FD",X"21",X"A8",X"E1",X"CD",X"CF",X"3F",X"FD",X"E1",X"CD",X"AE",
		X"3F",X"FD",X"E5",X"FD",X"21",X"08",X"E2",X"CD",X"CF",X"3F",X"FD",X"E1",X"CD",X"AE",X"3F",X"FD",
		X"E5",X"FD",X"21",X"68",X"E2",X"CD",X"CF",X"3F",X"FD",X"E1",X"CD",X"AE",X"3F",X"C9",X"3A",X"A4",
		X"E5",X"A7",X"CA",X"BB",X"3F",X"3A",X"A5",X"E5",X"FD",X"77",X"01",X"3A",X"B0",X"E5",X"A7",X"C8",
		X"D5",X"E1",X"01",X"01",X"E5",X"ED",X"42",X"D8",X"3E",X"01",X"12",X"CD",X"DB",X"38",X"C9",X"AF",
		X"32",X"A4",X"E5",X"32",X"B0",X"E5",X"32",X"AB",X"E5",X"DD",X"7E",X"03",X"FE",X"C0",X"DA",X"EE",
		X"3F",X"FD",X"7E",X"03",X"D6",X"20",X"FD",X"77",X"03",X"3E",X"0F",X"32",X"AB",X"E5",X"DD",X"7E",
		X"03",X"C6",X"20",X"DD",X"77",X"03",X"AF",X"CD",X"45",X"03",X"A7",X"C4",X"3B",X"40",X"DD",X"7E",
		X"03",X"D6",X"40",X"DD",X"77",X"03",X"AF",X"CD",X"45",X"03",X"A7",X"C4",X"3B",X"40",X"DD",X"7E",
		X"03",X"C6",X"20",X"DD",X"77",X"03",X"AF",X"CD",X"45",X"03",X"A7",X"CA",X"25",X"40",X"3A",X"B0",
		X"E5",X"3C",X"32",X"B0",X"E5",X"3A",X"A9",X"E5",X"C6",X"02",X"32",X"A9",X"E5",X"3A",X"AB",X"E5",
		X"A7",X"C8",X"FD",X"7E",X"03",X"C6",X"20",X"FD",X"77",X"03",X"C9",X"3A",X"A9",X"E5",X"21",X"52",
		X"40",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"1A",X"32",X"A5",X"E5",X"3E",X"0F",X"32",X"A4",
		X"E5",X"C9",X"01",X"E5",X"11",X"E5",X"21",X"E5",X"DD",X"21",X"F0",X"E1",X"FD",X"21",X"F8",X"E1",
		X"CD",X"C8",X"40",X"C4",X"28",X"41",X"DD",X"21",X"F0",X"E1",X"FD",X"21",X"00",X"E2",X"CD",X"C8",
		X"40",X"C4",X"4A",X"41",X"DD",X"21",X"F8",X"E1",X"FD",X"21",X"00",X"E2",X"CD",X"C8",X"40",X"C4",
		X"6C",X"41",X"3A",X"A6",X"E2",X"A7",X"C0",X"3A",X"96",X"E2",X"A7",X"C0",X"3A",X"B0",X"E2",X"A7",
		X"C0",X"DD",X"21",X"C0",X"E1",X"FD",X"21",X"F0",X"E1",X"CD",X"C8",X"40",X"C4",X"CA",X"42",X"C4",
		X"8E",X"41",X"DD",X"21",X"C0",X"E1",X"FD",X"21",X"F8",X"E1",X"CD",X"C8",X"40",X"C4",X"CA",X"42",
		X"C4",X"B7",X"41",X"DD",X"21",X"C0",X"E1",X"FD",X"21",X"00",X"E2",X"CD",X"C8",X"40",X"C4",X"CA",
		X"42",X"C4",X"E0",X"41",X"3E",X"F0",X"A7",X"C9",X"AF",X"32",X"AE",X"E5",X"32",X"AD",X"E5",X"DD",
		X"7E",X"02",X"FE",X"82",X"C8",X"FE",X"84",X"C8",X"DD",X"86",X"06",X"A7",X"C8",X"FD",X"7E",X"02",
		X"FE",X"82",X"C8",X"FE",X"84",X"C8",X"FD",X"86",X"06",X"A7",X"C8",X"3E",X"01",X"CD",X"45",X"03",
		X"A7",X"C8",X"DD",X"7E",X"03",X"FD",X"46",X"03",X"CD",X"08",X"41",X"DD",X"7E",X"00",X"FD",X"46",
		X"00",X"CD",X"18",X"41",X"3E",X"FF",X"A7",X"C9",X"90",X"D2",X"12",X"41",X"3E",X"10",X"32",X"AD",
		X"E5",X"C9",X"3E",X"F0",X"32",X"AD",X"E5",X"C9",X"90",X"D2",X"22",X"41",X"3E",X"10",X"32",X"AE",
		X"E5",X"C9",X"3E",X"F0",X"32",X"AE",X"E5",X"C9",X"DD",X"21",X"F0",X"E1",X"FD",X"21",X"30",X"E5",
		X"CD",X"09",X"42",X"DD",X"21",X"F8",X"E1",X"FD",X"21",X"40",X"E5",X"CD",X"6B",X"42",X"DD",X"21",
		X"30",X"E5",X"FD",X"21",X"40",X"E5",X"CD",X"F9",X"42",X"C9",X"DD",X"21",X"F0",X"E1",X"FD",X"21",
		X"30",X"E5",X"CD",X"09",X"42",X"DD",X"21",X"00",X"E2",X"FD",X"21",X"50",X"E5",X"CD",X"6B",X"42",
		X"DD",X"21",X"30",X"E5",X"FD",X"21",X"50",X"E5",X"CD",X"F9",X"42",X"C9",X"DD",X"21",X"F8",X"E1",
		X"FD",X"21",X"40",X"E5",X"CD",X"09",X"42",X"DD",X"21",X"00",X"E2",X"FD",X"21",X"50",X"E5",X"CD",
		X"6B",X"42",X"DD",X"21",X"40",X"E5",X"DD",X"21",X"50",X"E5",X"CD",X"F9",X"42",X"C9",X"DD",X"21",
		X"F0",X"E1",X"FD",X"21",X"30",X"E5",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"0E",X"01",X"FD",X"34",
		X"0B",X"06",X"03",X"3A",X"A7",X"E2",X"A7",X"CA",X"AC",X"41",X"06",X"01",X"FD",X"7E",X"0B",X"B8",
		X"D2",X"EA",X"42",X"CD",X"6B",X"42",X"C9",X"DD",X"21",X"F8",X"E1",X"FD",X"21",X"40",X"E5",X"FD",
		X"36",X"0A",X"00",X"FD",X"36",X"0E",X"01",X"FD",X"34",X"0B",X"06",X"03",X"3A",X"A7",X"E2",X"A7",
		X"CA",X"D5",X"41",X"06",X"01",X"FD",X"7E",X"0B",X"B8",X"D2",X"EA",X"42",X"CD",X"6B",X"42",X"C9",
		X"DD",X"21",X"00",X"E2",X"FD",X"21",X"50",X"E5",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"0E",X"01",
		X"FD",X"34",X"0B",X"06",X"03",X"3A",X"A7",X"E2",X"A7",X"CA",X"FE",X"41",X"06",X"01",X"FD",X"7E",
		X"0B",X"B8",X"D2",X"EA",X"42",X"CD",X"6B",X"42",X"C9",X"0E",X"06",X"3A",X"AE",X"E5",X"A7",X"CA",
		X"33",X"42",X"FE",X"10",X"CA",X"28",X"42",X"79",X"ED",X"44",X"FD",X"77",X"0D",X"DD",X"7E",X"00",
		X"C6",X"08",X"DD",X"77",X"00",X"C3",X"33",X"42",X"FD",X"71",X"0D",X"DD",X"7E",X"00",X"D6",X"08",
		X"DD",X"77",X"00",X"3A",X"AD",X"E5",X"A7",X"C8",X"FE",X"10",X"CA",X"4E",X"42",X"FD",X"66",X"04",
		X"FD",X"6E",X"05",X"01",X"08",X"00",X"09",X"FD",X"74",X"04",X"FD",X"75",X"05",X"C9",X"FD",X"66",
		X"04",X"FD",X"6E",X"05",X"01",X"08",X"00",X"ED",X"42",X"FD",X"74",X"04",X"FD",X"75",X"05",X"FD",
		X"35",X"01",X"FD",X"7E",X"01",X"A7",X"C0",X"FD",X"34",X"01",X"C9",X"0E",X"06",X"3A",X"AE",X"E5",
		X"A7",X"CA",X"95",X"42",X"FE",X"10",X"CA",X"87",X"42",X"FD",X"71",X"0D",X"DD",X"7E",X"00",X"D6",
		X"08",X"DD",X"77",X"00",X"C3",X"95",X"42",X"79",X"ED",X"44",X"FD",X"77",X"0D",X"DD",X"7E",X"00",
		X"C6",X"08",X"DD",X"77",X"00",X"3A",X"AD",X"E5",X"A7",X"C8",X"FE",X"10",X"C8",X"FD",X"66",X"04",
		X"FD",X"6E",X"05",X"01",X"08",X"00",X"ED",X"42",X"FD",X"74",X"04",X"FD",X"75",X"05",X"FD",X"35",
		X"01",X"FD",X"7E",X"01",X"A7",X"C0",X"FD",X"34",X"01",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"01",
		X"08",X"00",X"09",X"FD",X"74",X"04",X"FD",X"75",X"05",X"C9",X"3A",X"96",X"E2",X"A7",X"C2",X"D5",
		X"42",X"3C",X"32",X"96",X"E2",X"3E",X"01",X"32",X"A7",X"E5",X"FD",X"7E",X"00",X"32",X"AA",X"E2",
		X"FD",X"7E",X"03",X"32",X"AB",X"E2",X"3E",X"FF",X"A7",X"C9",X"FD",X"36",X"01",X"00",X"FD",X"7E",
		X"03",X"3C",X"32",X"BE",X"E5",X"FD",X"34",X"0F",X"C9",X"DD",X"7E",X"0E",X"A7",X"CA",X"0F",X"43",
		X"FD",X"36",X"0E",X"01",X"FD",X"36",X"0A",X"00",X"DD",X"34",X"0B",X"FD",X"34",X"0B",X"C9",X"FD",
		X"7E",X"0E",X"A7",X"C8",X"DD",X"36",X"0E",X"01",X"DD",X"36",X"0A",X"00",X"DD",X"34",X"0B",X"FD",
		X"34",X"0B",X"C9",X"DD",X"7E",X"02",X"DD",X"86",X"06",X"A7",X"C8",X"FD",X"E5",X"CD",X"7B",X"1F",
		X"FD",X"E1",X"D2",X"39",X"43",X"CD",X"DB",X"38",X"C9",X"DD",X"46",X"03",X"DD",X"36",X"03",X"E0",
		X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"70",X"03",X"D2",X"67",X"43",X"FD",X"7E",X"01",
		X"D6",X"04",X"3A",X"14",X"EC",X"DD",X"46",X"00",X"B8",X"D2",X"63",X"43",X"FD",X"36",X"02",X"10",
		X"C3",X"67",X"43",X"FD",X"36",X"02",X"F0",X"AF",X"32",X"B8",X"E5",X"DD",X"7E",X"00",X"47",X"C6",
		X"10",X"DD",X"77",X"00",X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"70",X"00",X"DA",X"95",
		X"43",X"DD",X"7E",X"00",X"47",X"D6",X"10",X"DD",X"77",X"00",X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",
		X"E1",X"DD",X"70",X"00",X"D0",X"3E",X"10",X"32",X"B8",X"E5",X"C9",X"3A",X"BF",X"E5",X"A7",X"C8",
		X"3A",X"83",X"E2",X"E6",X"03",X"FE",X"02",X"C0",X"3A",X"B6",X"E5",X"A7",X"C0",X"3A",X"BA",X"E5",
		X"3C",X"32",X"BA",X"E5",X"DD",X"21",X"D8",X"E1",X"FD",X"21",X"60",X"E5",X"CD",X"C0",X"43",X"C9",
		X"FD",X"7E",X"01",X"A7",X"CA",X"37",X"44",X"3A",X"C6",X"E2",X"A7",X"C2",X"09",X"44",X"CD",X"8C",
		X"35",X"CC",X"65",X"44",X"3A",X"C0",X"E5",X"A7",X"C8",X"CD",X"EE",X"44",X"CD",X"4F",X"44",X"DD",
		X"E5",X"FD",X"E5",X"CD",X"EF",X"45",X"CD",X"61",X"47",X"FD",X"E1",X"DD",X"E1",X"CD",X"A0",X"46",
		X"3E",X"02",X"32",X"BD",X"E5",X"06",X"01",X"CD",X"18",X"34",X"CD",X"1D",X"37",X"CD",X"0D",X"47",
		X"CD",X"64",X"38",X"06",X"06",X"CD",X"27",X"3F",X"C9",X"FD",X"7E",X"01",X"A7",X"C2",X"1F",X"44",
		X"CD",X"1D",X"37",X"CD",X"19",X"38",X"CD",X"64",X"38",X"06",X"06",X"CD",X"27",X"3F",X"C9",X"FD",
		X"36",X"01",X"0B",X"06",X"01",X"CD",X"18",X"34",X"CD",X"1D",X"37",X"CD",X"0D",X"47",X"CD",X"64",
		X"38",X"06",X"06",X"CD",X"27",X"3F",X"C9",X"CD",X"8C",X"35",X"CA",X"D1",X"43",X"CD",X"EB",X"34",
		X"CD",X"1D",X"37",X"CD",X"19",X"38",X"CD",X"64",X"38",X"06",X"06",X"CD",X"27",X"3F",X"C9",X"3A",
		X"C0",X"E5",X"A7",X"C8",X"FD",X"34",X"0A",X"FD",X"7E",X"0A",X"FE",X"05",X"D8",X"3E",X"16",X"D7",
		X"FD",X"36",X"0A",X"00",X"C9",X"AF",X"32",X"C0",X"E5",X"3A",X"A7",X"E2",X"A7",X"C0",X"3A",X"7E",
		X"E0",X"A7",X"C0",X"3A",X"BA",X"E5",X"FE",X"10",X"D0",X"FD",X"86",X"00",X"FD",X"77",X"00",X"CD",
		X"EB",X"1F",X"E6",X"03",X"21",X"EA",X"44",X"4F",X"06",X"00",X"09",X"7E",X"DD",X"77",X"00",X"3A",
		X"96",X"E2",X"A7",X"C0",X"AF",X"32",X"BB",X"E5",X"32",X"AC",X"E5",X"CD",X"EB",X"1F",X"E6",X"03",
		X"47",X"32",X"AC",X"E5",X"3A",X"82",X"E2",X"C6",X"02",X"FD",X"77",X"01",X"CD",X"C6",X"44",X"C0",
		X"FD",X"36",X"04",X"00",X"FD",X"36",X"05",X"D8",X"FD",X"36",X"0A",X"04",X"FD",X"36",X"0B",X"28",
		X"3E",X"01",X"32",X"C0",X"E5",X"C9",X"DD",X"E5",X"DD",X"21",X"A8",X"E1",X"CD",X"8C",X"35",X"DD",
		X"E1",X"C0",X"DD",X"E5",X"DD",X"21",X"08",X"E2",X"CD",X"8C",X"35",X"DD",X"E1",X"C0",X"DD",X"E5",
		X"DD",X"21",X"68",X"E2",X"CD",X"8C",X"35",X"DD",X"E1",X"C9",X"58",X"90",X"90",X"C8",X"FD",X"7E",
		X"04",X"FE",X"01",X"C0",X"3A",X"AC",X"E5",X"21",X"05",X"45",X"CB",X"27",X"06",X"00",X"4F",X"09",
		X"5E",X"23",X"56",X"EB",X"E9",X"0E",X"45",X"0E",X"45",X"88",X"45",X"88",X"45",X"C9",X"3A",X"C7",
		X"E1",X"C6",X"40",X"DD",X"4E",X"03",X"B9",X"D2",X"6A",X"45",X"3E",X"0F",X"32",X"BB",X"E5",X"3A",
		X"C4",X"E1",X"D6",X"10",X"DD",X"4E",X"00",X"B9",X"D2",X"35",X"45",X"3A",X"C4",X"E1",X"B9",X"DA",
		X"40",X"45",X"C3",X"48",X"45",X"DD",X"7E",X"00",X"C6",X"04",X"DD",X"77",X"00",X"C3",X"48",X"45",
		X"DD",X"7E",X"00",X"D6",X"04",X"DD",X"77",X"00",X"3A",X"82",X"E2",X"FD",X"77",X"01",X"FD",X"7E",
		X"0B",X"A7",X"CA",X"7F",X"45",X"FD",X"35",X"0B",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"01",X"02",
		X"00",X"ED",X"42",X"FD",X"74",X"04",X"FD",X"75",X"05",X"C9",X"3A",X"BB",X"E5",X"A7",X"C2",X"1A",
		X"45",X"FD",X"7E",X"01",X"A7",X"C8",X"3A",X"82",X"E2",X"3C",X"3C",X"FD",X"77",X"01",X"C9",X"3A",
		X"82",X"E2",X"C6",X"03",X"FD",X"77",X"01",X"C9",X"FD",X"35",X"0B",X"FD",X"7E",X"0B",X"A7",X"CA",
		X"E1",X"45",X"3A",X"C0",X"E1",X"DD",X"46",X"00",X"90",X"D2",X"9E",X"45",X"ED",X"44",X"FE",X"28",
		X"D2",X"E1",X"45",X"FE",X"04",X"DA",X"C1",X"45",X"3A",X"C0",X"E1",X"DD",X"46",X"00",X"B8",X"D2",
		X"BB",X"45",X"DD",X"35",X"00",X"DD",X"35",X"00",X"C3",X"C1",X"45",X"DD",X"34",X"00",X"DD",X"34",
		X"00",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"23",X"23",X"45",X"3A",X"C3",X"E1",X"90",X"FE",X"48",
		X"D8",X"FE",X"60",X"D0",X"3A",X"82",X"E2",X"FD",X"77",X"01",X"FD",X"74",X"04",X"FD",X"75",X"05",
		X"C9",X"3A",X"82",X"E2",X"C6",X"03",X"FD",X"77",X"01",X"C9",X"FD",X"36",X"01",X"00",X"C9",X"FD",
		X"21",X"D8",X"E1",X"3A",X"96",X"E2",X"A7",X"C2",X"03",X"46",X"CD",X"40",X"03",X"CA",X"03",X"46",
		X"32",X"96",X"E2",X"DD",X"21",X"F0",X"E1",X"AF",X"CD",X"45",X"03",X"CA",X"15",X"46",X"3A",X"31",
		X"E5",X"A7",X"CA",X"9B",X"46",X"DD",X"7E",X"00",X"FD",X"46",X"00",X"C6",X"10",X"90",X"DA",X"38",
		X"46",X"FE",X"30",X"D2",X"38",X"46",X"FE",X"18",X"D2",X"33",X"46",X"3E",X"08",X"32",X"3D",X"E5",
		X"C3",X"38",X"46",X"3E",X"F8",X"32",X"3D",X"E5",X"DD",X"21",X"F8",X"E1",X"AF",X"CD",X"45",X"03",
		X"CA",X"4A",X"46",X"3A",X"41",X"E5",X"A7",X"CA",X"9B",X"46",X"DD",X"7E",X"00",X"FD",X"46",X"00",
		X"C6",X"10",X"90",X"DA",X"6D",X"46",X"FE",X"30",X"D2",X"6D",X"46",X"FE",X"18",X"D2",X"68",X"46",
		X"3E",X"08",X"32",X"4D",X"E5",X"C3",X"6D",X"46",X"3E",X"F8",X"32",X"4D",X"E5",X"DD",X"21",X"00",
		X"E2",X"AF",X"CD",X"45",X"03",X"C8",X"3A",X"51",X"E5",X"A7",X"CA",X"9B",X"46",X"DD",X"7E",X"00",
		X"FD",X"46",X"00",X"C6",X"10",X"90",X"D8",X"FE",X"30",X"D0",X"FE",X"18",X"D2",X"95",X"46",X"3E",
		X"08",X"32",X"5D",X"E5",X"C9",X"3E",X"F8",X"32",X"5D",X"E5",X"C9",X"AF",X"32",X"61",X"E5",X"C9",
		X"DD",X"7E",X"03",X"47",X"C6",X"40",X"DD",X"77",X"03",X"DD",X"7E",X"00",X"4F",X"C6",X"08",X"DD",
		X"77",X"00",X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"71",X"00",X"DD",X"70",X"03",X"D2",
		X"CB",X"46",X"FD",X"36",X"01",X"00",X"FD",X"36",X"0B",X"00",X"C9",X"DD",X"7E",X"00",X"47",X"D6",
		X"10",X"DD",X"77",X"00",X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"70",X"00",X"D2",X"ED",
		X"46",X"DD",X"7E",X"00",X"C6",X"03",X"DD",X"77",X"00",X"FD",X"35",X"0B",X"C9",X"DD",X"7E",X"00",
		X"47",X"C6",X"10",X"DD",X"77",X"00",X"FD",X"E5",X"CD",X"7B",X"1F",X"FD",X"E1",X"DD",X"70",X"00",
		X"D0",X"DD",X"7E",X"00",X"D6",X"03",X"DD",X"77",X"00",X"FD",X"35",X"0B",X"C9",X"FD",X"34",X"03",
		X"FD",X"7E",X"03",X"CB",X"47",X"C0",X"FE",X"08",X"DA",X"1F",X"47",X"AF",X"FD",X"77",X"03",X"21",
		X"41",X"47",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",X"DD",X"E5",X"06",X"06",X"11",X"04",
		X"00",X"7E",X"DD",X"36",X"01",X"40",X"DD",X"77",X"02",X"23",X"DD",X"19",X"10",X"F3",X"DD",X"E1",
		X"C9",X"49",X"47",X"4F",X"47",X"55",X"47",X"5B",X"47",X"2F",X"2D",X"2E",X"2C",X"30",X"2B",X"41",
		X"3F",X"2E",X"2C",X"42",X"3D",X"2F",X"2D",X"40",X"3E",X"30",X"2B",X"41",X"3F",X"40",X"3E",X"42",
		X"3D",X"3A",X"01",X"E5",X"A7",X"CA",X"85",X"47",X"DD",X"21",X"A8",X"E1",X"FD",X"21",X"D8",X"E1",
		X"CD",X"0E",X"48",X"3A",X"B7",X"E5",X"A7",X"CA",X"85",X"47",X"DD",X"21",X"00",X"E5",X"FD",X"21",
		X"60",X"E5",X"CD",X"CA",X"47",X"3A",X"11",X"E5",X"A7",X"CA",X"A9",X"47",X"DD",X"21",X"08",X"E2",
		X"FD",X"21",X"D8",X"E1",X"CD",X"0E",X"48",X"3A",X"B7",X"E5",X"A7",X"CA",X"A9",X"47",X"DD",X"21",
		X"10",X"E5",X"FD",X"21",X"60",X"E5",X"CD",X"CA",X"47",X"3A",X"21",X"E5",X"A7",X"C8",X"DD",X"21",
		X"68",X"E2",X"FD",X"21",X"D8",X"E1",X"CD",X"0E",X"48",X"3A",X"B7",X"E5",X"A7",X"C8",X"DD",X"21",
		X"20",X"E5",X"FD",X"21",X"60",X"E5",X"CD",X"CA",X"47",X"C9",X"FD",X"7E",X"05",X"DD",X"46",X"05",
		X"B8",X"D2",X"F1",X"47",X"DD",X"7E",X"01",X"FE",X"02",X"D2",X"E4",X"47",X"AF",X"DD",X"77",X"01",
		X"FD",X"77",X"01",X"C9",X"FD",X"35",X"01",X"FD",X"35",X"01",X"DD",X"34",X"01",X"DD",X"34",X"01",
		X"C9",X"DD",X"7E",X"01",X"FE",X"02",X"D2",X"01",X"48",X"AF",X"DD",X"77",X"01",X"FD",X"77",X"01",
		X"C9",X"FD",X"34",X"01",X"FD",X"34",X"01",X"DD",X"35",X"01",X"DD",X"35",X"01",X"C9",X"AF",X"32",
		X"B7",X"E5",X"DD",X"7E",X"02",X"A7",X"C8",X"FD",X"7E",X"02",X"A7",X"C8",X"FD",X"7E",X"00",X"DD",
		X"46",X"00",X"90",X"D2",X"28",X"48",X"ED",X"44",X"FE",X"20",X"DA",X"33",X"48",X"FE",X"28",X"DA",
		X"45",X"48",X"C9",X"FD",X"7E",X"03",X"DD",X"46",X"03",X"90",X"D2",X"3F",X"48",X"ED",X"44",X"FE",
		X"40",X"DA",X"57",X"48",X"C9",X"FD",X"7E",X"03",X"DD",X"46",X"03",X"90",X"D2",X"51",X"48",X"ED",
		X"44",X"FE",X"40",X"DA",X"57",X"48",X"C9",X"3E",X"0F",X"32",X"B7",X"E5",X"C9",X"3A",X"B6",X"E5",
		X"A7",X"C2",X"93",X"48",X"3A",X"AF",X"E5",X"A7",X"C8",X"3A",X"7E",X"E0",X"A7",X"C0",X"3A",X"C0",
		X"E5",X"A7",X"C0",X"DD",X"21",X"A8",X"E1",X"CD",X"8C",X"35",X"C0",X"DD",X"21",X"08",X"E2",X"CD",
		X"8C",X"35",X"C0",X"DD",X"21",X"68",X"E2",X"CD",X"8C",X"35",X"C0",X"3E",X"01",X"32",X"B6",X"E5",
		X"C3",X"C0",X"48",X"3A",X"83",X"E2",X"E6",X"03",X"FE",X"03",X"C0",X"DD",X"21",X"D8",X"E1",X"CD",
		X"8C",X"35",X"C2",X"FC",X"48",X"DD",X"21",X"08",X"E2",X"CD",X"8C",X"35",X"C2",X"FC",X"48",X"AF",
		X"32",X"AF",X"E5",X"32",X"B6",X"E5",X"32",X"0B",X"E5",X"32",X"1B",X"E5",X"32",X"2B",X"E5",X"C9",
		X"3A",X"A7",X"E2",X"A7",X"C0",X"DD",X"21",X"D8",X"E1",X"FD",X"21",X"70",X"E5",X"CD",X"D1",X"36",
		X"E6",X"03",X"16",X"00",X"5F",X"21",X"E0",X"48",X"19",X"7E",X"DD",X"77",X"00",X"C3",X"E4",X"48",
		X"50",X"88",X"D0",X"88",X"3A",X"82",X"E2",X"C6",X"04",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",
		X"FD",X"36",X"04",X"00",X"FD",X"36",X"05",X"B8",X"FD",X"36",X"0A",X"02",X"DD",X"21",X"D8",X"E1",
		X"FD",X"21",X"70",X"E5",X"3E",X"03",X"32",X"BD",X"E5",X"06",X"01",X"CD",X"18",X"34",X"CD",X"35",
		X"49",X"CD",X"24",X"49",X"CD",X"97",X"49",X"CD",X"03",X"4A",X"CD",X"30",X"4A",X"CD",X"6A",X"4A",
		X"CD",X"81",X"4A",X"C9",X"FD",X"34",X"0A",X"FD",X"7E",X"0A",X"FE",X"03",X"D8",X"3E",X"16",X"D7",
		X"FD",X"36",X"0A",X"00",X"C9",X"DD",X"7E",X"02",X"A7",X"C8",X"DD",X"7E",X"03",X"FE",X"30",X"D8",
		X"FD",X"7E",X"02",X"A7",X"C2",X"62",X"49",X"3A",X"C4",X"E1",X"47",X"CD",X"EB",X"1F",X"FE",X"0A",
		X"D0",X"DD",X"7E",X"00",X"B8",X"D2",X"5D",X"49",X"FD",X"36",X"02",X"F0",X"C9",X"FD",X"36",X"02",
		X"10",X"C9",X"FD",X"7E",X"02",X"FE",X"10",X"CA",X"82",X"49",X"FE",X"F0",X"C0",X"DD",X"7E",X"00",
		X"C6",X"03",X"47",X"3A",X"C4",X"E1",X"B8",X"D2",X"7E",X"49",X"FD",X"36",X"02",X"80",X"DD",X"70",
		X"00",X"C9",X"DD",X"7E",X"00",X"D6",X"03",X"47",X"3A",X"C4",X"E1",X"B8",X"DA",X"93",X"49",X"FD",
		X"36",X"02",X"80",X"DD",X"70",X"00",X"C9",X"FD",X"21",X"08",X"E2",X"CD",X"A6",X"49",X"FD",X"21",
		X"D8",X"E1",X"CD",X"A6",X"49",X"C9",X"CD",X"40",X"03",X"CA",X"AF",X"49",X"32",X"96",X"E2",X"3A",
		X"31",X"E5",X"A7",X"CA",X"CC",X"49",X"DD",X"21",X"F0",X"E1",X"AF",X"CD",X"45",X"03",X"CA",X"CC",
		X"49",X"FD",X"E5",X"FD",X"21",X"30",X"E5",X"CD",X"DB",X"38",X"FD",X"E1",X"3A",X"41",X"E5",X"A7",
		X"CA",X"E9",X"49",X"DD",X"21",X"F8",X"E1",X"AF",X"CD",X"45",X"03",X"CA",X"E9",X"49",X"FD",X"E5",
		X"FD",X"21",X"40",X"E5",X"CD",X"DB",X"38",X"FD",X"E1",X"3A",X"51",X"E5",X"A7",X"C8",X"DD",X"21",
		X"00",X"E2",X"AF",X"CD",X"45",X"03",X"C8",X"FD",X"E5",X"FD",X"21",X"50",X"E5",X"CD",X"DB",X"38",
		X"FD",X"E1",X"C9",X"DD",X"21",X"D8",X"E1",X"FD",X"21",X"70",X"E5",X"CD",X"1D",X"37",X"DD",X"46",
		X"00",X"FD",X"66",X"08",X"FD",X"6E",X"09",X"DD",X"21",X"08",X"E2",X"FD",X"21",X"80",X"E5",X"11",
		X"10",X"00",X"19",X"DD",X"70",X"00",X"FD",X"74",X"04",X"FD",X"75",X"05",X"CD",X"1D",X"37",X"C9",
		X"FD",X"21",X"70",X"E5",X"FD",X"34",X"03",X"FD",X"7E",X"03",X"CB",X"47",X"C2",X"45",X"4A",X"21",
		X"94",X"4A",X"C3",X"48",X"4A",X"21",X"A0",X"4A",X"DD",X"21",X"D8",X"E1",X"CD",X"57",X"4A",X"DD",
		X"21",X"08",X"E2",X"CD",X"57",X"4A",X"C9",X"06",X"06",X"11",X"04",X"00",X"7E",X"DD",X"36",X"01",
		X"41",X"DD",X"77",X"02",X"23",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"21",X"D8",X"E1",X"FD",X"21",
		X"70",X"E5",X"CD",X"64",X"38",X"DD",X"21",X"08",X"E2",X"FD",X"21",X"80",X"E5",X"CD",X"64",X"38",
		X"C9",X"DD",X"21",X"D8",X"E1",X"06",X"06",X"CD",X"27",X"3F",X"DD",X"21",X"08",X"E2",X"06",X"06",
		X"CD",X"27",X"3F",X"C9",X"57",X"55",X"56",X"54",X"53",X"51",X"52",X"50",X"4F",X"4D",X"4E",X"4C",
		X"57",X"55",X"56",X"54",X"53",X"51",X"52",X"50",X"4F",X"4D",X"59",X"58",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"03",X"03",X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"03",X"03",
		X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"03",X"03",X"01",X"DD",X"DD",X"CD",X"CD",X"07",X"02",X"03",
		X"01",X"CD",X"CD",X"CD",X"CD",X"07",X"02",X"03",X"01",X"CD",X"CD",X"CD",X"CD",X"07",X"02",X"03",
		X"01",X"CD",X"CD",X"CD",X"CD",X"07",X"02",X"03",X"01",X"CD",X"CD",X"CD",X"CD",X"01",X"03",X"02",
		X"07",X"DD",X"DD",X"DD",X"DD",X"01",X"03",X"02",X"07",X"DD",X"DD",X"DD",X"DD",X"01",X"03",X"02",
		X"07",X"DD",X"DD",X"DD",X"DD",X"01",X"03",X"02",X"07",X"DD",X"DD",X"DD",X"DD",X"07",X"02",X"03",
		X"01",X"CD",X"CD",X"CD",X"CD",X"07",X"05",X"03",X"01",X"ED",X"ED",X"CD",X"CD",X"06",X"04",X"03",
		X"01",X"ED",X"ED",X"CD",X"CD",X"01",X"03",X"03",X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"03",X"03",
		X"01",X"DD",X"DD",X"CD",X"CD",X"06",X"04",X"03",X"01",X"CD",X"CD",X"CD",X"CD",X"07",X"05",X"03",
		X"01",X"CD",X"CD",X"CD",X"CD",X"07",X"02",X"03",X"01",X"CD",X"CD",X"CD",X"CD",X"01",X"03",X"02",
		X"07",X"DD",X"DD",X"DD",X"FD",X"01",X"03",X"05",X"07",X"DD",X"DD",X"FD",X"FD",X"01",X"03",X"04",
		X"06",X"DD",X"DD",X"FD",X"FD",X"01",X"03",X"03",X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"12",X"12",
		X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"10",X"10",X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"77",X"75",
		X"26",X"DD",X"ED",X"ED",X"ED",X"01",X"76",X"74",X"07",X"DD",X"ED",X"ED",X"ED",X"01",X"12",X"12",
		X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"10",X"10",X"01",X"DD",X"DD",X"CD",X"CD",X"26",X"75",X"77",
		X"01",X"FD",X"FD",X"FD",X"ED",X"07",X"74",X"76",X"01",X"FD",X"FD",X"FD",X"ED",X"7B",X"79",X"73",
		X"71",X"E8",X"E8",X"E8",X"E8",X"7A",X"78",X"72",X"70",X"E8",X"E8",X"E8",X"E8",X"0F",X"0D",X"0B",
		X"09",X"E8",X"E8",X"E8",X"E8",X"0E",X"0C",X"0A",X"08",X"E8",X"E8",X"E8",X"E8",X"14",X"16",X"1B",
		X"07",X"DD",X"DD",X"ED",X"ED",X"15",X"17",X"1A",X"18",X"DD",X"DD",X"ED",X"ED",X"18",X"1A",X"17",
		X"15",X"DD",X"DD",X"ED",X"ED",X"07",X"1B",X"16",X"14",X"DD",X"DD",X"ED",X"ED",X"07",X"1B",X"16",
		X"14",X"FD",X"FD",X"CD",X"CD",X"18",X"1A",X"17",X"15",X"FD",X"FD",X"CD",X"CD",X"15",X"17",X"1A",
		X"18",X"FD",X"FD",X"CD",X"CD",X"14",X"16",X"1B",X"07",X"FD",X"FD",X"CD",X"CD",X"5F",X"5D",X"57",
		X"55",X"E8",X"E8",X"E8",X"E8",X"5E",X"5C",X"56",X"54",X"E8",X"E8",X"E8",X"E8",X"5B",X"59",X"53",
		X"51",X"E8",X"E8",X"E8",X"E8",X"5A",X"58",X"52",X"50",X"E8",X"E8",X"E8",X"E8",X"F3",X"F1",X"07",
		X"27",X"ED",X"ED",X"ED",X"ED",X"F2",X"F0",X"25",X"28",X"ED",X"ED",X"ED",X"ED",X"29",X"25",X"F0",
		X"F4",X"ED",X"DD",X"DD",X"ED",X"07",X"07",X"F1",X"F3",X"DD",X"DD",X"DD",X"DD",X"01",X"03",X"21",
		X"22",X"FD",X"FD",X"FD",X"FD",X"01",X"03",X"21",X"22",X"FD",X"FD",X"FD",X"FD",X"1D",X"1F",X"20",
		X"22",X"FD",X"FD",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"24",X"2A",
		X"00",X"FD",X"FD",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"07",
		X"27",X"DD",X"CD",X"DD",X"CD",X"2C",X"2C",X"07",X"27",X"DD",X"CD",X"DD",X"CD",X"2C",X"2C",X"07",
		X"27",X"DD",X"CD",X"DD",X"CD",X"2C",X"2C",X"07",X"27",X"DD",X"CD",X"DD",X"CD",X"07",X"07",X"F1",
		X"F3",X"FD",X"FD",X"FD",X"FD",X"29",X"25",X"F0",X"F4",X"CD",X"FD",X"FD",X"CD",X"F2",X"F0",X"25",
		X"28",X"CD",X"CD",X"CD",X"CD",X"F3",X"F1",X"07",X"27",X"CD",X"CD",X"CD",X"CD",X"07",X"07",X"2C",
		X"2C",X"CD",X"CD",X"DD",X"CD",X"07",X"07",X"2C",X"2C",X"CD",X"CD",X"DD",X"CD",X"07",X"07",X"2C",
		X"2C",X"CD",X"CD",X"DD",X"CD",X"07",X"07",X"2C",X"2C",X"CD",X"CD",X"DD",X"CD",X"6F",X"6D",X"67",
		X"65",X"ED",X"ED",X"ED",X"ED",X"6E",X"6C",X"66",X"64",X"ED",X"ED",X"ED",X"ED",X"6B",X"69",X"63",
		X"61",X"ED",X"ED",X"ED",X"ED",X"6A",X"68",X"62",X"60",X"ED",X"ED",X"ED",X"ED",X"63",X"61",X"3B",
		X"39",X"A8",X"A8",X"A8",X"A8",X"62",X"60",X"3A",X"38",X"A8",X"A8",X"A8",X"A8",X"5F",X"5D",X"37",
		X"35",X"A8",X"A8",X"A8",X"A8",X"5E",X"5C",X"36",X"34",X"A8",X"A8",X"A8",X"A8",X"4F",X"4D",X"47",
		X"45",X"ED",X"ED",X"ED",X"ED",X"4E",X"4C",X"46",X"44",X"ED",X"ED",X"ED",X"ED",X"4B",X"49",X"43",
		X"41",X"ED",X"ED",X"ED",X"ED",X"4A",X"48",X"42",X"40",X"ED",X"ED",X"ED",X"ED",X"8B",X"89",X"83",
		X"81",X"ED",X"ED",X"ED",X"ED",X"8A",X"88",X"82",X"80",X"ED",X"ED",X"ED",X"ED",X"87",X"85",X"7F",
		X"7D",X"ED",X"ED",X"ED",X"ED",X"86",X"84",X"7E",X"7C",X"ED",X"ED",X"ED",X"ED",X"9B",X"99",X"93",
		X"91",X"ED",X"ED",X"ED",X"ED",X"9A",X"98",X"92",X"90",X"ED",X"ED",X"ED",X"ED",X"97",X"95",X"8F",
		X"8D",X"ED",X"ED",X"ED",X"ED",X"96",X"94",X"8E",X"8C",X"ED",X"ED",X"ED",X"ED",X"BB",X"B9",X"B3",
		X"B1",X"ED",X"ED",X"ED",X"ED",X"BA",X"B8",X"B2",X"B0",X"ED",X"ED",X"ED",X"ED",X"B7",X"B5",X"AF",
		X"AD",X"ED",X"ED",X"ED",X"ED",X"B6",X"B4",X"AE",X"AC",X"ED",X"ED",X"ED",X"ED",X"35",X"3D",X"37",
		X"35",X"ED",X"ED",X"ED",X"ED",X"35",X"3C",X"36",X"34",X"ED",X"ED",X"ED",X"ED",X"3B",X"39",X"33",
		X"31",X"ED",X"ED",X"ED",X"ED",X"3A",X"38",X"32",X"30",X"ED",X"ED",X"ED",X"ED",X"01",X"10",X"10",
		X"01",X"DD",X"FD",X"ED",X"CD",X"01",X"12",X"12",X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"12",X"12",
		X"01",X"DD",X"DD",X"CD",X"CD",X"01",X"10",X"10",X"01",X"DD",X"DD",X"CD",X"CD",X"E0",X"56",X"E0",
		X"56",X"E0",X"56",X"E0",X"56",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"41",
		X"65",X"A8",X"63",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"73",X"68",X"DA",
		X"66",X"A5",X"6B",X"12",X"5A",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"D1",X"7E",X"EA",X"7E",X"28",
		X"01",X"50",X"01",X"50",X"01",X"66",X"01",X"01",X"01",X"01",X"01",X"01",X"70",X"01",X"01",X"01",
		X"01",X"14",X"06",X"22",X"01",X"18",X"DD",X"5E",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",
		X"3E",X"6D",X"D7",X"6E",X"70",X"70",X"09",X"72",X"3E",X"6D",X"D7",X"6E",X"09",X"72",X"3E",X"6D",
		X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"44",X"5D",
		X"E0",X"56",X"44",X"5D",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",
		X"0C",X"6A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"47",X"55",X"E0",X"56",X"79",X"58",
		X"AE",X"53",X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",X"63",X"73",X"68",X"DA",X"66",X"A5",X"6B",
		X"06",X"7A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",
		X"AB",X"5B",X"44",X"5D",X"D1",X"7E",X"EA",X"7E",X"01",X"0A",X"01",X"01",X"14",X"41",X"01",X"28",
		X"01",X"1E",X"01",X"01",X"14",X"1E",X"01",X"01",X"0A",X"01",X"0A",X"08",X"03",X"08",X"0A",X"02",
		X"01",X"0A",X"01",X"01",X"0F",X"01",X"1E",X"01",X"01",X"14",X"01",X"3E",X"01",X"0A",X"01",X"01",
		X"01",X"01",X"01",X"01",X"0A",X"01",X"0A",X"01",X"01",X"0A",X"01",X"01",X"0F",X"01",X"18",X"9F",
		X"7B",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"A2",X"73",X"76",X"60",X"0F",
		X"62",X"76",X"60",X"0F",X"62",X"76",X"60",X"0F",X"62",X"76",X"60",X"0F",X"62",X"A2",X"73",X"76",
		X"60",X"0F",X"62",X"76",X"60",X"0F",X"62",X"A2",X"73",X"3B",X"75",X"D4",X"76",X"6D",X"78",X"73",
		X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"44",
		X"5D",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"0C",X"6A",X"A5",
		X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",X"63",X"73",
		X"68",X"DA",X"66",X"A5",X"6B",X"06",X"7A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"73",
		X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"D1",X"7E",X"EA",X"7E",X"01",X"0A",X"01",
		X"01",X"14",X"01",X"05",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"3C",X"01",X"01",X"01",
		X"01",X"03",X"01",X"50",X"01",X"01",X"01",X"1E",X"01",X"0A",X"08",X"0A",X"3F",X"0A",X"02",X"01",
		X"0A",X"01",X"01",X"0F",X"01",X"1E",X"01",X"01",X"1E",X"01",X"01",X"01",X"01",X"01",X"01",X"0A",
		X"01",X"12",X"01",X"01",X"0A",X"01",X"01",X"0F",X"01",X"18",X"DD",X"5E",X"41",X"65",X"A8",X"63",
		X"AE",X"53",X"47",X"55",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"12",X"5A",
		X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"0C",X"6A",
		X"A5",X"6B",X"06",X"7A",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"79",X"58",X"AE",X"53",
		X"73",X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",
		X"44",X"5D",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"0C",X"6A",X"A5",X"6B",
		X"AB",X"5B",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"41",X"65",X"A8",X"63",
		X"73",X"68",X"DA",X"66",X"A5",X"6B",X"06",X"7A",X"0C",X"6A",X"41",X"65",X"A8",X"63",X"73",X"68",
		X"DA",X"66",X"06",X"7A",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",
		X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",
		X"0C",X"6A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"47",X"55",X"E0",X"56",X"79",X"58",X"73",X"68",
		X"DA",X"66",X"41",X"65",X"A8",X"63",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"06",X"7A",X"41",X"65",
		X"A8",X"63",X"AE",X"53",X"47",X"55",X"E0",X"56",X"03",X"7F",X"1C",X"7F",X"01",X"01",X"01",X"0A",
		X"01",X"15",X"01",X"01",X"01",X"0E",X"06",X"18",X"01",X"01",X"14",X"01",X"01",X"04",X"01",X"04",
		X"01",X"0A",X"01",X"01",X"02",X"01",X"1E",X"01",X"01",X"0A",X"01",X"0A",X"08",X"03",X"08",X"0A",
		X"02",X"01",X"01",X"01",X"05",X"01",X"0A",X"01",X"1E",X"01",X"01",X"01",X"02",X"01",X"01",X"01",
		X"01",X"08",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0A",X"01",X"0A",X"08",X"03",X"32",X"03",
		X"08",X"0A",X"02",X"01",X"0A",X"01",X"01",X"01",X"0A",X"01",X"01",X"01",X"1E",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"0A",X"01",X"01",X"01",X"0F",X"01",X"1B",X"9F",X"7B",X"AE",X"53",X"AE",
		X"53",X"AE",X"53",X"47",X"55",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"12",
		X"5A",X"A5",X"6B",X"AB",X"5B",X"A2",X"73",X"76",X"60",X"0F",X"62",X"76",X"60",X"0F",X"62",X"76",
		X"60",X"0F",X"62",X"76",X"60",X"0F",X"62",X"A2",X"73",X"76",X"60",X"0F",X"62",X"76",X"60",X"0F",
		X"62",X"A2",X"73",X"E0",X"56",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",
		X"6B",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"79",
		X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"0C",X"6A",X"A5",X"6B",X"41",X"65",X"A8",
		X"63",X"AE",X"53",X"47",X"55",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",
		X"63",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"06",X"7A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",
		X"53",X"47",X"55",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",
		X"63",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"44",X"5D",X"03",X"7F",X"1C",X"7F",X"01",
		X"01",X"01",X"0A",X"01",X"15",X"01",X"01",X"01",X"0E",X"06",X"18",X"01",X"05",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"28",X"01",X"01",X"01",X"01",X"03",X"2C",X"11",X"01",X"14",X"01",
		X"01",X"0A",X"01",X"0A",X"08",X"03",X"08",X"0A",X"02",X"01",X"0A",X"01",X"01",X"0A",X"01",X"14",
		X"01",X"01",X"12",X"01",X"1E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"08",X"01",X"08",X"01",
		X"01",X"0F",X"01",X"2B",X"01",X"0A",X"01",X"01",X"01",X"01",X"01",X"01",X"0A",X"01",X"1B",X"9F",
		X"7B",X"AE",X"53",X"AE",X"53",X"AE",X"53",X"47",X"55",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",
		X"66",X"A5",X"6B",X"12",X"5A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"3E",X"6D",X"D7",
		X"6E",X"70",X"70",X"09",X"72",X"3E",X"6D",X"D7",X"6E",X"70",X"70",X"09",X"72",X"3E",X"6D",X"D7",
		X"6E",X"09",X"72",X"3E",X"6D",X"AE",X"53",X"73",X"68",X"DA",X"66",X"A5",X"6B",X"AB",X"5B",X"44",
		X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",
		X"68",X"DA",X"66",X"A5",X"6B",X"0C",X"6A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"47",
		X"55",X"E0",X"56",X"79",X"58",X"AE",X"53",X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",X"63",X"73",
		X"68",X"DA",X"66",X"A5",X"6B",X"06",X"7A",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"47",X"55",X"E0",
		X"56",X"03",X"7F",X"1C",X"7F",X"01",X"01",X"01",X"0A",X"01",X"15",X"01",X"01",X"01",X"0E",X"06",
		X"18",X"01",X"01",X"0F",X"28",X"01",X"1E",X"01",X"1E",X"01",X"14",X"01",X"0A",X"01",X"01",X"0A",
		X"1E",X"01",X"01",X"0A",X"01",X"0A",X"08",X"03",X"08",X"0A",X"02",X"01",X"0A",X"01",X"01",X"0F",
		X"01",X"1E",X"01",X"01",X"12",X"01",X"2A",X"01",X"08",X"01",X"01",X"01",X"01",X"01",X"01",X"08",
		X"01",X"09",X"01",X"01",X"01",X"1B",X"E0",X"56",X"79",X"58",X"73",X"68",X"DA",X"66",X"A5",X"6B",
		X"12",X"5A",X"A5",X"6B",X"A5",X"6B",X"41",X"65",X"A8",X"63",X"AE",X"53",X"73",X"68",X"DA",X"66",
		X"41",X"65",X"A8",X"63",X"47",X"55",X"E0",X"56",X"E0",X"56",X"E0",X"56",X"79",X"58",X"AE",X"53",
		X"73",X"68",X"DA",X"66",X"AB",X"5B",X"44",X"5D",X"E0",X"56",X"44",X"5D",X"E0",X"56",X"44",X"5D",
		X"E0",X"56",X"44",X"5D",X"79",X"58",X"73",X"68",X"DA",X"66",X"0C",X"6A",X"A5",X"6B",X"41",X"65",
		X"A8",X"63",X"47",X"55",X"79",X"58",X"47",X"55",X"E0",X"56",X"79",X"58",X"47",X"55",X"79",X"58",
		X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",X"63",X"73",X"68",X"DA",X"66",X"41",X"65",X"A8",X"63",
		X"73",X"68",X"DA",X"66",X"06",X"7A",X"41",X"65",X"A8",X"63",X"47",X"55",X"E0",X"56",X"E0",X"56",
		X"E0",X"56",X"E0",X"56",X"E0",X"56",X"E0",X"56",X"E0",X"56",X"79",X"58",X"AE",X"53",X"47",X"55",
		X"E0",X"56",X"38",X"7D",X"35",X"7F",X"4E",X"7F",X"35",X"7F",X"4E",X"7F",X"35",X"7F",X"19",X"01",
		X"01",X"01",X"0E",X"06",X"18",X"22",X"01",X"01",X"14",X"01",X"01",X"01",X"01",X"01",X"18",X"01",
		X"10",X"01",X"17",X"01",X"01",X"01",X"0A",X"08",X"03",X"08",X"03",X"08",X"0A",X"01",X"01",X"01",
		X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"15",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"15",X"01",X"15",X"01",X"15",X"01",X"49",
		X"01",X"1B",X"01",X"1A",X"01",X"02",X"43",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"70",X"F9",X"A2",
		X"F3",X"7B",X"79",X"80",X"95",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FD",X"F3",X"F3",X"A2",X"7A",X"78",X"96",X"94",X"FE",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A2",X"A2",
		X"F9",X"7F",X"7D",X"77",X"75",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F3",X"F9",X"7E",X"7C",X"76",X"74",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",
		X"F3",X"F3",X"F9",X"A2",X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"A2",X"F9",X"F3",X"F9",X"F3",X"F9",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",
		X"A2",X"F3",X"F9",X"F3",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"F3",X"F3",X"A2",X"F9",X"F3",X"A2",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"7B",
		X"79",X"80",X"95",X"F9",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"7A",X"78",X"96",X"94",X"F9",X"A2",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"7F",
		X"7D",X"77",X"75",X"F3",X"F9",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"7E",X"7C",X"76",X"74",X"F9",X"F3",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"A2",
		X"F3",X"F9",X"F3",X"A2",X"F9",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"F3",X"A2",X"F3",X"A2",X"F3",X"F3",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",
		X"F9",X"F3",X"F9",X"F3",X"A2",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FE",X"F3",X"F3",X"A2",X"F9",X"F9",X"F3",X"A2",X"FC",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"04",X"43",
		X"43",X"43",X"43",X"43",X"43",X"43",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"70",X"F3",X"F3",X"F3",X"F9",X"F9",X"F3",X"A2",X"FC",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"F3",
		X"F3",X"F9",X"A2",X"F9",X"F3",X"F4",X"FA",X"05",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"F9",X"F3",X"F9",X"F9",X"F9",X"F3",X"F5",X"FB",X"04",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",
		X"F3",X"F3",X"F9",X"F3",X"F9",X"F6",X"08",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",X"F9",X"F3",X"F9",X"F0",X"F7",X"07",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",
		X"F3",X"F3",X"F9",X"F9",X"F1",X"F8",X"06",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",X"F9",X"F3",X"EE",X"F2",X"0A",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",
		X"F3",X"F3",X"EC",X"EF",X"0B",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F3",X"E9",X"ED",X"0B",X"09",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"F9",
		X"E5",X"EA",X"0D",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"E6",X"EB",X"0C",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"E1",
		X"E7",X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"E2",X"E8",X"0E",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"E3",
		X"11",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"E4",X"10",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"01",X"60",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"70",
		X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",
		X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",
		X"91",X"69",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"91",X"92",X"69",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"92",
		X"51",X"69",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"51",X"51",X"69",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"51",
		X"51",X"69",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"51",X"51",X"69",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"51",
		X"93",X"69",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"93",X"91",X"69",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"69",X"91",
		X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",
		X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",X"90",X"2C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"2C",X"90",
		X"05",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"70",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"E4",X"10",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"E3",X"11",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"E2",X"E8",X"0E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"E1",X"E7",X"0F",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"A2",X"E6",X"EB",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"E5",X"EA",X"0D",X"09",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"F3",X"A2",X"E9",X"ED",X"0B",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"F9",X"F9",X"F3",X"EC",X"EF",X"0B",X"09",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"A2",X"F3",X"F9",X"F3",X"EE",X"F2",X"0A",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F3",X"A2",X"F9",X"A2",X"F1",X"F8",
		X"06",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"F9",X"F9",X"A2",X"F3",X"F9",X"F0",X"F7",X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F3",X"F3",X"A2",X"F3",X"F3",X"F6",
		X"F8",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FF",X"F9",X"A2",X"A2",X"F9",X"F9",X"F9",X"F5",X"FB",X"04",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"F3",X"F9",X"F3",X"F3",X"A2",X"F4",
		X"FA",X"05",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"FE",X"F3",X"A2",X"F3",X"F9",X"A2",X"F9",X"F3",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"09",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"51",X"51",X"51",X"51",X"51",X"00",X"A7",X"A7",X"FE",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"51",X"51",X"51",X"51",X"51",X"00",
		X"B5",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",X"B4",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",
		X"B3",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",X"B2",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",
		X"B1",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"51",X"51",X"51",X"51",X"51",X"00",X"B0",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"51",X"51",X"51",X"51",X"51",X"00",
		X"AF",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"51",X"51",X"51",X"6D",X"6C",X"00",X"A7",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5A",X"5B",X"59",X"6A",X"6B",X"00",
		X"AE",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"59",X"59",X"59",X"51",X"51",X"00",X"AD",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",
		X"AC",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",X"AB",X"A7",X"FF",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"51",X"51",X"51",X"51",X"51",X"00",
		X"AA",X"A7",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"51",X"51",X"51",X"51",X"51",X"00",X"A9",X"A7",X"FC",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"51",X"51",X"51",X"51",X"51",X"00",
		X"A8",X"A7",X"06",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"50",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"FD",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"F3",X"A2",X"F9",X"F9",
		X"A2",X"A2",X"F3",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"2D",X"01",X"01",X"01",X"01",
		X"01",X"01",X"05",X"FA",X"F4",X"F3",X"F3",X"F9",X"A2",X"F3",X"A2",X"FF",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"2E",X"34",X"01",X"01",X"01",X"01",X"01",X"04",X"FB",X"F5",X"F3",X"A2",X"F9",
		X"F3",X"F3",X"F9",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"2F",X"35",X"01",X"01",X"01",
		X"01",X"01",X"03",X"08",X"F6",X"A2",X"F9",X"F3",X"A2",X"F3",X"F9",X"FF",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"30",X"36",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"F7",X"F0",X"F3",X"F3",
		X"A2",X"F9",X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"31",X"37",X"3C",X"01",X"01",
		X"01",X"01",X"01",X"06",X"F8",X"F1",X"F3",X"A2",X"A2",X"F9",X"F3",X"FF",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"32",X"38",X"3D",X"42",X"01",X"01",X"01",X"01",X"01",X"0A",X"F2",X"EE",X"F3",
		X"F9",X"A2",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"30",X"39",X"3E",X"3D",X"42",
		X"01",X"01",X"01",X"01",X"09",X"0B",X"EF",X"EC",X"F3",X"F9",X"F9",X"FE",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"31",X"3A",X"39",X"3E",X"3D",X"42",X"01",X"01",X"01",X"01",X"09",X"0B",X"ED",
		X"E9",X"A2",X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"32",X"3F",X"3A",X"39",X"3E",
		X"43",X"01",X"01",X"01",X"01",X"01",X"09",X"0D",X"EA",X"E5",X"F9",X"FF",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"30",X"39",X"3F",X"3A",X"39",X"44",X"45",X"01",X"01",X"01",X"01",X"01",X"0C",
		X"EB",X"E6",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"31",X"3A",X"39",X"3F",X"3A",
		X"39",X"46",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"E7",X"E1",X"FF",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"32",X"3F",X"3A",X"39",X"3F",X"3A",X"47",X"49",X"01",X"01",X"01",X"01",X"01",
		X"0E",X"E8",X"E2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"30",X"39",X"3F",X"3A",X"39",
		X"3F",X"48",X"4A",X"01",X"01",X"01",X"01",X"01",X"01",X"11",X"E3",X"FF",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"31",X"3A",X"39",X"3F",X"3A",X"39",X"3F",X"4B",X"01",X"01",X"01",X"01",X"01",
		X"01",X"10",X"E4",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"33",X"3B",X"40",X"41",X"3B",
		X"40",X"41",X"33",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"1A",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"63",X"63",X"63",X"63",X"63",X"63",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8F",X"8A",X"8A",
		X"8A",X"8A",X"88",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8D",X"81",X"82",X"81",X"81",X"86",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8E",X"82",X"81",
		X"82",X"83",X"85",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8C",X"81",X"83",X"82",X"82",X"86",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8D",X"82",X"81",
		X"83",X"83",X"87",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8E",X"81",X"82",X"82",X"81",X"85",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FF",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8C",X"82",X"83",
		X"81",X"82",X"86",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"FC",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8D",X"83",X"82",X"82",X"83",X"87",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FC",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8E",X"81",X"82",
		X"83",X"81",X"85",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"FE",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8C",X"82",X"81",X"82",X"83",X"87",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FE",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8E",X"83",X"81",
		X"81",X"81",X"86",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8D",X"81",X"83",X"82",X"82",X"87",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8E",X"83",X"82",
		X"82",X"83",X"85",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8C",X"81",X"81",X"81",X"81",X"87",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"8C",X"81",X"83",
		X"82",X"82",X"85",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"8B",X"89",X"89",X"89",X"89",X"84",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"FF",X"07",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"53",X"53",X"53",
		X"53",X"53",X"53",X"53",X"53",X"53",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",X"A2",X"F3",X"F9",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"FC",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"05",X"FA",X"F4",
		X"F3",X"F9",X"A2",X"F3",X"4C",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"04",X"FB",X"F5",X"F9",X"F9",X"A2",X"F3",X"39",X"3A",X"09",X"01",
		X"01",X"01",X"01",X"01",X"01",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"08",X"F6",
		X"A2",X"F9",X"A2",X"A2",X"F3",X"39",X"3F",X"09",X"01",X"01",X"01",X"01",X"01",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"F7",X"F0",X"F3",X"A2",X"F9",X"F9",X"F3",X"39",X"3F",
		X"09",X"01",X"01",X"01",X"01",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"06",X"F8",
		X"F1",X"F9",X"F9",X"F3",X"A2",X"A2",X"A2",X"39",X"3F",X"09",X"01",X"01",X"01",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0A",X"F2",X"EE",X"F9",X"F9",X"F3",X"A2",X"F3",X"A2",
		X"39",X"4D",X"4E",X"4E",X"4E",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"09",
		X"0B",X"EF",X"EC",X"F9",X"F3",X"A2",X"F9",X"F3",X"A2",X"A2",X"F9",X"A2",X"F9",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"09",X"0B",X"ED",X"E9",X"F9",X"A2",X"F9",X"F3",
		X"A2",X"A2",X"F9",X"F3",X"F9",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"09",X"0D",X"EA",X"E5",X"A2",X"F9",X"F9",X"F3",X"F3",X"A2",X"F9",X"A2",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"EB",X"E6",X"F3",X"F3",X"F9",
		X"F9",X"A2",X"A2",X"F9",X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"0F",X"E7",X"E1",X"A2",X"F9",X"A2",X"A2",X"F9",X"F9",X"F3",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0E",X"E8",X"E2",X"F9",X"F3",
		X"F9",X"A2",X"F3",X"F3",X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"11",X"E3",X"F3",X"F9",X"A2",X"F9",X"F9",X"A2",X"F3",X"FE",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"10",X"F4",X"F9",X"A2",
		X"A2",X"A2",X"F9",X"F3",X"F3",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FC",X"A2",X"A2",X"F9",X"F3",X"F9",X"F9",X"F3",X"16",X"A4",X"A4",
		X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",
		X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"04",X"03",X"01",X"07",X"05",X"04",X"08",X"09",X"0A",X"0B",
		X"08",X"04",X"0A",X"09",X"0B",X"04",X"04",X"0B",X"0A",X"09",X"08",X"04",X"0B",X"03",X"08",X"FF",
		X"FD",X"FA",X"F8",X"09",X"0B",X"0A",X"04",X"09",X"04",X"08",X"04",X"0B",X"04",X"09",X"08",X"0A",
		X"08",X"04",X"09",X"0E",X"0C",X"FF",X"09",X"FE",X"FC",X"F7",X"F5",X"04",X"0B",X"09",X"08",X"04",
		X"08",X"09",X"0A",X"0B",X"0A",X"0A",X"09",X"04",X"0B",X"08",X"08",X"04",X"0B",X"FE",X"0A",X"02",
		X"F9",X"F6",X"06",X"0E",X"0C",X"04",X"0A",X"0B",X"08",X"04",X"0A",X"09",X"0B",X"04",X"04",X"0B",
		X"0A",X"03",X"01",X"07",X"05",X"02",X"03",X"01",X"07",X"05",X"03",X"01",X"07",X"05",X"09",X"04",
		X"08",X"04",X"0B",X"04",X"09",X"08",X"0A",X"08",X"04",X"FF",X"FD",X"FA",X"F8",X"08",X"FF",X"FD",
		X"FA",X"F8",X"FF",X"FD",X"FA",X"F8",X"0B",X"09",X"08",X"04",X"08",X"09",X"0A",X"0B",X"0A",X"0A",
		X"09",X"FE",X"FC",X"F7",X"F5",X"04",X"FE",X"FC",X"F7",X"F5",X"FE",X"FC",X"F7",X"F5",X"04",X"0A",
		X"0B",X"08",X"04",X"0A",X"09",X"0B",X"04",X"04",X"0B",X"02",X"F9",X"F6",X"06",X"0A",X"02",X"F9",
		X"F6",X"06",X"02",X"F9",X"F6",X"06",X"0E",X"0C",X"09",X"04",X"08",X"04",X"0B",X"04",X"09",X"03",
		X"01",X"07",X"05",X"09",X"08",X"04",X"04",X"03",X"01",X"07",X"05",X"0A",X"04",X"08",X"09",X"04",
		X"08",X"04",X"08",X"09",X"0A",X"0B",X"0A",X"FF",X"FD",X"FA",X"F8",X"04",X"08",X"0B",X"08",X"FF",
		X"FD",X"FA",X"F8",X"0B",X"0A",X"09",X"04",X"0B",X"0A",X"0B",X"08",X"04",X"0A",X"09",X"0B",X"FE",
		X"FC",X"F7",X"F5",X"08",X"0E",X"0C",X"09",X"FE",X"FC",X"F7",X"F5",X"04",X"09",X"0B",X"0A",X"08",
		X"04",X"08",X"04",X"0B",X"04",X"09",X"08",X"02",X"F9",X"F6",X"06",X"0A",X"0B",X"09",X"0A",X"02",
		X"F9",X"F6",X"06",X"08",X"09",X"0A",X"04",X"09",X"08",X"04",X"08",X"09",X"0A",X"0B",X"0A",X"04",
		X"04",X"0B",X"09",X"0E",X"0C",X"08",X"0C",X"04",X"0E",X"0C",X"08",X"09",X"08",X"0E",X"0C",X"0A",
		X"0B",X"08",X"04",X"0A",X"09",X"0B",X"09",X"04",X"0E",X"0C",X"08",X"0A",X"0B",X"0E",X"0E",X"0C",
		X"04",X"03",X"01",X"07",X"05",X"0E",X"0C",X"04",X"08",X"04",X"0B",X"04",X"09",X"08",X"0A",X"04",
		X"08",X"0A",X"0E",X"0C",X"09",X"08",X"01",X"07",X"05",X"FF",X"FD",X"FA",X"F8",X"09",X"0E",X"0C",
		X"08",X"04",X"08",X"09",X"0A",X"0B",X"0A",X"04",X"04",X"0B",X"09",X"0A",X"04",X"0E",X"FD",X"FA",
		X"F8",X"FE",X"FC",X"F7",X"F5",X"08",X"0E",X"0C",X"09",X"08",X"09",X"0A",X"0B",X"0A",X"04",X"04",
		X"0B",X"09",X"0E",X"0C",X"04",X"08",X"16",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",
		X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"FC",
		X"F7",X"F5",X"02",X"F9",X"F6",X"06",X"0E",X"0C",X"04",X"08",X"0A",X"0B",X"04",X"08",X"08",X"09",
		X"0A",X"04",X"08",X"09",X"0E",X"0C",X"04",X"F9",X"F6",X"03",X"01",X"07",X"05",X"0E",X"0C",X"09",
		X"0A",X"0B",X"04",X"09",X"09",X"04",X"04",X"08",X"0A",X"0B",X"08",X"04",X"09",X"09",X"0A",X"04",
		X"04",X"FF",X"FD",X"FA",X"F8",X"08",X"08",X"04",X"04",X"09",X"09",X"0A",X"0A",X"0B",X"0B",X"04",
		X"04",X"08",X"08",X"09",X"09",X"03",X"01",X"0C",X"09",X"FE",X"FC",X"F7",X"F5",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"04",X"04",X"04",X"09",X"09",X"09",X"03",X"03",X"03",X"09",X"FF",X"FD",X"0E",
		X"0C",X"02",X"F9",X"F6",X"06",X"04",X"08",X"0A",X"0B",X"04",X"08",X"08",X"09",X"0A",X"04",X"08",
		X"09",X"04",X"08",X"0A",X"0B",X"FE",X"FC",X"0C",X"09",X"0A",X"0B",X"04",X"09",X"09",X"04",X"04",
		X"08",X"0A",X"0B",X"08",X"04",X"09",X"09",X"0A",X"04",X"08",X"0B",X"09",X"04",X"02",X"F9",X"04",
		X"0E",X"0C",X"09",X"08",X"04",X"0A",X"0B",X"09",X"04",X"0B",X"0A",X"08",X"08",X"0E",X"0C",X"09",
		X"08",X"0A",X"04",X"04",X"03",X"01",X"07",X"0B",X"0A",X"0E",X"0C",X"09",X"0A",X"0B",X"04",X"09",
		X"09",X"04",X"04",X"08",X"03",X"01",X"07",X"05",X"08",X"09",X"04",X"08",X"FF",X"FD",X"FA",X"01",
		X"07",X"05",X"0B",X"04",X"04",X"08",X"0A",X"0B",X"04",X"08",X"04",X"09",X"FF",X"FD",X"FA",X"F8",
		X"08",X"04",X"0A",X"0B",X"FE",X"FC",X"F7",X"FD",X"FA",X"F8",X"0A",X"0B",X"0A",X"04",X"08",X"04",
		X"0A",X"0B",X"09",X"04",X"FE",X"FC",X"F7",X"F5",X"09",X"04",X"08",X"04",X"02",X"F9",X"F6",X"FC",
		X"F7",X"F5",X"09",X"0A",X"0B",X"04",X"09",X"09",X"04",X"08",X"0E",X"0C",X"02",X"F9",X"F6",X"06",
		X"0A",X"0B",X"04",X"03",X"01",X"07",X"05",X"F9",X"F6",X"06",X"08",X"0B",X"04",X"04",X"08",X"0A",
		X"0B",X"04",X"08",X"03",X"01",X"07",X"05",X"04",X"08",X"09",X"0A",X"FF",X"FD",X"FA",X"F8",X"04",
		X"08",X"0A",X"0B",X"0B",X"09",X"0A",X"08",X"03",X"01",X"07",X"05",X"FF",X"FD",X"FA",X"F8",X"0B",
		X"0B",X"0A",X"04",X"FE",X"FC",X"F7",X"F5",X"0B",X"0A",X"09",X"0A",X"04",X"08",X"0B",X"0B",X"FF",
		X"FD",X"FA",X"F8",X"FE",X"FC",X"F7",X"F5",X"04",X"08",X"09",X"0A",X"02",X"F9",X"F6",X"06",X"04",
		X"08",X"09",X"0A",X"0B",X"0A",X"0B",X"08",X"FE",X"FC",X"F7",X"F5",X"02",X"F9",X"F6",X"06",X"0A",
		X"09",X"0B",X"0B",X"0A",X"04",X"0E",X"0C",X"0E",X"0C",X"04",X"08",X"09",X"0A",X"0B",X"04",X"02",
		X"F9",X"F6",X"06",X"0A",X"0B",X"0E",X"0C",X"09",X"08",X"04",X"0A",X"0E",X"0C",X"0B",X"0A",X"0A",
		X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",
		X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"53",X"F3",X"F9",X"A2",X"B8",X"29",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"28",X"B9",X"BA",X"A2",X"F3",
		X"F9",X"F9",X"A2",X"B7",X"2A",X"2B",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"27",X"26",X"BB",X"F9",X"A2",X"A2",X"F3",X"F3",X"CA",X"CC",X"1F",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"25",X"BC",X"F3",X"F3",
		X"A2",X"A2",X"F9",X"CB",X"CD",X"1E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"17",X"BD",X"BF",X"F9",X"F3",X"F9",X"F9",X"A2",X"CE",X"1D",X"1C",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"22",X"BE",X"C0",X"F3",
		X"F9",X"A2",X"F3",X"F9",X"CF",X"D1",X"1B",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"24",X"23",X"C1",X"A2",X"F3",X"F3",X"F9",X"A2",X"D0",X"D2",X"1A",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"18",X"C2",X"F9",
		X"A2",X"A2",X"F3",X"F9",X"F3",X"D3",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"17",X"C3",X"C5",X"A2",X"F9",X"F9",X"F3",X"F9",X"D4",X"16",X"15",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"22",X"C4",X"C6",
		X"F9",X"F3",X"A2",X"A2",X"F3",X"D5",X"D7",X"19",X"01",X"01",X"01",X"01",X"01",X"24",X"19",X"01",
		X"01",X"01",X"01",X"01",X"01",X"21",X"20",X"C7",X"F3",X"A2",X"F9",X"F9",X"A2",X"D6",X"D8",X"18",
		X"01",X"01",X"01",X"01",X"01",X"01",X"18",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"C8",
		X"A2",X"A2",X"F3",X"F9",X"F3",X"F9",X"D9",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"17",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"C9",X"F9",X"F3",X"A2",X"F3",X"F9",X"A2",X"DA",X"16",
		X"15",X"01",X"01",X"01",X"01",X"01",X"22",X"15",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",
		X"F3",X"F3",X"F3",X"F3",X"F9",X"A2",X"DB",X"DE",X"14",X"01",X"01",X"01",X"01",X"01",X"21",X"14",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"A2",X"F3",X"F9",X"F9",X"A2",X"DC",X"DF",
		X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",
		X"F9",X"F3",X"F3",X"A2",X"F9",X"F9",X"DD",X"E0",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"12",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"0A",X"63",X"73",X"73",X"73",X"73",X"73",X"73",
		X"73",X"73",X"73",X"73",X"73",X"43",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"63",X"53",
		X"43",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"12",X"E0",X"DD",X"F3",X"F3",X"F9",X"A2",X"A2",X"F9",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"DF",X"DC",X"F9",X"A2",X"F3",X"F9",X"F9",
		X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"14",X"DE",X"DB",X"F9",X"F9",X"A2",X"F3",X"A2",X"A2",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"15",X"16",X"DA",X"A2",X"F3",X"F9",X"F9",X"A2",
		X"F3",X"C9",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"17",X"D9",X"F3",X"F3",X"A2",X"F9",X"A2",X"A2",X"C8",X"13",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"18",X"D8",X"D6",X"F9",X"F9",X"F3",X"F9",
		X"F3",X"C7",X"20",X"21",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"19",X"D7",X"D5",X"A2",X"F9",X"A2",X"F3",X"F3",X"C6",X"C4",X"22",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"15",X"16",X"D4",X"F9",X"F3",X"F9",X"F3",
		X"F3",X"C5",X"C3",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"17",X"D3",X"A2",X"A2",X"F9",X"F9",X"A2",X"F9",X"C2",X"18",X"01",X"01",X"01",X"01",
		X"01",X"01",X"15",X"22",X"01",X"01",X"01",X"01",X"01",X"01",X"1A",X"D2",X"D0",X"F3",X"F3",X"F3",
		X"F3",X"A2",X"C1",X"23",X"24",X"01",X"01",X"01",X"01",X"01",X"01",X"17",X"01",X"01",X"01",X"01",
		X"01",X"01",X"1B",X"D1",X"CF",X"F9",X"A2",X"F3",X"A2",X"F3",X"C0",X"BE",X"22",X"01",X"01",X"01",
		X"01",X"01",X"01",X"25",X"01",X"01",X"01",X"01",X"01",X"01",X"1C",X"1D",X"CE",X"F3",X"F9",X"F9",
		X"A2",X"F9",X"BF",X"BD",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"1B",X"27",X"01",X"01",X"01",
		X"01",X"01",X"01",X"1E",X"CD",X"CB",X"A2",X"F9",X"F3",X"F3",X"A2",X"BC",X"25",X"01",X"01",X"01",
		X"01",X"01",X"01",X"1C",X"28",X"01",X"01",X"01",X"01",X"01",X"01",X"1F",X"CC",X"CA",X"A2",X"F9",
		X"F9",X"A2",X"F9",X"BB",X"26",X"27",X"01",X"01",X"01",X"01",X"01",X"01",X"1E",X"01",X"01",X"01",
		X"01",X"01",X"01",X"2B",X"2A",X"B7",X"F9",X"A2",X"F9",X"F3",X"F9",X"BA",X"B9",X"28",X"01",X"01",
		X"01",X"01",X"01",X"01",X"1F",X"2B",X"01",X"01",X"01",X"01",X"01",X"01",X"29",X"B8",X"F9",X"F9",
		X"A2",X"0B",X"43",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",
		X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"43",X"53",X"73",X"F3",X"A2",X"BA",X"B9",X"28",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"29",X"B8",X"F3",
		X"F9",X"F9",X"F9",X"F3",X"BB",X"26",X"27",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"2B",X"2A",X"B7",X"F9",X"A2",X"F3",X"A2",X"F9",X"BC",X"25",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1F",X"CC",X"CA",X"F9",
		X"F3",X"F9",X"F9",X"BF",X"BD",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"1E",X"CD",X"CB",X"F3",X"A2",X"F9",X"F3",X"C0",X"BE",X"22",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1C",X"1D",X"CE",X"A2",X"F9",
		X"A2",X"F3",X"F3",X"C1",X"23",X"24",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"1B",X"D1",X"CF",X"F9",X"F3",X"F3",X"A2",X"A2",X"C2",X"18",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1A",X"D2",X"D0",X"F9",X"A2",
		X"A2",X"F9",X"C5",X"C3",X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"17",X"D3",X"F9",X"A2",X"F3",X"A2",X"F3",X"C6",X"C4",X"22",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"15",X"16",X"D4",X"A2",X"F3",X"F9",
		X"F9",X"F3",X"C7",X"20",X"21",X"01",X"01",X"01",X"01",X"01",X"01",X"19",X"24",X"01",X"01",X"01",
		X"01",X"01",X"19",X"D7",X"D5",X"F9",X"A2",X"F3",X"F9",X"A2",X"C8",X"13",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"18",X"01",X"01",X"01",X"01",X"01",X"01",X"18",X"D8",X"D6",X"F9",X"F3",X"F3",
		X"A2",X"F9",X"C9",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"17",X"01",X"01",X"01",X"01",
		X"01",X"01",X"17",X"D9",X"F3",X"F9",X"A2",X"F9",X"A2",X"F9",X"FC",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"15",X"22",X"01",X"01",X"01",X"01",X"01",X"15",X"16",X"DA",X"F3",X"A2",X"F3",X"F9",
		X"F9",X"A2",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"14",X"21",X"01",X"01",X"01",X"01",
		X"01",X"14",X"DE",X"DB",X"F9",X"F9",X"F3",X"A2",X"A2",X"F9",X"FE",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"DF",X"DC",X"F3",X"F3",X"A2",X"F3",
		X"F9",X"A2",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"01",
		X"01",X"12",X"E0",X"DD",X"A2",X"F3",X"F9",X"F9",X"A2",X"F3",X"0B",X"43",X"53",X"73",X"63",X"63",
		X"63",X"63",X"63",X"63",X"63",X"63",X"53",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",
		X"63",X"63",X"73",X"F3",X"A2",X"F9",X"F3",X"F3",X"A2",X"DD",X"E0",X"12",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"F9",X"F3",X"F3",X"A2",X"F9",
		X"F9",X"DC",X"DF",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"FE",X"A2",X"F9",X"A2",X"F9",X"F3",X"A2",X"DB",X"DE",X"14",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"A2",X"F3",X"F3",X"F9",
		X"A2",X"DA",X"16",X"15",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"FC",X"F9",X"F9",X"F9",X"A2",X"F9",X"F3",X"D9",X"17",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"C9",X"A2",X"F3",X"A2",X"F3",X"F9",
		X"D6",X"D8",X"18",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"13",X"C8",X"F9",X"F3",X"F9",X"F9",X"F3",X"D5",X"D7",X"19",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"20",X"C7",X"F3",X"A2",X"F9",X"F3",X"A2",
		X"D4",X"16",X"15",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"22",X"C4",X"C6",X"A2",X"F3",X"F3",X"F9",X"F9",X"D3",X"17",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"17",X"C3",X"C5",X"F3",X"A2",X"A2",X"F3",X"D0",
		X"D2",X"1A",X"01",X"01",X"01",X"01",X"01",X"01",X"22",X"15",X"01",X"01",X"01",X"01",X"01",X"01",
		X"18",X"C2",X"A2",X"A2",X"F3",X"F9",X"F9",X"CF",X"D1",X"1B",X"01",X"01",X"01",X"01",X"01",X"01",
		X"17",X"01",X"01",X"01",X"01",X"01",X"01",X"24",X"23",X"C1",X"F9",X"F3",X"F9",X"A2",X"F3",X"CE",
		X"1D",X"1C",X"01",X"01",X"01",X"01",X"01",X"01",X"25",X"01",X"01",X"01",X"01",X"01",X"01",X"22",
		X"BE",X"C0",X"F3",X"F9",X"A2",X"F3",X"CB",X"CD",X"1E",X"01",X"01",X"01",X"01",X"01",X"01",X"27",
		X"1B",X"01",X"01",X"01",X"01",X"01",X"01",X"17",X"BD",X"BF",X"F9",X"F3",X"A2",X"F9",X"CA",X"CC",
		X"1F",X"01",X"01",X"01",X"01",X"01",X"01",X"28",X"1C",X"01",X"01",X"01",X"01",X"01",X"01",X"25",
		X"BC",X"F3",X"A2",X"F9",X"F9",X"A2",X"B7",X"2A",X"2B",X"01",X"01",X"01",X"01",X"01",X"01",X"1E",
		X"01",X"01",X"01",X"01",X"01",X"01",X"27",X"26",X"BB",X"A2",X"F9",X"A2",X"F3",X"F3",X"B8",X"29",
		X"01",X"01",X"01",X"01",X"01",X"01",X"2B",X"1F",X"01",X"01",X"01",X"01",X"01",X"01",X"28",X"B9",
		X"BA",X"F9",X"F3",X"0E",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"72",X"72",X"76",X"76",X"76",X"76",X"76",X"FD",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"A1",X"9C",X"98",
		X"98",X"98",X"99",X"5C",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"FE",X"A0",X"9E",X"98",X"98",X"98",X"9A",X"5C",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A0",X"9C",X"98",
		X"98",X"9B",X"5C",X"5C",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"FF",X"9F",X"9D",X"98",X"98",X"9A",X"5C",X"5C",X"FF",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A1",X"9E",X"9A",
		X"9A",X"9A",X"5C",X"5D",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"FF",X"A0",X"9D",X"98",X"9B",X"5C",X"5C",X"5E",X"FE",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A0",X"9D",X"98",
		X"99",X"5C",X"5D",X"5E",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"FC",X"9F",X"9E",X"9B",X"5C",X"5C",X"5E",X"5F",X"B6",X"50",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"50",X"B6",X"A1",X"9C",X"99",
		X"5E",X"5E",X"5E",X"61",X"B6",X"52",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"52",X"B6",X"A0",X"9D",X"9A",X"5C",X"5C",X"5F",X"62",X"B6",X"4F",X"53",X"54",
		X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"53",X"4F",X"B6",X"A0",X"9E",X"99",
		X"5C",X"5C",X"60",X"64",X"B6",X"4F",X"4F",X"4F",X"55",X"56",X"00",X"00",X"00",X"00",X"00",X"56",
		X"55",X"4F",X"4F",X"4F",X"B6",X"9F",X"9C",X"9B",X"5C",X"5D",X"61",X"63",X"B6",X"57",X"58",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"B6",X"A1",X"9C",X"9A",
		X"5C",X"5E",X"60",X"62",X"B6",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"B6",X"A0",X"9E",X"9B",X"5C",X"5F",X"64",X"65",X"B6",X"4F",X"4F",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"B6",X"A0",X"9D",X"99",
		X"5C",X"61",X"63",X"65",X"B6",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"B6",X"9F",X"9C",X"99",X"5C",X"61",X"62",X"65",X"03",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"70",X"43",X"63",
		X"63",X"63",X"63",X"63",X"63",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FD",X"F9",X"7B",X"79",X"80",X"95",X"F3",X"F9",X"FE",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A2",X"7A",
		X"78",X"96",X"94",X"A2",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"7F",X"7D",X"77",X"75",X"F9",X"F9",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"7E",
		X"7C",X"76",X"74",X"A2",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"A2",X"F3",X"F9",X"A2",X"F3",X"A2",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"F9",
		X"A2",X"A2",X"F9",X"F9",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"F3",X"F3",X"F9",X"7B",X"79",X"80",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",
		X"A2",X"F9",X"7A",X"78",X"96",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"F3",X"F3",X"F9",X"7F",X"7D",X"77",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"F9",
		X"A2",X"F3",X"7E",X"7C",X"76",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"F3",X"F9",X"A2",X"F3",X"F3",X"F9",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"F9",
		X"A2",X"F9",X"F9",X"A2",X"F3",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",X"F9",X"F3",X"A2",X"A2",X"F3",X"F9",X"FF",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"A2",
		X"F9",X"F3",X"F9",X"A2",X"A2",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"FE",X"A2",X"F9",X"F9",X"A2",X"F3",X"F3",X"F9",X"FC",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"F9",X"F3",
		X"A2",X"A2",X"F9",X"F3",X"A2",X"12",X"01",X"21",X"11",X"31",X"01",X"31",X"21",X"31",X"11",X"01",
		X"21",X"02",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"11",X"21",X"31",X"11",X"62",X"63",
		X"99",X"62",X"99",X"62",X"63",X"99",X"63",X"63",X"72",X"6E",X"6F",X"82",X"83",X"82",X"85",X"81",
		X"83",X"8A",X"72",X"63",X"62",X"63",X"63",X"63",X"62",X"63",X"63",X"62",X"99",X"63",X"63",X"63",
		X"75",X"6E",X"6F",X"82",X"8A",X"81",X"82",X"8A",X"85",X"81",X"76",X"62",X"63",X"99",X"62",X"63",
		X"63",X"99",X"62",X"63",X"63",X"62",X"63",X"63",X"72",X"6E",X"6F",X"85",X"83",X"82",X"8A",X"81",
		X"8A",X"83",X"75",X"62",X"63",X"62",X"63",X"62",X"63",X"63",X"62",X"99",X"62",X"63",X"63",X"62",
		X"77",X"6E",X"6F",X"85",X"82",X"81",X"82",X"85",X"83",X"8A",X"72",X"63",X"99",X"99",X"63",X"63",
		X"62",X"63",X"99",X"62",X"63",X"99",X"62",X"63",X"76",X"6E",X"6F",X"81",X"85",X"82",X"8A",X"8A",
		X"83",X"82",X"77",X"63",X"99",X"63",X"63",X"63",X"63",X"63",X"63",X"62",X"99",X"63",X"63",X"63",
		X"72",X"6E",X"6F",X"82",X"83",X"82",X"85",X"8A",X"85",X"83",X"76",X"62",X"62",X"62",X"63",X"99",
		X"99",X"62",X"62",X"99",X"99",X"63",X"62",X"63",X"75",X"6E",X"6F",X"81",X"8A",X"82",X"85",X"83",
		X"82",X"81",X"75",X"63",X"99",X"99",X"63",X"62",X"63",X"63",X"99",X"62",X"62",X"63",X"63",X"63",
		X"76",X"6E",X"6F",X"82",X"82",X"83",X"8A",X"81",X"85",X"83",X"77",X"63",X"62",X"63",X"63",X"63",
		X"63",X"62",X"63",X"62",X"99",X"63",X"62",X"63",X"77",X"6E",X"6F",X"83",X"82",X"81",X"82",X"83",
		X"83",X"8A",X"72",X"99",X"62",X"62",X"63",X"63",X"63",X"63",X"99",X"63",X"62",X"63",X"63",X"63",
		X"75",X"6E",X"6F",X"82",X"82",X"85",X"85",X"83",X"82",X"8A",X"72",X"62",X"99",X"63",X"62",X"99",
		X"62",X"63",X"63",X"62",X"99",X"63",X"63",X"99",X"72",X"6E",X"6F",X"83",X"8A",X"82",X"82",X"82",
		X"81",X"81",X"76",X"99",X"63",X"99",X"63",X"63",X"63",X"99",X"62",X"63",X"63",X"63",X"62",X"63",
		X"72",X"6E",X"6F",X"8A",X"81",X"81",X"82",X"83",X"82",X"85",X"77",X"99",X"63",X"62",X"63",X"62",
		X"63",X"62",X"63",X"62",X"62",X"99",X"63",X"63",X"75",X"6E",X"6F",X"82",X"83",X"82",X"8A",X"81",
		X"85",X"83",X"75",X"62",X"99",X"63",X"62",X"63",X"99",X"63",X"63",X"99",X"99",X"62",X"63",X"63",
		X"76",X"6E",X"6F",X"82",X"85",X"8A",X"82",X"85",X"83",X"82",X"77",X"63",X"74",X"99",X"63",X"62",
		X"63",X"63",X"99",X"62",X"63",X"63",X"63",X"63",X"77",X"6E",X"6F",X"85",X"83",X"83",X"82",X"82",
		X"85",X"85",X"76",X"63",X"99",X"62",X"63",X"63",X"62",X"63",X"62",X"63",X"99",X"62",X"63",X"99",
		X"75",X"6E",X"6F",X"81",X"83",X"82",X"85",X"82",X"8A",X"81",X"72",X"62",X"63",X"99",X"11",X"21",
		X"11",X"11",X"11",X"21",X"12",X"22",X"22",X"22",X"22",X"22",X"22",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"11",X"11",X"11",X"11",X"11",X"99",X"63",X"63",X"74",X"99",X"7A",X"7B",X"7A",X"7B",
		X"7B",X"85",X"6E",X"6F",X"83",X"82",X"83",X"82",X"83",X"8A",X"77",X"63",X"75",X"99",X"76",X"63",
		X"74",X"75",X"99",X"63",X"7A",X"7B",X"7A",X"7B",X"7A",X"C0",X"6E",X"6F",X"82",X"81",X"83",X"8A",
		X"82",X"83",X"75",X"99",X"63",X"99",X"63",X"61",X"61",X"61",X"61",X"61",X"8A",X"8A",X"8A",X"8A",
		X"C3",X"BF",X"7E",X"7C",X"82",X"8A",X"82",X"81",X"83",X"82",X"77",X"74",X"99",X"74",X"99",X"E1",
		X"DE",X"DC",X"DA",X"EF",X"9C",X"CE",X"CB",X"C7",X"C1",X"91",X"70",X"7D",X"7F",X"86",X"83",X"82",
		X"8A",X"83",X"76",X"99",X"63",X"77",X"74",X"E0",X"DD",X"DB",X"D9",X"FB",X"9C",X"9C",X"9C",X"C6",
		X"BD",X"91",X"70",X"71",X"91",X"87",X"8B",X"8D",X"82",X"81",X"72",X"63",X"75",X"76",X"99",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"9C",X"9C",X"CA",X"C5",X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"8E",
		X"8F",X"AE",X"74",X"74",X"99",X"63",X"63",X"DF",X"FB",X"FB",X"D8",X"EF",X"D2",X"CD",X"C9",X"91",
		X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"91",X"90",X"B2",X"80",X"79",X"74",X"63",X"75",X"FB",
		X"FB",X"FB",X"D7",X"D5",X"D1",X"CC",X"C8",X"91",X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"91",
		X"9D",X"AD",X"B7",X"D3",X"74",X"63",X"63",X"D4",X"D6",X"EE",X"D6",X"D4",X"D0",X"C2",X"91",X"91",
		X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"A3",X"A4",X"9C",X"B9",X"EA",X"73",X"6D",X"99",X"61",
		X"61",X"61",X"78",X"78",X"CF",X"90",X"91",X"91",X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"A2",
		X"A5",X"9C",X"FB",X"FB",X"ED",X"6C",X"63",X"99",X"63",X"99",X"63",X"74",X"BE",X"8F",X"8E",X"91",
		X"91",X"91",X"70",X"71",X"91",X"91",X"AB",X"A1",X"A6",X"9C",X"BA",X"FB",X"FB",X"F5",X"69",X"75",
		X"63",X"63",X"99",X"72",X"8A",X"85",X"8D",X"8B",X"87",X"91",X"70",X"71",X"91",X"B1",X"AA",X"A0",
		X"AC",X"B3",X"FB",X"EB",X"FB",X"F6",X"68",X"74",X"63",X"99",X"75",X"75",X"82",X"83",X"82",X"81",
		X"86",X"7F",X"7D",X"71",X"91",X"B0",X"A9",X"9C",X"9C",X"B4",X"BB",X"EC",X"F1",X"FB",X"F7",X"74",
		X"99",X"63",X"74",X"77",X"8A",X"85",X"82",X"83",X"82",X"81",X"7C",X"7E",X"B6",X"AF",X"A8",X"9C",
		X"9C",X"9C",X"BC",X"FB",X"F2",X"FB",X"F8",X"99",X"63",X"99",X"99",X"76",X"82",X"81",X"8A",X"85",
		X"82",X"83",X"6E",X"6F",X"B5",X"88",X"A7",X"9F",X"9C",X"9C",X"C4",X"FB",X"F3",X"FB",X"F9",X"74",
		X"63",X"99",X"63",X"75",X"8A",X"85",X"82",X"83",X"82",X"81",X"6E",X"6F",X"85",X"89",X"8C",X"9E",
		X"9C",X"9C",X"FB",X"FB",X"F4",X"FB",X"FA",X"10",X"11",X"11",X"11",X"11",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"02",X"12",X"21",X"11",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"99",X"63",X"63",X"72",X"8A",X"81",X"82",X"83",X"82",X"85",X"8A",X"6E",X"6F",X"72",X"75",X"8A",
		X"E5",X"FB",X"E2",X"E3",X"FB",X"E9",X"FB",X"E6",X"62",X"63",X"62",X"76",X"81",X"83",X"82",X"85",
		X"8A",X"82",X"81",X"6E",X"6F",X"75",X"72",X"8A",X"E5",X"FB",X"E2",X"FB",X"E9",X"E7",X"FB",X"E6",
		X"99",X"63",X"62",X"75",X"85",X"82",X"81",X"82",X"81",X"82",X"82",X"6E",X"6F",X"72",X"76",X"8A",
		X"E4",X"FB",X"E3",X"E2",X"E7",X"FB",X"FB",X"E8",X"63",X"99",X"63",X"72",X"82",X"83",X"82",X"8A",
		X"82",X"8A",X"82",X"6E",X"6F",X"77",X"77",X"8A",X"E4",X"FB",X"E2",X"FB",X"FB",X"E3",X"FB",X"E8",
		X"62",X"99",X"63",X"77",X"83",X"85",X"81",X"81",X"83",X"82",X"81",X"6E",X"6F",X"76",X"76",X"8A",
		X"E5",X"FB",X"E7",X"FB",X"FB",X"FB",X"FB",X"E6",X"99",X"62",X"62",X"76",X"82",X"8A",X"8A",X"85",
		X"83",X"82",X"83",X"6E",X"6F",X"72",X"75",X"8A",X"E4",X"FB",X"FB",X"FB",X"FB",X"E2",X"FB",X"E8",
		X"63",X"99",X"63",X"75",X"85",X"83",X"83",X"82",X"82",X"8A",X"81",X"6E",X"6F",X"75",X"77",X"8A",
		X"E5",X"FB",X"E2",X"E2",X"E7",X"FB",X"FB",X"E6",X"62",X"62",X"63",X"77",X"8A",X"8A",X"83",X"82",
		X"81",X"82",X"81",X"6E",X"6F",X"76",X"72",X"8A",X"E5",X"FB",X"E2",X"FB",X"FB",X"E9",X"FB",X"E6",
		X"63",X"62",X"99",X"72",X"81",X"82",X"83",X"81",X"8A",X"85",X"82",X"6E",X"6F",X"77",X"72",X"8A",
		X"E4",X"FB",X"E9",X"E3",X"E9",X"E7",X"FB",X"E8",X"63",X"63",X"62",X"72",X"83",X"83",X"82",X"82",
		X"83",X"82",X"81",X"6E",X"6F",X"75",X"76",X"8A",X"E5",X"FB",X"E2",X"E2",X"E7",X"E9",X"FB",X"E6",
		X"99",X"63",X"99",X"76",X"82",X"81",X"82",X"8A",X"83",X"83",X"82",X"6E",X"6F",X"72",X"77",X"8A",
		X"E4",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E6",X"62",X"99",X"99",X"77",X"85",X"85",X"82",X"83",
		X"85",X"82",X"82",X"6E",X"6F",X"72",X"75",X"8A",X"E4",X"FB",X"E3",X"FB",X"FB",X"E3",X"FB",X"E6",
		X"63",X"99",X"62",X"75",X"81",X"82",X"81",X"82",X"8A",X"8A",X"82",X"6E",X"6F",X"75",X"77",X"8A",
		X"E4",X"FB",X"E9",X"FB",X"E9",X"E2",X"FB",X"E8",X"99",X"74",X"63",X"77",X"83",X"81",X"82",X"82",
		X"81",X"83",X"85",X"6E",X"6F",X"76",X"76",X"8A",X"E5",X"FB",X"E2",X"E2",X"FB",X"FB",X"FB",X"E8",
		X"62",X"99",X"63",X"76",X"81",X"82",X"83",X"82",X"81",X"82",X"85",X"6E",X"6F",X"77",X"75",X"8A",
		X"E5",X"FB",X"E3",X"E3",X"E7",X"E9",X"FB",X"E6",X"99",X"63",X"62",X"72",X"85",X"8A",X"83",X"82",
		X"81",X"8A",X"81",X"6E",X"6F",X"75",X"72",X"8A",X"E4",X"FB",X"E2",X"FB",X"FB",X"E7",X"FB",X"E8",
		X"0D",X"01",X"31",X"31",X"31",X"01",X"32",X"02",X"02",X"02",X"02",X"02",X"02",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"31",X"31",X"31",X"31",X"31",X"74",X"63",X"99",X"63",X"75",X"8A",X"85",
		X"82",X"83",X"82",X"81",X"6E",X"6F",X"85",X"89",X"8C",X"9E",X"9C",X"9C",X"FB",X"FB",X"F4",X"FB",
		X"FA",X"99",X"63",X"99",X"99",X"76",X"82",X"81",X"8A",X"85",X"82",X"83",X"6E",X"6F",X"B5",X"88",
		X"A7",X"9F",X"9C",X"9C",X"C4",X"FB",X"F3",X"FB",X"F9",X"74",X"99",X"63",X"74",X"77",X"8A",X"85",
		X"82",X"83",X"82",X"81",X"7C",X"7E",X"B6",X"AF",X"A8",X"9C",X"9C",X"9C",X"BC",X"FB",X"F2",X"FB",
		X"F8",X"74",X"63",X"99",X"75",X"72",X"82",X"83",X"82",X"81",X"86",X"7F",X"7D",X"71",X"91",X"B0",
		X"A9",X"9C",X"9C",X"B4",X"BB",X"EC",X"F1",X"FB",X"F7",X"75",X"63",X"63",X"99",X"75",X"8A",X"8A",
		X"8D",X"8B",X"87",X"91",X"70",X"71",X"91",X"B1",X"AA",X"A0",X"AC",X"B3",X"FB",X"EB",X"FB",X"F6",
		X"68",X"99",X"63",X"99",X"63",X"74",X"BE",X"8F",X"8E",X"91",X"91",X"91",X"70",X"71",X"91",X"91",
		X"AB",X"A1",X"A6",X"9C",X"BA",X"FB",X"FB",X"F5",X"69",X"61",X"61",X"61",X"78",X"78",X"CF",X"90",
		X"91",X"91",X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"A2",X"A5",X"9C",X"FB",X"FB",X"ED",X"6C",
		X"63",X"D4",X"D6",X"EE",X"D6",X"D4",X"D0",X"C2",X"91",X"91",X"91",X"91",X"70",X"71",X"91",X"91",
		X"91",X"A3",X"A4",X"9C",X"B9",X"EA",X"73",X"6D",X"99",X"FB",X"FB",X"FB",X"D7",X"D5",X"D1",X"CC",
		X"C8",X"91",X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"91",X"9D",X"AD",X"B7",X"D3",X"74",X"99",
		X"63",X"DF",X"FB",X"FB",X"D8",X"EF",X"D2",X"CD",X"C9",X"91",X"91",X"91",X"70",X"71",X"91",X"91",
		X"91",X"91",X"90",X"B2",X"80",X"79",X"74",X"63",X"75",X"FB",X"FB",X"FB",X"FB",X"FB",X"9C",X"9C",
		X"CA",X"C5",X"91",X"91",X"70",X"71",X"91",X"91",X"91",X"8E",X"8F",X"AE",X"74",X"74",X"99",X"63",
		X"63",X"E0",X"DD",X"DB",X"D9",X"FB",X"9C",X"9C",X"9C",X"C6",X"BD",X"91",X"70",X"71",X"91",X"87",
		X"8B",X"8D",X"8A",X"85",X"72",X"63",X"75",X"76",X"99",X"E1",X"DE",X"DC",X"DA",X"EF",X"9C",X"CE",
		X"CB",X"C7",X"C1",X"91",X"70",X"7D",X"7F",X"86",X"83",X"8A",X"82",X"83",X"76",X"99",X"63",X"77",
		X"74",X"61",X"61",X"61",X"61",X"61",X"8A",X"8A",X"8A",X"8A",X"C3",X"BF",X"7E",X"7C",X"82",X"8A",
		X"82",X"81",X"83",X"82",X"77",X"74",X"99",X"74",X"99",X"63",X"74",X"75",X"99",X"63",X"7A",X"7B",
		X"7A",X"7B",X"7A",X"C0",X"6E",X"6F",X"82",X"81",X"83",X"8A",X"82",X"83",X"75",X"99",X"63",X"99",
		X"63",X"99",X"63",X"63",X"74",X"99",X"7A",X"7B",X"7A",X"7B",X"7B",X"85",X"6E",X"6F",X"83",X"82",
		X"83",X"82",X"83",X"8A",X"77",X"63",X"75",X"99",X"76",X"15",X"84",X"94",X"A4",X"B4",X"84",X"94",
		X"A4",X"B4",X"84",X"94",X"A4",X"B4",X"84",X"94",X"A4",X"B4",X"84",X"94",X"A4",X"B4",X"84",X"94",
		X"A4",X"B4",X"04",X"08",X"09",X"0A",X"0B",X"04",X"09",X"0A",X"08",X"0B",X"09",X"09",X"08",X"04",
		X"0A",X"0A",X"0B",X"08",X"08",X"09",X"04",X"0B",X"0B",X"04",X"09",X"0A",X"0B",X"04",X"08",X"0A",
		X"0B",X"08",X"04",X"04",X"0A",X"04",X"09",X"0B",X"0A",X"08",X"08",X"0A",X"0B",X"04",X"0A",X"0B",
		X"09",X"08",X"04",X"08",X"09",X"04",X"09",X"0B",X"04",X"08",X"04",X"08",X"0A",X"0A",X"0A",X"09",
		X"04",X"0B",X"0B",X"0A",X"08",X"09",X"04",X"08",X"0B",X"0B",X"08",X"0A",X"09",X"0A",X"0B",X"04",
		X"09",X"0A",X"08",X"0B",X"09",X"09",X"08",X"04",X"0A",X"0A",X"0B",X"08",X"08",X"09",X"04",X"0B",
		X"0B",X"04",X"0A",X"0B",X"04",X"08",X"0A",X"0B",X"08",X"04",X"04",X"0A",X"04",X"09",X"0B",X"0A",
		X"08",X"08",X"0A",X"0B",X"04",X"0A",X"0B",X"09",X"08",X"04",X"09",X"04",X"09",X"0B",X"04",X"08",
		X"04",X"08",X"0A",X"0A",X"0A",X"09",X"04",X"0B",X"0B",X"0A",X"08",X"09",X"04",X"08",X"0B",X"0B",
		X"04",X"09",X"08",X"09",X"0A",X"0B",X"04",X"09",X"0A",X"08",X"0B",X"09",X"09",X"08",X"04",X"0A",
		X"0A",X"0B",X"0A",X"08",X"09",X"04",X"08",X"0B",X"0B",X"0A",X"0B",X"04",X"08",X"0A",X"0B",X"08",
		X"04",X"04",X"0A",X"04",X"09",X"0B",X"0A",X"08",X"08",X"0A",X"0B",X"04",X"0A",X"0B",X"09",X"08",
		X"04",X"04",X"09",X"0B",X"04",X"08",X"04",X"08",X"0A",X"0B",X"0A",X"09",X"04",X"0A",X"0B",X"0A",
		X"08",X"09",X"04",X"08",X"0B",X"0B",X"04",X"09",X"08",X"04",X"09",X"0A",X"0B",X"04",X"09",X"0A",
		X"08",X"0B",X"09",X"09",X"08",X"04",X"0A",X"0A",X"0B",X"0A",X"08",X"09",X"04",X"08",X"0B",X"0B",
		X"04",X"09",X"0A",X"0B",X"08",X"04",X"04",X"0A",X"04",X"09",X"0B",X"0A",X"08",X"08",X"0A",X"0B",
		X"04",X"0A",X"0B",X"09",X"08",X"04",X"04",X"09",X"0A",X"0B",X"08",X"0B",X"09",X"0B",X"0A",X"04",
		X"09",X"04",X"09",X"0B",X"0A",X"04",X"08",X"09",X"09",X"0A",X"08",X"0B",X"0A",X"09",X"08",X"04",
		X"04",X"09",X"04",X"08",X"0A",X"0B",X"08",X"04",X"04",X"0A",X"04",X"09",X"0B",X"0A",X"08",X"08",
		X"0A",X"0B",X"04",X"0A",X"0B",X"09",X"08",X"04",X"08",X"0A",X"0A",X"0B",X"04",X"09",X"0A",X"08",
		X"0B",X"09",X"09",X"08",X"04",X"0A",X"0A",X"0B",X"0A",X"08",X"09",X"04",X"08",X"0B",X"0B",X"04",
		X"09",X"04",X"04",X"08",X"04",X"08",X"0A",X"0B",X"0A",X"09",X"0A",X"0B",X"04",X"0A",X"08",X"09",
		X"04",X"08",X"0B",X"0B",X"04",X"09",X"08",X"04",X"09",X"08",X"0A",X"0B",X"04",X"09",X"04",X"09",
		X"04",X"09",X"0B",X"0A",X"04",X"08",X"09",X"09",X"0A",X"08",X"0B",X"0A",X"09",X"08",X"04",X"04",
		X"09",X"0A",X"17",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"63",X"53",X"53",X"61",X"5D",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",
		X"F3",X"F9",X"F3",X"60",X"5E",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"99",X"F3",X"F9",X"F9",X"62",X"61",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",
		X"F9",X"F3",X"A2",X"63",X"60",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"9A",X"F9",X"F3",X"F9",X"65",X"63",X"60",X"5E",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"99",
		X"F3",X"F9",X"BA",X"65",X"65",X"63",X"61",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",X"F3",X"A2",X"BB",X"65",X"65",X"62",X"5F",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",
		X"F9",X"A2",X"BC",X"65",X"64",X"60",X"5E",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"9A",X"F3",X"BF",X"BD",X"65",X"65",X"63",X"5F",X"5E",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"99",
		X"F9",X"C0",X"BE",X"65",X"65",X"64",X"60",X"5E",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"F9",X"C1",X"23",X"65",X"65",X"65",X"63",X"60",
		X"5E",X"5D",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"99",X"98",
		X"F9",X"C2",X"18",X"65",X"65",X"65",X"65",X"63",X"60",X"5E",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"C5",X"C3",X"17",X"65",X"65",X"65",X"65",X"63",
		X"62",X"5F",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",X"98",X"98",
		X"C6",X"C4",X"22",X"65",X"65",X"65",X"65",X"64",X"60",X"5E",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"98",X"C7",X"20",X"21",X"65",X"65",X"65",X"65",X"65",
		X"63",X"61",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"9A",X"98",X"98",
		X"C8",X"13",X"01",X"65",X"65",X"65",X"65",X"65",X"64",X"60",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"98",X"98",X"C9",X"12",X"01",X"17",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"62",
		X"62",X"70",X"60",X"60",X"97",X"66",X"65",X"65",X"65",X"65",X"63",X"60",X"5E",X"5D",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",X"98",X"9D",X"A1",X"FD",X"02",X"01",X"97",X"97",X"68",X"65",
		X"65",X"65",X"65",X"63",X"60",X"5E",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"9B",X"98",X"9E",
		X"A0",X"FE",X"02",X"01",X"97",X"97",X"97",X"67",X"65",X"65",X"65",X"65",X"62",X"61",X"5C",X"5C",
		X"5C",X"5D",X"5C",X"5C",X"5C",X"99",X"98",X"9C",X"A0",X"FF",X"02",X"01",X"97",X"97",X"68",X"65",
		X"65",X"65",X"65",X"64",X"60",X"5E",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"9A",X"98",X"9C",
		X"9F",X"FF",X"02",X"01",X"97",X"97",X"67",X"65",X"65",X"65",X"65",X"62",X"5F",X"5D",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"99",X"98",X"9D",X"A1",X"FF",X"02",X"01",X"97",X"66",X"65",X"65",
		X"65",X"65",X"62",X"60",X"5E",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",X"98",X"9E",
		X"A0",X"FF",X"02",X"01",X"97",X"97",X"68",X"65",X"65",X"65",X"65",X"63",X"60",X"5E",X"5C",X"5C",
		X"5C",X"5D",X"5C",X"5C",X"5C",X"9B",X"98",X"9C",X"A0",X"FF",X"02",X"01",X"97",X"97",X"97",X"67",
		X"65",X"65",X"65",X"65",X"63",X"61",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"99",X"98",X"9D",
		X"9F",X"FF",X"02",X"01",X"97",X"97",X"66",X"65",X"65",X"65",X"65",X"62",X"5F",X"5E",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"9C",X"A1",X"FF",X"02",X"01",X"97",X"67",X"65",X"65",
		X"65",X"65",X"62",X"5F",X"5E",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",X"98",X"9E",
		X"A0",X"FF",X"02",X"01",X"68",X"65",X"65",X"65",X"65",X"62",X"5F",X"5E",X"5D",X"5C",X"5C",X"5C",
		X"5D",X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"9D",X"A0",X"FF",X"02",X"01",X"67",X"65",X"65",X"65",
		X"64",X"60",X"5E",X"5E",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"5C",X"5C",X"99",X"98",X"9D",
		X"9F",X"FF",X"02",X"01",X"66",X"65",X"65",X"65",X"65",X"63",X"60",X"5E",X"5D",X"5C",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"9B",X"98",X"9C",X"A1",X"FF",X"02",X"01",X"97",X"68",X"65",X"65",
		X"65",X"65",X"63",X"60",X"5E",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"99",X"98",X"9E",
		X"A0",X"FF",X"02",X"01",X"97",X"97",X"67",X"65",X"65",X"65",X"65",X"63",X"61",X"5C",X"5D",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"9A",X"98",X"9D",X"A0",X"FE",X"02",X"01",X"97",X"97",X"66",X"65",
		X"65",X"65",X"65",X"64",X"60",X"5C",X"5C",X"5C",X"5C",X"5D",X"5C",X"5C",X"5C",X"99",X"98",X"9C",
		X"9F",X"FC",X"02",X"01",X"17",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"43",X"43",X"43",X"43",X"43",X"43",X"97",X"67",X"65",
		X"65",X"65",X"65",X"97",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"F9",
		X"F9",X"F3",X"FC",X"02",X"01",X"66",X"65",X"65",X"65",X"65",X"62",X"97",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"F3",X"F9",X"F4",X"FA",X"05",X"01",X"65",X"65",X"65",
		X"65",X"62",X"5F",X"97",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"A2",
		X"A2",X"F5",X"FB",X"04",X"01",X"65",X"65",X"65",X"62",X"5F",X"5E",X"97",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"F3",X"F9",X"56",X"08",X"03",X"01",X"65",X"65",X"62",
		X"5F",X"5E",X"5E",X"97",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"A2",
		X"F0",X"F7",X"07",X"01",X"01",X"65",X"64",X"60",X"5E",X"5D",X"5D",X"97",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"A2",X"F1",X"F8",X"06",X"01",X"01",X"65",X"62",X"61",
		X"5D",X"5C",X"5C",X"97",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"97",X"EE",
		X"F2",X"0A",X"01",X"01",X"01",X"62",X"60",X"5F",X"5C",X"5C",X"5C",X"97",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"01",X"EF",X"0B",X"09",X"01",X"01",X"01",X"60",X"5E",X"5C",
		X"5C",X"5C",X"5C",X"97",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"01",X"01",X"0D",
		X"09",X"01",X"01",X"01",X"01",X"5F",X"5D",X"5C",X"5C",X"5C",X"9A",X"97",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5E",X"5C",X"5C",
		X"5C",X"99",X"98",X"97",X"51",X"51",X"51",X"51",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"5C",X"5C",X"5C",X"9B",X"98",X"98",X"97",X"51",X"51",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5C",X"5C",X"9A",
		X"98",X"98",X"98",X"97",X"51",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"5C",X"99",X"98",X"98",X"98",X"98",X"97",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"9A",X"98",X"98",
		X"98",X"98",X"98",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"98",X"98",X"98",X"98",X"98",X"98",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"4F",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"52",
		X"52",X"56",X"56",X"56",X"56",X"56",X"B6",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"B6",X"9F",X"9C",X"99",X"5C",X"61",X"62",X"65",X"B6",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"B6",X"A0",
		X"9D",X"99",X"5C",X"61",X"63",X"65",X"B6",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"B6",X"A0",X"9E",X"9B",X"5C",X"5F",X"64",X"65",X"B6",X"4F",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"B6",X"A1",
		X"9C",X"9A",X"5C",X"5E",X"60",X"62",X"B6",X"4F",X"4F",X"4F",X"55",X"56",X"00",X"00",X"00",X"00",
		X"00",X"56",X"55",X"4F",X"4F",X"4F",X"B6",X"9F",X"9C",X"9B",X"5C",X"5D",X"61",X"63",X"B6",X"4F",
		X"53",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"53",X"4F",X"B6",X"A0",
		X"9E",X"99",X"5C",X"5C",X"60",X"64",X"B6",X"52",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"52",X"B6",X"A0",X"9D",X"9A",X"5C",X"5C",X"5F",X"62",X"B6",X"50",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"50",X"B6",X"A1",
		X"9C",X"99",X"5E",X"5E",X"5E",X"61",X"FD",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"9F",X"9E",X"9B",X"5C",X"5C",X"5E",X"5F",X"FE",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A0",
		X"9D",X"98",X"99",X"5C",X"5D",X"5E",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A0",X"9D",X"98",X"9B",X"5C",X"5C",X"5E",X"FF",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A1",
		X"9E",X"9A",X"9A",X"9A",X"5C",X"5D",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"9F",X"9D",X"98",X"98",X"9A",X"5C",X"5C",X"FF",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A0",
		X"9C",X"98",X"98",X"9B",X"5C",X"5C",X"FE",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A0",X"9E",X"98",X"98",X"98",X"9A",X"5C",X"FC",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"A1",
		X"9C",X"98",X"98",X"98",X"99",X"5C",X"08",X"63",X"73",X"73",X"73",X"73",X"73",X"73",X"43",X"43",
		X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"FC",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"F3",X"F3",X"F9",X"A2",X"F9",X"FC",X"02",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"4C",
		X"A2",X"F3",X"F9",X"F9",X"F4",X"FA",X"05",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"01",
		X"01",X"01",X"01",X"01",X"01",X"09",X"3A",X"39",X"F9",X"F3",X"A2",X"F3",X"F5",X"FB",X"04",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"01",X"01",X"01",X"01",X"01",X"09",X"3F",X"39",X"F3",
		X"A2",X"F9",X"F3",X"F9",X"F6",X"08",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"01",
		X"01",X"01",X"01",X"09",X"3F",X"39",X"F3",X"F9",X"F3",X"F9",X"A2",X"F0",X"F7",X"07",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"01",X"01",X"01",X"09",X"3F",X"39",X"A2",X"F3",X"A2",
		X"F3",X"A2",X"F9",X"F1",X"F8",X"06",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"4E",
		X"4E",X"4E",X"4D",X"39",X"F9",X"F3",X"F9",X"A2",X"F9",X"F3",X"EE",X"F2",X"0A",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A2",X"F9",X"A2",X"F9",X"A2",X"F3",X"F9",X"A2",X"A2",
		X"F9",X"EC",X"EF",X"0B",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",
		X"F9",X"F3",X"F9",X"A2",X"F3",X"A2",X"F3",X"A2",X"E9",X"ED",X"0B",X"09",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"A2",X"F3",X"F9",X"F3",X"A2",X"A2",X"F9",X"E5",
		X"EA",X"0D",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",
		X"F9",X"A2",X"F9",X"F3",X"F3",X"F9",X"A2",X"E6",X"EB",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F3",X"A2",X"F3",X"A2",X"F3",X"F9",X"A2",X"E1",X"E7",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",
		X"F9",X"F9",X"F3",X"F9",X"A2",X"F9",X"E2",X"E8",X"0E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"A2",X"F9",X"A2",X"F3",X"F3",X"F9",X"F3",X"E3",X"11",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FF",X"F9",
		X"F3",X"A2",X"F9",X"F3",X"A2",X"A2",X"E4",X"10",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"FE",X"A2",X"F9",X"F3",X"A2",X"F3",X"F9",X"F3",X"FD",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FD",X"18",
		X"F8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",
		X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"E8",X"FB",X"2E",X"83",X"83",X"86",X"84",X"83",X"83",
		X"2F",X"83",X"83",X"86",X"84",X"83",X"83",X"2F",X"83",X"83",X"86",X"84",X"83",X"83",X"2E",X"FB",
		X"FF",X"2E",X"1A",X"1A",X"82",X"80",X"1A",X"1A",X"2F",X"1A",X"1A",X"82",X"80",X"1A",X"1A",X"2F",
		X"1A",X"1A",X"82",X"80",X"1A",X"1A",X"2E",X"FF",X"FC",X"2E",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"2F",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"2F",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"2E",X"FC",
		X"FD",X"1B",X"67",X"79",X"79",X"79",X"79",X"65",X"1B",X"67",X"79",X"79",X"79",X"79",X"65",X"1B",
		X"67",X"79",X"79",X"79",X"79",X"65",X"1B",X"FD",X"FC",X"1B",X"66",X"78",X"78",X"78",X"78",X"64",
		X"1B",X"66",X"78",X"78",X"78",X"78",X"64",X"1B",X"66",X"78",X"78",X"78",X"78",X"64",X"1B",X"FC",
		X"FD",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"FD",X"FE",X"1B",X"6F",X"6F",X"81",X"6F",X"6F",X"81",
		X"6F",X"6F",X"81",X"6F",X"6F",X"81",X"6F",X"6F",X"81",X"6F",X"6F",X"81",X"6F",X"6F",X"1B",X"FE",
		X"00",X"1B",X"00",X"69",X"73",X"7F",X"7D",X"7B",X"33",X"77",X"75",X"71",X"27",X"77",X"75",X"31",
		X"7F",X"7D",X"6D",X"6B",X"69",X"00",X"1B",X"00",X"00",X"1B",X"00",X"68",X"72",X"7E",X"7C",X"7A",
		X"32",X"76",X"74",X"70",X"26",X"76",X"74",X"30",X"7E",X"7C",X"6C",X"6A",X"68",X"00",X"1B",X"00",
		X"00",X"1B",X"6E",X"6E",X"81",X"6E",X"6E",X"81",X"6E",X"6E",X"81",X"6E",X"6E",X"81",X"6E",X"6E",
		X"81",X"6E",X"6E",X"81",X"6E",X"6E",X"1B",X"00",X"00",X"16",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"14",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"2B",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"29",
		X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"1B",
		X"2A",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"28",X"1B",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"16",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"14",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9A",X"40",X"42",X"B9",X"CF",X"40",X"42",X"BE",X"BF",X"40",X"42",
		X"C3",X"AF",X"40",X"42",X"CF",X"9F",X"40",X"42",X"DB",X"8F",X"40",X"42",X"E7",X"7F",X"50",X"42",
		X"BA",X"CF",X"50",X"42",X"BF",X"BF",X"50",X"42",X"C4",X"AF",X"50",X"42",X"D0",X"9F",X"50",X"42",
		X"DC",X"8F",X"50",X"42",X"E8",X"7F",X"60",X"42",X"BB",X"CF",X"60",X"42",X"C0",X"BF",X"60",X"42",
		X"C5",X"AF",X"60",X"42",X"D1",X"9F",X"60",X"42",X"DD",X"8F",X"60",X"42",X"E9",X"7F",X"70",X"42",
		X"C6",X"AF",X"70",X"42",X"D2",X"9F",X"70",X"42",X"DE",X"8F",X"70",X"42",X"EA",X"7F",X"80",X"42",
		X"C7",X"AF",X"80",X"42",X"D3",X"9F",X"80",X"42",X"DF",X"8F",X"80",X"42",X"EB",X"7F",X"90",X"42",
		X"C8",X"AF",X"90",X"42",X"D4",X"9F",X"90",X"42",X"E0",X"8F",X"90",X"42",X"EC",X"7F",X"A0",X"42",
		X"C9",X"AF",X"A0",X"42",X"D5",X"9F",X"A0",X"42",X"E1",X"8F",X"A0",X"42",X"ED",X"7F",X"B0",X"42",
		X"CA",X"AF",X"B0",X"42",X"D6",X"9F",X"B0",X"42",X"E2",X"8F",X"B0",X"42",X"EE",X"7F",X"C0",X"42",
		X"CB",X"AF",X"C0",X"42",X"D7",X"9F",X"C0",X"42",X"E3",X"8F",X"C0",X"42",X"EF",X"7F",X"D0",X"42",
		X"CC",X"AF",X"D0",X"42",X"D8",X"9F",X"D0",X"42",X"E4",X"8F",X"D0",X"42",X"F0",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
