library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3A",X"00",X"40",X"FE",X"55",X"CA",X"01",X"40",X"3A",X"00",X"88",X"31",X"00",X"88",X"C3",X"B1",
		X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"3A",X"FE",X"83",X"B7",X"C8",X"E5",X"21",
		X"00",X"83",X"34",X"7E",X"6F",X"71",X"E1",X"C9",X"1A",X"77",X"7D",X"D6",X"20",X"6F",X"30",X"01",
		X"25",X"13",X"10",X"F4",X"C9",X"FF",X"FF",X"FF",X"11",X"10",X"20",X"21",X"00",X"A8",X"06",X"20",
		X"73",X"23",X"10",X"FC",X"0E",X"15",X"10",X"FE",X"0D",X"20",X"FB",X"15",X"20",X"F0",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"E5",X"D5",X"C5",X"DD",X"E5",X"FD",X"E5",X"3A",X"00",
		X"88",X"AF",X"32",X"08",X"B8",X"CD",X"00",X"3E",X"21",X"07",X"80",X"11",X"07",X"B0",X"7E",X"12",
		X"2C",X"1C",X"06",X"1C",X"7E",X"0F",X"0F",X"0F",X"0F",X"12",X"2C",X"1C",X"7E",X"12",X"2C",X"1C",
		X"10",X"F2",X"0E",X"08",X"3A",X"2F",X"84",X"B7",X"28",X"05",X"0E",X"06",X"1E",X"48",X"6B",X"7E",
		X"0F",X"0F",X"0F",X"0F",X"12",X"2C",X"1C",X"06",X"03",X"7E",X"12",X"2C",X"1C",X"10",X"FA",X"0D",
		X"20",X"ED",X"21",X"7F",X"83",X"7E",X"B7",X"28",X"07",X"35",X"20",X"04",X"AF",X"32",X"1C",X"B8",
		X"21",X"7E",X"83",X"7E",X"B7",X"28",X"07",X"35",X"20",X"04",X"AF",X"32",X"18",X"B8",X"3A",X"04",
		X"E0",X"E6",X"08",X"CA",X"FC",X"00",X"3A",X"FE",X"83",X"A7",X"CA",X"FC",X"00",X"3A",X"FD",X"83",
		X"A7",X"28",X"19",X"3D",X"28",X"16",X"0E",X"02",X"21",X"43",X"80",X"11",X"43",X"B0",X"7E",X"81",
		X"12",X"0E",X"02",X"21",X"47",X"80",X"11",X"47",X"B0",X"7E",X"81",X"12",X"3A",X"FE",X"83",X"B7",
		X"CA",X"22",X"01",X"CD",X"BF",X"07",X"3A",X"EA",X"83",X"B7",X"CA",X"53",X"02",X"2A",X"D2",X"83",
		X"7C",X"B5",X"CA",X"7F",X"01",X"2B",X"22",X"D2",X"83",X"CD",X"40",X"25",X"CD",X"8B",X"28",X"C3",
		X"53",X"02",X"3A",X"86",X"83",X"A7",X"CA",X"30",X"01",X"3D",X"32",X"86",X"83",X"C3",X"53",X"02",
		X"3A",X"D6",X"83",X"FE",X"02",X"D2",X"66",X"01",X"B7",X"CC",X"D4",X"0D",X"CD",X"CA",X"33",X"AF",
		X"32",X"CD",X"83",X"32",X"CF",X"83",X"32",X"B5",X"83",X"67",X"6F",X"22",X"93",X"82",X"21",X"5C",
		X"82",X"11",X"5D",X"82",X"01",X"0B",X"00",X"70",X"ED",X"B0",X"21",X"AF",X"83",X"36",X"80",X"2C",
		X"77",X"2C",X"77",X"C3",X"53",X"02",X"21",X"D8",X"83",X"7E",X"B7",X"CA",X"53",X"02",X"35",X"C2",
		X"53",X"02",X"2D",X"7E",X"B7",X"C2",X"53",X"02",X"21",X"D6",X"83",X"35",X"C3",X"53",X"02",X"2A",
		X"82",X"83",X"7C",X"B5",X"28",X"12",X"2B",X"22",X"82",X"83",X"7C",X"B5",X"20",X"0A",X"3E",X"0F",
		X"DF",X"3E",X"B0",X"DF",X"AF",X"32",X"71",X"83",X"3A",X"FD",X"83",X"3D",X"C2",X"82",X"02",X"3A",
		X"5C",X"82",X"FE",X"05",X"CA",X"6C",X"02",X"3A",X"98",X"82",X"A7",X"28",X"07",X"3D",X"32",X"98",
		X"82",X"C3",X"F0",X"01",X"3A",X"97",X"82",X"A7",X"C2",X"65",X"02",X"2A",X"9D",X"82",X"7C",X"B5",
		X"20",X"2E",X"CD",X"93",X"08",X"CD",X"DE",X"2A",X"3A",X"B5",X"83",X"B7",X"20",X"22",X"3C",X"32",
		X"B5",X"83",X"3E",X"FF",X"32",X"84",X"83",X"3A",X"80",X"83",X"B7",X"28",X"13",X"AF",X"32",X"80",
		X"83",X"21",X"40",X"00",X"22",X"82",X"83",X"11",X"11",X"10",X"21",X"51",X"AA",X"06",X"07",X"EF",
		X"3A",X"84",X"83",X"B7",X"28",X"0A",X"3D",X"32",X"84",X"83",X"21",X"50",X"A8",X"CC",X"6B",X"2A",
		X"CD",X"8E",X"30",X"CD",X"8B",X"28",X"3A",X"07",X"81",X"A7",X"28",X"07",X"3A",X"09",X"81",X"3D",
		X"32",X"09",X"81",X"3A",X"08",X"81",X"A7",X"28",X"07",X"3A",X"24",X"81",X"3D",X"32",X"24",X"81",
		X"CD",X"48",X"22",X"3A",X"07",X"81",X"A7",X"28",X"07",X"3A",X"09",X"81",X"3C",X"32",X"09",X"81",
		X"3A",X"08",X"81",X"A7",X"28",X"07",X"3A",X"24",X"81",X"3C",X"32",X"24",X"81",X"CD",X"81",X"27",
		X"CD",X"40",X"25",X"CD",X"00",X"1C",X"CD",X"50",X"30",X"CD",X"A0",X"02",X"3A",X"97",X"82",X"A7",
		X"C4",X"B5",X"06",X"3A",X"00",X"88",X"FD",X"E1",X"DD",X"E1",X"C1",X"D1",X"E1",X"3E",X"01",X"32",
		X"08",X"B8",X"F1",X"ED",X"45",X"3D",X"32",X"97",X"82",X"C3",X"F0",X"01",X"21",X"5E",X"82",X"11",
		X"5F",X"82",X"01",X"04",X"00",X"70",X"ED",X"B0",X"AF",X"32",X"5C",X"82",X"CD",X"E6",X"05",X"C3",
		X"53",X"02",X"3A",X"5D",X"82",X"FE",X"05",X"C2",X"A7",X"01",X"21",X"63",X"82",X"11",X"64",X"82",
		X"01",X"04",X"00",X"70",X"ED",X"B0",X"AF",X"32",X"5D",X"82",X"CD",X"E6",X"05",X"C3",X"53",X"02",
		X"2A",X"9D",X"82",X"7C",X"B5",X"C8",X"2B",X"22",X"9D",X"82",X"7C",X"B5",X"C0",X"32",X"AE",X"83",
		X"C9",X"AF",X"32",X"08",X"B8",X"32",X"05",X"88",X"32",X"10",X"B8",X"32",X"0C",X"B8",X"21",X"00",
		X"80",X"11",X"01",X"80",X"01",X"FF",X"07",X"75",X"ED",X"B0",X"21",X"00",X"B0",X"01",X"00",X"00",
		X"71",X"2C",X"10",X"FC",X"3A",X"02",X"E0",X"11",X"D6",X"0E",X"E6",X"03",X"83",X"5F",X"30",X"01",
		X"14",X"1A",X"32",X"E4",X"83",X"3A",X"04",X"E0",X"67",X"CB",X"5C",X"28",X"05",X"3E",X"01",X"32",
		X"C2",X"83",X"7C",X"E6",X"06",X"32",X"D4",X"83",X"21",X"E0",X"0E",X"11",X"EB",X"83",X"01",X"12",
		X"00",X"ED",X"B0",X"CD",X"BC",X"20",X"3E",X"01",X"32",X"70",X"83",X"32",X"08",X"B8",X"FF",X"AF",
		X"32",X"01",X"B0",X"3E",X"06",X"32",X"03",X"B0",X"21",X"00",X"01",X"22",X"C7",X"83",X"3E",X"15",
		X"32",X"81",X"83",X"21",X"87",X"0F",X"11",X"00",X"84",X"01",X"20",X"00",X"ED",X"B0",X"21",X"06",
		X"E0",X"36",X"9B",X"21",X"06",X"D0",X"36",X"88",X"3E",X"18",X"32",X"D9",X"83",X"32",X"02",X"D0",
		X"AF",X"CD",X"A7",X"07",X"3A",X"D9",X"83",X"E6",X"EF",X"32",X"D9",X"83",X"32",X"02",X"D0",X"3E",
		X"FF",X"CD",X"A7",X"07",X"3A",X"D6",X"83",X"FE",X"02",X"D4",X"74",X"0C",X"CD",X"42",X"0B",X"3A",
		X"D6",X"83",X"3D",X"C4",X"8A",X"0B",X"CD",X"98",X"33",X"3E",X"02",X"21",X"54",X"82",X"77",X"23",
		X"77",X"3E",X"09",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"2A",X"C7",X"83",X"7C",X"B5",
		X"2B",X"20",X"FB",X"3A",X"FE",X"83",X"B7",X"C2",X"1E",X"04",X"3A",X"B3",X"83",X"B7",X"20",X"C4",
		X"3A",X"02",X"E0",X"07",X"30",X"07",X"07",X"38",X"BB",X"0E",X"02",X"18",X"02",X"0E",X"01",X"3A",
		X"E1",X"83",X"B9",X"38",X"AF",X"91",X"27",X"32",X"E1",X"83",X"79",X"32",X"70",X"83",X"21",X"00",
		X"85",X"11",X"01",X"85",X"01",X"FF",X"01",X"75",X"ED",X"B0",X"32",X"FE",X"83",X"3E",X"01",X"32",
		X"FD",X"83",X"32",X"B3",X"83",X"67",X"6F",X"32",X"B7",X"83",X"22",X"B8",X"83",X"CD",X"2D",X"0B",
		X"3E",X"03",X"32",X"3D",X"80",X"CD",X"EC",X"07",X"AF",X"32",X"71",X"80",X"DF",X"3E",X"09",X"DF",
		X"3E",X"0A",X"DF",X"3E",X"0B",X"DF",X"21",X"20",X"00",X"22",X"9D",X"82",X"21",X"A0",X"01",X"22",
		X"82",X"83",X"21",X"00",X"00",X"22",X"D2",X"83",X"CD",X"F9",X"07",X"FF",X"CD",X"C6",X"32",X"AF",
		X"67",X"6F",X"32",X"2F",X"84",X"32",X"2D",X"84",X"22",X"93",X"82",X"21",X"40",X"84",X"11",X"41",
		X"84",X"01",X"4F",X"00",X"70",X"ED",X"B0",X"32",X"04",X"80",X"3C",X"32",X"5A",X"82",X"3A",X"EA",
		X"83",X"B7",X"C2",X"6A",X"04",X"3A",X"CD",X"83",X"B7",X"20",X"0D",X"3A",X"FE",X"83",X"3D",X"28",
		X"04",X"FF",X"CD",X"01",X"07",X"CD",X"42",X"0B",X"3A",X"6D",X"82",X"A7",X"C4",X"03",X"06",X"CD",
		X"65",X"09",X"32",X"EA",X"83",X"CD",X"39",X"0A",X"21",X"9E",X"83",X"36",X"20",X"2D",X"36",X"10",
		X"2D",X"36",X"20",X"3A",X"FE",X"83",X"3D",X"C4",X"D4",X"07",X"AF",X"32",X"6D",X"82",X"3A",X"CD",
		X"83",X"32",X"B6",X"83",X"CD",X"6B",X"0A",X"C3",X"7B",X"03",X"CD",X"42",X"0B",X"3A",X"CE",X"83",
		X"B7",X"CA",X"7B",X"03",X"CD",X"17",X"08",X"CD",X"F9",X"07",X"AF",X"21",X"9A",X"83",X"77",X"2C",
		X"77",X"32",X"CC",X"83",X"32",X"EA",X"83",X"21",X"A0",X"83",X"11",X"A1",X"83",X"01",X"0D",X"00",
		X"77",X"ED",X"B0",X"3E",X"80",X"DF",X"3A",X"CF",X"83",X"B7",X"20",X"06",X"CD",X"45",X"08",X"C3",
		X"7B",X"03",X"CD",X"35",X"08",X"3E",X"0C",X"DF",X"3E",X"0D",X"DF",X"2A",X"C5",X"83",X"2B",X"22",
		X"C5",X"83",X"7C",X"B5",X"20",X"F8",X"3A",X"FE",X"83",X"3D",X"CA",X"5A",X"05",X"3A",X"FD",X"83",
		X"3D",X"C2",X"06",X"05",X"21",X"C9",X"83",X"36",X"01",X"23",X"7E",X"B7",X"C2",X"47",X"05",X"FF",
		X"CD",X"45",X"08",X"3E",X"01",X"32",X"FE",X"83",X"32",X"5C",X"82",X"21",X"5E",X"82",X"11",X"5F",
		X"82",X"01",X"04",X"00",X"36",X"00",X"ED",X"B0",X"21",X"00",X"86",X"11",X"FF",X"80",X"01",X"B7",
		X"00",X"ED",X"B0",X"21",X"C0",X"85",X"11",X"0C",X"80",X"01",X"2B",X"00",X"ED",X"B0",X"3E",X"01",
		X"32",X"3F",X"80",X"C3",X"7B",X"03",X"21",X"CA",X"83",X"36",X"01",X"2B",X"7E",X"B7",X"C2",X"6A",
		X"05",X"FF",X"CD",X"45",X"08",X"3E",X"01",X"32",X"FE",X"83",X"32",X"5D",X"82",X"21",X"63",X"82",
		X"11",X"64",X"82",X"01",X"04",X"00",X"70",X"ED",X"B0",X"21",X"C0",X"86",X"11",X"0C",X"80",X"01",
		X"2B",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"3F",X"80",X"21",X"00",X"85",X"11",X"FF",X"80",X"01",
		X"B7",X"00",X"ED",X"B0",X"C3",X"7B",X"03",X"AF",X"32",X"5C",X"82",X"21",X"5E",X"82",X"11",X"5F",
		X"82",X"01",X"04",X"00",X"70",X"ED",X"B0",X"C3",X"7A",X"05",X"AF",X"32",X"5C",X"82",X"21",X"5E",
		X"82",X"11",X"5F",X"82",X"01",X"04",X"00",X"70",X"ED",X"B0",X"AF",X"32",X"5D",X"82",X"21",X"63",
		X"82",X"11",X"64",X"82",X"01",X"04",X"00",X"70",X"ED",X"B0",X"FF",X"CD",X"F9",X"07",X"CD",X"8A",
		X"0B",X"CD",X"B3",X"0E",X"CD",X"42",X"0B",X"21",X"00",X"81",X"11",X"01",X"81",X"01",X"5F",X"01",
		X"75",X"ED",X"B0",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"04",X"00",X"70",X"ED",X"B0",X"21",
		X"0C",X"80",X"11",X"0D",X"80",X"01",X"2E",X"00",X"70",X"ED",X"B0",X"AF",X"32",X"C3",X"83",X"32",
		X"FE",X"83",X"32",X"BF",X"83",X"21",X"C9",X"83",X"77",X"2C",X"77",X"67",X"6F",X"32",X"10",X"B8",
		X"32",X"0C",X"B8",X"22",X"93",X"82",X"32",X"BB",X"83",X"32",X"CB",X"83",X"32",X"D8",X"83",X"32",
		X"C4",X"83",X"32",X"BA",X"83",X"32",X"95",X"82",X"32",X"5B",X"82",X"3E",X"03",X"32",X"D6",X"83",
		X"CD",X"FE",X"07",X"C3",X"7B",X"03",X"3E",X"01",X"32",X"6D",X"82",X"32",X"5A",X"82",X"32",X"CD",
		X"83",X"AF",X"32",X"5B",X"82",X"32",X"EA",X"83",X"3E",X"FF",X"32",X"97",X"82",X"3E",X"40",X"32",
		X"98",X"82",X"C9",X"3E",X"10",X"DF",X"3E",X"30",X"DF",X"3A",X"FD",X"83",X"3D",X"20",X"0C",X"21",
		X"93",X"82",X"34",X"7E",X"D6",X"05",X"20",X"0D",X"77",X"18",X"0A",X"21",X"94",X"82",X"34",X"7E",
		X"D6",X"05",X"20",X"01",X"77",X"CD",X"3C",X"06",X"CD",X"5E",X"06",X"CD",X"C6",X"32",X"CD",X"8B",
		X"2A",X"3E",X"01",X"32",X"80",X"83",X"11",X"00",X"01",X"C3",X"03",X"09",X"CD",X"F9",X"07",X"21",
		X"9A",X"83",X"AF",X"77",X"2C",X"77",X"3C",X"32",X"CC",X"83",X"3E",X"20",X"21",X"06",X"A8",X"CD",
		X"8C",X"07",X"2C",X"2C",X"CD",X"8C",X"07",X"0E",X"0A",X"09",X"3D",X"20",X"F2",X"C9",X"21",X"0C",
		X"80",X"11",X"0D",X"80",X"01",X"2B",X"00",X"70",X"ED",X"B0",X"21",X"0C",X"80",X"11",X"0C",X"B0",
		X"01",X"2B",X"00",X"ED",X"B0",X"21",X"00",X"81",X"11",X"01",X"81",X"01",X"62",X"00",X"36",X"00",
		X"ED",X"B0",X"C9",X"21",X"64",X"AB",X"CD",X"A8",X"06",X"21",X"A4",X"AA",X"CD",X"A8",X"06",X"21",
		X"E4",X"A9",X"CD",X"A8",X"06",X"21",X"24",X"A9",X"CD",X"A8",X"06",X"21",X"64",X"A8",X"CD",X"A8",
		X"06",X"AF",X"32",X"2F",X"84",X"C3",X"82",X"0A",X"3E",X"10",X"77",X"23",X"77",X"01",X"1F",X"00",
		X"09",X"77",X"23",X"77",X"C9",X"FE",X"C0",X"CA",X"D4",X"06",X"FE",X"90",X"CA",X"DA",X"06",X"FE",
		X"70",X"CA",X"E0",X"06",X"FE",X"50",X"CA",X"E6",X"06",X"FE",X"30",X"CA",X"EC",X"06",X"FE",X"10",
		X"CA",X"83",X"06",X"C9",X"21",X"64",X"AB",X"C3",X"F2",X"06",X"21",X"A4",X"AA",X"C3",X"F2",X"06",
		X"21",X"E4",X"A9",X"C3",X"F2",X"06",X"21",X"24",X"A9",X"C3",X"F2",X"06",X"21",X"64",X"A8",X"C3",
		X"F2",X"06",X"36",X"FC",X"23",X"36",X"FD",X"01",X"1F",X"00",X"09",X"36",X"FE",X"23",X"36",X"FF",
		X"C9",X"3A",X"FD",X"83",X"3D",X"20",X"32",X"21",X"0C",X"80",X"11",X"C0",X"85",X"01",X"2B",X"00",
		X"ED",X"B0",X"21",X"FF",X"80",X"11",X"00",X"86",X"01",X"B7",X"00",X"ED",X"B0",X"21",X"C0",X"86",
		X"11",X"0C",X"80",X"01",X"2B",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"3F",X"80",X"21",X"00",X"85",
		X"11",X"FF",X"80",X"01",X"B7",X"00",X"ED",X"B0",X"C9",X"21",X"FF",X"80",X"11",X"00",X"85",X"01",
		X"B7",X"00",X"ED",X"B0",X"21",X"0C",X"80",X"11",X"C0",X"86",X"01",X"2B",X"00",X"ED",X"B0",X"21",
		X"00",X"86",X"11",X"FF",X"80",X"01",X"B7",X"00",X"ED",X"B0",X"21",X"C0",X"85",X"11",X"0C",X"80",
		X"01",X"2B",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"3F",X"80",X"3A",X"95",X"82",X"A7",X"C0",X"AF",
		X"32",X"5B",X"82",X"3E",X"01",X"32",X"95",X"82",X"C9",X"21",X"02",X"A8",X"11",X"10",X"20",X"0E",
		X"04",X"06",X"1C",X"73",X"23",X"10",X"FC",X"09",X"15",X"20",X"F6",X"C9",X"01",X"10",X"0A",X"71",
		X"23",X"10",X"FC",X"C9",X"21",X"08",X"A8",X"11",X"10",X"20",X"0E",X"0A",X"06",X"16",X"73",X"23",
		X"10",X"FC",X"09",X"15",X"20",X"F6",X"C9",X"32",X"00",X"D0",X"3A",X"D9",X"83",X"E6",X"F7",X"32",
		X"02",X"D0",X"00",X"00",X"00",X"00",X"3A",X"D9",X"83",X"F6",X"08",X"32",X"02",X"D0",X"C9",X"21",
		X"00",X"83",X"7E",X"B7",X"C8",X"35",X"4F",X"2C",X"7E",X"CD",X"A7",X"07",X"54",X"5D",X"2C",X"06",
		X"00",X"ED",X"B0",X"C9",X"3A",X"FD",X"83",X"3D",X"CA",X"E1",X"07",X"3E",X"01",X"32",X"5B",X"82",
		X"C9",X"3A",X"6D",X"82",X"A7",X"C8",X"3E",X"01",X"32",X"5B",X"82",X"C9",X"21",X"00",X"83",X"11",
		X"01",X"83",X"01",X"2F",X"00",X"70",X"ED",X"B0",X"C9",X"3A",X"FE",X"83",X"3D",X"C8",X"AF",X"21",
		X"44",X"80",X"11",X"45",X"80",X"01",X"1F",X"00",X"70",X"ED",X"B0",X"21",X"20",X"84",X"11",X"21",
		X"84",X"0E",X"0B",X"77",X"ED",X"B0",X"C9",X"21",X"44",X"80",X"AF",X"36",X"01",X"2C",X"77",X"2C",
		X"2C",X"77",X"3A",X"FE",X"83",X"FE",X"02",X"C0",X"21",X"40",X"00",X"22",X"D2",X"83",X"21",X"40",
		X"00",X"22",X"DA",X"83",X"C9",X"21",X"50",X"A8",X"CD",X"6B",X"2A",X"21",X"70",X"AA",X"11",X"D6",
		X"0F",X"06",X"09",X"EF",X"C9",X"AF",X"32",X"71",X"83",X"3A",X"FE",X"83",X"3D",X"C8",X"3A",X"FD",
		X"83",X"EE",X"03",X"32",X"FD",X"83",X"21",X"B8",X"83",X"3D",X"28",X"01",X"2C",X"7E",X"32",X"B7",
		X"83",X"AF",X"32",X"B6",X"83",X"3C",X"32",X"5A",X"82",X"3A",X"C2",X"83",X"B7",X"C8",X"3A",X"CB",
		X"83",X"EE",X"01",X"32",X"CB",X"83",X"67",X"32",X"10",X"B8",X"32",X"0C",X"B8",X"C9",X"21",X"51",
		X"AA",X"11",X"04",X"10",X"06",X"04",X"EF",X"11",X"DA",X"0F",X"06",X"05",X"EF",X"3E",X"01",X"32",
		X"04",X"80",X"C9",X"3A",X"CD",X"83",X"B7",X"C0",X"3A",X"04",X"80",X"B7",X"C0",X"3A",X"AE",X"83",
		X"B7",X"20",X"07",X"3C",X"32",X"AE",X"83",X"3E",X"06",X"DF",X"CD",X"DD",X"0A",X"3A",X"DF",X"83",
		X"B7",X"20",X"35",X"21",X"DC",X"83",X"35",X"C0",X"36",X"20",X"23",X"7E",X"B7",X"CA",X"7E",X"08",
		X"3D",X"77",X"2C",X"7E",X"3D",X"27",X"77",X"2D",X"FE",X"10",X"20",X"07",X"3E",X"05",X"DF",X"AF",
		X"32",X"3F",X"80",X"66",X"7C",X"E6",X"03",X"4F",X"AC",X"07",X"07",X"6F",X"26",X"00",X"29",X"11",
		X"DF",X"A8",X"19",X"3E",X"10",X"91",X"77",X"C9",X"3A",X"E0",X"83",X"B7",X"C0",X"3C",X"32",X"E0",
		X"83",X"21",X"51",X"AA",X"11",X"04",X"10",X"06",X"05",X"EF",X"3A",X"DE",X"83",X"5F",X"16",X"00",
		X"CD",X"C3",X"0B",X"3A",X"FE",X"83",X"B7",X"C8",X"3A",X"FD",X"83",X"3D",X"28",X"05",X"21",X"EB",
		X"83",X"18",X"03",X"21",X"ED",X"83",X"7B",X"86",X"27",X"77",X"5F",X"23",X"7A",X"8E",X"27",X"77",
		X"57",X"3A",X"FD",X"83",X"3D",X"20",X"09",X"01",X"E7",X"83",X"0A",X"B7",X"20",X"2B",X"18",X"07",
		X"01",X"E8",X"83",X"0A",X"B7",X"20",X"22",X"2A",X"DE",X"0E",X"ED",X"52",X"28",X"02",X"30",X"19",
		X"32",X"CF",X"83",X"3C",X"02",X"0D",X"0D",X"0A",X"3C",X"02",X"21",X"DE",X"AB",X"01",X"E0",X"FF",
		X"09",X"3D",X"20",X"FC",X"36",X"4D",X"3E",X"07",X"DF",X"2A",X"EF",X"83",X"B7",X"ED",X"52",X"D0",
		X"ED",X"53",X"EF",X"83",X"C9",X"AF",X"32",X"CE",X"83",X"3A",X"CD",X"83",X"B7",X"20",X"04",X"AF",
		X"32",X"CF",X"83",X"3A",X"FE",X"83",X"B7",X"28",X"74",X"3A",X"FD",X"83",X"3D",X"20",X"05",X"21",
		X"E5",X"83",X"18",X"03",X"21",X"E6",X"83",X"3A",X"CD",X"83",X"B7",X"20",X"08",X"35",X"20",X"05",
		X"3E",X"01",X"32",X"CF",X"83",X"CD",X"DB",X"29",X"3A",X"CD",X"83",X"B7",X"20",X"0A",X"3C",X"32",
		X"B5",X"83",X"21",X"50",X"A8",X"CD",X"6B",X"2A",X"3A",X"6C",X"82",X"EE",X"01",X"32",X"B5",X"83",
		X"3A",X"FD",X"83",X"3D",X"C2",X"F5",X"09",X"21",X"5E",X"82",X"CD",X"FE",X"09",X"3A",X"5A",X"82",
		X"A7",X"28",X"0A",X"CD",X"C6",X"32",X"CD",X"23",X"20",X"AF",X"32",X"5A",X"82",X"21",X"44",X"80",
		X"36",X"80",X"2C",X"36",X"1E",X"2C",X"36",X"03",X"2C",X"36",X"E0",X"AF",X"32",X"CD",X"83",X"32",
		X"2D",X"84",X"32",X"2C",X"84",X"32",X"69",X"82",X"3C",X"32",X"C3",X"83",X"C9",X"3A",X"CD",X"83",
		X"B7",X"C8",X"C3",X"CD",X"09",X"21",X"63",X"82",X"CD",X"FE",X"09",X"C3",X"BD",X"09",X"AF",X"B6",
		X"11",X"64",X"AB",X"C4",X"28",X"0A",X"23",X"AF",X"B6",X"11",X"A4",X"AA",X"C4",X"28",X"0A",X"23",
		X"AF",X"B6",X"11",X"E4",X"A9",X"C4",X"28",X"0A",X"23",X"AF",X"B6",X"11",X"24",X"A9",X"C4",X"28",
		X"0A",X"23",X"AF",X"B6",X"11",X"64",X"A8",X"C8",X"EB",X"36",X"6C",X"23",X"36",X"6D",X"01",X"1F",
		X"00",X"09",X"36",X"6E",X"23",X"36",X"6F",X"EB",X"C9",X"3A",X"E4",X"83",X"3C",X"C8",X"3A",X"FE",
		X"83",X"B7",X"20",X"05",X"21",X"E4",X"83",X"18",X"0E",X"3A",X"FD",X"83",X"3D",X"20",X"05",X"21",
		X"E5",X"83",X"18",X"03",X"21",X"E6",X"83",X"46",X"78",X"B7",X"3E",X"4D",X"11",X"E0",X"FF",X"21",
		X"BE",X"AB",X"28",X"04",X"77",X"19",X"10",X"FC",X"36",X"10",X"C9",X"3A",X"B7",X"83",X"21",X"7E",
		X"A8",X"11",X"20",X"00",X"FE",X"0F",X"38",X"02",X"3E",X"0F",X"47",X"0E",X"4C",X"71",X"19",X"10",
		X"FC",X"C9",X"AF",X"32",X"CC",X"83",X"21",X"B8",X"83",X"3A",X"FD",X"83",X"3D",X"28",X"01",X"2C",
		X"34",X"7E",X"32",X"B7",X"83",X"FE",X"10",X"D0",X"26",X"00",X"11",X"5E",X"A8",X"87",X"87",X"87",
		X"87",X"6F",X"29",X"19",X"36",X"4C",X"C9",X"06",X"05",X"21",X"F2",X"83",X"7A",X"BE",X"38",X"27",
		X"28",X"19",X"78",X"3D",X"28",X"0F",X"87",X"4F",X"06",X"00",X"D5",X"11",X"FA",X"83",X"21",X"F8",
		X"83",X"ED",X"B8",X"EB",X"D1",X"72",X"2D",X"73",X"87",X"3C",X"C9",X"2D",X"7E",X"2C",X"BB",X"38",
		X"E1",X"20",X"04",X"78",X"3D",X"28",X"F1",X"2C",X"2C",X"10",X"D1",X"AF",X"C9",X"3A",X"2D",X"84",
		X"B7",X"C0",X"3C",X"32",X"2D",X"84",X"3E",X"03",X"32",X"3F",X"80",X"AF",X"32",X"E0",X"83",X"21",
		X"BF",X"A8",X"11",X"04",X"10",X"06",X"04",X"EF",X"21",X"DF",X"A8",X"11",X"20",X"00",X"01",X"0C",
		X"0F",X"71",X"19",X"10",X"FC",X"21",X"20",X"3C",X"22",X"DC",X"83",X"3E",X"60",X"32",X"DE",X"83",
		X"C9",X"E5",X"D5",X"21",X"00",X"84",X"35",X"20",X"02",X"36",X"1F",X"54",X"5E",X"7B",X"C6",X"0D",
		X"FE",X"20",X"38",X"02",X"D6",X"1F",X"6F",X"1A",X"AE",X"77",X"D1",X"E1",X"C9",X"21",X"00",X"00",
		X"22",X"ED",X"83",X"22",X"EB",X"83",X"22",X"E7",X"83",X"3A",X"E4",X"83",X"67",X"6F",X"22",X"E5",
		X"83",X"C9",X"11",X"AA",X"0F",X"21",X"60",X"AA",X"06",X"08",X"EF",X"21",X"41",X"AA",X"ED",X"5B",
		X"EF",X"83",X"CD",X"B8",X"0B",X"3E",X"01",X"21",X"20",X"AB",X"CD",X"CC",X"0B",X"11",X"A7",X"0F",
		X"06",X"03",X"EF",X"21",X"41",X"AB",X"ED",X"5B",X"ED",X"83",X"CD",X"B8",X"0B",X"3A",X"70",X"83",
		X"3D",X"C8",X"3E",X"02",X"21",X"00",X"A9",X"CD",X"CC",X"0B",X"11",X"A7",X"0F",X"06",X"03",X"EF",
		X"21",X"21",X"A9",X"ED",X"5B",X"EB",X"83",X"C3",X"B8",X"0B",X"3A",X"B4",X"83",X"B7",X"20",X"11",
		X"3C",X"32",X"B4",X"83",X"21",X"1F",X"A8",X"11",X"20",X"00",X"01",X"10",X"20",X"71",X"19",X"10",
		X"FC",X"11",X"FE",X"0F",X"21",X"7F",X"A9",X"06",X"06",X"EF",X"3E",X"01",X"32",X"3F",X"80",X"21",
		X"9F",X"A8",X"3A",X"E1",X"83",X"C3",X"C3",X"0B",X"CD",X"BE",X"0B",X"AF",X"18",X"0E",X"7A",X"CD",
		X"C3",X"0B",X"7B",X"4F",X"0F",X"0F",X"0F",X"0F",X"CD",X"CC",X"0B",X"79",X"E6",X"0F",X"77",X"7D",
		X"D6",X"20",X"6F",X"D0",X"25",X"C9",X"21",X"D8",X"83",X"35",X"2D",X"AF",X"77",X"32",X"B3",X"83",
		X"CD",X"79",X"07",X"3E",X"03",X"32",X"19",X"80",X"21",X"1F",X"80",X"06",X"05",X"AF",X"77",X"2C",
		X"2C",X"2C",X"2C",X"10",X"F9",X"CD",X"60",X"0C",X"21",X"AC",X"AA",X"11",X"AD",X"0F",X"06",X"0D",
		X"EF",X"3E",X"01",X"26",X"AA",X"ED",X"47",X"87",X"C6",X"CD",X"6F",X"ED",X"57",X"CD",X"CC",X"0B",
		X"ED",X"57",X"08",X"06",X"03",X"EF",X"D9",X"21",X"EF",X"83",X"08",X"47",X"2C",X"2C",X"10",X"FC",
		X"5E",X"2C",X"56",X"26",X"A9",X"87",X"C6",X"ED",X"6F",X"CD",X"B8",X"0B",X"11",X"4B",X"10",X"06",
		X"04",X"EF",X"ED",X"57",X"D9",X"3C",X"FE",X"06",X"20",X"C9",X"11",X"DF",X"0F",X"21",X"3C",X"AB",
		X"06",X"13",X"AF",X"32",X"39",X"80",X"EF",X"C9",X"7A",X"CD",X"4D",X"0C",X"7B",X"4F",X"E6",X"0F",
		X"CD",X"58",X"0C",X"79",X"0F",X"0F",X"0F",X"0F",X"77",X"7D",X"D6",X"20",X"6F",X"D0",X"25",X"C9",
		X"26",X"80",X"ED",X"4B",X"FB",X"83",X"11",X"04",X"30",X"CD",X"6D",X"0C",X"48",X"7A",X"91",X"BA",
		X"C8",X"6F",X"73",X"C9",X"3A",X"D8",X"83",X"B7",X"C0",X"3A",X"D6",X"83",X"FE",X"03",X"CA",X"D6",
		X"0B",X"3A",X"E1",X"83",X"B7",X"C2",X"A6",X"0C",X"3A",X"D6",X"83",X"FE",X"04",X"CA",X"00",X"18",
		X"FE",X"02",X"CA",X"9B",X"3E",X"FE",X"05",X"C0",X"21",X"D8",X"83",X"36",X"30",X"2D",X"AF",X"77",
		X"32",X"15",X"80",X"C3",X"3A",X"0C",X"CD",X"F9",X"07",X"3A",X"BA",X"83",X"B7",X"C0",X"67",X"6F",
		X"22",X"93",X"82",X"22",X"B3",X"81",X"32",X"5B",X"82",X"32",X"9A",X"82",X"3C",X"32",X"BA",X"83",
		X"CD",X"C6",X"32",X"CD",X"17",X"08",X"CD",X"79",X"07",X"CD",X"5E",X"06",X"3E",X"04",X"32",X"1B",
		X"80",X"3E",X"06",X"32",X"29",X"80",X"21",X"28",X"AA",X"11",X"0D",X"10",X"06",X"04",X"EF",X"21",
		X"AD",X"AA",X"13",X"06",X"0C",X"EF",X"CD",X"13",X"0D",X"21",X"74",X"AB",X"11",X"1E",X"10",X"06",
		X"03",X"EF",X"11",X"39",X"10",X"06",X"06",X"EF",X"11",X"3F",X"10",X"06",X"05",X"EF",X"13",X"06",
		X"07",X"EF",X"21",X"94",X"A9",X"ED",X"5B",X"DE",X"0E",X"CD",X"B8",X"0B",X"11",X"4B",X"10",X"06",
		X"04",X"EF",X"C9",X"3A",X"E1",X"83",X"11",X"1E",X"10",X"3D",X"28",X"11",X"3E",X"03",X"32",X"23",
		X"80",X"21",X"11",X"AB",X"06",X"04",X"EF",X"06",X"0D",X"EF",X"36",X"23",X"C9",X"21",X"F1",X"AA",
		X"06",X"04",X"EF",X"11",X"29",X"10",X"06",X"0B",X"EF",X"C9",X"3E",X"03",X"32",X"0D",X"80",X"32",
		X"0F",X"80",X"3A",X"BC",X"83",X"3D",X"32",X"BC",X"83",X"C0",X"3E",X"20",X"32",X"BC",X"83",X"3A",
		X"D7",X"83",X"87",X"16",X"00",X"5F",X"21",X"59",X"0D",X"19",X"E9",X"18",X"46",X"18",X"3A",X"18",
		X"2E",X"18",X"22",X"18",X"16",X"18",X"0A",X"21",X"06",X"AB",X"11",X"40",X"80",X"3E",X"D4",X"18",
		X"3A",X"21",X"A6",X"AA",X"11",X"44",X"80",X"3E",X"D8",X"18",X"30",X"21",X"46",X"AA",X"11",X"48",
		X"80",X"3E",X"DC",X"18",X"26",X"21",X"E6",X"A9",X"11",X"4C",X"80",X"3E",X"F4",X"18",X"1C",X"21",
		X"86",X"A9",X"11",X"50",X"80",X"3E",X"F4",X"18",X"12",X"21",X"26",X"A9",X"11",X"54",X"80",X"3E",
		X"F8",X"18",X"08",X"21",X"C6",X"A8",X"11",X"58",X"80",X"3E",X"D8",X"01",X"1F",X"00",X"77",X"3C",
		X"2C",X"77",X"3C",X"09",X"77",X"3C",X"2C",X"77",X"EB",X"01",X"00",X"04",X"71",X"2C",X"10",X"FC",
		X"21",X"D7",X"83",X"35",X"C0",X"36",X"07",X"AF",X"32",X"BF",X"83",X"32",X"BB",X"83",X"3E",X"05",
		X"32",X"D6",X"83",X"C9",X"3A",X"E1",X"83",X"B7",X"20",X"F4",X"21",X"BF",X"83",X"7E",X"B7",X"20",
		X"2D",X"CD",X"79",X"07",X"CD",X"5E",X"06",X"21",X"40",X"80",X"01",X"03",X"07",X"11",X"00",X"81",
		X"73",X"2C",X"2C",X"71",X"2C",X"72",X"2C",X"10",X"F7",X"21",X"04",X"05",X"22",X"BD",X"83",X"21",
		X"D7",X"83",X"36",X"07",X"21",X"BC",X"83",X"36",X"20",X"21",X"BF",X"83",X"34",X"C9",X"3D",X"20",
		X"5F",X"3A",X"D7",X"83",X"87",X"16",X"00",X"5F",X"21",X"1B",X"0E",X"19",X"E9",X"18",X"34",X"18",
		X"2B",X"18",X"22",X"18",X"19",X"18",X"10",X"18",X"07",X"21",X"40",X"80",X"06",X"31",X"18",X"28",
		X"21",X"44",X"80",X"06",X"49",X"18",X"21",X"21",X"48",X"80",X"06",X"61",X"18",X"1A",X"21",X"4C",
		X"80",X"06",X"79",X"18",X"13",X"21",X"50",X"80",X"06",X"91",X"18",X"0C",X"21",X"54",X"80",X"06",
		X"A9",X"18",X"05",X"21",X"58",X"80",X"06",X"C1",X"CD",X"98",X"0E",X"4F",X"35",X"35",X"35",X"35",
		X"7E",X"2C",X"71",X"B8",X"D0",X"36",X"1E",X"21",X"D7",X"83",X"35",X"C0",X"36",X"14",X"18",X"99",
		X"3D",X"C2",X"3A",X"0D",X"CD",X"98",X"0E",X"D6",X"03",X"4F",X"3A",X"D7",X"83",X"B7",X"CA",X"FF",
		X"0D",X"06",X"07",X"11",X"06",X"00",X"21",X"43",X"80",X"35",X"35",X"35",X"35",X"2D",X"2D",X"71",
		X"19",X"10",X"F6",X"3D",X"32",X"D7",X"83",X"C9",X"E5",X"21",X"BD",X"83",X"35",X"20",X"11",X"36",
		X"08",X"2C",X"35",X"20",X"02",X"36",X"04",X"7E",X"21",X"F1",X"0E",X"85",X"6F",X"7E",X"E1",X"C9",
		X"F1",X"F1",X"C9",X"ED",X"5B",X"ED",X"83",X"2A",X"EB",X"83",X"44",X"4D",X"B7",X"ED",X"52",X"38",
		X"05",X"D5",X"C5",X"D1",X"18",X"01",X"C5",X"CD",X"A7",X"0A",X"D1",X"F5",X"CD",X"A7",X"0A",X"67",
		X"F1",X"6F",X"22",X"FB",X"83",X"C9",X"03",X"05",X"07",X"FF",X"00",X"02",X"04",X"06",X"00",X"20",
		X"00",X"00",X"58",X"01",X"63",X"04",X"63",X"04",X"05",X"02",X"97",X"01",X"58",X"01",X"27",X"01",
		X"05",X"00",X"1F",X"20",X"21",X"20",X"25",X"26",X"27",X"26",X"2C",X"2D",X"2E",X"2D",X"2F",X"30",
		X"31",X"30",X"2C",X"2E",X"30",X"2E",X"2D",X"2F",X"31",X"2F",X"25",X"26",X"27",X"2C",X"2D",X"2E",
		X"2F",X"30",X"31",X"2C",X"2E",X"30",X"2D",X"2F",X"31",X"04",X"04",X"04",X"08",X"08",X"08",X"08",
		X"08",X"08",X"10",X"10",X"10",X"02",X"03",X"03",X"05",X"05",X"06",X"08",X"09",X"54",X"58",X"5A",
		X"5E",X"56",X"5C",X"03",X"03",X"06",X"08",X"10",X"18",X"30",X"50",X"60",X"80",X"C0",X"E0",X"05",
		X"02",X"02",X"02",X"08",X"08",X"05",X"08",X"02",X"08",X"08",X"08",X"0E",X"08",X"08",X"0E",X"08",
		X"0E",X"08",X"0E",X"08",X"0E",X"08",X"05",X"05",X"08",X"05",X"02",X"0B",X"05",X"08",X"FF",X"C0",
		X"02",X"00",X"03",X"00",X"03",X"80",X"01",X"80",X"02",X"80",X"02",X"00",X"02",X"00",X"02",X"80",
		X"03",X"E0",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"00",X"03",X"80",X"02",X"C0",X"02",X"C0",
		X"02",X"80",X"03",X"20",X"02",X"20",X"02",X"10",X"3B",X"8C",X"D9",X"AF",X"7F",X"3C",X"30",X"70",
		X"A9",X"47",X"E7",X"A7",X"FF",X"BC",X"36",X"10",X"F9",X"40",X"D2",X"D7",X"C4",X"37",X"A6",X"9B",
		X"A1",X"00",X"C7",X"AC",X"8D",X"C5",X"06",X"2B",X"25",X"20",X"18",X"19",X"2B",X"23",X"13",X"1F",
		X"22",X"15",X"10",X"22",X"11",X"1E",X"1B",X"19",X"1E",X"17",X"10",X"23",X"24",X"10",X"1E",X"14",
		X"10",X"22",X"14",X"10",X"24",X"18",X"10",X"24",X"18",X"2B",X"20",X"1F",X"19",X"1E",X"24",X"10",
		X"24",X"11",X"12",X"1C",X"15",X"2B",X"17",X"11",X"1D",X"15",X"10",X"1F",X"26",X"15",X"22",X"10",
		X"10",X"10",X"23",X"15",X"17",X"11",X"10",X"10",X"4E",X"10",X"10",X"01",X"09",X"08",X"01",X"10",
		X"10",X"10",X"19",X"1E",X"23",X"15",X"22",X"24",X"10",X"13",X"1F",X"19",X"1E",X"23",X"13",X"22",
		X"15",X"14",X"19",X"24",X"24",X"19",X"1D",X"15",X"10",X"10",X"20",X"15",X"22",X"20",X"25",X"23",
		X"18",X"10",X"23",X"24",X"11",X"22",X"24",X"10",X"12",X"25",X"24",X"24",X"1F",X"1E",X"1F",X"1E",
		X"15",X"10",X"1F",X"22",X"10",X"24",X"27",X"1F",X"10",X"20",X"1C",X"11",X"29",X"15",X"22",X"10",
		X"1F",X"1E",X"1C",X"29",X"12",X"1F",X"1E",X"25",X"23",X"10",X"15",X"28",X"24",X"22",X"11",X"10",
		X"16",X"22",X"1F",X"17",X"23",X"10",X"11",X"16",X"24",X"15",X"22",X"10",X"20",X"24",X"23",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"86",X"83",X"A7",X"C2",X"B0",X"19",X"21",X"D8",X"83",X"7E",X"B7",X"C0",X"36",X"80",X"2D",
		X"7E",X"34",X"21",X"1F",X"18",X"07",X"4F",X"06",X"00",X"09",X"46",X"23",X"66",X"68",X"E9",X"3B",
		X"18",X"68",X"18",X"7A",X"18",X"97",X"18",X"B4",X"18",X"D7",X"18",X"DD",X"18",X"21",X"19",X"38",
		X"19",X"49",X"19",X"5A",X"19",X"77",X"19",X"88",X"19",X"A5",X"19",X"3E",X"06",X"32",X"17",X"80",
		X"32",X"19",X"80",X"32",X"1B",X"80",X"32",X"1D",X"80",X"3E",X"03",X"32",X"21",X"80",X"32",X"23",
		X"80",X"32",X"25",X"80",X"32",X"27",X"80",X"3E",X"01",X"32",X"2B",X"80",X"32",X"2D",X"80",X"32",
		X"31",X"80",X"32",X"2F",X"80",X"C3",X"15",X"19",X"11",X"B5",X"19",X"06",X"18",X"21",X"88",X"AB",
		X"EF",X"06",X"1B",X"21",X"89",X"AB",X"EF",X"C3",X"15",X"19",X"11",X"E8",X"19",X"06",X"14",X"21",
		X"8B",X"AB",X"EF",X"06",X"1A",X"21",X"8C",X"AB",X"EF",X"06",X"15",X"21",X"8D",X"AB",X"EF",X"06",
		X"1A",X"21",X"8E",X"AB",X"EF",X"18",X"7E",X"11",X"45",X"1A",X"06",X"16",X"21",X"90",X"AB",X"EF",
		X"06",X"15",X"21",X"91",X"AB",X"EF",X"06",X"14",X"21",X"92",X"AB",X"EF",X"06",X"0A",X"21",X"93",
		X"AB",X"EF",X"18",X"61",X"11",X"8E",X"1A",X"06",X"15",X"21",X"95",X"AB",X"EF",X"06",X"19",X"21",
		X"96",X"AB",X"EF",X"06",X"14",X"21",X"97",X"AB",X"EF",X"06",X"0E",X"21",X"98",X"AB",X"EF",X"3E",
		X"A0",X"32",X"86",X"83",X"C3",X"1B",X"19",X"21",X"D8",X"83",X"36",X"C0",X"C9",X"CD",X"79",X"07",
		X"3E",X"06",X"32",X"0F",X"80",X"32",X"15",X"80",X"32",X"1B",X"80",X"32",X"25",X"80",X"32",X"2B",
		X"80",X"32",X"33",X"80",X"3E",X"03",X"32",X"0D",X"80",X"32",X"13",X"80",X"32",X"19",X"80",X"32",
		X"21",X"80",X"32",X"23",X"80",X"32",X"29",X"80",X"32",X"2F",X"80",X"32",X"31",X"80",X"AF",X"32",
		X"0B",X"80",X"32",X"1F",X"80",X"21",X"D8",X"83",X"36",X"80",X"C9",X"21",X"D8",X"83",X"36",X"F0",
		X"C9",X"11",X"DE",X"1A",X"06",X"12",X"21",X"85",X"AB",X"EF",X"06",X"13",X"21",X"86",X"AB",X"EF",
		X"06",X"0B",X"21",X"87",X"AB",X"EF",X"18",X"DD",X"11",X"0E",X"1B",X"06",X"15",X"21",X"89",X"AB",
		X"EF",X"06",X"0B",X"21",X"8A",X"AB",X"EF",X"18",X"CC",X"11",X"2E",X"1B",X"06",X"1A",X"21",X"8C",
		X"AB",X"EF",X"06",X"1A",X"21",X"8D",X"AB",X"EF",X"18",X"BB",X"11",X"62",X"1B",X"06",X"18",X"21",
		X"8F",X"AB",X"EF",X"06",X"12",X"21",X"90",X"AB",X"EF",X"06",X"0C",X"21",X"91",X"AB",X"EF",X"06",
		X"0C",X"21",X"92",X"AB",X"EF",X"18",X"9E",X"11",X"A4",X"1B",X"06",X"13",X"21",X"94",X"AB",X"EF",
		X"06",X"0C",X"21",X"95",X"AB",X"EF",X"18",X"8D",X"11",X"C3",X"1B",X"06",X"13",X"21",X"97",X"AB",
		X"EF",X"06",X"14",X"21",X"98",X"AB",X"EF",X"06",X"0D",X"21",X"99",X"AB",X"EF",X"3E",X"A0",X"32",
		X"86",X"83",X"C3",X"1B",X"19",X"3E",X"03",X"32",X"D6",X"83",X"21",X"D8",X"83",X"36",X"C0",X"C9",
		X"21",X"86",X"83",X"35",X"C9",X"1D",X"1F",X"26",X"15",X"10",X"16",X"22",X"1F",X"17",X"10",X"26",
		X"15",X"22",X"24",X"19",X"13",X"11",X"1C",X"1C",X"29",X"10",X"1F",X"22",X"10",X"18",X"1F",X"22",
		X"19",X"2A",X"1F",X"1E",X"24",X"11",X"1C",X"1C",X"29",X"10",X"25",X"23",X"19",X"1E",X"17",X"10",
		X"1A",X"1F",X"29",X"23",X"24",X"19",X"13",X"1B",X"1F",X"12",X"1A",X"15",X"13",X"24",X"10",X"19",
		X"23",X"10",X"24",X"1F",X"10",X"23",X"11",X"16",X"15",X"1C",X"29",X"10",X"1D",X"11",X"1E",X"15",
		X"25",X"26",X"15",X"22",X"10",X"16",X"22",X"1F",X"17",X"10",X"24",X"1F",X"10",X"19",X"24",X"23",
		X"10",X"18",X"1F",X"1D",X"15",X"10",X"27",X"19",X"24",X"18",X"19",X"1E",X"10",X"11",X"1C",X"1C",
		X"1F",X"24",X"24",X"15",X"14",X"10",X"24",X"19",X"1D",X"15",X"10",X"2B",X"23",X"19",X"28",X"24",
		X"29",X"10",X"12",X"15",X"11",X"24",X"23",X"10",X"1F",X"1E",X"10",X"24",X"18",X"15",X"10",X"24",
		X"19",X"1D",X"15",X"22",X"2B",X"13",X"22",X"1F",X"23",X"23",X"10",X"18",X"19",X"17",X"18",X"27",
		X"11",X"29",X"10",X"27",X"19",X"24",X"18",X"1F",X"25",X"24",X"10",X"17",X"15",X"24",X"24",X"19",
		X"1E",X"17",X"10",X"22",X"25",X"1E",X"10",X"1F",X"26",X"15",X"22",X"10",X"11",X"1E",X"14",X"10",
		X"13",X"22",X"1F",X"23",X"23",X"10",X"22",X"19",X"26",X"15",X"22",X"10",X"27",X"19",X"24",X"18",
		X"1F",X"25",X"24",X"10",X"16",X"11",X"1C",X"1C",X"19",X"1E",X"17",X"10",X"19",X"1E",X"11",X"26",
		X"1F",X"19",X"14",X"10",X"24",X"22",X"11",X"16",X"16",X"19",X"13",X"10",X"14",X"15",X"11",X"14",
		X"1C",X"29",X"10",X"23",X"1E",X"11",X"1B",X"15",X"23",X"10",X"1F",X"24",X"24",X"15",X"22",X"23",
		X"10",X"13",X"22",X"1F",X"13",X"1F",X"14",X"19",X"1C",X"15",X"23",X"10",X"11",X"1E",X"14",X"10",
		X"24",X"18",X"15",X"10",X"24",X"22",X"15",X"11",X"13",X"18",X"15",X"22",X"1F",X"25",X"23",X"10",
		X"14",X"19",X"26",X"19",X"1E",X"17",X"10",X"24",X"25",X"22",X"24",X"1C",X"15",X"23",X"20",X"1F",
		X"19",X"1E",X"24",X"23",X"10",X"11",X"22",X"15",X"10",X"23",X"13",X"1F",X"22",X"15",X"14",X"10",
		X"16",X"1F",X"22",X"10",X"15",X"11",X"13",X"18",X"10",X"23",X"11",X"16",X"15",X"10",X"1A",X"25",
		X"1D",X"20",X"10",X"2B",X"01",X"00",X"10",X"20",X"1F",X"19",X"1E",X"24",X"23",X"2B",X"23",X"11",
		X"16",X"15",X"1C",X"29",X"10",X"11",X"22",X"22",X"19",X"26",X"19",X"1E",X"17",X"10",X"18",X"1F",
		X"1D",X"15",X"10",X"2B",X"05",X"00",X"10",X"20",X"1F",X"19",X"1E",X"24",X"23",X"2B",X"11",X"1E",
		X"14",X"10",X"16",X"1F",X"22",X"10",X"12",X"15",X"11",X"24",X"19",X"1E",X"17",X"10",X"24",X"18",
		X"15",X"10",X"24",X"19",X"1D",X"15",X"22",X"10",X"2B",X"01",X"00",X"10",X"20",X"1F",X"19",X"1E",
		X"24",X"23",X"10",X"20",X"15",X"22",X"10",X"12",X"15",X"11",X"24",X"10",X"23",X"11",X"26",X"15",
		X"14",X"2B",X"12",X"1F",X"1E",X"25",X"23",X"10",X"20",X"1F",X"19",X"1E",X"24",X"23",X"10",X"11",
		X"22",X"15",X"10",X"23",X"13",X"1F",X"22",X"15",X"14",X"10",X"12",X"29",X"10",X"15",X"23",X"13",
		X"1F",X"22",X"24",X"19",X"1E",X"17",X"10",X"18",X"1F",X"1D",X"15",X"10",X"11",X"10",X"1C",X"11",
		X"14",X"29",X"10",X"16",X"22",X"1F",X"17",X"10",X"2B",X"02",X"00",X"00",X"10",X"20",X"1F",X"19",
		X"1E",X"24",X"23",X"2B",X"17",X"1F",X"12",X"12",X"1C",X"19",X"1E",X"17",X"10",X"11",X"1E",X"10",
		X"19",X"1E",X"23",X"15",X"13",X"24",X"10",X"2B",X"02",X"00",X"00",X"10",X"20",X"1F",X"19",X"1E",
		X"24",X"23",X"2B",X"11",X"1E",X"14",X"10",X"23",X"11",X"16",X"15",X"1C",X"29",X"10",X"17",X"15",
		X"24",X"24",X"19",X"1E",X"17",X"10",X"11",X"1C",X"1C",X"10",X"16",X"19",X"26",X"15",X"10",X"16",
		X"22",X"1F",X"17",X"23",X"10",X"18",X"1F",X"1D",X"15",X"10",X"2B",X"01",X"00",X"00",X"00",X"10",
		X"20",X"1F",X"19",X"1E",X"24",X"23",X"2B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"B7",X"83",X"FE",X"03",X"38",X"2A",X"3A",X"FD",X"83",X"3D",X"20",X"06",X"DD",X"21",X"40",
		X"84",X"18",X"04",X"DD",X"21",X"60",X"84",X"FD",X"21",X"48",X"80",X"CD",X"49",X"1C",X"3A",X"B7",
		X"83",X"FE",X"06",X"38",X"07",X"11",X"10",X"00",X"DD",X"19",X"FD",X"21",X"50",X"80",X"CD",X"49",
		X"1C",X"3A",X"FD",X"83",X"3D",X"20",X"06",X"DD",X"21",X"80",X"84",X"18",X"04",X"DD",X"21",X"90",
		X"84",X"FD",X"21",X"58",X"80",X"CD",X"13",X"1E",X"C9",X"CD",X"FA",X"1C",X"CD",X"59",X"1C",X"CD",
		X"89",X"1C",X"CD",X"83",X"1D",X"CD",X"E8",X"1D",X"C9",X"DD",X"35",X"08",X"C0",X"DD",X"36",X"08",
		X"0C",X"DD",X"7E",X"06",X"B7",X"C8",X"3D",X"20",X"02",X"3E",X"04",X"DD",X"77",X"06",X"6F",X"26",
		X"00",X"11",X"65",X"1F",X"19",X"7E",X"DD",X"B6",X"05",X"FD",X"77",X"01",X"3C",X"FD",X"77",X"05",
		X"FD",X"36",X"02",X"04",X"FD",X"36",X"06",X"04",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",X"3A",X"2C",
		X"84",X"B7",X"C0",X"DD",X"35",X"09",X"C0",X"DD",X"36",X"09",X"08",X"FD",X"7E",X"03",X"FE",X"60",
		X"30",X"2A",X"DD",X"36",X"07",X"01",X"DD",X"7E",X"05",X"B7",X"C2",X"BD",X"1C",X"3A",X"14",X"80",
		X"DD",X"96",X"00",X"D8",X"FD",X"BE",X"00",X"30",X"2A",X"DD",X"34",X"02",X"C9",X"3A",X"14",X"80",
		X"DD",X"96",X"01",X"FD",X"BE",X"00",X"38",X"1B",X"DD",X"35",X"02",X"C9",X"DD",X"36",X"07",X"01",
		X"DD",X"7E",X"05",X"B7",X"28",X"04",X"3E",X"02",X"18",X"02",X"3E",X"FE",X"DD",X"86",X"03",X"DD",
		X"77",X"03",X"C9",X"DD",X"7E",X"05",X"EE",X"80",X"DD",X"77",X"05",X"FD",X"7E",X"04",X"FD",X"77",
		X"00",X"FD",X"7E",X"01",X"EE",X"80",X"FD",X"77",X"01",X"C9",X"3A",X"B7",X"83",X"FE",X"03",X"D8",
		X"4F",X"DD",X"35",X"0A",X"C0",X"DD",X"7E",X"06",X"B7",X"C0",X"CD",X"11",X"0B",X"47",X"79",X"87",
		X"87",X"87",X"C6",X"80",X"B8",X"D8",X"CD",X"11",X"0B",X"E6",X"03",X"28",X"1D",X"0E",X"40",X"21",
		X"76",X"82",X"7E",X"0F",X"0F",X"C6",X"24",X"57",X"2C",X"2C",X"46",X"3A",X"14",X"80",X"D6",X"10",
		X"38",X"08",X"91",X"38",X"19",X"92",X"38",X"02",X"10",X"F8",X"DD",X"36",X"04",X"7E",X"CD",X"11",
		X"0B",X"0F",X"38",X"1E",X"DD",X"36",X"05",X"00",X"DD",X"36",X"03",X"F0",X"18",X"1C",X"81",X"47",
		X"3A",X"14",X"80",X"DD",X"77",X"02",X"90",X"DD",X"77",X"01",X"81",X"DD",X"77",X"00",X"DD",X"36",
		X"04",X"4E",X"DD",X"36",X"05",X"80",X"DD",X"36",X"03",X"00",X"DD",X"36",X"06",X"01",X"DD",X"36",
		X"08",X"0B",X"DD",X"36",X"09",X"08",X"3A",X"71",X"83",X"B7",X"C0",X"3C",X"32",X"71",X"83",X"3E",
		X"90",X"DF",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",X"CD",X"76",X"1D",X"DD",X"7E",X"04",X"FE",X"60",
		X"30",X"0C",X"3A",X"14",X"80",X"DD",X"96",X"02",X"4F",X"FD",X"77",X"00",X"18",X"06",X"DD",X"4E",
		X"03",X"FD",X"71",X"00",X"DD",X"7E",X"04",X"FD",X"77",X"03",X"FD",X"77",X"07",X"DD",X"7E",X"05",
		X"B7",X"20",X"0A",X"3E",X"0F",X"81",X"FD",X"77",X"04",X"3C",X"C0",X"18",X"09",X"3E",X"F1",X"81",
		X"FD",X"77",X"04",X"79",X"B7",X"C0",X"DD",X"7E",X"07",X"B7",X"C8",X"DD",X"E5",X"E1",X"54",X"5D",
		X"1C",X"01",X"0F",X"00",X"70",X"ED",X"B0",X"01",X"07",X"00",X"FD",X"E5",X"E1",X"54",X"5D",X"1C",
		X"70",X"ED",X"B0",X"DD",X"36",X"0A",X"20",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",X"DD",X"7E",X"04",
		X"C6",X"02",X"21",X"47",X"80",X"BE",X"C0",X"DD",X"7E",X"05",X"B7",X"FD",X"7E",X"00",X"21",X"44",
		X"80",X"28",X"02",X"C6",X"10",X"96",X"D8",X"FE",X"10",X"D0",X"3E",X"01",X"32",X"04",X"80",X"32",
		X"2C",X"84",X"C9",X"CD",X"A3",X"1E",X"CD",X"3B",X"1E",X"CD",X"23",X"1E",X"CD",X"38",X"1F",X"CD",
		X"8B",X"1E",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",X"DD",X"6E",X"0B",X"26",X"80",X"7E",X"DD",X"96",
		X"02",X"FD",X"77",X"00",X"DD",X"7E",X"04",X"FD",X"77",X"03",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",
		X"DD",X"35",X"09",X"C0",X"DD",X"36",X"09",X"08",X"DD",X"6E",X"0B",X"26",X"80",X"DD",X"7E",X"05",
		X"B7",X"28",X"0D",X"7E",X"DD",X"96",X"00",X"FD",X"BE",X"00",X"30",X"11",X"DD",X"34",X"02",X"C9",
		X"7E",X"DD",X"96",X"01",X"FD",X"BE",X"00",X"38",X"04",X"DD",X"35",X"02",X"C9",X"3A",X"04",X"80",
		X"B7",X"C0",X"DD",X"E5",X"E1",X"54",X"5D",X"1C",X"01",X"0F",X"00",X"70",X"ED",X"B0",X"21",X"58",
		X"80",X"11",X"59",X"80",X"01",X"03",X"00",X"70",X"ED",X"B0",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",
		X"21",X"69",X"1F",X"4F",X"06",X"00",X"09",X"7E",X"DD",X"B6",X"05",X"FD",X"77",X"01",X"FD",X"36",
		X"02",X"02",X"C9",X"3A",X"B7",X"83",X"FE",X"03",X"D8",X"4F",X"DD",X"7E",X"06",X"B7",X"C0",X"CD",
		X"11",X"0B",X"47",X"79",X"87",X"87",X"87",X"C6",X"80",X"B8",X"D8",X"0E",X"40",X"CD",X"11",X"0B",
		X"E6",X"07",X"FE",X"05",X"D0",X"4F",X"0F",X"0F",X"0F",X"0F",X"C6",X"30",X"DD",X"77",X"04",X"CD",
		X"11",X"0B",X"47",X"79",X"87",X"5F",X"16",X"00",X"21",X"76",X"1F",X"19",X"5E",X"2C",X"6E",X"26",
		X"80",X"DD",X"75",X"0B",X"7E",X"57",X"79",X"87",X"4F",X"06",X"00",X"21",X"6C",X"1F",X"09",X"4E",
		X"2C",X"66",X"69",X"7E",X"0F",X"0F",X"D6",X"10",X"4F",X"2C",X"2C",X"46",X"7A",X"93",X"D8",X"91",
		X"38",X"02",X"10",X"F9",X"81",X"47",X"DD",X"6E",X"0B",X"26",X"80",X"7E",X"DD",X"77",X"02",X"90",
		X"DD",X"77",X"01",X"81",X"DD",X"77",X"00",X"CD",X"11",X"0B",X"0F",X"38",X"0A",X"DD",X"36",X"05",
		X"80",X"DD",X"36",X"03",X"F0",X"18",X"08",X"DD",X"36",X"05",X"00",X"DD",X"36",X"03",X"00",X"DD",
		X"36",X"06",X"01",X"DD",X"36",X"09",X"08",X"C9",X"DD",X"7E",X"06",X"B7",X"C8",X"DD",X"7E",X"04",
		X"21",X"47",X"80",X"BE",X"C0",X"DD",X"7E",X"05",X"B7",X"FD",X"7E",X"00",X"21",X"44",X"80",X"20",
		X"04",X"C6",X"14",X"18",X"02",X"D6",X"04",X"96",X"D8",X"FE",X"10",X"D0",X"3E",X"01",X"32",X"04",
		X"80",X"DD",X"36",X"06",X"02",X"C9",X"2C",X"2E",X"30",X"2E",X"27",X"38",X"70",X"82",X"73",X"82",
		X"76",X"82",X"79",X"82",X"7C",X"82",X"50",X"0C",X"30",X"10",X"70",X"14",X"40",X"18",X"40",X"1C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"18",X"81",X"A7",X"C8",X"11",X"06",X"A8",X"06",X"08",X"21",X"9C",X"24",X"7E",X"12",X"23",
		X"13",X"7E",X"12",X"23",X"C5",X"01",X"1F",X"00",X"EB",X"09",X"EB",X"C1",X"10",X"EF",X"AF",X"32",
		X"18",X"81",X"C9",X"2A",X"00",X"80",X"01",X"32",X"20",X"26",X"00",X"29",X"09",X"4E",X"23",X"66",
		X"69",X"E9",X"48",X"20",X"E1",X"20",X"04",X"21",X"24",X"21",X"44",X"21",X"64",X"21",X"81",X"21",
		X"A1",X"21",X"C1",X"21",X"E1",X"21",X"01",X"22",X"21",X"70",X"82",X"7E",X"23",X"46",X"23",X"4E",
		X"2A",X"76",X"24",X"11",X"8C",X"24",X"DD",X"21",X"00",X"81",X"FD",X"21",X"00",X"81",X"32",X"B1",
		X"81",X"ED",X"53",X"01",X"80",X"E5",X"C5",X"D5",X"CD",X"21",X"22",X"3A",X"5B",X"82",X"A7",X"20",
		X"0B",X"79",X"2F",X"3C",X"DD",X"77",X"01",X"DD",X"23",X"FD",X"34",X"00",X"D1",X"C1",X"E1",X"78",
		X"32",X"03",X"80",X"1A",X"77",X"23",X"13",X"1A",X"77",X"2B",X"D5",X"11",X"20",X"00",X"19",X"D1",
		X"10",X"1A",X"3A",X"B1",X"81",X"5F",X"16",X"00",X"19",X"0D",X"C2",X"B0",X"20",X"21",X"00",X"80",
		X"34",X"7E",X"FE",X"0B",X"DA",X"23",X"20",X"AF",X"77",X"C3",X"BB",X"20",X"13",X"C3",X"83",X"20",
		X"ED",X"5B",X"01",X"80",X"3A",X"03",X"80",X"47",X"C3",X"65",X"20",X"C9",X"01",X"FF",X"03",X"21",
		X"00",X"A8",X"3A",X"00",X"88",X"36",X"28",X"23",X"0B",X"78",X"A7",X"20",X"F5",X"79",X"A7",X"20",
		X"F1",X"01",X"FF",X"EF",X"3A",X"00",X"88",X"0B",X"78",X"A7",X"20",X"F8",X"79",X"A7",X"20",X"F4",
		X"C9",X"CD",X"00",X"20",X"21",X"73",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"78",X"24",X"11",
		X"AC",X"24",X"DD",X"21",X"09",X"81",X"FD",X"21",X"09",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",
		X"80",X"C3",X"65",X"20",X"21",X"76",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"7A",X"24",X"11",
		X"C4",X"24",X"DD",X"21",X"12",X"81",X"FD",X"21",X"12",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",
		X"80",X"C3",X"65",X"20",X"21",X"79",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"7C",X"24",X"11",
		X"DC",X"24",X"DD",X"21",X"1B",X"81",X"FD",X"21",X"1B",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",
		X"80",X"C3",X"65",X"20",X"21",X"7C",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"7E",X"24",X"11",
		X"E8",X"24",X"DD",X"21",X"24",X"81",X"FD",X"21",X"24",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",
		X"80",X"C3",X"65",X"20",X"C3",X"9D",X"20",X"11",X"24",X"25",X"01",X"04",X"02",X"DD",X"21",X"2D",
		X"81",X"FD",X"21",X"2D",X"81",X"3E",X"80",X"32",X"B1",X"81",X"ED",X"53",X"01",X"80",X"C3",X"65",
		X"20",X"21",X"82",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"82",X"24",X"11",X"28",X"25",X"DD",
		X"21",X"36",X"81",X"FD",X"21",X"36",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",X"80",X"C3",X"65",
		X"20",X"21",X"85",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"84",X"24",X"11",X"30",X"25",X"DD",
		X"21",X"3F",X"81",X"FD",X"21",X"3F",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",X"80",X"C3",X"65",
		X"20",X"21",X"88",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"86",X"24",X"11",X"34",X"25",X"DD",
		X"21",X"48",X"81",X"FD",X"21",X"48",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",X"80",X"C3",X"65",
		X"20",X"21",X"8B",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"88",X"24",X"11",X"38",X"25",X"DD",
		X"21",X"51",X"81",X"FD",X"21",X"51",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",X"80",X"C3",X"65",
		X"20",X"21",X"8E",X"82",X"7E",X"23",X"46",X"23",X"4E",X"2A",X"8A",X"24",X"11",X"3C",X"25",X"DD",
		X"21",X"5A",X"81",X"FD",X"21",X"5A",X"81",X"32",X"B1",X"81",X"ED",X"53",X"01",X"80",X"C3",X"65",
		X"20",X"11",X"00",X"A8",X"ED",X"52",X"7D",X"01",X"00",X"06",X"E6",X"E0",X"6F",X"7C",X"E6",X"04",
		X"CA",X"39",X"22",X"CB",X"01",X"0C",X"C3",X"3B",X"22",X"CB",X"01",X"CB",X"05",X"CB",X"14",X"10",
		X"EC",X"CB",X"01",X"CB",X"01",X"CB",X"01",X"C9",X"3A",X"CD",X"83",X"B7",X"C0",X"3A",X"04",X"80",
		X"A7",X"C0",X"21",X"47",X"80",X"7E",X"4F",X"E6",X"0F",X"FE",X"09",X"D2",X"92",X"22",X"79",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"6F",X"26",X"00",X"01",X"72",X"22",X"29",X"09",X"4E",X"23",X"66",
		X"69",X"E9",X"92",X"22",X"95",X"22",X"98",X"22",X"9B",X"22",X"A3",X"22",X"AB",X"22",X"B3",X"22",
		X"BB",X"22",X"C3",X"22",X"CB",X"22",X"D3",X"22",X"DB",X"22",X"E3",X"22",X"EB",X"22",X"F3",X"22",
		X"F6",X"22",X"C3",X"6D",X"23",X"C3",X"6D",X"23",X"C3",X"6D",X"23",X"21",X"00",X"81",X"0E",X"3C",
		X"C3",X"F9",X"22",X"21",X"09",X"81",X"0E",X"1F",X"C3",X"F9",X"22",X"21",X"12",X"81",X"0E",X"5C",
		X"C3",X"F9",X"22",X"21",X"1B",X"81",X"0E",X"2C",X"C3",X"F9",X"22",X"21",X"24",X"81",X"0E",X"2F",
		X"C3",X"F9",X"22",X"C3",X"6D",X"23",X"0E",X"17",X"C3",X"F9",X"22",X"21",X"36",X"81",X"0E",X"22",
		X"C3",X"F9",X"22",X"21",X"3F",X"81",X"0E",X"12",X"C3",X"F9",X"22",X"21",X"48",X"81",X"0E",X"12",
		X"C3",X"F9",X"22",X"21",X"51",X"81",X"0E",X"12",X"C3",X"F9",X"22",X"21",X"5A",X"81",X"0E",X"12",
		X"C3",X"F9",X"22",X"C3",X"6D",X"23",X"C3",X"6D",X"23",X"3A",X"47",X"80",X"FE",X"80",X"DA",X"22",
		X"23",X"3A",X"44",X"80",X"C6",X"03",X"57",X"81",X"5F",X"46",X"DA",X"2A",X"23",X"23",X"7E",X"BA",
		X"DA",X"3F",X"23",X"BB",X"D2",X"3F",X"23",X"3A",X"47",X"80",X"FE",X"80",X"DA",X"6D",X"23",X"C3",
		X"59",X"23",X"3A",X"44",X"80",X"C6",X"0C",X"C3",X"06",X"23",X"23",X"7E",X"BA",X"D2",X"34",X"23",
		X"BB",X"D2",X"4C",X"23",X"3A",X"47",X"80",X"FE",X"80",X"DA",X"6D",X"23",X"C3",X"59",X"23",X"10",
		X"CC",X"3A",X"47",X"80",X"FE",X"80",X"DA",X"59",X"23",X"C3",X"6D",X"23",X"10",X"DC",X"3A",X"47",
		X"80",X"FE",X"80",X"DA",X"59",X"23",X"C3",X"6D",X"23",X"3E",X"01",X"32",X"04",X"80",X"3A",X"47",
		X"80",X"FE",X"80",X"D0",X"FE",X"30",X"D8",X"3E",X"01",X"32",X"9C",X"82",X"C9",X"3A",X"04",X"80",
		X"A7",X"C0",X"21",X"47",X"80",X"7E",X"C6",X"0F",X"4F",X"E6",X"0F",X"FE",X"05",X"DA",X"B4",X"23",
		X"79",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"6F",X"26",X"00",X"01",X"94",X"23",X"29",X"09",X"4E",
		X"23",X"66",X"69",X"E9",X"B4",X"23",X"B7",X"23",X"BA",X"23",X"BD",X"23",X"C5",X"23",X"CD",X"23",
		X"D5",X"23",X"DD",X"23",X"E5",X"23",X"ED",X"23",X"F5",X"23",X"FD",X"23",X"05",X"24",X"0D",X"24",
		X"15",X"24",X"15",X"24",X"C3",X"6A",X"24",X"C3",X"6A",X"24",X"C3",X"6A",X"24",X"21",X"00",X"81",
		X"0E",X"3C",X"C3",X"18",X"24",X"21",X"09",X"81",X"0E",X"1F",X"C3",X"18",X"24",X"21",X"12",X"81",
		X"0E",X"5C",X"C3",X"18",X"24",X"21",X"1B",X"81",X"0E",X"2C",X"C3",X"18",X"24",X"21",X"24",X"81",
		X"0E",X"2F",X"C3",X"18",X"24",X"C3",X"6A",X"24",X"0E",X"17",X"C3",X"18",X"24",X"21",X"36",X"81",
		X"0E",X"22",X"C3",X"18",X"24",X"21",X"3F",X"81",X"0E",X"12",X"C3",X"18",X"24",X"21",X"48",X"81",
		X"0E",X"12",X"C3",X"18",X"24",X"21",X"51",X"81",X"0E",X"12",X"C3",X"18",X"24",X"21",X"5A",X"81",
		X"0E",X"12",X"C3",X"18",X"24",X"C3",X"6A",X"24",X"3A",X"2F",X"80",X"FE",X"80",X"DA",X"42",X"24",
		X"3A",X"44",X"80",X"C6",X"03",X"57",X"81",X"5F",X"46",X"DA",X"4A",X"24",X"23",X"7E",X"BA",X"DA",
		X"60",X"24",X"BB",X"D2",X"60",X"24",X"3A",X"47",X"80",X"FE",X"80",X"D8",X"3E",X"01",X"32",X"04",
		X"80",X"C9",X"3A",X"44",X"80",X"C6",X"0C",X"C3",X"25",X"24",X"23",X"7E",X"BA",X"D2",X"54",X"24",
		X"BB",X"D2",X"6B",X"24",X"3A",X"47",X"80",X"FE",X"80",X"D8",X"3E",X"01",X"32",X"04",X"80",X"C9",
		X"10",X"CA",X"3A",X"47",X"80",X"FE",X"80",X"DA",X"59",X"23",X"C9",X"10",X"DD",X"3A",X"47",X"80",
		X"FE",X"80",X"DA",X"59",X"23",X"C9",X"06",X"A8",X"08",X"A8",X"0A",X"A8",X"0C",X"A8",X"0E",X"A8",
		X"10",X"A8",X"12",X"A8",X"14",X"A8",X"16",X"A8",X"18",X"A8",X"1A",X"A8",X"5C",X"5D",X"5E",X"5F",
		X"58",X"59",X"5A",X"5B",X"58",X"59",X"5A",X"5B",X"54",X"55",X"56",X"57",X"10",X"10",X"10",X"10",
		X"D0",X"D1",X"D2",X"D3",X"CC",X"CD",X"CE",X"CF",X"C8",X"C9",X"CA",X"CB",X"34",X"35",X"36",X"37",
		X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",
		X"3C",X"3D",X"3E",X"3F",X"5C",X"5D",X"5E",X"5F",X"58",X"59",X"5A",X"5B",X"58",X"59",X"5A",X"5B",
		X"58",X"59",X"5A",X"5B",X"58",X"59",X"5A",X"5B",X"54",X"55",X"56",X"57",X"5C",X"5D",X"5E",X"5F",
		X"58",X"59",X"5A",X"5B",X"54",X"55",X"56",X"57",X"34",X"35",X"36",X"37",X"34",X"35",X"36",X"37",
		X"34",X"35",X"36",X"37",X"34",X"35",X"36",X"37",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",
		X"38",X"39",X"3A",X"3B",X"38",X"39",X"3A",X"3B",X"38",X"39",X"3A",X"3B",X"38",X"39",X"3A",X"3B",
		X"3C",X"3D",X"3E",X"3F",X"3C",X"3D",X"3E",X"3F",X"3C",X"3D",X"3E",X"3F",X"3C",X"3D",X"3E",X"3F",
		X"3C",X"3D",X"3E",X"3F",X"47",X"47",X"47",X"47",X"AC",X"AD",X"AE",X"AF",X"A8",X"A9",X"AA",X"AB",
		X"A0",X"A1",X"A2",X"A3",X"30",X"31",X"32",X"33",X"A4",X"A5",X"A6",X"A7",X"50",X"51",X"52",X"53",
		X"3A",X"FF",X"80",X"01",X"50",X"25",X"26",X"00",X"87",X"6F",X"09",X"4E",X"23",X"66",X"69",X"E9",
		X"66",X"25",X"77",X"25",X"88",X"25",X"99",X"25",X"AA",X"25",X"BB",X"25",X"CC",X"25",X"DD",X"25",
		X"EE",X"25",X"FF",X"25",X"10",X"26",X"21",X"9B",X"81",X"11",X"00",X"81",X"DD",X"21",X"0C",X"80",
		X"FD",X"21",X"A6",X"81",X"C3",X"21",X"26",X"21",X"9C",X"81",X"11",X"09",X"81",X"DD",X"21",X"10",
		X"80",X"FD",X"21",X"A7",X"81",X"C3",X"C7",X"26",X"21",X"9D",X"81",X"11",X"12",X"81",X"DD",X"21",
		X"14",X"80",X"FD",X"21",X"A8",X"81",X"C3",X"21",X"26",X"21",X"9E",X"81",X"11",X"1B",X"81",X"DD",
		X"21",X"18",X"80",X"FD",X"21",X"A9",X"81",X"C3",X"21",X"26",X"21",X"9F",X"81",X"11",X"24",X"81",
		X"DD",X"21",X"1C",X"80",X"FD",X"21",X"AA",X"81",X"C3",X"C7",X"26",X"C3",X"67",X"26",X"11",X"2D",
		X"81",X"DD",X"21",X"20",X"80",X"FD",X"21",X"AB",X"81",X"C3",X"21",X"26",X"21",X"A1",X"81",X"11",
		X"36",X"81",X"DD",X"21",X"24",X"80",X"FD",X"21",X"AC",X"81",X"C3",X"C7",X"26",X"21",X"A2",X"81",
		X"11",X"3F",X"81",X"DD",X"21",X"28",X"80",X"FD",X"21",X"AD",X"81",X"C3",X"21",X"26",X"21",X"A3",
		X"81",X"11",X"48",X"81",X"DD",X"21",X"2C",X"80",X"FD",X"21",X"AE",X"81",X"C3",X"C7",X"26",X"21",
		X"A4",X"81",X"11",X"51",X"81",X"DD",X"21",X"30",X"80",X"FD",X"21",X"AF",X"81",X"C3",X"21",X"26",
		X"21",X"A5",X"81",X"11",X"5A",X"81",X"DD",X"21",X"34",X"80",X"FD",X"21",X"B0",X"81",X"C3",X"C7",
		X"26",X"FD",X"7E",X"00",X"4F",X"A7",X"C2",X"5D",X"27",X"7E",X"47",X"E6",X"0F",X"4F",X"78",X"E6",
		X"10",X"C2",X"5D",X"27",X"1A",X"47",X"13",X"1A",X"81",X"12",X"10",X"FA",X"DD",X"7E",X"00",X"81",
		X"DD",X"77",X"00",X"DD",X"77",X"02",X"3A",X"47",X"80",X"FE",X"30",X"DA",X"63",X"26",X"3A",X"47",
		X"80",X"FE",X"73",X"D2",X"63",X"26",X"47",X"E6",X"0F",X"FE",X"03",X"DA",X"74",X"26",X"FE",X"0C",
		X"D2",X"A8",X"26",X"FD",X"36",X"00",X"00",X"21",X"FF",X"80",X"34",X"7E",X"FE",X"0B",X"DA",X"40",
		X"25",X"36",X"00",X"C9",X"78",X"E6",X"F0",X"08",X"08",X"D6",X"30",X"0F",X"0F",X"0F",X"0F",X"47",
		X"3A",X"FF",X"80",X"B8",X"C2",X"63",X"26",X"3A",X"47",X"80",X"FE",X"30",X"DA",X"63",X"26",X"3A",
		X"44",X"80",X"81",X"32",X"44",X"80",X"FE",X"08",X"DA",X"A0",X"26",X"FE",X"E7",X"DA",X"63",X"26",
		X"3E",X"01",X"32",X"04",X"80",X"C3",X"63",X"26",X"78",X"E6",X"F0",X"C6",X"10",X"08",X"08",X"D6",
		X"30",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"FF",X"80",X"B8",X"C2",X"63",X"26",X"3A",X"44",X"80",
		X"81",X"32",X"44",X"80",X"C3",X"63",X"26",X"FD",X"7E",X"00",X"4F",X"A7",X"C2",X"6F",X"27",X"7E",
		X"47",X"E6",X"0F",X"4F",X"78",X"E6",X"10",X"C2",X"6F",X"27",X"1A",X"47",X"13",X"1A",X"91",X"12",
		X"10",X"FA",X"DD",X"7E",X"00",X"91",X"DD",X"77",X"00",X"DD",X"77",X"02",X"3A",X"47",X"80",X"FE",
		X"73",X"D2",X"01",X"27",X"47",X"E6",X"0F",X"FE",X"03",X"DA",X"12",X"27",X"FE",X"0C",X"D2",X"3E",
		X"27",X"FD",X"36",X"00",X"00",X"21",X"FF",X"80",X"34",X"7E",X"FE",X"0B",X"DA",X"40",X"25",X"36",
		X"00",X"C9",X"78",X"E6",X"F0",X"08",X"08",X"D6",X"30",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"FF",
		X"80",X"B8",X"C2",X"01",X"27",X"3A",X"44",X"80",X"91",X"32",X"44",X"80",X"FE",X"08",X"DA",X"36",
		X"27",X"FE",X"E7",X"DA",X"01",X"27",X"3E",X"01",X"32",X"04",X"80",X"C3",X"01",X"27",X"78",X"E6",
		X"F0",X"C6",X"10",X"08",X"08",X"D6",X"30",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"FF",X"80",X"B8",
		X"C2",X"01",X"27",X"3A",X"44",X"80",X"91",X"32",X"44",X"80",X"C3",X"01",X"27",X"79",X"FE",X"01",
		X"C2",X"68",X"27",X"0E",X"01",X"C3",X"34",X"26",X"0D",X"FD",X"71",X"00",X"C3",X"67",X"26",X"79",
		X"FE",X"01",X"C2",X"7A",X"27",X"0E",X"01",X"C3",X"DA",X"26",X"0D",X"FD",X"71",X"00",X"C3",X"05",
		X"27",X"3A",X"04",X"80",X"A7",X"C8",X"3A",X"50",X"81",X"CB",X"47",X"28",X"05",X"3E",X"01",X"32",
		X"18",X"81",X"3A",X"20",X"81",X"A7",X"28",X"03",X"32",X"21",X"81",X"CD",X"57",X"36",X"CD",X"3C",
		X"38",X"3A",X"47",X"82",X"3C",X"32",X"47",X"82",X"D6",X"10",X"C0",X"32",X"47",X"82",X"3E",X"07",
		X"32",X"46",X"80",X"21",X"44",X"80",X"3A",X"B2",X"81",X"3C",X"32",X"B2",X"81",X"4F",X"3A",X"9C",
		X"82",X"A7",X"C2",X"06",X"28",X"79",X"FE",X"06",X"20",X"44",X"CD",X"17",X"08",X"AF",X"32",X"B2",
		X"81",X"32",X"04",X"80",X"32",X"47",X"82",X"32",X"69",X"82",X"32",X"9C",X"82",X"21",X"48",X"82",
		X"11",X"49",X"82",X"01",X"0B",X"00",X"77",X"ED",X"B0",X"3C",X"32",X"CE",X"83",X"3A",X"D6",X"83",
		X"3D",X"20",X"12",X"3A",X"FE",X"83",X"A7",X"20",X"0C",X"32",X"D6",X"83",X"32",X"99",X"82",X"32",
		X"9A",X"82",X"32",X"5B",X"82",X"C9",X"79",X"FE",X"05",X"20",X"03",X"C3",X"CA",X"27",X"3A",X"9C",
		X"82",X"A7",X"C2",X"4D",X"28",X"23",X"3A",X"B2",X"81",X"3D",X"28",X"0B",X"3D",X"28",X"15",X"3D",
		X"28",X"15",X"3D",X"28",X"15",X"18",X"16",X"36",X"39",X"AF",X"67",X"6F",X"22",X"82",X"83",X"DF",
		X"3E",X"03",X"DF",X"C9",X"36",X"39",X"C9",X"36",X"3A",X"C9",X"36",X"3B",X"C9",X"36",X"3C",X"AF",
		X"32",X"AE",X"83",X"CD",X"DF",X"38",X"21",X"D8",X"00",X"22",X"82",X"83",X"C9",X"23",X"3A",X"B2",
		X"81",X"3D",X"28",X"08",X"3D",X"28",X"12",X"3D",X"28",X"12",X"18",X"13",X"36",X"22",X"AF",X"67",
		X"6F",X"22",X"82",X"83",X"DF",X"3E",X"02",X"DF",X"C9",X"36",X"23",X"C9",X"36",X"24",X"C9",X"36",
		X"3C",X"AF",X"32",X"AE",X"83",X"32",X"10",X"81",X"32",X"07",X"81",X"32",X"1A",X"81",X"32",X"19",
		X"81",X"CD",X"DF",X"38",X"21",X"D8",X"00",X"22",X"82",X"83",X"C9",X"3A",X"4F",X"81",X"A7",X"C0",
		X"3A",X"5B",X"81",X"A7",X"C0",X"3A",X"B4",X"81",X"A7",X"C2",X"BB",X"28",X"67",X"3A",X"B3",X"81",
		X"6F",X"11",X"CA",X"28",X"29",X"19",X"4E",X"23",X"66",X"69",X"EB",X"21",X"B3",X"81",X"34",X"7E",
		X"23",X"36",X"15",X"D6",X"0A",X"C2",X"C0",X"28",X"2B",X"77",X"C9",X"21",X"B4",X"81",X"35",X"C9",
		X"EB",X"11",X"9B",X"81",X"01",X"0B",X"00",X"ED",X"B0",X"C9",X"F4",X"28",X"FF",X"28",X"0A",X"29",
		X"15",X"29",X"20",X"29",X"2B",X"29",X"36",X"29",X"41",X"29",X"4C",X"29",X"57",X"29",X"62",X"29",
		X"6D",X"29",X"78",X"29",X"83",X"29",X"8E",X"29",X"99",X"29",X"A4",X"29",X"AF",X"29",X"BA",X"29",
		X"C5",X"29",X"D0",X"29",X"13",X"12",X"11",X"16",X"12",X"00",X"12",X"13",X"14",X"15",X"16",X"12",
		X"13",X"12",X"15",X"01",X"00",X"13",X"02",X"12",X"13",X"12",X"12",X"12",X"13",X"14",X"12",X"00",
		X"12",X"01",X"13",X"12",X"13",X"12",X"01",X"12",X"13",X"13",X"00",X"12",X"02",X"12",X"01",X"14",
		X"13",X"12",X"01",X"12",X"12",X"00",X"12",X"01",X"01",X"12",X"13",X"13",X"01",X"12",X"13",X"13",
		X"00",X"01",X"02",X"12",X"13",X"12",X"12",X"12",X"13",X"12",X"12",X"00",X"12",X"01",X"13",X"12",
		X"13",X"13",X"13",X"12",X"13",X"01",X"00",X"13",X"02",X"12",X"01",X"12",X"12",X"12",X"13",X"12",
		X"12",X"00",X"12",X"01",X"01",X"12",X"13",X"13",X"01",X"12",X"01",X"13",X"00",X"01",X"02",X"12",
		X"13",X"13",X"12",X"12",X"01",X"12",X"12",X"00",X"01",X"01",X"13",X"12",X"12",X"01",X"13",X"01",
		X"13",X"01",X"00",X"12",X"01",X"12",X"01",X"01",X"12",X"12",X"01",X"12",X"12",X"00",X"01",X"02",
		X"13",X"12",X"01",X"01",X"12",X"01",X"12",X"01",X"00",X"01",X"03",X"12",X"01",X"12",X"12",X"12",
		X"01",X"12",X"12",X"00",X"01",X"02",X"13",X"12",X"12",X"01",X"01",X"12",X"01",X"12",X"00",X"01",
		X"01",X"12",X"01",X"01",X"01",X"01",X"12",X"01",X"12",X"00",X"01",X"01",X"12",X"01",X"01",X"12",
		X"01",X"13",X"12",X"01",X"00",X"12",X"02",X"01",X"12",X"12",X"01",X"12",X"14",X"01",X"12",X"00",
		X"01",X"03",X"12",X"13",X"01",X"12",X"01",X"13",X"12",X"13",X"00",X"12",X"02",X"13",X"12",X"12",
		X"13",X"12",X"12",X"13",X"12",X"00",X"13",X"01",X"14",X"13",X"14",X"21",X"43",X"A8",X"0E",X"05",
		X"11",X"7F",X"2A",X"06",X"04",X"1A",X"77",X"13",X"C5",X"01",X"20",X"00",X"09",X"C1",X"10",X"F5",
		X"11",X"40",X"00",X"19",X"0D",X"C2",X"E0",X"29",X"21",X"A4",X"A8",X"0E",X"04",X"11",X"83",X"2A",
		X"06",X"04",X"1A",X"77",X"13",X"C5",X"01",X"20",X"00",X"09",X"C1",X"10",X"F5",X"11",X"40",X"00",
		X"19",X"0D",X"C2",X"FD",X"29",X"21",X"A5",X"A8",X"0E",X"04",X"11",X"87",X"2A",X"06",X"04",X"1A",
		X"77",X"13",X"C5",X"01",X"20",X"00",X"09",X"C1",X"10",X"F5",X"11",X"40",X"00",X"19",X"0D",X"C2",
		X"1A",X"2A",X"21",X"C3",X"A8",X"06",X"04",X"36",X"47",X"11",X"20",X"00",X"19",X"36",X"47",X"11",
		X"A0",X"00",X"19",X"10",X"F2",X"21",X"44",X"A8",X"36",X"41",X"23",X"36",X"42",X"01",X"5F",X"03",
		X"09",X"36",X"45",X"23",X"36",X"46",X"21",X"5C",X"A8",X"CD",X"6B",X"2A",X"21",X"07",X"80",X"3E",
		X"01",X"77",X"2C",X"2C",X"77",X"2C",X"2C",X"77",X"C3",X"8B",X"2A",X"06",X"0E",X"36",X"48",X"23",
		X"36",X"49",X"11",X"1F",X"00",X"19",X"36",X"4A",X"23",X"36",X"4B",X"19",X"10",X"EF",X"C9",X"40",
		X"43",X"43",X"44",X"45",X"47",X"47",X"41",X"46",X"43",X"43",X"42",X"3E",X"05",X"32",X"25",X"80",
		X"32",X"27",X"80",X"3E",X"04",X"32",X"2D",X"80",X"32",X"2F",X"80",X"3E",X"07",X"32",X"35",X"80",
		X"32",X"37",X"80",X"3E",X"06",X"32",X"21",X"80",X"32",X"23",X"80",X"32",X"39",X"80",X"32",X"3B",
		X"80",X"3E",X"05",X"06",X"0A",X"21",X"0D",X"80",X"77",X"23",X"23",X"10",X"FB",X"32",X"29",X"80",
		X"32",X"2B",X"80",X"32",X"31",X"80",X"32",X"33",X"80",X"3E",X"02",X"32",X"0D",X"80",X"32",X"0F",
		X"80",X"32",X"15",X"80",X"32",X"17",X"80",X"32",X"19",X"80",X"32",X"1B",X"80",X"C9",X"3A",X"FE",
		X"83",X"B7",X"28",X"34",X"CD",X"44",X"39",X"CD",X"A6",X"39",X"CD",X"73",X"38",X"CD",X"2F",X"37",
		X"CD",X"8F",X"39",X"3A",X"40",X"83",X"A7",X"C4",X"28",X"2B",X"CD",X"74",X"34",X"3A",X"B7",X"83",
		X"CB",X"47",X"CA",X"36",X"2B",X"3A",X"22",X"81",X"3C",X"32",X"22",X"81",X"A7",X"CC",X"83",X"34",
		X"3A",X"22",X"81",X"FE",X"70",X"CC",X"57",X"36",X"3A",X"47",X"80",X"FE",X"31",X"DA",X"88",X"2D",
		X"3A",X"FE",X"83",X"B7",X"C8",X"C3",X"54",X"2B",X"3D",X"32",X"40",X"83",X"FE",X"01",X"C0",X"CD",
		X"23",X"37",X"CD",X"67",X"38",X"C9",X"3A",X"22",X"81",X"3C",X"32",X"22",X"81",X"A7",X"CC",X"1F",
		X"35",X"3A",X"22",X"81",X"FE",X"50",X"CC",X"BB",X"35",X"3A",X"22",X"81",X"FE",X"B0",X"CC",X"57",
		X"36",X"C3",X"18",X"2B",X"3A",X"6C",X"82",X"A7",X"C0",X"3A",X"68",X"82",X"A7",X"28",X"08",X"3D",
		X"32",X"68",X"82",X"CD",X"74",X"34",X"C9",X"3A",X"04",X"80",X"A7",X"C0",X"21",X"44",X"80",X"11",
		X"47",X"80",X"3A",X"04",X"E0",X"CB",X"5F",X"28",X"07",X"3A",X"FD",X"83",X"3D",X"C2",X"FD",X"2B",
		X"3A",X"00",X"E0",X"4F",X"3A",X"48",X"82",X"A7",X"C2",X"43",X"2C",X"3A",X"04",X"E0",X"CB",X"5F",
		X"28",X"07",X"3A",X"FD",X"83",X"3D",X"C2",X"04",X"2C",X"3A",X"04",X"E0",X"CB",X"77",X"CA",X"14",
		X"2C",X"AF",X"32",X"4C",X"82",X"32",X"50",X"82",X"3A",X"49",X"82",X"A7",X"C2",X"96",X"2C",X"3A",
		X"4A",X"82",X"47",X"3A",X"4B",X"82",X"80",X"20",X"1D",X"3A",X"04",X"E0",X"CB",X"5F",X"28",X"07",
		X"3A",X"FD",X"83",X"3D",X"C2",X"0C",X"2C",X"3A",X"04",X"E0",X"CB",X"67",X"CA",X"6D",X"2C",X"AF",
		X"32",X"4D",X"82",X"32",X"51",X"82",X"3A",X"4A",X"82",X"A7",X"C2",X"FF",X"2C",X"CB",X"61",X"CA",
		X"CA",X"2C",X"AF",X"32",X"4E",X"82",X"32",X"52",X"82",X"3A",X"4B",X"82",X"A7",X"C2",X"5E",X"2D",
		X"CB",X"69",X"CA",X"29",X"2D",X"AF",X"32",X"4F",X"82",X"32",X"53",X"82",X"C9",X"3A",X"02",X"E0",
		X"4F",X"C3",X"84",X"2B",X"3A",X"04",X"E0",X"CB",X"47",X"C3",X"9E",X"2B",X"3A",X"00",X"E0",X"CB",
		X"47",X"C3",X"CC",X"2B",X"3A",X"47",X"80",X"FE",X"F0",X"D0",X"3A",X"50",X"82",X"A7",X"20",X"10",
		X"3E",X"04",X"DF",X"23",X"7E",X"2B",X"FE",X"DE",X"CA",X"3D",X"2C",X"3E",X"DE",X"32",X"45",X"80",
		X"3A",X"50",X"82",X"3C",X"32",X"50",X"82",X"B7",X"C8",X"AF",X"32",X"50",X"82",X"3A",X"56",X"82",
		X"32",X"50",X"82",X"3A",X"4C",X"82",X"A7",X"C0",X"3C",X"32",X"48",X"82",X"3A",X"50",X"82",X"3D",
		X"32",X"50",X"82",X"C2",X"61",X"2C",X"32",X"48",X"82",X"3C",X"32",X"4C",X"82",X"23",X"36",X"DE",
		X"C9",X"EB",X"3A",X"54",X"82",X"86",X"77",X"EB",X"23",X"3E",X"DC",X"77",X"C9",X"3A",X"51",X"82",
		X"A7",X"20",X"10",X"3E",X"04",X"DF",X"23",X"7E",X"2B",X"FE",X"1E",X"CA",X"90",X"2C",X"3E",X"1E",
		X"32",X"45",X"80",X"3A",X"51",X"82",X"3C",X"32",X"51",X"82",X"B7",X"C8",X"AF",X"32",X"51",X"82",
		X"3A",X"57",X"82",X"32",X"51",X"82",X"CD",X"74",X"34",X"3A",X"4D",X"82",X"A7",X"C0",X"3C",X"32",
		X"49",X"82",X"3A",X"51",X"82",X"3D",X"32",X"51",X"82",X"C2",X"BC",X"2C",X"32",X"49",X"82",X"3C",
		X"32",X"4D",X"82",X"23",X"36",X"1E",X"D5",X"CD",X"5F",X"30",X"D1",X"C9",X"EB",X"3A",X"54",X"82",
		X"47",X"7E",X"90",X"77",X"EB",X"23",X"3E",X"1C",X"77",X"C9",X"3A",X"47",X"80",X"FE",X"30",X"D8",
		X"3A",X"44",X"80",X"FE",X"E0",X"D0",X"3A",X"52",X"82",X"A7",X"20",X"10",X"3E",X"04",X"DF",X"23",
		X"7E",X"2B",X"FE",X"A1",X"CA",X"F9",X"2C",X"3E",X"A1",X"32",X"45",X"80",X"3A",X"52",X"82",X"3C",
		X"32",X"52",X"82",X"B7",X"C8",X"AF",X"32",X"52",X"82",X"3A",X"58",X"82",X"32",X"52",X"82",X"3A",
		X"4E",X"82",X"A7",X"C0",X"3C",X"32",X"4A",X"82",X"3A",X"52",X"82",X"3D",X"32",X"52",X"82",X"C2",
		X"1D",X"2D",X"32",X"4A",X"82",X"3C",X"32",X"4E",X"82",X"23",X"36",X"A1",X"C9",X"3A",X"55",X"82",
		X"47",X"7E",X"80",X"77",X"23",X"3E",X"9F",X"77",X"C9",X"3A",X"47",X"80",X"FE",X"30",X"D8",X"3A",
		X"44",X"80",X"FE",X"20",X"D8",X"3A",X"53",X"82",X"A7",X"20",X"10",X"3E",X"04",X"DF",X"23",X"7E",
		X"2B",X"FE",X"21",X"CA",X"58",X"2D",X"3E",X"21",X"32",X"45",X"80",X"3A",X"53",X"82",X"3C",X"32",
		X"53",X"82",X"B7",X"C8",X"AF",X"32",X"53",X"82",X"3A",X"59",X"82",X"32",X"53",X"82",X"3A",X"4F",
		X"82",X"A7",X"C0",X"3C",X"32",X"4B",X"82",X"3A",X"53",X"82",X"3D",X"32",X"53",X"82",X"C2",X"7C",
		X"2D",X"32",X"4B",X"82",X"3C",X"32",X"4F",X"82",X"23",X"36",X"21",X"C9",X"3A",X"55",X"82",X"47",
		X"7E",X"90",X"77",X"23",X"3E",X"1F",X"77",X"C9",X"3A",X"44",X"80",X"FE",X"15",X"DA",X"00",X"2E",
		X"FE",X"1C",X"CA",X"10",X"2E",X"DA",X"10",X"2E",X"FE",X"2E",X"DA",X"00",X"2E",X"FE",X"35",X"CA",
		X"00",X"2E",X"DA",X"00",X"2E",X"FE",X"45",X"DA",X"00",X"2E",X"FE",X"4C",X"CA",X"61",X"2E",X"DA",
		X"61",X"2E",X"FE",X"5E",X"DA",X"00",X"2E",X"FE",X"65",X"CA",X"00",X"2E",X"DA",X"00",X"2E",X"FE",
		X"75",X"DA",X"00",X"2E",X"FE",X"7C",X"CA",X"B2",X"2E",X"DA",X"B2",X"2E",X"FE",X"8E",X"DA",X"00",
		X"2E",X"FE",X"95",X"CA",X"00",X"2E",X"DA",X"00",X"2E",X"FE",X"A5",X"DA",X"00",X"2E",X"FE",X"AC",
		X"CA",X"03",X"2F",X"DA",X"03",X"2F",X"FE",X"BE",X"DA",X"00",X"2E",X"FE",X"C5",X"CA",X"00",X"2E",
		X"DA",X"00",X"2E",X"FE",X"D5",X"DA",X"00",X"2E",X"FE",X"DC",X"CA",X"54",X"2F",X"DA",X"54",X"2F",
		X"3A",X"47",X"80",X"FE",X"2A",X"D2",X"54",X"2B",X"3E",X"01",X"32",X"04",X"80",X"C3",X"54",X"2B",
		X"3A",X"FD",X"83",X"3D",X"20",X"3C",X"3A",X"5E",X"82",X"A7",X"C0",X"3A",X"47",X"80",X"FE",X"2A",
		X"D2",X"54",X"2B",X"06",X"18",X"3A",X"21",X"81",X"D6",X"01",X"CC",X"FC",X"36",X"21",X"64",X"AB",
		X"CD",X"A5",X"2F",X"3A",X"34",X"81",X"A7",X"28",X"09",X"06",X"18",X"CD",X"54",X"38",X"AF",X"32",
		X"34",X"81",X"3A",X"FD",X"83",X"3D",X"20",X"0F",X"3E",X"01",X"32",X"5E",X"82",X"21",X"5C",X"82",
		X"34",X"C9",X"3A",X"63",X"82",X"18",X"C2",X"3E",X"01",X"32",X"63",X"82",X"21",X"5D",X"82",X"34",
		X"C9",X"3A",X"FD",X"83",X"3D",X"20",X"3C",X"3A",X"5F",X"82",X"A7",X"C0",X"3A",X"47",X"80",X"FE",
		X"2A",X"D2",X"54",X"2B",X"06",X"48",X"3A",X"21",X"81",X"D6",X"02",X"CC",X"FC",X"36",X"21",X"A4",
		X"AA",X"CD",X"A5",X"2F",X"3A",X"34",X"81",X"A7",X"28",X"09",X"06",X"48",X"CD",X"54",X"38",X"AF",
		X"32",X"34",X"81",X"3A",X"FD",X"83",X"3D",X"20",X"0F",X"3E",X"01",X"32",X"5F",X"82",X"21",X"5C",
		X"82",X"34",X"C9",X"3A",X"64",X"82",X"18",X"C2",X"3E",X"01",X"32",X"64",X"82",X"21",X"5D",X"82",
		X"34",X"C9",X"3A",X"FD",X"83",X"3D",X"20",X"3C",X"3A",X"60",X"82",X"A7",X"C0",X"3A",X"47",X"80",
		X"FE",X"2A",X"D2",X"54",X"2B",X"06",X"78",X"3A",X"21",X"81",X"D6",X"03",X"CC",X"FC",X"36",X"21",
		X"E4",X"A9",X"CD",X"A5",X"2F",X"3A",X"34",X"81",X"A7",X"28",X"09",X"06",X"78",X"CD",X"54",X"38",
		X"AF",X"32",X"34",X"81",X"3A",X"FD",X"83",X"3D",X"20",X"0F",X"3E",X"01",X"32",X"60",X"82",X"21",
		X"5C",X"82",X"34",X"C9",X"3A",X"65",X"82",X"18",X"C2",X"3E",X"01",X"32",X"65",X"82",X"21",X"5D",
		X"82",X"34",X"C9",X"3A",X"FD",X"83",X"3D",X"20",X"3C",X"3A",X"61",X"82",X"A7",X"C0",X"3A",X"47",
		X"80",X"FE",X"2A",X"D2",X"54",X"2B",X"06",X"A8",X"3A",X"21",X"81",X"D6",X"04",X"CC",X"FC",X"36",
		X"21",X"24",X"A9",X"CD",X"A5",X"2F",X"3A",X"34",X"81",X"A7",X"28",X"09",X"06",X"A8",X"CD",X"54",
		X"38",X"AF",X"32",X"34",X"81",X"3A",X"FD",X"83",X"3D",X"20",X"0F",X"3E",X"01",X"32",X"61",X"82",
		X"21",X"5C",X"82",X"34",X"C9",X"3A",X"66",X"82",X"18",X"C2",X"3E",X"01",X"32",X"66",X"82",X"21",
		X"5D",X"82",X"34",X"C9",X"3A",X"FD",X"83",X"3D",X"20",X"3C",X"3A",X"62",X"82",X"A7",X"C0",X"3A",
		X"47",X"80",X"FE",X"2A",X"D2",X"54",X"2B",X"06",X"D8",X"3A",X"21",X"81",X"D6",X"05",X"CC",X"FC",
		X"36",X"21",X"64",X"A8",X"CD",X"A5",X"2F",X"3A",X"34",X"81",X"A7",X"28",X"09",X"06",X"D8",X"CD",
		X"54",X"38",X"AF",X"32",X"34",X"81",X"3A",X"FD",X"83",X"3D",X"20",X"0F",X"3E",X"01",X"32",X"62",
		X"82",X"21",X"5C",X"82",X"34",X"C9",X"3A",X"67",X"82",X"18",X"C2",X"3E",X"01",X"32",X"67",X"82",
		X"21",X"5D",X"82",X"34",X"C9",X"3A",X"34",X"81",X"A7",X"28",X"09",X"11",X"20",X"00",X"CD",X"03",
		X"09",X"CD",X"45",X"38",X"36",X"6C",X"23",X"36",X"6D",X"01",X"1F",X"00",X"09",X"36",X"6E",X"23",
		X"36",X"6F",X"E5",X"D5",X"11",X"05",X"00",X"CD",X"03",X"09",X"CD",X"E8",X"08",X"3A",X"FE",X"83",
		X"B7",X"28",X"4A",X"AF",X"67",X"6F",X"22",X"82",X"83",X"DF",X"3E",X"F0",X"DF",X"3A",X"FD",X"83",
		X"21",X"5C",X"82",X"3D",X"28",X"01",X"2C",X"7E",X"FE",X"04",X"28",X"1E",X"3E",X"08",X"DF",X"3E",
		X"0E",X"DF",X"21",X"81",X"83",X"35",X"20",X"02",X"36",X"14",X"7E",X"21",X"5D",X"0F",X"87",X"85",
		X"6F",X"7E",X"2C",X"66",X"6F",X"22",X"82",X"83",X"18",X"13",X"32",X"2F",X"84",X"CD",X"F9",X"07",
		X"21",X"40",X"B0",X"01",X"00",X"18",X"71",X"2C",X"10",X"FC",X"CD",X"45",X"38",X"3E",X"20",X"32",
		X"6A",X"82",X"3E",X"80",X"DF",X"21",X"44",X"80",X"AF",X"77",X"23",X"77",X"23",X"77",X"23",X"36",
		X"F0",X"D1",X"E1",X"AF",X"32",X"9B",X"82",X"32",X"EA",X"83",X"32",X"4D",X"82",X"32",X"49",X"82",
		X"32",X"51",X"82",X"3C",X"32",X"6C",X"82",X"32",X"CD",X"83",X"3E",X"10",X"32",X"68",X"82",X"C9",
		X"3A",X"6C",X"82",X"A7",X"C8",X"21",X"6A",X"82",X"35",X"C0",X"AF",X"32",X"6C",X"82",X"C9",X"3A",
		X"47",X"80",X"FE",X"30",X"D8",X"FE",X"D0",X"4F",X"28",X"17",X"D0",X"3A",X"69",X"82",X"B9",X"D8",
		X"C8",X"79",X"32",X"69",X"82",X"11",X"01",X"00",X"FE",X"80",X"C8",X"E5",X"CD",X"03",X"09",X"E1",
		X"C9",X"3A",X"69",X"82",X"A7",X"20",X"E4",X"3E",X"E0",X"32",X"69",X"82",X"18",X"DD",X"DD",X"21",
		X"73",X"82",X"DD",X"7E",X"02",X"32",X"1A",X"81",X"3A",X"10",X"81",X"3C",X"32",X"10",X"81",X"FE",
		X"50",X"D4",X"84",X"31",X"DD",X"21",X"7C",X"82",X"DD",X"7E",X"02",X"32",X"19",X"81",X"3A",X"11",
		X"81",X"3C",X"3C",X"32",X"11",X"81",X"FE",X"A0",X"DC",X"25",X"32",X"3A",X"6E",X"82",X"3C",X"32",
		X"6E",X"82",X"FE",X"10",X"CA",X"D2",X"30",X"FE",X"20",X"CA",X"F8",X"30",X"FE",X"30",X"CA",X"1E",
		X"31",X"C9",X"21",X"73",X"82",X"7E",X"23",X"46",X"21",X"1A",X"81",X"4E",X"11",X"AC",X"24",X"32",
		X"B1",X"81",X"CD",X"55",X"31",X"21",X"7C",X"82",X"7E",X"23",X"46",X"21",X"19",X"81",X"4E",X"11",
		X"E8",X"24",X"32",X"B1",X"81",X"C3",X"48",X"31",X"21",X"73",X"82",X"7E",X"23",X"46",X"21",X"1A",
		X"81",X"4E",X"11",X"B4",X"24",X"32",X"B1",X"81",X"CD",X"55",X"31",X"21",X"7C",X"82",X"7E",X"23",
		X"46",X"21",X"19",X"81",X"4E",X"11",X"FC",X"24",X"32",X"B1",X"81",X"C3",X"48",X"31",X"21",X"73",
		X"82",X"7E",X"23",X"46",X"21",X"1A",X"81",X"4E",X"11",X"BC",X"24",X"32",X"B1",X"81",X"AF",X"32",
		X"6E",X"82",X"CD",X"55",X"31",X"21",X"7C",X"82",X"7E",X"23",X"46",X"21",X"19",X"81",X"4E",X"11",
		X"10",X"25",X"32",X"B1",X"81",X"C3",X"48",X"31",X"2A",X"7E",X"24",X"ED",X"53",X"01",X"80",X"78",
		X"32",X"03",X"80",X"18",X"0B",X"2A",X"78",X"24",X"ED",X"53",X"01",X"80",X"78",X"32",X"03",X"80",
		X"1A",X"77",X"23",X"13",X"1A",X"77",X"2B",X"D5",X"11",X"20",X"00",X"19",X"D1",X"13",X"10",X"F0",
		X"3A",X"B1",X"81",X"5F",X"16",X"00",X"19",X"3A",X"03",X"80",X"47",X"ED",X"5B",X"01",X"80",X"0D",
		X"C2",X"60",X"31",X"C9",X"DD",X"21",X"73",X"82",X"AF",X"67",X"DD",X"46",X"01",X"C6",X"20",X"10",
		X"FC",X"4F",X"DD",X"6E",X"00",X"09",X"5D",X"54",X"AF",X"6F",X"67",X"DD",X"46",X"02",X"05",X"19",
		X"10",X"FD",X"11",X"08",X"A8",X"19",X"0E",X"02",X"3A",X"10",X"81",X"FE",X"50",X"CA",X"C7",X"31",
		X"FE",X"80",X"CA",X"D5",X"31",X"FE",X"A0",X"CA",X"EE",X"31",X"FE",X"B0",X"CA",X"D5",X"31",X"FE",
		X"D0",X"CA",X"C7",X"31",X"C3",X"11",X"32",X"06",X"02",X"11",X"19",X"32",X"CD",X"01",X"32",X"0D",
		X"20",X"F5",X"C3",X"11",X"32",X"06",X"02",X"11",X"1D",X"32",X"CD",X"01",X"32",X"0D",X"20",X"F5",
		X"3A",X"07",X"81",X"A7",X"CA",X"11",X"32",X"AF",X"32",X"07",X"81",X"C3",X"11",X"32",X"06",X"02",
		X"11",X"21",X"32",X"CD",X"01",X"32",X"0D",X"20",X"F5",X"3E",X"01",X"32",X"07",X"81",X"C3",X"11",
		X"32",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"D5",X"11",X"1F",X"00",X"19",X"D1",X"10",X"F1",
		X"C9",X"DD",X"7E",X"02",X"3D",X"32",X"1A",X"81",X"C9",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",
		X"9B",X"10",X"10",X"10",X"10",X"DD",X"21",X"7C",X"82",X"AF",X"67",X"DD",X"46",X"01",X"C6",X"20",
		X"10",X"FC",X"4F",X"DD",X"6E",X"00",X"09",X"5D",X"54",X"AF",X"6F",X"67",X"DD",X"46",X"02",X"05",
		X"19",X"10",X"FD",X"11",X"0E",X"A8",X"19",X"0E",X"03",X"3A",X"11",X"81",X"FE",X"00",X"CA",X"68",
		X"32",X"FE",X"30",X"CA",X"76",X"32",X"FE",X"50",X"CA",X"8F",X"32",X"FE",X"60",X"CA",X"76",X"32",
		X"FE",X"70",X"CA",X"68",X"32",X"C3",X"B2",X"32",X"06",X"02",X"11",X"BA",X"32",X"CD",X"A2",X"32",
		X"0D",X"20",X"F5",X"C3",X"B2",X"32",X"06",X"02",X"11",X"BE",X"32",X"CD",X"A2",X"32",X"0D",X"20",
		X"F5",X"3A",X"08",X"81",X"A7",X"CA",X"B2",X"32",X"AF",X"32",X"08",X"81",X"C3",X"B2",X"32",X"06",
		X"02",X"11",X"C2",X"32",X"CD",X"A2",X"32",X"0D",X"20",X"F5",X"3E",X"01",X"32",X"08",X"81",X"C3",
		X"B2",X"32",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"D5",X"11",X"1F",X"00",X"19",X"D1",X"10",
		X"F1",X"C9",X"DD",X"7E",X"02",X"3D",X"32",X"19",X"81",X"C9",X"94",X"95",X"96",X"97",X"98",X"99",
		X"9A",X"9B",X"10",X"10",X"10",X"10",X"D9",X"21",X"93",X"82",X"3A",X"FD",X"83",X"3D",X"28",X"01",
		X"2C",X"7E",X"01",X"E9",X"32",X"26",X"00",X"6F",X"85",X"6F",X"09",X"5E",X"23",X"56",X"EB",X"11",
		X"70",X"82",X"01",X"21",X"00",X"ED",X"B0",X"D9",X"C9",X"F3",X"32",X"14",X"33",X"35",X"33",X"56",
		X"33",X"77",X"33",X"60",X"08",X"03",X"60",X"04",X"04",X"80",X"0C",X"02",X"80",X"06",X"03",X"40",
		X"06",X"04",X"80",X"02",X"04",X"E0",X"04",X"02",X"60",X"02",X"01",X"C0",X"02",X"03",X"C0",X"02",
		X"03",X"E0",X"02",X"03",X"60",X"08",X"03",X"40",X"04",X"05",X"80",X"0C",X"01",X"60",X"06",X"03",
		X"C0",X"06",X"03",X"80",X"02",X"04",X"E0",X"04",X"03",X"60",X"02",X"02",X"E0",X"02",X"04",X"C0",
		X"02",X"04",X"E0",X"02",X"04",X"60",X"08",X"02",X"80",X"04",X"04",X"80",X"0C",X"01",X"C0",X"06",
		X"03",X"60",X"06",X"03",X"80",X"02",X"04",X"A0",X"04",X"03",X"E0",X"02",X"02",X"A0",X"02",X"05",
		X"E0",X"02",X"04",X"C0",X"02",X"04",X"60",X"08",X"02",X"A0",X"04",X"03",X"80",X"0C",X"01",X"E0",
		X"06",X"02",X"80",X"06",X"03",X"80",X"02",X"04",X"80",X"04",X"04",X"C0",X"02",X"03",X"E0",X"02",
		X"04",X"A0",X"02",X"04",X"E0",X"02",X"04",X"60",X"08",X"01",X"E0",X"04",X"03",X"80",X"0C",X"01",
		X"A0",X"06",X"02",X"E0",X"06",X"02",X"80",X"02",X"04",X"60",X"04",X"03",X"A0",X"02",X"04",X"80",
		X"02",X"05",X"C0",X"02",X"04",X"A0",X"02",X"05",X"3A",X"D6",X"83",X"3D",X"C0",X"3A",X"9B",X"82",
		X"A7",X"C0",X"32",X"B4",X"83",X"CD",X"DD",X"0A",X"CD",X"3C",X"06",X"CD",X"C6",X"32",X"AF",X"32",
		X"5B",X"82",X"CD",X"DB",X"29",X"21",X"50",X"A8",X"CD",X"6B",X"2A",X"CD",X"CD",X"09",X"CD",X"23",
		X"20",X"3E",X"01",X"32",X"5B",X"82",X"32",X"9B",X"82",X"C9",X"3A",X"D6",X"83",X"3D",X"C0",X"3A",
		X"9B",X"82",X"A7",X"C8",X"CD",X"F6",X"33",X"CD",X"DE",X"2A",X"CD",X"40",X"34",X"CD",X"65",X"09",
		X"CD",X"93",X"08",X"CD",X"8E",X"30",X"CD",X"8B",X"28",X"CD",X"48",X"22",X"CD",X"81",X"27",X"CD",
		X"50",X"30",X"CD",X"40",X"25",X"C9",X"3A",X"6C",X"82",X"B7",X"C0",X"3A",X"04",X"80",X"A7",X"C0",
		X"3A",X"99",X"82",X"A7",X"C2",X"6F",X"34",X"11",X"47",X"80",X"3E",X"30",X"32",X"99",X"82",X"21",
		X"9A",X"82",X"34",X"4E",X"06",X"00",X"21",X"3E",X"0F",X"09",X"4E",X"0C",X"CA",X"35",X"34",X"21",
		X"25",X"34",X"09",X"E5",X"21",X"44",X"80",X"C9",X"C3",X"29",X"2D",X"C3",X"CA",X"2C",X"C3",X"6D",
		X"2C",X"C3",X"14",X"2C",X"C9",X"AF",X"32",X"9A",X"82",X"32",X"99",X"82",X"32",X"5B",X"82",X"C9",
		X"21",X"44",X"80",X"11",X"47",X"80",X"3A",X"48",X"82",X"A7",X"C2",X"43",X"2C",X"32",X"4C",X"82",
		X"3A",X"49",X"82",X"A7",X"C2",X"96",X"2C",X"32",X"4D",X"82",X"3A",X"4A",X"82",X"A7",X"C2",X"FF",
		X"2C",X"32",X"4E",X"82",X"3A",X"4B",X"82",X"A7",X"C2",X"5E",X"2D",X"32",X"4F",X"82",X"C9",X"3D",
		X"32",X"99",X"82",X"C9",X"3A",X"23",X"81",X"3C",X"32",X"23",X"81",X"FE",X"06",X"D8",X"AF",X"32",
		X"23",X"81",X"C9",X"3A",X"FD",X"83",X"4F",X"3A",X"23",X"81",X"32",X"21",X"81",X"FE",X"01",X"CA",
		X"A7",X"34",X"FE",X"02",X"CA",X"BC",X"34",X"FE",X"03",X"CA",X"D1",X"34",X"FE",X"04",X"CA",X"E6",
		X"34",X"FE",X"05",X"CA",X"FB",X"34",X"C9",X"0D",X"20",X"0B",X"3A",X"5E",X"82",X"A7",X"C0",X"21",
		X"64",X"AB",X"C3",X"10",X"35",X"3A",X"63",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",
		X"5F",X"82",X"A7",X"C0",X"21",X"A4",X"AA",X"C3",X"10",X"35",X"3A",X"64",X"82",X"A7",X"C0",X"18",
		X"F3",X"0D",X"20",X"0B",X"3A",X"60",X"82",X"A7",X"C0",X"21",X"E4",X"A9",X"C3",X"10",X"35",X"3A",
		X"65",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"61",X"82",X"A7",X"C0",X"21",X"24",
		X"A9",X"C3",X"10",X"35",X"3A",X"66",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"62",
		X"82",X"A7",X"C0",X"21",X"64",X"A8",X"C3",X"10",X"35",X"3A",X"67",X"82",X"A7",X"C0",X"18",X"F3",
		X"36",X"2C",X"23",X"36",X"2D",X"01",X"1F",X"00",X"09",X"36",X"2E",X"23",X"36",X"2F",X"C9",X"3A",
		X"FD",X"83",X"4F",X"3A",X"23",X"81",X"32",X"20",X"81",X"FE",X"01",X"CA",X"43",X"35",X"FE",X"02",
		X"CA",X"58",X"35",X"FE",X"03",X"CA",X"6D",X"35",X"FE",X"04",X"CA",X"82",X"35",X"FE",X"05",X"CA",
		X"97",X"35",X"C9",X"0D",X"20",X"0B",X"3A",X"5E",X"82",X"A7",X"C0",X"21",X"64",X"AB",X"C3",X"AC",
		X"35",X"3A",X"63",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"5F",X"82",X"A7",X"C0",
		X"21",X"A4",X"AA",X"C3",X"AC",X"35",X"3A",X"64",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",
		X"3A",X"60",X"82",X"A7",X"C0",X"21",X"E4",X"A9",X"C3",X"AC",X"35",X"3A",X"65",X"82",X"A7",X"C0",
		X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"61",X"82",X"A7",X"C0",X"21",X"24",X"A9",X"C3",X"AC",X"35",
		X"3A",X"66",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"62",X"82",X"A7",X"C0",X"21",
		X"64",X"A8",X"C3",X"AC",X"35",X"3A",X"67",X"82",X"A7",X"C0",X"18",X"F3",X"36",X"10",X"23",X"36",
		X"10",X"01",X"1F",X"00",X"09",X"36",X"D0",X"23",X"36",X"D1",X"C9",X"3A",X"FD",X"83",X"4F",X"3A",
		X"20",X"81",X"32",X"21",X"81",X"FE",X"01",X"CA",X"DF",X"35",X"FE",X"02",X"CA",X"F4",X"35",X"FE",
		X"03",X"CA",X"09",X"36",X"FE",X"04",X"CA",X"1E",X"36",X"FE",X"05",X"CA",X"33",X"36",X"C9",X"0D",
		X"20",X"0B",X"3A",X"5E",X"82",X"A7",X"C0",X"21",X"64",X"AB",X"C3",X"48",X"36",X"3A",X"63",X"82",
		X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"5F",X"82",X"A7",X"C0",X"21",X"A4",X"AA",X"C3",
		X"48",X"36",X"3A",X"64",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"60",X"82",X"A7",
		X"C0",X"21",X"E4",X"A9",X"C3",X"48",X"36",X"3A",X"65",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",
		X"0B",X"3A",X"61",X"82",X"A7",X"C0",X"21",X"24",X"A9",X"C3",X"48",X"36",X"3A",X"66",X"82",X"A7",
		X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"62",X"82",X"A7",X"C0",X"21",X"64",X"A8",X"C3",X"48",
		X"36",X"3A",X"67",X"82",X"A7",X"C0",X"18",X"F3",X"36",X"D0",X"23",X"36",X"D1",X"01",X"1F",X"00",
		X"09",X"36",X"D2",X"23",X"36",X"D3",X"C9",X"3A",X"FD",X"83",X"4F",X"3A",X"21",X"81",X"FE",X"01",
		X"CA",X"78",X"36",X"FE",X"02",X"CA",X"8D",X"36",X"FE",X"03",X"CA",X"A2",X"36",X"FE",X"04",X"CA",
		X"B7",X"36",X"FE",X"05",X"CA",X"CC",X"36",X"C9",X"0D",X"20",X"0B",X"3A",X"5E",X"82",X"A7",X"C0",
		X"21",X"64",X"AB",X"C3",X"E1",X"36",X"3A",X"63",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",
		X"3A",X"5F",X"82",X"A7",X"C0",X"21",X"A4",X"AA",X"C3",X"E1",X"36",X"3A",X"64",X"82",X"A7",X"C0",
		X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"60",X"82",X"A7",X"C0",X"21",X"E4",X"A9",X"C3",X"E1",X"36",
		X"3A",X"65",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",X"61",X"82",X"A7",X"C0",X"21",
		X"24",X"A9",X"C3",X"E1",X"36",X"3A",X"66",X"82",X"A7",X"C0",X"18",X"F3",X"0D",X"20",X"0B",X"3A",
		X"62",X"82",X"A7",X"C0",X"21",X"64",X"A8",X"C3",X"E1",X"36",X"3A",X"67",X"82",X"A7",X"C0",X"18",
		X"F3",X"36",X"10",X"23",X"36",X"10",X"01",X"1F",X"00",X"09",X"36",X"10",X"23",X"36",X"10",X"3A",
		X"04",X"80",X"A7",X"C0",X"AF",X"32",X"21",X"81",X"32",X"20",X"81",X"C9",X"3A",X"20",X"81",X"A7",
		X"C2",X"1C",X"37",X"21",X"5C",X"80",X"70",X"23",X"36",X"19",X"23",X"36",X"03",X"23",X"36",X"20",
		X"3E",X"A0",X"32",X"40",X"83",X"11",X"20",X"00",X"CD",X"03",X"09",X"C9",X"3E",X"01",X"32",X"04",
		X"80",X"E1",X"C9",X"21",X"5C",X"80",X"AF",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"C9",X"3A",
		X"34",X"81",X"A7",X"C2",X"79",X"37",X"DD",X"21",X"1B",X"81",X"DD",X"7E",X"01",X"A7",X"CC",X"96",
		X"37",X"3A",X"3D",X"81",X"CB",X"47",X"C2",X"3C",X"38",X"3A",X"35",X"81",X"A7",X"20",X"01",X"C9",
		X"3A",X"34",X"81",X"A7",X"20",X"23",X"CD",X"B8",X"37",X"3A",X"47",X"80",X"FE",X"5A",X"D8",X"FE",
		X"68",X"D0",X"3A",X"40",X"80",X"47",X"3A",X"44",X"80",X"C6",X"04",X"B8",X"D8",X"D6",X"08",X"B8",
		X"D0",X"3E",X"01",X"32",X"34",X"81",X"3E",X"18",X"DF",X"DD",X"21",X"44",X"80",X"FD",X"21",X"40",
		X"80",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"DD",X"7E",X"03",
		X"C6",X"02",X"FD",X"77",X"03",X"C9",X"3A",X"35",X"81",X"A7",X"C0",X"21",X"3D",X"81",X"34",X"21",
		X"41",X"80",X"36",X"1E",X"23",X"36",X"04",X"23",X"36",X"60",X"3E",X"01",X"32",X"35",X"81",X"32",
		X"3D",X"83",X"3E",X"3C",X"32",X"3E",X"83",X"C9",X"21",X"3E",X"83",X"7E",X"A7",X"28",X"2B",X"35",
		X"3E",X"3C",X"CB",X"3F",X"BE",X"20",X"0F",X"2B",X"7E",X"A7",X"3E",X"21",X"32",X"41",X"80",X"F0",
		X"3E",X"A1",X"32",X"41",X"80",X"C9",X"2B",X"7E",X"E6",X"7F",X"21",X"28",X"38",X"3C",X"CD",X"23",
		X"38",X"7E",X"21",X"1C",X"81",X"86",X"32",X"40",X"80",X"C9",X"2B",X"7E",X"A7",X"F2",X"F2",X"37",
		X"35",X"35",X"34",X"7E",X"E6",X"7F",X"21",X"28",X"38",X"CD",X"23",X"38",X"7E",X"FE",X"01",X"38",
		X"0A",X"28",X"1A",X"21",X"1C",X"81",X"86",X"32",X"40",X"80",X"C9",X"21",X"3D",X"83",X"7E",X"EE",
		X"80",X"77",X"3E",X"3C",X"32",X"3E",X"83",X"3E",X"1E",X"32",X"41",X"80",X"C9",X"3E",X"3C",X"32",
		X"3E",X"83",X"C9",X"85",X"6F",X"D0",X"24",X"C9",X"00",X"EE",X"EC",X"EA",X"E8",X"E6",X"E4",X"E2",
		X"E0",X"01",X"DE",X"DC",X"DA",X"D8",X"D6",X"D4",X"D2",X"D0",X"00",X"D0",X"3A",X"35",X"81",X"A7",
		X"C8",X"AF",X"32",X"34",X"81",X"21",X"40",X"80",X"AF",X"77",X"23",X"77",X"23",X"77",X"23",X"77",
		X"32",X"35",X"81",X"C9",X"21",X"40",X"80",X"70",X"23",X"36",X"19",X"23",X"36",X"03",X"23",X"36",
		X"10",X"3E",X"A0",X"32",X"40",X"83",X"C9",X"21",X"40",X"80",X"AF",X"77",X"23",X"77",X"23",X"77",
		X"23",X"77",X"C9",X"3A",X"B7",X"83",X"FE",X"02",X"DA",X"FC",X"38",X"FE",X"05",X"D2",X"FD",X"38",
		X"3A",X"01",X"81",X"A7",X"CC",X"15",X"39",X"3A",X"4F",X"81",X"A7",X"C8",X"21",X"46",X"81",X"7E",
		X"23",X"BE",X"C2",X"39",X"39",X"35",X"11",X"06",X"A8",X"3A",X"50",X"81",X"CB",X"47",X"CA",X"F6",
		X"38",X"21",X"9C",X"24",X"AF",X"47",X"3A",X"4E",X"81",X"4F",X"3C",X"3C",X"32",X"4E",X"81",X"09",
		X"06",X"00",X"EB",X"3A",X"45",X"81",X"4F",X"09",X"EB",X"0E",X"20",X"3A",X"45",X"81",X"81",X"32",
		X"45",X"81",X"7E",X"12",X"23",X"13",X"7E",X"12",X"3A",X"4E",X"81",X"FE",X"10",X"D8",X"AF",X"32",
		X"4F",X"81",X"32",X"4E",X"81",X"32",X"45",X"81",X"32",X"46",X"81",X"32",X"47",X"81",X"C9",X"3A",
		X"FE",X"83",X"FE",X"02",X"C0",X"AF",X"32",X"4F",X"81",X"32",X"4E",X"81",X"32",X"45",X"81",X"32",
		X"46",X"81",X"32",X"47",X"81",X"C9",X"21",X"8C",X"24",X"C3",X"A4",X"38",X"C9",X"3A",X"01",X"81",
		X"A7",X"CC",X"07",X"39",X"C3",X"87",X"38",X"3A",X"4F",X"81",X"A7",X"C0",X"3E",X"01",X"32",X"50",
		X"81",X"CD",X"25",X"39",X"C9",X"3A",X"4F",X"81",X"A7",X"C0",X"3A",X"50",X"81",X"3C",X"32",X"50",
		X"81",X"CD",X"25",X"39",X"C9",X"3A",X"9B",X"81",X"E6",X"0F",X"87",X"87",X"87",X"21",X"46",X"81",
		X"77",X"23",X"77",X"3E",X"01",X"32",X"4F",X"81",X"C9",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"3A",
		X"46",X"81",X"77",X"C9",X"3A",X"50",X"81",X"CB",X"47",X"C8",X"3A",X"B7",X"83",X"FE",X"02",X"D8",
		X"3A",X"47",X"80",X"C6",X"08",X"FE",X"2A",X"D8",X"FE",X"3B",X"D0",X"3A",X"44",X"80",X"C6",X"08",
		X"47",X"3A",X"01",X"81",X"4F",X"C6",X"08",X"B8",X"D8",X"79",X"D6",X"20",X"B8",X"D0",X"79",X"D6",
		X"08",X"B8",X"30",X"04",X"CD",X"59",X"23",X"C9",X"3E",X"01",X"32",X"04",X"80",X"21",X"46",X"A8",
		X"36",X"68",X"23",X"36",X"69",X"01",X"1F",X"00",X"09",X"36",X"6A",X"23",X"36",X"6B",X"C9",X"3A",
		X"FE",X"83",X"A7",X"C8",X"3A",X"A2",X"81",X"FE",X"0F",X"D0",X"FE",X"02",X"D8",X"3A",X"40",X"81",
		X"A7",X"C0",X"3E",X"D0",X"DF",X"C9",X"3A",X"01",X"81",X"A7",X"20",X"05",X"AF",X"32",X"3F",X"83",
		X"C9",X"3A",X"50",X"81",X"CB",X"47",X"C8",X"3A",X"4F",X"81",X"A7",X"C0",X"21",X"3F",X"83",X"34",
		X"7E",X"FE",X"40",X"28",X"05",X"FE",X"70",X"28",X"13",X"C9",X"21",X"46",X"A8",X"36",X"68",X"23",
		X"36",X"69",X"01",X"1F",X"00",X"09",X"36",X"6A",X"23",X"36",X"6B",X"C9",X"21",X"46",X"A8",X"36",
		X"D0",X"23",X"36",X"D1",X"01",X"1F",X"00",X"09",X"36",X"D2",X"23",X"36",X"D3",X"AF",X"32",X"3F",
		X"83",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"E2",X"83",X"7E",X"B7",X"3A",X"00",X"E0",X"2F",X"20",X"04",X"E6",X"C4",X"77",X"C9",X"E6",
		X"C4",X"C0",X"3C",X"CD",X"A7",X"07",X"AF",X"32",X"86",X"83",X"ED",X"5B",X"D4",X"83",X"CB",X"76",
		X"C2",X"3E",X"3E",X"CB",X"56",X"77",X"20",X"09",X"3C",X"32",X"18",X"B8",X"3E",X"04",X"32",X"7E",
		X"83",X"21",X"36",X"3E",X"19",X"E9",X"18",X"24",X"18",X"1B",X"18",X"19",X"18",X"1E",X"77",X"3C",
		X"32",X"1C",X"B8",X"3E",X"04",X"32",X"7F",X"83",X"21",X"4D",X"3E",X"19",X"E9",X"18",X"0D",X"18",
		X"04",X"18",X"11",X"18",X"13",X"21",X"E3",X"83",X"34",X"CB",X"46",X"C0",X"0E",X"01",X"18",X"0A",
		X"0E",X"02",X"18",X"06",X"0E",X"03",X"18",X"02",X"0E",X"06",X"3A",X"E1",X"83",X"81",X"27",X"30",
		X"02",X"3E",X"99",X"32",X"E1",X"83",X"3A",X"FE",X"83",X"B7",X"C0",X"3A",X"D6",X"83",X"FE",X"05",
		X"CC",X"13",X"0D",X"3E",X"05",X"32",X"D6",X"83",X"AF",X"32",X"D8",X"83",X"21",X"40",X"80",X"11",
		X"41",X"80",X"01",X"1F",X"00",X"70",X"ED",X"B0",X"C3",X"8A",X"0B",X"21",X"D8",X"83",X"36",X"FF",
		X"CD",X"79",X"07",X"AF",X"32",X"9B",X"82",X"32",X"21",X"80",X"3E",X"05",X"32",X"1B",X"80",X"3E",
		X"03",X"32",X"2B",X"80",X"11",X"F2",X"0F",X"21",X"8D",X"AA",X"06",X"0B",X"EF",X"3A",X"E4",X"83",
		X"FE",X"0A",X"D0",X"21",X"15",X"AB",X"CD",X"CC",X"0B",X"11",X"3F",X"10",X"06",X"07",X"EF",X"11",
		X"09",X"10",X"06",X"04",X"EF",X"11",X"28",X"10",X"06",X"07",X"EF",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
