library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tcs_rom4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tcs_rom4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"58",X"49",X"58",X"49",X"58",X"49",X"FD",X"60",X"00",X"DC",X"08",X"83",X"00",X"01",X"DD",X"08",
		X"10",X"26",X"FE",X"36",X"10",X"9E",X"12",X"EC",X"A9",X"00",X"0F",X"10",X"26",X"00",X"5E",X"0F",
		X"03",X"0F",X"04",X"10",X"BE",X"E1",X"00",X"10",X"9F",X"12",X"10",X"9F",X"14",X"0F",X"01",X"0F",
		X"02",X"EC",X"A1",X"DD",X"08",X"DD",X"0A",X"A6",X"A0",X"97",X"1C",X"97",X"3C",X"EC",X"A1",X"DD",
		X"1F",X"DD",X"3F",X"A6",X"A0",X"97",X"24",X"97",X"44",X"EC",X"A1",X"DD",X"27",X"DD",X"47",X"A6",
		X"A0",X"97",X"2C",X"97",X"4C",X"EC",X"A1",X"DD",X"2F",X"DD",X"4F",X"A6",X"A0",X"97",X"34",X"97",
		X"54",X"EC",X"A4",X"DD",X"37",X"DD",X"57",X"CC",X"00",X"00",X"DD",X"1D",X"DD",X"25",X"DD",X"2D",
		X"DD",X"35",X"DD",X"3D",X"DD",X"45",X"DD",X"4D",X"DD",X"55",X"7E",X"DE",X"4A",X"10",X"83",X"FF",
		X"F8",X"27",X"15",X"31",X"A9",X"00",X"0F",X"10",X"9F",X"12",X"31",X"22",X"DD",X"08",X"EC",X"A1",
		X"DD",X"1F",X"44",X"56",X"DD",X"57",X"20",X"15",X"31",X"A9",X"00",X"11",X"EC",X"A1",X"DD",X"08",
		X"10",X"9F",X"12",X"EC",X"A1",X"DD",X"1F",X"EC",X"A9",X"00",X"0D",X"DD",X"57",X"A6",X"A0",X"97",
		X"24",X"97",X"2C",X"EC",X"A1",X"DD",X"27",X"EC",X"A1",X"DD",X"2F",X"EC",X"A1",X"DD",X"37",X"EC",
		X"A1",X"DD",X"3F",X"EC",X"A1",X"DD",X"47",X"86",X"C5",X"97",X"1C",X"97",X"54",X"86",X"D6",X"97",
		X"34",X"97",X"3C",X"97",X"44",X"7E",X"DE",X"4A",X"00",X"08",X"00",X"35",X"00",X"0A",X"00",X"55",
		X"00",X"0C",X"00",X"75",X"00",X"0E",X"00",X"95",X"00",X"10",X"00",X"B5",X"00",X"12",X"00",X"03",
		X"00",X"14",X"00",X"04",X"00",X"16",X"00",X"05",X"00",X"18",X"00",X"06",X"00",X"1A",X"00",X"07",
		X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",
		X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"F5",X"14",X"E9",X"61",X"E3",X"DA",X"EE",X"FA",
		X"E1",X"AA",X"E1",X"BA",X"E1",X"CA",X"E1",X"DA",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",
		X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",
		X"E1",X"EA",X"E1",X"FA",X"E2",X"0A",X"E2",X"1A",X"E2",X"2A",X"E2",X"3A",X"E1",X"9A",X"E1",X"9A",
		X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",
		X"E2",X"4A",X"E2",X"5A",X"E2",X"6A",X"E2",X"7A",X"E2",X"8A",X"E2",X"9A",X"E2",X"AA",X"E2",X"BA",
		X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",X"E1",X"9A",
		X"E2",X"CA",X"E2",X"DA",X"E2",X"EA",X"E2",X"FA",X"E3",X"0A",X"E3",X"1A",X"E3",X"2A",X"E3",X"3A",
		X"E3",X"4A",X"E3",X"5A",X"E3",X"6A",X"E3",X"7A",X"E3",X"8A",X"0F",X"F8",X"C1",X"00",X"00",X"C1",
		X"00",X"00",X"C1",X"00",X"00",X"C1",X"00",X"00",X"E1",X"9A",X"00",X"90",X"C0",X"F8",X"40",X"CB",
		X"01",X"50",X"C2",X"02",X"00",X"C2",X"00",X"02",X"E1",X"AA",X"00",X"70",X"C0",X"F4",X"40",X"CB",
		X"01",X"40",X"C2",X"02",X"00",X"C2",X"00",X"02",X"E1",X"BA",X"00",X"50",X"C0",X"F0",X"40",X"CB",
		X"01",X"40",X"C2",X"02",X"00",X"C2",X"00",X"02",X"E1",X"CA",X"00",X"30",X"C0",X"EC",X"40",X"CB",
		X"01",X"60",X"C2",X"02",X"30",X"C2",X"00",X"02",X"E1",X"DA",X"00",X"90",X"C0",X"01",X"60",X"CB",
		X"01",X"60",X"CD",X"06",X"20",X"C2",X"00",X"02",X"E1",X"EA",X"00",X"58",X"C0",X"02",X"60",X"CB",
		X"01",X"60",X"CD",X"06",X"20",X"C2",X"00",X"02",X"E1",X"FA",X"00",X"38",X"C0",X"04",X"60",X"CB",
		X"01",X"60",X"CD",X"06",X"20",X"C2",X"00",X"02",X"E2",X"0A",X"00",X"28",X"C0",X"08",X"60",X"CB",
		X"01",X"60",X"CD",X"06",X"20",X"C2",X"00",X"02",X"E2",X"1A",X"00",X"20",X"C0",X"FB",X"00",X"CB",
		X"04",X"00",X"C2",X"FF",X"FB",X"C2",X"00",X"04",X"E2",X"2A",X"00",X"20",X"C0",X"FB",X"00",X"CB",
		X"02",X"00",X"C2",X"FF",X"F6",X"C2",X"00",X"02",X"E2",X"3A",X"00",X"C0",X"C8",X"90",X"00",X"D4",
		X"30",X"22",X"C2",X"FF",X"00",X"C2",X"01",X"40",X"00",X"00",X"00",X"A0",X"C8",X"20",X"00",X"D4",
		X"04",X"09",X"C2",X"00",X"00",X"C2",X"01",X"90",X"00",X"00",X"01",X"90",X"C8",X"8F",X"E0",X"D4",
		X"01",X"00",X"C2",X"00",X"00",X"C2",X"00",X"A0",X"00",X"00",X"02",X"80",X"C1",X"06",X"0B",X"C1",
		X"03",X"20",X"C1",X"00",X"00",X"C2",X"00",X"60",X"00",X"00",X"00",X"C0",X"C8",X"A0",X"00",X"D4",
		X"08",X"40",X"C2",X"FF",X"1F",X"C2",X"01",X"40",X"00",X"00",X"01",X"90",X"C8",X"A0",X"00",X"D4",
		X"33",X"12",X"C2",X"FE",X"7F",X"C2",X"00",X"A0",X"00",X"00",X"00",X"C0",X"C8",X"FF",X"00",X"D4",
		X"70",X"31",X"C2",X"FF",X"7F",X"C2",X"01",X"40",X"00",X"00",X"01",X"90",X"C8",X"F0",X"00",X"D4",
		X"10",X"10",X"C0",X"FF",X"FB",X"C2",X"00",X"A0",X"00",X"00",X"04",X"00",X"CA",X"A0",X"11",X"C1",
		X"21",X"43",X"C1",X"00",X"00",X"C2",X"00",X"40",X"00",X"00",X"04",X"00",X"CA",X"67",X"70",X"C8",
		X"E4",X"55",X"C1",X"00",X"00",X"C2",X"00",X"40",X"00",X"00",X"00",X"80",X"D0",X"AE",X"55",X"C5",
		X"08",X"55",X"C1",X"00",X"00",X"C2",X"02",X"00",X"00",X"00",X"00",X"80",X"C0",X"01",X"00",X"C1",
		X"00",X"40",X"C1",X"00",X"00",X"C2",X"02",X"00",X"00",X"00",X"04",X"00",X"C0",X"E0",X"00",X"C0",
		X"40",X"10",X"C1",X"00",X"00",X"C2",X"00",X"40",X"00",X"00",X"07",X"F8",X"C1",X"0F",X"A0",X"C1",
		X"00",X"00",X"C1",X"00",X"00",X"C2",X"00",X"04",X"00",X"00",X"04",X"00",X"C0",X"80",X"00",X"C6",
		X"00",X"10",X"C1",X"00",X"00",X"C2",X"00",X"40",X"00",X"00",X"04",X"00",X"C0",X"E0",X"00",X"C8",
		X"00",X"80",X"C1",X"00",X"00",X"C2",X"00",X"40",X"00",X"00",X"04",X"00",X"C0",X"E0",X"00",X"C8",
		X"00",X"04",X"C1",X"00",X"00",X"C2",X"00",X"40",X"00",X"00",X"02",X"00",X"C0",X"FC",X"00",X"C1",
		X"00",X"20",X"C1",X"00",X"00",X"C2",X"00",X"80",X"00",X"00",X"02",X"00",X"C0",X"00",X"00",X"C1",
		X"00",X"A0",X"C1",X"00",X"00",X"C2",X"00",X"80",X"00",X"00",X"02",X"00",X"C0",X"01",X"40",X"C0",
		X"74",X"0A",X"C6",X"00",X"10",X"C2",X"00",X"80",X"00",X"00",X"02",X"00",X"C0",X"F9",X"12",X"C0",
		X"20",X"0F",X"C6",X"00",X"10",X"C2",X"00",X"80",X"00",X"00",X"20",X"20",X"44",X"45",X"4D",X"4F",
		X"20",X"42",X"55",X"59",X"49",X"4E",X"2C",X"20",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",
		X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"2C",X"20",X"4E",X"45",X"49",X"4C",X"20",X"46",X"41",
		X"4C",X"43",X"4F",X"4E",X"45",X"52",X"20",X"46",X"4F",X"52",X"20",X"42",X"41",X"4C",X"4C",X"59",
		X"20",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"20",X"20",X"02",X"C0",X"03",X"BA",X"D6",X"0F",
		X"03",X"0E",X"C9",X"03",X"BA",X"05",X"94",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",
		X"0E",X"C9",X"00",X"00",X"05",X"94",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",
		X"C9",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"03",
		X"BA",X"06",X"44",X"07",X"72",X"02",X"C0",X"00",X"00",X"D7",X"0F",X"03",X"0E",X"C9",X"00",X"00",
		X"06",X"44",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D8",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"00",
		X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D9",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"14",X"08",X"13",X"BC",X"03",X"BA",X"06",X"A2",X"07",
		X"72",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"06",X"A2",X"00",X"00",
		X"02",X"C0",X"03",X"BA",X"D6",X"10",X"D8",X"10",X"98",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",
		X"C0",X"00",X"00",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"00",X"00",X"07",X"72",X"02",X"C0",
		X"03",X"84",X"D6",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"06",X"44",X"07",X"72",X"02",X"C0",X"00",
		X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"06",X"44",X"07",X"72",X"02",X"C0",X"03",X"52",
		X"D6",X"0D",X"5F",X"0D",X"2D",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",
		X"0D",X"5F",X"0D",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"0B",
		X"3D",X"0B",X"13",X"02",X"CA",X"04",X"2E",X"09",X"F2",X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",
		X"0B",X"13",X"00",X"00",X"04",X"2E",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",
		X"13",X"02",X"CA",X"00",X"00",X"08",X"5C",X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",
		X"00",X"00",X"00",X"00",X"08",X"5C",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",
		X"CA",X"04",X"B2",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",
		X"04",X"B2",X"07",X"72",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"00",
		X"00",X"06",X"A2",X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"00",X"00",
		X"06",X"A2",X"02",X"C0",X"02",X"CA",X"D6",X"0A",X"9C",X"0A",X"74",X"02",X"CA",X"04",X"F8",X"05",
		X"94",X"02",X"C0",X"00",X"00",X"D7",X"0A",X"05",X"09",X"DF",X"00",X"00",X"04",X"F8",X"05",X"94",
		X"02",X"C0",X"02",X"CA",X"D8",X"09",X"74",X"09",X"50",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",
		X"C0",X"00",X"00",X"D9",X"08",X"ED",X"08",X"CB",X"00",X"00",X"00",X"00",X"05",X"94",X"02",X"C0",
		X"02",X"F4",X"DA",X"08",X"6C",X"08",X"4C",X"02",X"CA",X"04",X"B2",X"05",X"94",X"02",X"C0",X"00",
		X"00",X"DB",X"07",X"F3",X"07",X"D5",X"00",X"00",X"04",X"B2",X"02",X"F4",X"02",X"C0",X"03",X"22",
		X"DC",X"07",X"80",X"07",X"64",X"02",X"CA",X"00",X"00",X"06",X"44",X"02",X"C0",X"00",X"00",X"DD",
		X"07",X"15",X"06",X"FB",X"00",X"00",X"00",X"00",X"06",X"A2",X"02",X"C0",X"03",X"BA",X"D6",X"0F",
		X"03",X"0E",X"C9",X"03",X"BA",X"05",X"94",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",
		X"0E",X"C9",X"00",X"00",X"05",X"94",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",
		X"C9",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"03",
		X"BA",X"06",X"44",X"07",X"72",X"02",X"C0",X"00",X"00",X"DB",X"0F",X"03",X"0E",X"C9",X"00",X"00",
		X"06",X"44",X"00",X"00",X"02",X"C0",X"03",X"BA",X"DC",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"00",
		X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"DD",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"16",X"7D",X"16",X"27",X"03",X"BA",X"06",X"A2",X"07",
		X"72",X"02",X"C0",X"00",X"00",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"06",X"A2",X"07",X"72",
		X"02",X"C0",X"03",X"BA",X"D6",X"14",X"08",X"13",X"BC",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",
		X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"07",X"72",X"02",X"C0",
		X"03",X"84",X"D6",X"10",X"D8",X"10",X"98",X"03",X"BA",X"06",X"44",X"07",X"72",X"02",X"C0",X"00",
		X"00",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"06",X"44",X"07",X"72",X"02",X"C0",X"03",X"52",
		X"D6",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",
		X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"0D",
		X"5F",X"0D",X"2D",X"02",X"CA",X"04",X"2E",X"0B",X"28",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",
		X"0D",X"2D",X"00",X"00",X"04",X"2E",X"0B",X"28",X"02",X"C0",X"02",X"CA",X"D6",X"0D",X"5F",X"0D",
		X"2D",X"02",X"CA",X"00",X"00",X"09",X"F2",X"02",X"C0",X"00",X"00",X"D6",X"0E",X"2B",X"0D",X"F5",
		X"00",X"00",X"00",X"00",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"D7",X"0F",X"03",X"0E",X"C9",X"02",
		X"CA",X"04",X"B2",X"08",X"5C",X"02",X"C0",X"00",X"00",X"D8",X"0F",X"E6",X"0F",X"AA",X"00",X"00",
		X"04",X"B2",X"08",X"5C",X"02",X"C0",X"02",X"CA",X"D9",X"10",X"D8",X"10",X"98",X"02",X"CA",X"00",
		X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"DA",X"11",X"DA",X"11",X"96",X"00",X"00",X"00",X"00",
		X"07",X"72",X"02",X"C0",X"02",X"CA",X"D6",X"1E",X"06",X"1D",X"92",X"02",X"CA",X"04",X"F8",X"06",
		X"A2",X"02",X"C0",X"00",X"00",X"D6",X"1C",X"54",X"1B",X"E8",X"00",X"00",X"02",X"7C",X"07",X"08",
		X"02",X"C0",X"02",X"CA",X"D6",X"1A",X"BD",X"1A",X"57",X"02",X"CA",X"00",X"00",X"06",X"A2",X"02",
		X"C0",X"00",X"00",X"D6",X"19",X"3E",X"18",X"DE",X"00",X"00",X"00",X"00",X"06",X"44",X"02",X"C0",
		X"02",X"CA",X"D6",X"17",X"D4",X"17",X"78",X"02",X"CA",X"04",X"B2",X"05",X"EA",X"02",X"C0",X"00",
		X"00",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"04",X"B2",X"05",X"94",X"02",X"C0",X"02",X"CA",
		X"D6",X"15",X"3B",X"14",X"E9",X"02",X"CA",X"00",X"00",X"05",X"44",X"02",X"C0",X"00",X"00",X"D6",
		X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"04",X"F8",X"02",X"C0",X"04",X"2E",X"D6",X"16",
		X"7D",X"16",X"27",X"04",X"2E",X"06",X"44",X"08",X"5C",X"02",X"C0",X"00",X"00",X"D6",X"1A",X"BD",
		X"1A",X"57",X"00",X"00",X"06",X"44",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"1E",X"06",X"1D",
		X"92",X"04",X"2E",X"00",X"00",X"08",X"5C",X"02",X"C0",X"00",X"00",X"D6",X"1A",X"BD",X"1A",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"16",X"7D",X"16",X"27",X"04",
		X"2E",X"07",X"08",X"0B",X"28",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",
		X"07",X"08",X"0D",X"46",X"02",X"C0",X"04",X"2E",X"D6",X"16",X"7D",X"16",X"27",X"04",X"2E",X"00",
		X"00",X"0E",X"E6",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",
		X"0D",X"46",X"02",X"C0",X"04",X"2E",X"D6",X"10",X"D8",X"10",X"98",X"04",X"2E",X"07",X"72",X"0B",
		X"28",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"07",X"72",X"09",X"F2",
		X"02",X"C0",X"04",X"2E",X"D6",X"0D",X"5F",X"0D",X"2D",X"04",X"2E",X"00",X"00",X"0B",X"28",X"02",
		X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"09",X"F2",X"02",X"C0",
		X"04",X"2E",X"D6",X"10",X"D8",X"10",X"98",X"04",X"2E",X"07",X"08",X"08",X"5C",X"02",X"C0",X"00",
		X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"07",X"08",X"07",X"72",X"02",X"C0",X"04",X"2E",
		X"D6",X"0D",X"5F",X"0D",X"2D",X"04",X"2E",X"00",X"00",X"06",X"A2",X"02",X"C0",X"00",X"00",X"D6",
		X"0B",X"3D",X"0B",X"13",X"00",X"00",X"00",X"00",X"05",X"94",X"02",X"C0",X"02",X"CA",X"D6",X"15",
		X"3B",X"14",X"E9",X"0A",X"88",X"08",X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"D6",X"16",X"7D",
		X"16",X"27",X"0B",X"28",X"08",X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"D7",X"16",X"7D",X"16",
		X"27",X"0B",X"28",X"08",X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"D8",X"16",X"7D",X"16",X"27",
		X"0B",X"28",X"08",X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"D9",X"16",X"7D",X"16",X"27",X"0B",
		X"28",X"08",X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"DA",X"16",X"7D",X"16",X"27",X"0B",X"28",
		X"08",X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"DB",X"16",X"7D",X"16",X"27",X"00",X"00",X"08",
		X"5C",X"09",X"F2",X"02",X"C0",X"02",X"CA",X"DC",X"16",X"7D",X"16",X"27",X"00",X"00",X"08",X"5C",
		X"00",X"00",X"02",X"C0",X"02",X"CA",X"DD",X"16",X"7D",X"16",X"27",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"00",X"00",X"D6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"44",X"45",X"4D",X"4F",X"20",X"53",X"54",X"41",X"52",X"54",X"2C",X"20",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"2C",X"20",
		X"4E",X"45",X"49",X"4C",X"20",X"46",X"41",X"4C",X"43",X"4F",X"4E",X"45",X"52",X"20",X"46",X"4F",
		X"52",X"20",X"42",X"41",X"4C",X"4C",X"59",X"20",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"20",
		X"20",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"04",X"2E",X"05",X"94",
		X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"04",X"2E",X"00",X"00",X"02",
		X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",
		X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",
		X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"04",X"B2",X"05",X"94",X"02",X"C0",X"00",X"00",
		X"DB",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"04",X"B2",X"00",X"00",X"02",X"C0",X"02",X"CA",X"DC",
		X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",X"00",X"00",X"DD",X"0B",
		X"3D",X"0B",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"16",X"7D",
		X"16",X"27",X"02",X"CA",X"04",X"F8",X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"16",X"7D",X"16",
		X"27",X"00",X"00",X"04",X"F8",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"14",X"08",X"13",X"BC",
		X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"52",X"D6",X"10",X"D8",X"10",X"98",X"03",X"52",
		X"04",X"B2",X"06",X"A2",X"02",X"C0",X"00",X"00",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"04",
		X"B2",X"00",X"00",X"02",X"C0",X"03",X"84",X"D6",X"0D",X"5F",X"0D",X"2D",X"03",X"84",X"00",X"00",
		X"07",X"08",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",X"0D",X"2D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"05",X"94",X"07",X"72",
		X"02",X"C0",X"00",X"00",X"D6",X"0E",X"2B",X"0D",X"F5",X"00",X"00",X"05",X"94",X"00",X"00",X"02",
		X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",
		X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",
		X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"06",X"44",X"07",X"72",X"02",X"C0",X"00",X"00",
		X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"06",X"44",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D7",
		X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D8",X"0E",
		X"2B",X"0D",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"10",X"D8",
		X"10",X"98",X"03",X"BA",X"06",X"A2",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"10",X"D8",X"10",
		X"98",X"00",X"00",X"06",X"A2",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0D",X"5F",X"0D",X"2D",
		X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",X"0D",X"2D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"84",X"D6",X"0B",X"3D",X"0B",X"13",X"03",X"BA",
		X"06",X"44",X"07",X"08",X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"06",
		X"44",X"00",X"00",X"02",X"C0",X"03",X"52",X"D6",X"0A",X"05",X"09",X"DF",X"03",X"BA",X"00",X"00",
		X"06",X"A2",X"02",X"C0",X"00",X"00",X"D6",X"0A",X"05",X"09",X"DF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"04",X"2E",X"05",X"94",
		X"02",X"C0",X"00",X"00",X"D6",X"0A",X"9C",X"0A",X"74",X"00",X"00",X"04",X"2E",X"00",X"00",X"02",
		X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",
		X"00",X"00",X"D6",X"0A",X"05",X"09",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",
		X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"04",X"B2",X"05",X"94",X"02",X"C0",X"00",X"00",
		X"D6",X"09",X"74",X"09",X"50",X"00",X"00",X"04",X"B2",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",
		X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"08",
		X"ED",X"08",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"1A",X"BD",
		X"1A",X"57",X"02",X"CA",X"04",X"F8",X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"1A",X"BD",X"1A",
		X"57",X"00",X"00",X"04",X"F8",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"16",X"7D",X"16",X"27",
		X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"16",X"7D",X"16",X"27",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"14",X"08",X"13",X"BC",X"02",X"CA",
		X"04",X"B2",X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"04",
		X"B2",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"0D",X"5F",X"0D",X"2D",X"02",X"CA",X"00",X"00",
		X"05",X"94",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",X"0D",X"2D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"03",X"BA",X"D6",X"16",X"7D",X"16",X"27",X"03",X"BA",X"05",X"94",X"07",X"72",
		X"02",X"C0",X"00",X"00",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"05",X"94",X"00",X"00",X"02",
		X"C0",X"03",X"BA",X"D6",X"14",X"08",X"13",X"BC",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",
		X"00",X"00",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",
		X"BA",X"D6",X"10",X"D8",X"10",X"98",X"03",X"BA",X"06",X"44",X"07",X"72",X"02",X"C0",X"00",X"00",
		X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"06",X"44",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",
		X"0F",X"03",X"0E",X"C9",X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"0F",
		X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"14",X"08",
		X"13",X"BC",X"03",X"BA",X"06",X"A2",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",X"13",
		X"BC",X"00",X"00",X"06",X"A2",X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"16",X"7D",X"16",X"27",
		X"03",X"BA",X"00",X"00",X"07",X"72",X"02",X"C0",X"00",X"00",X"D6",X"16",X"7D",X"16",X"27",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"84",X"D6",X"10",X"D8",X"10",X"98",X"03",X"84",
		X"06",X"44",X"07",X"08",X"02",X"C0",X"00",X"00",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"06",
		X"44",X"00",X"00",X"02",X"C0",X"03",X"52",X"D6",X"0A",X"05",X"09",X"DF",X"03",X"52",X"00",X"00",
		X"06",X"A2",X"02",X"C0",X"00",X"00",X"D6",X"0A",X"05",X"09",X"DF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"04",X"2E",X"05",X"94",
		X"02",X"C0",X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"04",X"2E",X"00",X"00",X"02",
		X"C0",X"02",X"CA",X"D6",X"0B",X"3D",X"0B",X"13",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",
		X"00",X"00",X"D6",X"0B",X"3D",X"0B",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",
		X"CA",X"D6",X"0B",X"E9",X"0B",X"BB",X"02",X"CA",X"04",X"B2",X"05",X"94",X"02",X"C0",X"00",X"00",
		X"D7",X"0C",X"9E",X"0C",X"6E",X"00",X"00",X"04",X"B2",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D8",
		X"0D",X"5F",X"0D",X"2D",X"02",X"CA",X"00",X"00",X"05",X"94",X"02",X"C0",X"00",X"00",X"DD",X"0D",
		X"5F",X"0D",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"F8",X"D6",X"1A",X"BD",
		X"1A",X"57",X"04",X"F8",X"04",X"F8",X"09",X"F2",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",X"0D",
		X"2D",X"00",X"00",X"04",X"F8",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"19",X"3E",X"18",X"DE",
		X"04",X"2E",X"00",X"00",X"08",X"5C",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"03",X"52",X"D6",X"16",X"7D",X"16",X"27",X"03",X"52",
		X"04",X"B2",X"06",X"A2",X"02",X"C0",X"00",X"00",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"04",
		X"B2",X"00",X"00",X"02",X"C0",X"03",X"22",X"D6",X"14",X"08",X"13",X"BC",X"03",X"22",X"00",X"00",
		X"06",X"44",X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"F8",X"02",X"C0",X"02",X"CA",X"D6",X"16",X"7D",X"16",X"27",X"0D",X"46",X"07",X"08",
		X"0B",X"28",X"09",X"F2",X"FF",X"F8",X"02",X"C0",X"02",X"CA",X"D7",X"16",X"7D",X"16",X"27",X"0D",
		X"46",X"07",X"08",X"0B",X"28",X"09",X"F2",X"FF",X"F8",X"02",X"C0",X"02",X"CA",X"D8",X"16",X"7D",
		X"16",X"27",X"0D",X"46",X"07",X"08",X"0B",X"28",X"09",X"F2",X"FF",X"F8",X"02",X"C0",X"02",X"CA",
		X"D9",X"16",X"7D",X"16",X"27",X"0D",X"46",X"07",X"08",X"0B",X"28",X"09",X"F2",X"FF",X"F8",X"02",
		X"C0",X"02",X"CA",X"DA",X"16",X"7D",X"16",X"27",X"0D",X"46",X"07",X"08",X"0B",X"28",X"09",X"F2",
		X"FF",X"F8",X"02",X"C0",X"02",X"CA",X"DB",X"16",X"7D",X"16",X"27",X"00",X"00",X"07",X"08",X"0B",
		X"28",X"09",X"F2",X"FF",X"F8",X"02",X"C0",X"02",X"CA",X"DC",X"16",X"7D",X"16",X"27",X"00",X"00",
		X"07",X"08",X"00",X"00",X"00",X"00",X"FF",X"F8",X"02",X"C0",X"02",X"CA",X"DD",X"16",X"7D",X"16",
		X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"00",X"00",X"D6",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"44",X"45",X"4D",X"4F",
		X"20",X"54",X"52",X"4F",X"50",X"48",X"59",X"2C",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",
		X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"2C",X"20",X"4E",X"45",X"49",X"4C",X"20",X"46",X"41",
		X"4C",X"43",X"4F",X"4E",X"45",X"52",X"20",X"46",X"4F",X"52",X"20",X"42",X"41",X"4C",X"4C",X"59",
		X"20",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"20",X"20",X"02",X"C0",X"02",X"CA",X"D6",X"05",
		X"9E",X"05",X"8A",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"02",X"CA",X"D6",X"05",X"9E",
		X"05",X"8A",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",X"05",X"9E",X"05",
		X"8A",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",X"05",X"9E",X"05",X"8A",
		X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"02",X"CA",X"D6",X"05",X"4E",X"05",X"3A",X"06",
		X"A2",X"09",X"62",X"0C",X"86",X"02",X"C0",X"02",X"CA",X"D6",X"05",X"01",X"04",X"EF",X"06",X"44",
		X"08",X"DC",X"0B",X"D2",X"02",X"C0",X"03",X"84",X"D6",X"04",X"BB",X"04",X"A9",X"05",X"EA",X"08",
		X"5C",X"0B",X"28",X"02",X"C0",X"03",X"84",X"D6",X"04",X"76",X"04",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"04",X"36",X"04",X"26",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"04",X"2E",X"D6",X"04",X"36",X"04",X"26",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"C0",X"04",X"B2",X"DC",X"04",X"36",X"04",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"C0",X"04",X"B2",X"DD",X"04",X"36",X"04",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",
		X"04",X"F8",X"D6",X"0F",X"E6",X"0F",X"AA",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"04",
		X"F8",X"D6",X"10",X"D8",X"10",X"98",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"00",X"00",
		X"D6",X"10",X"D8",X"10",X"98",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"00",X"00",X"D6",
		X"10",X"D8",X"10",X"98",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"04",X"F8",X"D6",X"14",
		X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",
		X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"F8",X"D6",X"0F",X"03",X"0E",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"F8",X"D6",X"0F",X"03",X"0E",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"B2",X"D6",X"10",X"D8",X"10",X"98",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"B2",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"0E",
		X"E6",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"0E",X"E6",
		X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"0E",X"E6",X"02",
		X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"0E",X"E6",X"02",X"C0",
		X"03",X"BA",X"D6",X"0E",X"2B",X"0D",X"F5",X"08",X"DC",X"0A",X"88",X"0E",X"10",X"02",X"C0",X"03",
		X"BA",X"D6",X"0D",X"5F",X"0D",X"2D",X"08",X"5C",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"04",X"B2",
		X"D6",X"0C",X"9E",X"0C",X"6E",X"07",X"E4",X"09",X"62",X"0C",X"86",X"02",X"C0",X"04",X"B2",X"D9",
		X"0B",X"E9",X"0B",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"DA",X"0B",
		X"3D",X"0B",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"DB",X"0B",X"3D",
		X"0B",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",X"44",X"DC",X"0B",X"3D",X"0B",
		X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",X"44",X"DD",X"0B",X"3D",X"0B",X"13",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",X"A2",X"D6",X"16",X"7D",X"16",X"27",X"09",
		X"62",X"0B",X"28",X"0D",X"46",X"02",X"C0",X"06",X"A2",X"D6",X"16",X"7D",X"16",X"27",X"09",X"62",
		X"0B",X"28",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",X"1A",X"BD",X"1A",X"57",X"09",X"62",X"0B",
		X"28",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",X"1A",X"BD",X"1A",X"57",X"09",X"62",X"0B",X"28",
		X"0D",X"46",X"02",X"C0",X"06",X"A2",X"D6",X"19",X"3E",X"18",X"DE",X"00",X"00",X"00",X"00",X"0C",
		X"86",X"02",X"C0",X"00",X"00",X"D6",X"19",X"3E",X"18",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"C0",X"06",X"A2",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"C0",X"06",X"A2",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",
		X"06",X"44",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",
		X"44",X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",
		X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"D6",
		X"10",X"D8",X"10",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"0D",
		X"5F",X"0D",X"2D",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"02",X"CA",X"D6",X"0D",X"5F",
		X"0D",X"2D",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",X"0D",
		X"2D",X"07",X"08",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"00",X"00",X"D6",X"0D",X"5F",X"0D",X"2D",
		X"06",X"A2",X"09",X"F2",X"0B",X"28",X"02",X"C0",X"02",X"CA",X"D6",X"0C",X"9E",X"0C",X"6E",X"06",
		X"44",X"09",X"62",X"0A",X"88",X"02",X"C0",X"02",X"CA",X"D6",X"0B",X"E9",X"0B",X"BB",X"05",X"EA",
		X"08",X"DC",X"09",X"F2",X"02",X"C0",X"03",X"84",X"D6",X"0B",X"3D",X"0B",X"13",X"05",X"94",X"08",
		X"5C",X"09",X"62",X"02",X"C0",X"03",X"84",X"D6",X"0B",X"E9",X"0B",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"0C",X"9E",X"0C",X"6E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"C0",X"04",X"2E",X"D7",X"0D",X"5F",X"0D",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"C0",X"04",X"B2",X"D8",X"0E",X"2B",X"0D",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"C0",X"04",X"B2",X"D9",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",
		X"04",X"F8",X"D6",X"15",X"3B",X"14",X"E9",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"04",
		X"F8",X"D6",X"16",X"7D",X"16",X"27",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"00",X"00",
		X"D6",X"16",X"7D",X"16",X"27",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",
		X"16",X"7D",X"16",X"27",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"04",X"F8",X"D6",X"14",
		X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"00",X"00",X"D6",X"14",X"08",
		X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"D6",X"0F",X"03",X"0E",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"D6",X"0F",X"03",X"0E",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"F8",X"D6",X"10",X"D8",X"10",X"98",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"F8",X"D6",X"10",X"D8",X"10",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"0D",X"5F",X"0D",X"2D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"C0",X"04",X"2E",X"D6",X"0D",X"5F",X"0D",X"2D",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"C0",X"03",X"BA",X"D6",X"0E",X"2B",X"0D",X"F5",X"09",X"62",X"0B",X"28",X"07",
		X"72",X"02",X"C0",X"03",X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"07",X"72",
		X"02",X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"07",X"72",X"02",
		X"C0",X"00",X"00",X"D6",X"0F",X"03",X"0E",X"C9",X"09",X"62",X"0B",X"28",X"07",X"72",X"02",X"C0",
		X"03",X"BA",X"D6",X"0E",X"2B",X"0D",X"F5",X"00",X"00",X"00",X"00",X"07",X"08",X"02",X"C0",X"03",
		X"BA",X"D6",X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"B2",
		X"D6",X"0E",X"2B",X"0D",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"04",X"B2",X"D6",
		X"0F",X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"D6",X"0F",
		X"03",X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"DB",X"0F",X"03",
		X"0E",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",X"44",X"DC",X"0F",X"03",X"0E",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",X"44",X"DD",X"0F",X"03",X"0E",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",X"A2",X"D6",X"1F",X"CD",X"1F",X"53",X"09",
		X"62",X"0B",X"28",X"0D",X"46",X"02",X"C0",X"06",X"A2",X"D6",X"21",X"B3",X"21",X"31",X"09",X"62",
		X"0B",X"28",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",X"1E",X"06",X"1D",X"92",X"09",X"62",X"0B",
		X"28",X"0D",X"46",X"02",X"C0",X"00",X"00",X"D6",X"1E",X"06",X"1D",X"92",X"09",X"62",X"0B",X"28",
		X"0D",X"46",X"02",X"C0",X"06",X"A2",X"D6",X"1A",X"BD",X"1A",X"57",X"08",X"DC",X"0A",X"88",X"0C",
		X"86",X"02",X"C0",X"00",X"00",X"D6",X"1A",X"BD",X"1A",X"57",X"08",X"5C",X"09",X"F2",X"0B",X"D2",
		X"02",X"C0",X"07",X"72",X"D6",X"1E",X"06",X"1D",X"92",X"07",X"E4",X"09",X"62",X"0B",X"28",X"02",
		X"C0",X"07",X"72",X"D6",X"1A",X"BD",X"1A",X"57",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",
		X"06",X"A2",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"06",
		X"A2",X"D6",X"16",X"7D",X"16",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",
		X"D6",X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"05",X"94",X"D6",
		X"14",X"08",X"13",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"02",X"CA",X"D6",X"15",
		X"3B",X"14",X"E9",X"07",X"08",X"09",X"F2",X"0D",X"46",X"16",X"00",X"02",X"CA",X"D6",X"16",X"7D",
		X"16",X"27",X"07",X"08",X"09",X"F2",X"0D",X"46",X"02",X"C0",X"02",X"A2",X"D6",X"15",X"3B",X"14",
		X"E9",X"06",X"A2",X"09",X"62",X"0C",X"86",X"02",X"C0",X"02",X"7C",X"D6",X"14",X"08",X"13",X"BC",
		X"06",X"44",X"08",X"DC",X"0B",X"D2",X"02",X"C0",X"02",X"58",X"D6",X"12",X"E8",X"12",X"A0",X"05",
		X"EA",X"08",X"5C",X"0B",X"28",X"02",X"C0",X"02",X"36",X"D6",X"11",X"DA",X"11",X"96",X"05",X"94",
		X"07",X"E4",X"0A",X"88",X"02",X"C0",X"02",X"18",X"D6",X"10",X"D8",X"10",X"98",X"06",X"44",X"07",
		X"72",X"09",X"F2",X"02",X"C0",X"00",X"00",X"D6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"02",X"36",X"D6",X"08",X"ED",X"08",X"CB",X"04",X"6E",X"04",
		X"6E",X"04",X"6E",X"05",X"80",X"00",X"00",X"D6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"80",X"02",X"7C",X"D6",X"0A",X"05",X"09",X"DF",X"04",X"F8",X"04",X"F8",X"04",
		X"F8",X"0B",X"00",X"02",X"A2",X"D6",X"0A",X"9C",X"0A",X"74",X"05",X"44",X"05",X"44",X"05",X"44",
		X"0B",X"00",X"02",X"36",X"D6",X"08",X"ED",X"08",X"CB",X"04",X"6E",X"04",X"6E",X"04",X"6E",X"02",
		X"C0",X"00",X"00",X"D6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"2C",X"20",
		X"42",X"41",X"4C",X"4C",X"59",X"20",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"4D",X"46",X"47",
		X"2E",X"20",X"43",X"4F",X"2E",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",
		X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"D5",X"41",X"35",X"39",X"2D",X"30",X"58",
		X"58",X"2D",X"55",X"34",X"20",X"20",X"00",X"00",X"FF",X"34",X"76",X"B6",X"60",X"00",X"F6",X"60",
		X"01",X"C4",X"0F",X"34",X"04",X"86",X"3E",X"B7",X"60",X"02",X"B6",X"60",X"02",X"2A",X"FB",X"B6",
		X"60",X"01",X"F6",X"60",X"00",X"C6",X"3D",X"F7",X"60",X"02",X"48",X"48",X"48",X"48",X"AB",X"E0",
		X"27",X"7E",X"81",X"4D",X"10",X"24",X"03",X"4B",X"8E",X"E1",X"00",X"10",X"8E",X"00",X"1C",X"1F",
		X"89",X"81",X"03",X"23",X"55",X"81",X"0C",X"10",X"25",X"03",X"38",X"81",X"10",X"10",X"25",X"01",
		X"27",X"0D",X"02",X"27",X"0D",X"81",X"44",X"27",X"07",X"81",X"45",X"27",X"03",X"7E",X"F9",X"33",
		X"0F",X"02",X"58",X"3A",X"AE",X"84",X"81",X"14",X"10",X"25",X"01",X"72",X"81",X"20",X"10",X"25",
		X"03",X"11",X"81",X"24",X"10",X"25",X"01",X"BD",X"81",X"30",X"10",X"25",X"03",X"05",X"81",X"38",
		X"25",X"0F",X"81",X"40",X"10",X"25",X"02",X"FB",X"81",X"4D",X"10",X"25",X"01",X"FA",X"7E",X"F9",
		X"33",X"81",X"34",X"10",X"25",X"02",X"A1",X"16",X"02",X"AC",X"10",X"27",X"01",X"37",X"0D",X"02",
		X"10",X"26",X"02",X"DF",X"81",X"02",X"10",X"27",X"01",X"87",X"81",X"01",X"10",X"27",X"01",X"2A",
		X"BE",X"E1",X"00",X"9F",X"12",X"9F",X"14",X"9F",X"16",X"9F",X"18",X"9F",X"1A",X"EC",X"81",X"DD",
		X"08",X"DD",X"0A",X"DD",X"0C",X"DD",X"0E",X"DD",X"10",X"A6",X"80",X"97",X"1C",X"97",X"3C",X"97",
		X"5C",X"97",X"7C",X"97",X"9C",X"EC",X"81",X"DD",X"1F",X"DD",X"3F",X"DD",X"5F",X"DD",X"7F",X"DD",
		X"9F",X"A6",X"80",X"97",X"24",X"97",X"44",X"97",X"64",X"97",X"84",X"97",X"A4",X"EC",X"81",X"DD",
		X"27",X"DD",X"47",X"DD",X"67",X"DD",X"87",X"DD",X"A7",X"A6",X"80",X"97",X"2C",X"97",X"4C",X"97",
		X"6C",X"97",X"8C",X"97",X"AC",X"EC",X"81",X"DD",X"2F",X"DD",X"4F",X"DD",X"6F",X"DD",X"8F",X"DD",
		X"AF",X"A6",X"80",X"97",X"34",X"97",X"54",X"97",X"74",X"97",X"94",X"97",X"B4",X"EC",X"81",X"DD",
		X"37",X"DD",X"57",X"DD",X"77",X"DD",X"97",X"DD",X"B7",X"CC",X"00",X"00",X"97",X"03",X"97",X"04",
		X"97",X"05",X"97",X"06",X"97",X"07",X"DD",X"1D",X"DD",X"25",X"DD",X"2D",X"DD",X"35",X"DD",X"3D",
		X"DD",X"45",X"DD",X"4D",X"DD",X"55",X"DD",X"5D",X"DD",X"65",X"DD",X"6D",X"DD",X"75",X"DD",X"7D",
		X"DD",X"85",X"DD",X"8D",X"DD",X"95",X"DD",X"9D",X"DD",X"A5",X"DD",X"AD",X"DD",X"B5",X"DD",X"3A",
		X"DD",X"5A",X"DD",X"7A",X"DD",X"9A",X"DD",X"BA",X"97",X"01",X"97",X"02",X"10",X"CE",X"04",X"00",
		X"FC",X"60",X"00",X"1C",X"EF",X"7E",X"DE",X"4A",X"C6",X"FF",X"D7",X"01",X"D7",X"02",X"97",X"03",
		X"1F",X"89",X"58",X"8E",X"E1",X"00",X"3A",X"AE",X"84",X"9F",X"12",X"EC",X"81",X"DD",X"08",X"EC",
		X"81",X"DD",X"1F",X"44",X"56",X"DD",X"57",X"A6",X"80",X"97",X"24",X"97",X"2C",X"EC",X"81",X"DD",
		X"27",X"EC",X"81",X"DD",X"2F",X"EC",X"81",X"DD",X"37",X"EC",X"81",X"DD",X"3F",X"EC",X"81",X"DD",
		X"47",X"86",X"C5",X"97",X"1C",X"97",X"54",X"86",X"D6",X"97",X"34",X"97",X"3C",X"97",X"44",X"CC",
		X"00",X"00",X"DD",X"1D",X"DD",X"25",X"DD",X"2D",X"DD",X"35",X"DD",X"3D",X"DD",X"45",X"DD",X"4D",
		X"DD",X"55",X"7E",X"F9",X"33",X"0F",X"02",X"7E",X"F9",X"33",X"4F",X"BE",X"E1",X"00",X"10",X"8E",
		X"00",X"1C",X"97",X"03",X"9F",X"12",X"EC",X"81",X"DD",X"08",X"0D",X"01",X"10",X"27",X"01",X"62",
		X"0F",X"01",X"BE",X"E1",X"00",X"9F",X"14",X"EC",X"81",X"DD",X"0A",X"A6",X"80",X"97",X"3C",X"EC",
		X"81",X"DD",X"3F",X"A6",X"80",X"97",X"44",X"EC",X"81",X"DD",X"47",X"A6",X"80",X"97",X"4C",X"EC",
		X"81",X"DD",X"4F",X"A6",X"80",X"97",X"54",X"EC",X"84",X"DD",X"57",X"CC",X"00",X"00",X"DD",X"3D",
		X"DD",X"45",X"DD",X"4D",X"DD",X"55",X"DD",X"5A",X"97",X"04",X"9E",X"12",X"30",X"02",X"16",X"01",
		X"21",X"4F",X"BE",X"E1",X"00",X"10",X"8E",X"00",X"3C",X"97",X"04",X"9F",X"14",X"EC",X"81",X"DD",
		X"0A",X"0D",X"01",X"10",X"27",X"01",X"0B",X"0F",X"01",X"BE",X"E1",X"00",X"9F",X"12",X"EC",X"81",
		X"DD",X"08",X"A6",X"80",X"97",X"1C",X"EC",X"81",X"DD",X"1F",X"A6",X"80",X"97",X"24",X"EC",X"81",
		X"DD",X"27",X"A6",X"80",X"97",X"2C",X"EC",X"81",X"DD",X"2F",X"A6",X"80",X"97",X"34",X"EC",X"84",
		X"DD",X"37",X"CC",X"00",X"00",X"DD",X"1D",X"DD",X"25",X"DD",X"2D",X"DD",X"35",X"DD",X"3A",X"97",
		X"03",X"9E",X"14",X"30",X"02",X"16",X"00",X"CA",X"0D",X"01",X"10",X"27",X"00",X"9C",X"97",X"05",
		X"9F",X"16",X"BE",X"E1",X"00",X"9F",X"12",X"9F",X"14",X"9F",X"18",X"9F",X"1A",X"EC",X"81",X"DD",
		X"08",X"DD",X"0A",X"DD",X"0E",X"DD",X"10",X"A6",X"80",X"97",X"1C",X"97",X"3C",X"97",X"7C",X"97",
		X"9C",X"EC",X"81",X"DD",X"1F",X"DD",X"3F",X"DD",X"7F",X"DD",X"9F",X"A6",X"80",X"97",X"24",X"97",
		X"44",X"97",X"84",X"97",X"A4",X"EC",X"81",X"DD",X"27",X"DD",X"47",X"DD",X"87",X"DD",X"A7",X"A6",
		X"80",X"97",X"2C",X"97",X"4C",X"97",X"8C",X"97",X"AC",X"EC",X"81",X"DD",X"2F",X"DD",X"4F",X"DD",
		X"8F",X"DD",X"AF",X"A6",X"80",X"97",X"34",X"97",X"54",X"97",X"94",X"97",X"B4",X"EC",X"81",X"DD",
		X"37",X"DD",X"57",X"DD",X"97",X"DD",X"B7",X"CC",X"00",X"00",X"97",X"03",X"97",X"04",X"97",X"06",
		X"97",X"07",X"DD",X"1D",X"DD",X"25",X"DD",X"2D",X"DD",X"35",X"DD",X"3D",X"DD",X"45",X"DD",X"4D",
		X"DD",X"55",X"DD",X"7D",X"DD",X"85",X"DD",X"8D",X"DD",X"95",X"DD",X"9D",X"DD",X"A5",X"DD",X"AD",
		X"DD",X"B5",X"97",X"01",X"97",X"02",X"96",X"05",X"9E",X"16",X"10",X"8E",X"00",X"5C",X"97",X"05",
		X"9F",X"16",X"EC",X"81",X"DD",X"0C",X"20",X"1A",X"10",X"8E",X"00",X"7C",X"97",X"06",X"9F",X"18",
		X"EC",X"81",X"DD",X"0E",X"20",X"0C",X"10",X"8E",X"00",X"9C",X"97",X"07",X"9F",X"1A",X"EC",X"81",
		X"DD",X"10",X"CE",X"00",X"00",X"A6",X"80",X"A7",X"A0",X"EF",X"A1",X"EC",X"81",X"ED",X"A4",X"31",
		X"25",X"A6",X"80",X"A7",X"A0",X"EF",X"A1",X"EC",X"81",X"ED",X"A4",X"31",X"25",X"A6",X"80",X"A7",
		X"A0",X"EF",X"A1",X"EC",X"81",X"ED",X"A4",X"31",X"25",X"A6",X"80",X"A7",X"A0",X"EF",X"A1",X"EC",
		X"81",X"ED",X"A4",X"35",X"76",X"3B",X"34",X"76",X"86",X"44",X"7E",X"F5",X"E0",X"CC",X"FF",X"C0",
		X"B7",X"60",X"00",X"CC",X"3D",X"34",X"FD",X"60",X"02",X"86",X"3C",X"B7",X"60",X"03",X"8E",X"F5",
		X"A9",X"E6",X"0C",X"27",X"11",X"C1",X"20",X"22",X"0B",X"4F",X"8E",X"E0",X"00",X"AB",X"84",X"30",
		X"01",X"26",X"FA",X"4C",X"26",X"FE",X"CC",X"FF",X"FF",X"83",X"00",X"01",X"26",X"FB",X"86",X"34",
		X"B7",X"60",X"03",X"CC",X"FF",X"FF",X"83",X"00",X"01",X"26",X"FB",X"86",X"3C",X"B7",X"60",X"03",
		X"8E",X"DE",X"3A",X"E6",X"0C",X"27",X"12",X"C1",X"20",X"22",X"0C",X"4F",X"8E",X"C0",X"00",X"AB",
		X"80",X"8C",X"E0",X"00",X"26",X"F9",X"4C",X"26",X"FE",X"CC",X"FF",X"FF",X"83",X"00",X"01",X"26",
		X"FB",X"86",X"34",X"B7",X"60",X"03",X"CC",X"FF",X"FF",X"83",X"00",X"01",X"26",X"FB",X"86",X"3C",
		X"B7",X"60",X"03",X"8E",X"04",X"00",X"86",X"80",X"A7",X"84",X"A1",X"84",X"26",X"FE",X"44",X"26",
		X"F7",X"A7",X"84",X"30",X"1F",X"8C",X"FF",X"FF",X"26",X"EC",X"CC",X"FF",X"FF",X"83",X"00",X"01",
		X"26",X"FB",X"86",X"34",X"B7",X"60",X"03",X"CC",X"FF",X"FF",X"83",X"00",X"01",X"26",X"FB",X"86",
		X"3C",X"B7",X"60",X"03",X"86",X"80",X"B7",X"60",X"00",X"B1",X"60",X"00",X"26",X"FE",X"44",X"26",
		X"F5",X"CC",X"FF",X"FF",X"83",X"00",X"01",X"26",X"FB",X"86",X"34",X"B7",X"60",X"03",X"86",X"3D",
		X"B7",X"60",X"02",X"8E",X"00",X"00",X"10",X"8E",X"04",X"00",X"CC",X"00",X"00",X"ED",X"81",X"31",
		X"3F",X"26",X"FA",X"12",X"BE",X"E1",X"00",X"9F",X"12",X"9F",X"14",X"9F",X"16",X"9F",X"18",X"9F",
		X"1A",X"EC",X"81",X"DD",X"08",X"DD",X"0A",X"DD",X"0C",X"DD",X"0E",X"DD",X"10",X"A6",X"80",X"97",
		X"1C",X"97",X"3C",X"97",X"5C",X"97",X"7C",X"97",X"9C",X"EC",X"81",X"DD",X"1F",X"DD",X"3F",X"DD",
		X"5F",X"DD",X"7F",X"DD",X"9F",X"A6",X"80",X"97",X"24",X"97",X"44",X"97",X"64",X"97",X"84",X"97",
		X"A4",X"EC",X"81",X"DD",X"27",X"DD",X"47",X"DD",X"67",X"DD",X"87",X"DD",X"A7",X"A6",X"80",X"97",
		X"2C",X"97",X"4C",X"97",X"6C",X"97",X"8C",X"97",X"AC",X"EC",X"81",X"DD",X"2F",X"DD",X"4F",X"DD",
		X"6F",X"DD",X"8F",X"DD",X"AF",X"A6",X"80",X"97",X"34",X"97",X"54",X"97",X"74",X"97",X"94",X"97",
		X"B4",X"EC",X"81",X"DD",X"37",X"DD",X"57",X"DD",X"77",X"DD",X"97",X"DD",X"B7",X"CC",X"00",X"00",
		X"DD",X"03",X"DD",X"04",X"DD",X"05",X"DD",X"06",X"DD",X"07",X"DD",X"1D",X"DD",X"25",X"DD",X"2D",
		X"DD",X"35",X"DD",X"3D",X"DD",X"45",X"DD",X"4D",X"DD",X"55",X"DD",X"5D",X"DD",X"65",X"DD",X"6D",
		X"DD",X"75",X"DD",X"7D",X"DD",X"85",X"DD",X"8D",X"DD",X"95",X"DD",X"9D",X"DD",X"A5",X"DD",X"AD",
		X"DD",X"B5",X"10",X"CE",X"04",X"00",X"FC",X"60",X"00",X"1C",X"EF",X"7E",X"DE",X"4A",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F9",X"35",X"F9",X"35",X"F9",X"35",X"F9",X"35",X"F5",X"B9",X"F9",X"35",X"F9",X"36",X"F9",X"3D");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
